

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO router 
  PIN localRouterAddress[3] 
    ANTENNAPARTIALMETALAREA 0.72 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.664 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 40.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 150.664 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.48 LAYER M3 ; 
    ANTENNAMAXAREACAR 205.109 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 763.537 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.5641 LAYER VL ;
  END localRouterAddress[3]
  PIN localRouterAddress[2] 
    ANTENNAPARTIALMETALAREA 8.68 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 32.264 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 53.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 198.912 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.48 LAYER M3 ; 
    ANTENNAMAXAREACAR 130.444 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 489.233 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.08333 LAYER VL ;
  END localRouterAddress[2]
  PIN localRouterAddress[1] 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 52.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 196.84 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.96 LAYER M3 ; 
    ANTENNAMAXAREACAR 150.315 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 554.524 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.78571 LAYER VL ;
  END localRouterAddress[1]
  PIN localRouterAddress[0] 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 65.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 244.2 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.96 LAYER M3 ; 
    ANTENNAMAXAREACAR 103.625 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 380.8 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.78571 LAYER VL ;
  END localRouterAddress[0]
  PIN destinationAddressIn_NORTH[11] 
    ANTENNAPARTIALMETALAREA 7.56 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 27.972 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 13.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 50.912 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3168 LAYER M3 ; 
    ANTENNAMAXAREACAR 185.32 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 701.63 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER VL ;
  END destinationAddressIn_NORTH[11]
  PIN destinationAddressIn_NORTH[10] 
    ANTENNAPARTIALMETALAREA 8.42 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 31.154 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 14.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 56.24 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3168 LAYER M3 ; 
    ANTENNAMAXAREACAR 184.867 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 696.141 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.5641 LAYER VL ;
  END destinationAddressIn_NORTH[10]
  PIN destinationAddressIn_NORTH[9] 
    ANTENNAPARTIALMETALAREA 2.42 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.954 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 24.62 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 92.278 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3264 LAYER M3 ; 
    ANTENNAMAXAREACAR 79.7879 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 300.702 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.28205 LAYER VL ;
  END destinationAddressIn_NORTH[9]
  PIN destinationAddressIn_NORTH[8] 
    ANTENNAPARTIALMETALAREA 9.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 33.966 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 29.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 111.888 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3264 LAYER M3 ; 
    ANTENNAMAXAREACAR 103.806 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 386.467 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.28205 LAYER VL ;
  END destinationAddressIn_NORTH[8]
  PIN destinationAddressIn_NORTH[7] 
    ANTENNAPARTIALMETALAREA 2.54 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.546 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 43.141 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 161.481 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END destinationAddressIn_NORTH[7]
  PIN destinationAddressIn_NORTH[6] 
    ANTENNAPARTIALMETALAREA 1.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.81 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.768 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 63.9744 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 240.936 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.28205 LAYER VL ;
  END destinationAddressIn_NORTH[6]
  PIN destinationAddressIn_NORTH[5] 
    ANTENNAPARTIALMETALAREA 2.34 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.658 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.06 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.07 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.6282 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 96.0192 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.28205 LAYER VL ;
  END destinationAddressIn_NORTH[5]
  PIN destinationAddressIn_NORTH[4] 
    ANTENNAPARTIALMETALAREA 2.82 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.434 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 47.6282 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 175.712 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END destinationAddressIn_NORTH[4]
  PIN destinationAddressIn_NORTH[3] 
    ANTENNAPARTIALMETALAREA 2.52 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.324 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 42.8205 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 157.923 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END destinationAddressIn_NORTH[3]
  PIN destinationAddressIn_NORTH[2] 
    ANTENNAPARTIALMETALAREA 2.58 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.546 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 43.7821 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 161.481 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END destinationAddressIn_NORTH[2]
  PIN destinationAddressIn_NORTH[1] 
    ANTENNAPARTIALMETALAREA 2.52 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.324 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 42.8205 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 157.923 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END destinationAddressIn_NORTH[1]
  PIN destinationAddressIn_NORTH[0] 
    ANTENNAPARTIALMETALAREA 2.62 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.694 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 44.4231 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 163.853 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END destinationAddressIn_NORTH[0]
  PIN requesterAddressIn_NORTH[3] 
    ANTENNAPARTIALMETALAREA 2.54 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.546 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 43.141 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 161.481 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END requesterAddressIn_NORTH[3]
  PIN requesterAddressIn_NORTH[2] 
    ANTENNAPARTIALMETALAREA 2.54 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.546 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 43.141 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 161.481 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END requesterAddressIn_NORTH[2]
  PIN requesterAddressIn_NORTH[1] 
    ANTENNAPARTIALMETALAREA 2.7 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.138 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 45.7051 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 170.968 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END requesterAddressIn_NORTH[1]
  PIN requesterAddressIn_NORTH[0] 
    ANTENNAPARTIALMETALAREA 2.42 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.954 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.14 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 59.8462 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 227.538 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.28205 LAYER VL ;
  END requesterAddressIn_NORTH[0]
  PIN dataIn_NORTH[5] 
    ANTENNAPARTIALMETALAREA 2.54 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.546 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 43.141 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 161.481 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END dataIn_NORTH[5]
  PIN dataIn_NORTH[4] 
    ANTENNAPARTIALMETALAREA 3.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.174 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 50.8333 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 187.571 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END dataIn_NORTH[4]
  PIN dataIn_NORTH[3] 
    ANTENNAPARTIALMETALAREA 2.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.25 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.5 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.998 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 15.5513 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 63.0833 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.28205 LAYER VL ;
  END dataIn_NORTH[3]
  PIN dataIn_NORTH[2] 
    ANTENNAPARTIALMETALAREA 2.9 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.73 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 48.9103 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 180.455 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END dataIn_NORTH[2]
  PIN dataIn_NORTH[1] 
    ANTENNAPARTIALMETALAREA 2.54 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.546 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 43.141 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 161.481 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END dataIn_NORTH[1]
  PIN dataIn_NORTH[0] 
    ANTENNAPARTIALMETALAREA 2.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.25 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.368 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 15.2564 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 60.6795 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.28205 LAYER VL ;
  END dataIn_NORTH[0]
  PIN destinationAddressOut_NORTH[11] 
    ANTENNAPARTIALMETALAREA 8.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 30.266 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 24.272 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 5.89677 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 23.0302 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END destinationAddressOut_NORTH[11]
  PIN destinationAddressOut_NORTH[10] 
    ANTENNAPARTIALMETALAREA 2.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.25 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 24.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 92.056 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 14.4079 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 54.6746 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END destinationAddressOut_NORTH[10]
  PIN destinationAddressOut_NORTH[9] 
    ANTENNAPARTIALMETALAREA 5.98 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.274 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.208 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 11.8969 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 45.2306 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END destinationAddressOut_NORTH[9]
  PIN destinationAddressOut_NORTH[8] 
    ANTENNAPARTIALMETALAREA 3.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.838 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 23.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 88.8 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 15.8244 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 58.906 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.252177 LAYER VL ;
  END destinationAddressOut_NORTH[8]
  PIN destinationAddressOut_NORTH[7] 
    ANTENNAPARTIALMETALAREA 6.28 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.384 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.76 LAYER M2 ; 
    ANTENNAMAXAREACAR 3.73 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 13.9548 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.0454545 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.144 LAYER M3 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 4.28877 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 16.0988 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END destinationAddressOut_NORTH[7]
  PIN destinationAddressOut_NORTH[6] 
    ANTENNAPARTIALMETALAREA 3.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.322 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 25.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 93.832 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 15.1813 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 57.3064 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END destinationAddressOut_NORTH[6]
  PIN destinationAddressOut_NORTH[5] 
    ANTENNAPARTIALMETALAREA 3.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.322 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.76 LAYER M2 ; 
    ANTENNAMAXAREACAR 1.87773 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 7.10136 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.0454545 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.584 LAYER M3 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 8.37408 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 32.0431 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END destinationAddressOut_NORTH[5]
  PIN destinationAddressOut_NORTH[4] 
    ANTENNAPARTIALMETALAREA 3.82 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.282 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.76 LAYER M2 ; 
    ANTENNAMAXAREACAR 2.33227 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 8.78318 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.0454545 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.808 LAYER M3 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.95907 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 15.7075 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END destinationAddressOut_NORTH[4]
  PIN destinationAddressOut_NORTH[3] 
    ANTENNAPARTIALMETALAREA 0.42 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.554 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 25.3 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 93.906 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 22.2289 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 82.5539 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END destinationAddressOut_NORTH[3]
  PIN destinationAddressOut_NORTH[2] 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 27.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 101.824 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 16.6584 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 63.1543 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END destinationAddressOut_NORTH[2]
  PIN destinationAddressOut_NORTH[1] 
    ANTENNAPARTIALMETALAREA 4.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.354 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 8.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 32.856 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 8.4239 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 32.6103 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END destinationAddressOut_NORTH[1]
  PIN destinationAddressOut_NORTH[0] 
    ANTENNAPARTIALMETALAREA 9.82 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 36.482 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.064 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 5.38904 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 21.0611 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END destinationAddressOut_NORTH[0]
  PIN requesterAddressOut_NORTH[3] 
    ANTENNAPARTIALMETALAREA 10.54 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 39.146 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.88 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 5.13334 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 20.2055 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END requesterAddressOut_NORTH[3]
  PIN requesterAddressOut_NORTH[2] 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.37 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 23.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 88.504 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 14.8165 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 56.2628 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END requesterAddressOut_NORTH[2]
  PIN requesterAddressOut_NORTH[1] 
    ANTENNAPARTIALMETALAREA 5.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 18.722 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.384 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 4.76389 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 19.1448 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END requesterAddressOut_NORTH[1]
  PIN requesterAddressOut_NORTH[0] 
    ANTENNAPARTIALMETALAREA 8.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 30.266 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 12.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 45.584 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 7.81531 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 29.502 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.252177 LAYER VL ;
  END requesterAddressOut_NORTH[0]
  PIN dataOut_NORTH[5] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 27.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 102.12 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 28.2324 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 106.132 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END dataOut_NORTH[5]
  PIN dataOut_NORTH[4] 
    ANTENNAPARTIALMETALAREA 4.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.466 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 22.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 82.88 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 16.2828 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 61.9178 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END dataOut_NORTH[4]
  PIN dataOut_NORTH[3] 
    ANTENNAPARTIALMETALAREA 0.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.85 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 23.14 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 87.246 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 14.5371 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 55.6119 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END dataOut_NORTH[3]
  PIN dataOut_NORTH[2] 
    ANTENNAPARTIALMETALAREA 13.96 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 51.8 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 7.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 26.936 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 5.36896 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 21.14 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END dataOut_NORTH[2]
  PIN dataOut_NORTH[1] 
    ANTENNAPARTIALMETALAREA 12.58 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 46.842 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 26.344 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 6.2121 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 24.2596 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END dataOut_NORTH[1]
  PIN dataOut_NORTH[0] 
    ANTENNAPARTIALMETALAREA 6.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 25.826 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 18.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 68.08 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 12.5112 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 47.5661 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END dataOut_NORTH[0]
  PIN destinationAddressIn_SOUTH[11] 
    ANTENNAPARTIALMETALAREA 3.96 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.652 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 11.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 42.92 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3168 LAYER M3 ; 
    ANTENNAMAXAREACAR 42.7701 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 161.531 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.28205 LAYER VL ;
  END destinationAddressIn_SOUTH[11]
  PIN destinationAddressIn_SOUTH[10] 
    ANTENNAPARTIALMETALAREA 3.86 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.282 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 11.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 42.328 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3168 LAYER M3 ; 
    ANTENNAMAXAREACAR 40.3438 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 151.598 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.28205 LAYER VL ;
  END destinationAddressIn_SOUTH[10]
  PIN destinationAddressIn_SOUTH[9] 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 8.22 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 30.71 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3264 LAYER M3 ; 
    ANTENNAMAXAREACAR 37.8066 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 140.002 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.28205 LAYER VL ;
  END destinationAddressIn_SOUTH[9]
  PIN destinationAddressIn_SOUTH[8] 
    ANTENNAPARTIALMETALAREA 3.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.838 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 9.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 36.408 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3264 LAYER M3 ; 
    ANTENNAMAXAREACAR 34.3835 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 129.531 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.28205 LAYER VL ;
  END destinationAddressIn_SOUTH[8]
  PIN destinationAddressIn_SOUTH[7] 
    ANTENNAPARTIALMETALAREA 2.4 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.028 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 40.8974 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 153.179 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END destinationAddressIn_SOUTH[7]
  PIN destinationAddressIn_SOUTH[6] 
    ANTENNAPARTIALMETALAREA 2.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.954 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 40.5769 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 151.994 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END destinationAddressIn_SOUTH[6]
  PIN destinationAddressIn_SOUTH[5] 
    ANTENNAPARTIALMETALAREA 2.7 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.138 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 45.7051 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 170.968 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END destinationAddressIn_SOUTH[5]
  PIN destinationAddressIn_SOUTH[4] 
    ANTENNAPARTIALMETALAREA 2.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.954 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 42.7308 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 160.712 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END destinationAddressIn_SOUTH[4]
  PIN destinationAddressIn_SOUTH[3] 
    ANTENNAPARTIALMETALAREA 2.54 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.546 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 45.2949 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 170.199 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END destinationAddressIn_SOUTH[3]
  PIN destinationAddressIn_SOUTH[2] 
    ANTENNAPARTIALMETALAREA 2.34 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.658 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.48 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 13.3077 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 54.7821 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.28205 LAYER VL ;
  END destinationAddressIn_SOUTH[2]
  PIN destinationAddressIn_SOUTH[1] 
    ANTENNAPARTIALMETALAREA 2.4 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.88 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 43.9231 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 163.231 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END destinationAddressIn_SOUTH[1]
  PIN destinationAddressIn_SOUTH[0] 
    ANTENNAPARTIALMETALAREA 2.46 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.102 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 41.859 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 154.365 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END destinationAddressIn_SOUTH[0]
  PIN requesterAddressIn_SOUTH[3] 
    ANTENNAPARTIALMETALAREA 2.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.954 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 40.5769 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 151.994 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END requesterAddressIn_SOUTH[3]
  PIN requesterAddressIn_SOUTH[2] 
    ANTENNAPARTIALMETALAREA 1.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.178 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.624 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 33.2051 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 127.09 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.28205 LAYER VL ;
  END requesterAddressIn_SOUTH[2]
  PIN requesterAddressIn_SOUTH[1] 
    ANTENNAPARTIALMETALAREA 2.54 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.546 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 43.141 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 161.481 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END requesterAddressIn_SOUTH[1]
  PIN requesterAddressIn_SOUTH[0] 
    ANTENNAPARTIALMETALAREA 2.54 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.546 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 43.141 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 161.481 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END requesterAddressIn_SOUTH[0]
  PIN dataIn_SOUTH[5] 
    ANTENNAPARTIALMETALAREA 3.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.618 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 54.2692 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 203.404 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END dataIn_SOUTH[5]
  PIN dataIn_SOUTH[4] 
    ANTENNAPARTIALMETALAREA 2.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.954 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 40.5769 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 151.994 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END dataIn_SOUTH[4]
  PIN dataIn_SOUTH[3] 
    ANTENNAPARTIALMETALAREA 2.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.954 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 40.5769 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 151.994 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END dataIn_SOUTH[3]
  PIN dataIn_SOUTH[2] 
    ANTENNAPARTIALMETALAREA 2.44 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.176 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 41.5385 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 155.551 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END dataIn_SOUTH[2]
  PIN dataIn_SOUTH[1] 
    ANTENNAPARTIALMETALAREA 2.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.026 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 49.5513 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 185.199 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END dataIn_SOUTH[1]
  PIN dataIn_SOUTH[0] 
    ANTENNAPARTIALMETALAREA 2.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.954 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 40.5769 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 151.994 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END dataIn_SOUTH[0]
  PIN destinationAddressOut_SOUTH[11] 
    ANTENNAPARTIALMETALAREA 6.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.458 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 9.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 34.04 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 6.0355 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 22.8402 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.252177 LAYER VL ;
  END destinationAddressOut_SOUTH[11]
  PIN destinationAddressOut_SOUTH[10] 
    ANTENNAPARTIALMETALAREA 1.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.178 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 15.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 58.312 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 9.6158 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 36.0873 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.252177 LAYER VL ;
  END destinationAddressOut_SOUTH[10]
  PIN destinationAddressOut_SOUTH[9] 
    ANTENNAPARTIALMETALAREA 17.56 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 65.416 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.536 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 9.46818 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 36.1539 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END destinationAddressOut_SOUTH[9]
  PIN destinationAddressOut_SOUTH[8] 
    ANTENNAPARTIALMETALAREA 3.86 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.43 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 25.16 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 5.03293 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 20.0637 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END destinationAddressOut_SOUTH[8]
  PIN destinationAddressOut_SOUTH[7] 
    ANTENNAPARTIALMETALAREA 2.62 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.842 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.76 LAYER M2 ; 
    ANTENNAMAXAREACAR 1.65045 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 6.26045 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.0454545 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.664 LAYER M3 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 8.00923 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 30.6931 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END destinationAddressOut_SOUTH[7]
  PIN destinationAddressOut_SOUTH[6] 
    ANTENNAPARTIALMETALAREA 3.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.322 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.76 LAYER M2 ; 
    ANTENNAMAXAREACAR 1.87773 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 7.10136 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.0454545 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.848 LAYER M3 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.39511 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 9.09226 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END destinationAddressOut_SOUTH[6]
  PIN destinationAddressOut_SOUTH[5] 
    ANTENNAPARTIALMETALAREA 1.04 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.848 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 10.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 38.776 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 7.48265 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 28.8213 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END destinationAddressOut_SOUTH[5]
  PIN destinationAddressOut_SOUTH[4] 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.37 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 8.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 32.708 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 8.94895 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 34.2467 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END destinationAddressOut_SOUTH[4]
  PIN destinationAddressOut_SOUTH[3] 
    ANTENNAPARTIALMETALAREA 7.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 26.64 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.76 LAYER M2 ; 
    ANTENNAMAXAREACAR 4.23 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 15.8048 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.0454545 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.848 LAYER M3 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 4.74738 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 17.7957 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END destinationAddressOut_SOUTH[3]
  PIN destinationAddressOut_SOUTH[2] 
    ANTENNAPARTIALMETALAREA 4.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 18.426 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.76 LAYER M2 ; 
    ANTENNAMAXAREACAR 2.96864 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 11.1377 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.0454545 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.624 LAYER M3 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 13.0528 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 49.3542 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END destinationAddressOut_SOUTH[2]
  PIN destinationAddressOut_SOUTH[1] 
    ANTENNAPARTIALMETALAREA 1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.84 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 4.79378 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 18.0161 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.252177 LAYER VL ;
  END destinationAddressOut_SOUTH[1]
  PIN destinationAddressOut_SOUTH[0] 
    ANTENNAPARTIALMETALAREA 5.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 18.87 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.584 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 13.0037 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 49.1727 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END destinationAddressOut_SOUTH[0]
  PIN requesterAddressOut_SOUTH[3] 
    ANTENNAPARTIALMETALAREA 7.34 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 27.306 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.76 LAYER M2 ; 
    ANTENNAMAXAREACAR 4.33227 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 16.1832 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.0454545 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.368 LAYER M3 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 4.6427 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 17.4083 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END requesterAddressOut_SOUTH[3]
  PIN requesterAddressOut_SOUTH[2] 
    ANTENNAPARTIALMETALAREA 6.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.162 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.76 LAYER M2 ; 
    ANTENNAMAXAREACAR 3.69591 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 13.8286 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.0454545 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.736 LAYER M3 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 8.80822 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 33.6355 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END requesterAddressOut_SOUTH[2]
  PIN requesterAddressOut_SOUTH[1] 
    ANTENNAPARTIALMETALAREA 3.42 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.802 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.24 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 13.5472 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 51.26 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END requesterAddressOut_SOUTH[1]
  PIN requesterAddressOut_SOUTH[0] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.46 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 9.20726 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 35.279 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END requesterAddressOut_SOUTH[0]
  PIN dataOut_SOUTH[5] 
    ANTENNAPARTIALMETALAREA 4.32 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.984 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.92 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.05537 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 11.5839 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.252177 LAYER VL ;
  END dataOut_SOUTH[5]
  PIN dataOut_SOUTH[4] 
    ANTENNAPARTIALMETALAREA 6.82 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 25.234 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M2 ; 
    ANTENNAMAXAREACAR 4.473 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 16.676 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.231481 LAYER V2 ;
  END dataOut_SOUTH[4]
  PIN dataOut_SOUTH[3] 
    ANTENNAPARTIALMETALAREA 4.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.762 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.104 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.55868 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 9.7462 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.252177 LAYER VL ;
  END dataOut_SOUTH[3]
  PIN dataOut_SOUTH[2] 
    ANTENNAPARTIALMETALAREA 4.86 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.982 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.76 LAYER M2 ; 
    ANTENNAMAXAREACAR 2.92318 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 10.8855 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.0454545 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.848 LAYER M3 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 8.68405 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 33.1761 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END dataOut_SOUTH[2]
  PIN dataOut_SOUTH[1] 
    ANTENNAPARTIALMETALAREA 2.64 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.768 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.104 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.45471 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 13.0894 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END dataOut_SOUTH[1]
  PIN dataOut_SOUTH[0] 
    ANTENNAPARTIALMETALAREA 1.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.178 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.912 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 4.95735 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 19.5404 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END dataOut_SOUTH[0]
  PIN destinationAddressIn_EAST[11] 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.37 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 37.42 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 139.046 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3168 LAYER M3 ; 
    ANTENNAMAXAREACAR 142.99 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 532.792 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER VL ;
  END destinationAddressIn_EAST[11]
  PIN destinationAddressIn_EAST[10] 
    ANTENNAPARTIALMETALAREA 1.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.514 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 37.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 139.712 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3168 LAYER M3 ; 
    ANTENNAMAXAREACAR 148.687 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 553.869 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.28205 LAYER VL ;
  END destinationAddressIn_EAST[10]
  PIN destinationAddressIn_EAST[9] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 25.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 95.904 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3264 LAYER M3 ; 
    ANTENNAMAXAREACAR 101.352 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 378.221 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER VL ;
  END destinationAddressIn_EAST[9]
  PIN destinationAddressIn_EAST[8] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 19.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 73.704 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3264 LAYER M3 ; 
    ANTENNAMAXAREACAR 140.662 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 523.668 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.92308 LAYER VL ;
  END destinationAddressIn_EAST[8]
  PIN destinationAddressIn_EAST[7] 
    ANTENNAPARTIALMETALAREA 0.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.518 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.54 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.246 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 63.2436 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 238.981 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.28205 LAYER VL ;
  END destinationAddressIn_EAST[7]
  PIN destinationAddressIn_EAST[6] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.7 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.838 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 64.9359 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 244.494 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.28205 LAYER VL ;
  END destinationAddressIn_EAST[6]
  PIN destinationAddressIn_EAST[5] 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.58 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 17.094 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 77.7564 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 291.929 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.28205 LAYER VL ;
  END destinationAddressIn_EAST[5]
  PIN destinationAddressIn_EAST[4] 
    ANTENNAPARTIALMETALAREA 0.98 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.626 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 57.0641 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 231.596 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END destinationAddressIn_EAST[4]
  PIN destinationAddressIn_EAST[3] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.248 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 84.4872 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 316.833 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.28205 LAYER VL ;
  END destinationAddressIn_EAST[3]
  PIN destinationAddressIn_EAST[2] 
    ANTENNAPARTIALMETALAREA 1.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.922 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 58.3462 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 236.34 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END destinationAddressIn_EAST[2]
  PIN destinationAddressIn_EAST[1] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 56.9359 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 237.75 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END destinationAddressIn_EAST[1]
  PIN destinationAddressIn_EAST[0] 
    ANTENNAPARTIALMETALAREA 0.12 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.444 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 59.6923 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 250.346 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END destinationAddressIn_EAST[0]
  PIN requesterAddressIn_EAST[3] 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.58 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.394 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 109.167 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 408.147 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.28205 LAYER VL ;
  END requesterAddressIn_EAST[3]
  PIN requesterAddressIn_EAST[2] 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.768 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 83.9231 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 315.41 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.28205 LAYER VL ;
  END requesterAddressIn_EAST[2]
  PIN requesterAddressIn_EAST[1] 
    ANTENNAPARTIALMETALAREA 2.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.398 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 56.8077 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 219.481 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END requesterAddressIn_EAST[1]
  PIN requesterAddressIn_EAST[0] 
    ANTENNAPARTIALMETALAREA 0.12 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.444 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 40.9744 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 170.795 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END requesterAddressIn_EAST[0]
  PIN dataIn_EAST[5] 
    ANTENNAPARTIALMETALAREA 0.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.518 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.064 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 84.4872 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 316.833 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.28205 LAYER VL ;
  END dataIn_EAST[5]
  PIN dataIn_EAST[4] 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.84 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 71.7692 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 272.218 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.28205 LAYER VL ;
  END dataIn_EAST[4]
  PIN dataIn_EAST[3] 
    ANTENNAPARTIALMETALAREA 1.42 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.402 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 57.9615 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 233.904 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END dataIn_EAST[3]
  PIN dataIn_EAST[2] 
    ANTENNAPARTIALMETALAREA 0.12 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.444 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.472 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 46.8974 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 178.5 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.28205 LAYER VL ;
  END dataIn_EAST[2]
  PIN dataIn_EAST[1] 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.37 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 31.6795 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 131.468 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END dataIn_EAST[1]
  PIN dataIn_EAST[0] 
    ANTENNAPARTIALMETALAREA 1.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.178 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 60.141 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 236.212 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END dataIn_EAST[0]
  PIN destinationAddressOut_EAST[11] 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.332 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 20.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 75.776 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 18.675 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 70.2331 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END destinationAddressOut_EAST[11]
  PIN destinationAddressOut_EAST[10] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 17.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 65.712 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 14.027 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 53.0354 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END destinationAddressOut_EAST[10]
  PIN destinationAddressOut_EAST[9] 
    ANTENNAPARTIALMETALAREA 0.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.518 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 15.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 58.904 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 13.075 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 49.513 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END destinationAddressOut_EAST[9]
  PIN destinationAddressOut_EAST[8] 
    ANTENNAPARTIALMETALAREA 0.12 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.444 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 13.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 49.432 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 13.1857 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 49.9087 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END destinationAddressOut_EAST[8]
  PIN destinationAddressOut_EAST[7] 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.37 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 8.5 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 31.598 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 11.5922 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 43.9502 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END destinationAddressOut_EAST[7]
  PIN destinationAddressOut_EAST[6] 
    ANTENNAPARTIALMETALAREA 0.08 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.296 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 22.2 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 7.06291 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 27.2544 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END destinationAddressOut_EAST[6]
  PIN destinationAddressOut_EAST[5] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.128 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 9.52781 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 36.3468 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END destinationAddressOut_EAST[5]
  PIN destinationAddressOut_EAST[4] 
    ANTENNAPARTIALMETALAREA 0.12 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.444 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.72 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 12.8282 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 48.5998 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END destinationAddressOut_EAST[4]
  PIN destinationAddressOut_EAST[3] 
    ANTENNAPARTIALMETALAREA 0.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.258 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 12.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 47.952 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 11.5435 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 43.8466 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END destinationAddressOut_EAST[3]
  PIN destinationAddressOut_EAST[2] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 12.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 45.88 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 12.1797 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 46.2005 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END destinationAddressOut_EAST[2]
  PIN destinationAddressOut_EAST[1] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 10.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 40.848 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 10.5295 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 40.1711 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END destinationAddressOut_EAST[1]
  PIN destinationAddressOut_EAST[0] 
    ANTENNAPARTIALMETALAREA 0.12 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.444 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 9.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 35.816 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 14.4761 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 54.6973 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END destinationAddressOut_EAST[0]
  PIN requesterAddressOut_EAST[3] 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 17.82 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 66.082 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 10.8587 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 41.2361 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END requesterAddressOut_EAST[3]
  PIN requesterAddressOut_EAST[2] 
    ANTENNAPARTIALMETALAREA 0.08 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.296 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 12.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 47.36 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 8.22001 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 31.5496 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END requesterAddressOut_EAST[2]
  PIN requesterAddressOut_EAST[1] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 18.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 67.488 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 18.442 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 69.3709 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END requesterAddressOut_EAST[1]
  PIN requesterAddressOut_EAST[0] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 19.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 73.704 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 18.406 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 69.1611 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END requesterAddressOut_EAST[0]
  PIN dataOut_EAST[5] 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.37 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 23.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 87.024 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 13.9618 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 52.0144 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.252177 LAYER VL ;
  END dataOut_EAST[5]
  PIN dataOut_EAST[4] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 27.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 101.824 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 16.6791 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 63.1543 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END dataOut_EAST[4]
  PIN dataOut_EAST[3] 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 26.38 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 98.198 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 15.2875 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 57.8524 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END dataOut_EAST[3]
  PIN dataOut_EAST[2] 
    ANTENNAPARTIALMETALAREA 0.12 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.444 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 23.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 87.616 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 15.2173 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 57.5163 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END dataOut_EAST[2]
  PIN dataOut_EAST[1] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 22.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 82.88 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 21.4995 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 80.7604 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END dataOut_EAST[1]
  PIN dataOut_EAST[0] 
    ANTENNAPARTIALMETALAREA 0.28 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.184 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 19.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 71.336 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 13.8668 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 52.5192 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END dataOut_EAST[0]
  PIN destinationAddressIn_WEST[11] 
    ANTENNAPARTIALMETALAREA 0.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.518 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.984 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3168 LAYER M3 ; 
    ANTENNAMAXAREACAR 60.4183 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 226.682 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.13854 LAYER VL ;
  END destinationAddressIn_WEST[11]
  PIN destinationAddressIn_WEST[10] 
    ANTENNAPARTIALMETALAREA 0.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.518 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 9.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 35.816 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3168 LAYER M3 ; 
    ANTENNAMAXAREACAR 85.1235 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 321.799 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.28205 LAYER VL ;
  END destinationAddressIn_WEST[10]
  PIN destinationAddressIn_WEST[9] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.288 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3264 LAYER M3 ; 
    ANTENNAMAXAREACAR 38.3499 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 144.081 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.763575 LAYER VL ;
  END destinationAddressIn_WEST[9]
  PIN destinationAddressIn_WEST[8] 
    ANTENNAPARTIALMETALAREA 6.92 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 25.9 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3264 LAYER M2 ; 
    ANTENNAMAXAREACAR 26.6625 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 100.274 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END destinationAddressIn_WEST[8]
  PIN destinationAddressIn_WEST[7] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.32 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 78.0769 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 293.115 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.28205 LAYER VL ;
  END destinationAddressIn_WEST[7]
  PIN destinationAddressIn_WEST[6] 
    ANTENNAPARTIALMETALAREA 2.52 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.472 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 67.3846 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 264.256 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END destinationAddressIn_WEST[6]
  PIN destinationAddressIn_WEST[5] 
    ANTENNAPARTIALMETALAREA 3.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.618 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 65.3974 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 250.699 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END destinationAddressIn_WEST[5]
  PIN destinationAddressIn_WEST[4] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.248 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 55 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 207.731 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.28205 LAYER VL ;
  END destinationAddressIn_WEST[4]
  PIN destinationAddressIn_WEST[3] 
    ANTENNAPARTIALMETALAREA 0.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.518 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.472 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 57.5641 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 217.218 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.28205 LAYER VL ;
  END destinationAddressIn_WEST[3]
  PIN destinationAddressIn_WEST[2] 
    ANTENNAPARTIALMETALAREA 0.82 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.034 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 40.141 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 161.083 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END destinationAddressIn_WEST[2]
  PIN destinationAddressIn_WEST[1] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.84 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 66.5385 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 250.423 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.28205 LAYER VL ;
  END destinationAddressIn_WEST[1]
  PIN destinationAddressIn_WEST[0] 
    ANTENNAPARTIALMETALAREA 0.52 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.924 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.768 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 47.3077 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 179.269 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.28205 LAYER VL ;
  END destinationAddressIn_WEST[0]
  PIN requesterAddressIn_WEST[3] 
    ANTENNAPARTIALMETALAREA 2.34 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.806 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 63.4744 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 249.224 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END requesterAddressIn_WEST[3]
  PIN requesterAddressIn_WEST[2] 
    ANTENNAPARTIALMETALAREA 0.98 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.626 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 49.8846 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 201.083 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END requesterAddressIn_WEST[2]
  PIN requesterAddressIn_WEST[1] 
    ANTENNAPARTIALMETALAREA 1.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.514 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 47.9615 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 193.519 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END requesterAddressIn_WEST[1]
  PIN requesterAddressIn_WEST[0] 
    ANTENNAPARTIALMETALAREA 2.88 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.804 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 57.7692 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 220.218 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END requesterAddressIn_WEST[0]
  PIN dataIn_WEST[5] 
    ANTENNAPARTIALMETALAREA 0.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.518 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.472 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 47.3077 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 179.269 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.28205 LAYER VL ;
  END dataIn_WEST[5]
  PIN dataIn_WEST[4] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.992 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 119.103 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 444.91 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.28205 LAYER VL ;
  END dataIn_WEST[4]
  PIN dataIn_WEST[3] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.472 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 51.1538 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 193.5 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.28205 LAYER VL ;
  END dataIn_WEST[3]
  PIN dataIn_WEST[2] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.88 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 115.718 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 433.615 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.28205 LAYER VL ;
  END dataIn_WEST[2]
  PIN dataIn_WEST[1] 
    ANTENNAPARTIALMETALAREA 0.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.518 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 32.3205 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 133.84 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END dataIn_WEST[1]
  PIN dataIn_WEST[0] 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.4 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 66.7436 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 252.974 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.28205 LAYER VL ;
  END dataIn_WEST[0]
  PIN destinationAddressOut_WEST[11] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 26.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 99.456 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 18.642 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 70.494 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END destinationAddressOut_WEST[11]
  PIN destinationAddressOut_WEST[10] 
    ANTENNAPARTIALMETALAREA 0.08 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.296 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 32.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 120.472 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 22.5274 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 84.7933 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END destinationAddressOut_WEST[10]
  PIN destinationAddressOut_WEST[9] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 27.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 102.12 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 19.4775 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 73.5853 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END destinationAddressOut_WEST[9]
  PIN destinationAddressOut_WEST[8] 
    ANTENNAPARTIALMETALAREA 0.12 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.444 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 26.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 100.344 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 16.4867 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 61.5094 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.252177 LAYER VL ;
  END destinationAddressOut_WEST[8]
  PIN destinationAddressOut_WEST[7] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 25.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 95.904 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 17.7238 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 66.9433 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END destinationAddressOut_WEST[7]
  PIN destinationAddressOut_WEST[6] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 26.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 97.088 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 14.8103 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 55.3836 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.252177 LAYER VL ;
  END destinationAddressOut_WEST[6]
  PIN destinationAddressOut_WEST[5] 
    ANTENNAPARTIALMETALAREA 0.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.518 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 23.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 89.392 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 16.7718 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 63.5741 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END destinationAddressOut_WEST[5]
  PIN destinationAddressOut_WEST[4] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 17.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 65.12 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 14.3658 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 54.4421 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END destinationAddressOut_WEST[4]
  PIN destinationAddressOut_WEST[3] 
    ANTENNAPARTIALMETALAREA 0.62 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.442 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.384 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 19.7312 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 73.3124 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END destinationAddressOut_WEST[3]
  PIN destinationAddressOut_WEST[2] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.424 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 8.84206 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 33.0991 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END destinationAddressOut_WEST[2]
  PIN destinationAddressOut_WEST[1] 
    ANTENNAPARTIALMETALAREA 0.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.518 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.384 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 4.82597 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 19.1448 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END destinationAddressOut_WEST[1]
  PIN destinationAddressOut_WEST[0] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.536 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 4.33419 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 17.3113 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END destinationAddressOut_WEST[0]
  PIN requesterAddressOut_WEST[3] 
    ANTENNAPARTIALMETALAREA 20.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 74.37 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 9.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 34.928 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 6.90471 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 25.8265 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.252177 LAYER VL ;
  END requesterAddressOut_WEST[3]
  PIN requesterAddressOut_WEST[2] 
    ANTENNAPARTIALMETALAREA 5.72 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 21.312 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 17.464 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 4.01886 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 16.0819 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END requesterAddressOut_WEST[2]
  PIN requesterAddressOut_WEST[1] 
    ANTENNAPARTIALMETALAREA 24.98 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 92.574 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.584 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.81852 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 11.4875 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END requesterAddressOut_WEST[1]
  PIN requesterAddressOut_WEST[0] 
    ANTENNAPARTIALMETALAREA 27.44 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 101.676 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.688 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.8582 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 15.3204 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END requesterAddressOut_WEST[0]
  PIN dataOut_WEST[5] 
    ANTENNAPARTIALMETALAREA 15.92 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 59.052 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 23.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 89.096 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 14.0817 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 53.3006 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END dataOut_WEST[5]
  PIN dataOut_WEST[4] 
    ANTENNAPARTIALMETALAREA 0.08 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.296 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 14.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 52.688 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 25.1481 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 94.2599 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END dataOut_WEST[4]
  PIN dataOut_WEST[3] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 13.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 51.8 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 15.7439 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 59.5412 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END dataOut_WEST[3]
  PIN dataOut_WEST[2] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 23.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 87.912 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 27.213 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 102.206 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END dataOut_WEST[2]
  PIN dataOut_WEST[1] 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.37 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 20.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 76.072 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 13.5203 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 51.5436 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END dataOut_WEST[1]
  PIN dataOut_WEST[0] 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 19.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 71.928 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 17.1696 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 64.8163 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END dataOut_WEST[0]
  PIN cacheDataIn_A[5] 
    ANTENNAPARTIALMETALAREA 2.9 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.878 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.76 LAYER M2 ; 
    ANTENNAMAXAREACAR 1.80955 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 6.84909 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.0454545 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.624 LAYER M3 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 8.94628 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 33.3056 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END cacheDataIn_A[5]
  PIN cacheDataIn_A[4] 
    ANTENNAPARTIALMETALAREA 0.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.518 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 16.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 62.752 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 12.2844 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 45.7331 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END cacheDataIn_A[4]
  PIN cacheDataIn_A[3] 
    ANTENNAPARTIALMETALAREA 5.4 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.128 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.312 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 8.36221 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 31.1445 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END cacheDataIn_A[3]
  PIN cacheDataIn_A[2] 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 20.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 75.184 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 17.7265 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 65.8307 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END cacheDataIn_A[2]
  PIN cacheDataIn_A[1] 
    ANTENNAPARTIALMETALAREA 4.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.762 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 20.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 74.888 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 13.0141 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 48.5861 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END cacheDataIn_A[1]
  PIN cacheDataIn_A[0] 
    ANTENNAPARTIALMETALAREA 7.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 26.714 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 18.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 68.376 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 12.6078 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 46.9299 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END cacheDataIn_A[0]
  PIN cacheAddressIn_A[7] 
    ANTENNAPARTIALMETALAREA 3.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.986 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.952 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 4.13576 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 15.5067 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END cacheAddressIn_A[7]
  PIN cacheAddressIn_A[6] 
    ANTENNAPARTIALMETALAREA 3.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.654 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M2 ; 
    ANTENNAMAXAREACAR 3.67931 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 12.9613 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.231481 LAYER V2 ;
  END cacheAddressIn_A[6]
  PIN cacheAddressIn_A[5] 
    ANTENNAPARTIALMETALAREA 2.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.324 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.76 LAYER M2 ; 
    ANTENNAMAXAREACAR 1.57091 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 5.96614 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.0454545 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.584 LAYER M3 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 6.11945 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 22.8463 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END cacheAddressIn_A[5]
  PIN cacheAddressIn_A[4] 
    ANTENNAPARTIALMETALAREA 4.66 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.538 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.76 LAYER M2 ; 
    ANTENNAMAXAREACAR 2.80955 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 10.6332 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.0454545 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.472 LAYER M3 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 12.7251 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 47.2872 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END cacheAddressIn_A[4]
  PIN cacheAddressIn_A[3] 
    ANTENNAPARTIALMETALAREA 3.58 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.394 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 10.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 38.776 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 9.833 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 36.3013 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.252177 LAYER VL ;
  END cacheAddressIn_A[3]
  PIN cacheAddressIn_A[2] 
    ANTENNAPARTIALMETALAREA 5.58 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.794 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 11.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 41.736 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 14.4175 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 53.7023 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END cacheAddressIn_A[2]
  PIN cacheAddressIn_A[1] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 17.62 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 65.49 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 11.7413 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 43.7238 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END cacheAddressIn_A[1]
  PIN cacheAddressIn_A[0] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 10.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 39.368 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 15.0123 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 55.9031 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END cacheAddressIn_A[0]
  PIN cacheDataOut_A[5] 
    ANTENNAPARTIALMETALAREA 1.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.178 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.1 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.762 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1152 LAYER M3 ; 
    ANTENNAMAXAREACAR 41.5382 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 159.944 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END cacheDataOut_A[5]
  PIN cacheDataOut_A[4] 
    ANTENNAPARTIALMETALAREA 1.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.178 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.472 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1152 LAYER M3 ; 
    ANTENNAMAXAREACAR 60.4618 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 226.108 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END cacheDataOut_A[4]
  PIN cacheDataOut_A[3] 
    ANTENNAPARTIALMETALAREA 7.82 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 29.082 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.552 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1488 LAYER M3 ; 
    ANTENNAMAXAREACAR 8.6371 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 35.8038 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.537634 LAYER VL ;
  END cacheDataOut_A[3]
  PIN cacheDataOut_A[2] 
    ANTENNAPARTIALMETALAREA 3.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.986 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.368 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1152 LAYER M3 ; 
    ANTENNAMAXAREACAR 21.9201 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 84.7882 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END cacheDataOut_A[2]
  PIN cacheDataOut_A[1] 
    ANTENNAPARTIALMETALAREA 8.44 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 31.228 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.4 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1152 LAYER M3 ; 
    ANTENNAMAXAREACAR 21.2257 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 82.151 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END cacheDataOut_A[1]
  PIN cacheDataOut_A[0] 
    ANTENNAPARTIALMETALAREA 3.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.618 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 17.76 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1656 LAYER M3 ; 
    ANTENNAMAXAREACAR 36.5266 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 136.744 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.483092 LAYER VL ;
  END cacheDataOut_A[0]
  PIN cacheDataIn_B[5] 
    ANTENNAPARTIALMETALAREA 3.26 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.21 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.76 LAYER M2 ; 
    ANTENNAMAXAREACAR 2.01409 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 7.60591 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.0454545 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M3 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 5.24154 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 19.736 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END cacheDataIn_B[5]
  PIN cacheDataIn_B[4] 
    ANTENNAPARTIALMETALAREA 5.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 19.018 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M2 ; 
    ANTENNAMAXAREACAR 7.41889 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 28.1382 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER V2 ;
  END cacheDataIn_B[4]
  PIN cacheDataIn_B[3] 
    ANTENNAPARTIALMETALAREA 6.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.458 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.584 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.78394 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 14.2815 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END cacheDataIn_B[3]
  PIN cacheDataIn_B[2] 
    ANTENNAPARTIALMETALAREA 6.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 25.826 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M2 ; 
    ANTENNAMAXAREACAR 42.0926 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 155.87 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M3 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 42.3202 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 156.789 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END cacheDataIn_B[2]
  PIN cacheDataIn_B[1] 
    ANTENNAPARTIALMETALAREA 5.26 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 19.61 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 13.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 49.728 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 19.7017 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 73.2539 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END cacheDataIn_B[1]
  PIN cacheDataIn_B[0] 
    ANTENNAPARTIALMETALAREA 10.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 38.554 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M2 ; 
    ANTENNAMAXAREACAR 62 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 229.528 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.256 LAYER M3 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 62.4346 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 231.212 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END cacheDataIn_B[0]
  PIN cacheAddressIn_B[7] 
    ANTENNAPARTIALMETALAREA 3.88 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.504 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M2 ; 
    ANTENNAMAXAREACAR 24.3843 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 90.3495 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.96 LAYER M3 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.7568 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 91.881 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END cacheAddressIn_B[7]
  PIN cacheAddressIn_B[6] 
    ANTENNAPARTIALMETALAREA 3.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.098 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 22.2 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 6.17157 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 23.0392 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END cacheAddressIn_B[6]
  PIN cacheAddressIn_B[5] 
    ANTENNAPARTIALMETALAREA 3.66 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.69 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M2 ; 
    ANTENNAMAXAREACAR 23.1111 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 85.6389 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.104 LAYER M3 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.0838 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 89.3144 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END cacheAddressIn_B[5]
  PIN cacheAddressIn_B[4] 
    ANTENNAPARTIALMETALAREA 6.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.754 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.832 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 7.6923 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 28.6659 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END cacheAddressIn_B[4]
  PIN cacheAddressIn_B[3] 
    ANTENNAPARTIALMETALAREA 6.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.866 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.84 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 4.23924 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 15.9661 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END cacheAddressIn_B[3]
  PIN cacheAddressIn_B[2] 
    ANTENNAPARTIALMETALAREA 1.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.514 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 21.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 79.032 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 14.3271 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 52.5112 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.252177 LAYER VL ;
  END cacheAddressIn_B[2]
  PIN cacheAddressIn_B[1] 
    ANTENNAPARTIALMETALAREA 3.58 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.394 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 19.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 73.408 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 16.9945 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 63.2371 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END cacheAddressIn_B[1]
  PIN cacheAddressIn_B[0] 
    ANTENNAPARTIALMETALAREA 6.62 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 24.642 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 LAYER M2 ; 
    ANTENNAMAXAREACAR 40.2407 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 149.019 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.624 LAYER M3 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 41.0065 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 151.928 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END cacheAddressIn_B[0]
  PIN cacheDataOut_B[5] 
    ANTENNAPARTIALMETALAREA 2.58 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.546 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.86 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.478 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1152 LAYER M3 ; 
    ANTENNAMAXAREACAR 12.6215 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 50.2847 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END cacheDataOut_B[5]
  PIN cacheDataOut_B[4] 
    ANTENNAPARTIALMETALAREA 4.54 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.798 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.36 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1152 LAYER M3 ; 
    ANTENNAMAXAREACAR 26.4167 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 101.425 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END cacheDataOut_B[4]
  PIN cacheDataOut_B[3] 
    ANTENNAPARTIALMETALAREA 1.86 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.882 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.62 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 17.538 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1584 LAYER M3 ; 
    ANTENNAMAXAREACAR 34.5025 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 131.227 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.505051 LAYER VL ;
  END cacheDataOut_B[3]
  PIN cacheDataOut_B[2] 
    ANTENNAPARTIALMETALAREA 5.62 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.794 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 18.056 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1152 LAYER M3 ; 
    ANTENNAMAXAREACAR 43.4479 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 167.01 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END cacheDataOut_B[2]
  PIN cacheDataOut_B[1] 
    ANTENNAPARTIALMETALAREA 1.86 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.882 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.42 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.394 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 46.491 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 182.523 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END cacheDataOut_B[1]
  PIN cacheDataOut_B[0] 
    ANTENNAPARTIALMETALAREA 1.86 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.882 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.332 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1656 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.3043 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 91.3092 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.483092 LAYER VL ;
  END cacheDataOut_B[0]
  PIN clk 
    ANTENNAPARTIALMETALAREA 41.7 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 155.474 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.7016 LAYER M3 ; 
    ANTENNAMAXAREACAR 25.0983 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 93.8138 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0470146 LAYER VL ;
  END clk
  PIN reset 
    ANTENNAPARTIALMETALAREA 7.06 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 26.122 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1152 LAYER M3 ; 
    ANTENNAMAXAREACAR 89.4549 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 332.097 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END reset
  PIN readIn_NORTH 
    ANTENNAPARTIALMETALAREA 2.62 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.842 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 44.4231 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 166.224 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END readIn_NORTH
  PIN writeIn_NORTH 
    ANTENNAPARTIALMETALAREA 2.54 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.546 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 47.3462 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 178.917 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END writeIn_NORTH
  PIN readIn_SOUTH 
    ANTENNAPARTIALMETALAREA 2.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.954 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 40.5769 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 151.994 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END readIn_SOUTH
  PIN writeIn_SOUTH 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.37 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.06 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.47 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 88.0128 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 329.878 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.28205 LAYER VL ;
  END writeIn_SOUTH
  PIN readIn_EAST 
    ANTENNAPARTIALMETALAREA 0.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.924 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 35.7179 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 147.654 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END readIn_EAST
  PIN writeIn_EAST 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.544 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 71.2564 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 268.628 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.28205 LAYER VL ;
  END writeIn_EAST
  PIN readIn_WEST 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.176 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M3 ; 
    ANTENNAMAXAREACAR 81.9231 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 307.346 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.28205 LAYER VL ;
  END readIn_WEST
  PIN writeIn_WEST 
    ANTENNAPARTIALMETALAREA 1.46 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.55 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 LAYER M2 ; 
    ANTENNAMAXAREACAR 50.3974 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 201.404 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.641026 LAYER V2 ;
  END writeIn_WEST
  PIN portA_writtenTo 
  END portA_writtenTo
  PIN portB_writtenTo 
  END portB_writtenTo
  PIN readOut_NORTH 
    ANTENNAPARTIALMETALAREA 8.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 29.97 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.848 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.15627 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 9.03719 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END readOut_NORTH
  PIN writeOut_NORTH 
    ANTENNAPARTIALMETALAREA 2.78 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.434 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 18 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 67.192 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 13.2666 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 50.3752 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END writeOut_NORTH
  PIN readOut_SOUTH 
    ANTENNAPARTIALMETALAREA 5.42 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.202 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.664 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.93782 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 7.44901 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.252177 LAYER VL ;
  END readOut_SOUTH
  PIN writeOut_SOUTH 
    ANTENNAPARTIALMETALAREA 7 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 26.048 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.328 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 6.5092 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 25.2196 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END writeOut_SOUTH
  PIN readOut_EAST 
    ANTENNAPARTIALMETALAREA 0.12 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.444 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.24 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 5.23452 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 20.4267 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END readOut_EAST
  PIN writeOut_EAST 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.37 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 8.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 30.784 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 5.6216 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 21.079 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.252177 LAYER VL ;
  END writeOut_EAST
  PIN readOut_WEST 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 10.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 40.552 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 9.60844 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 36.7495 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END readOut_WEST
  PIN writeOut_WEST 
    ANTENNAPARTIALMETALAREA 0.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.518 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 13.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 51.8 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9328 LAYER M3 ; 
    ANTENNAMAXAREACAR 24.1236 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 90.532 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.462963 LAYER VL ;
  END writeOut_WEST
  PIN memWrite_A 
    ANTENNAPARTIALMETALAREA 3.12 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.692 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.76 LAYER M2 ; 
    ANTENNAMAXAREACAR 1.93455 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 7.31159 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.0454545 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.96 LAYER M3 ;
    ANTENNAGATEAREA 1.8248 LAYER M3 ; 
    ANTENNAMAXAREACAR 14.5214 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 55.9554 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.23457 LAYER VL ;
  END memWrite_A
  PIN memWrite_B 
    ANTENNAPARTIALMETALAREA 13.34 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 49.506 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.76 LAYER M2 ; 
    ANTENNAMAXAREACAR 7.74136 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 28.7968 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAMAXCUTCAR 0.0454545 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M3 ;
    ANTENNAGATEAREA 1.8272 LAYER M3 ; 
    ANTENNAMAXAREACAR 7.98217 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 29.7688 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.19048 LAYER VL ;
  END memWrite_B
END router

END LIBRARY
