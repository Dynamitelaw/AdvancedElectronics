
module outputPortArbiter ( clk, reset, selectBit_NORTH, 
        destinationAddressIn_NORTH, requesterAddressIn_NORTH, readIn_NORTH, 
        writeIn_NORTH, dataIn_NORTH, selectBit_SOUTH, 
        destinationAddressIn_SOUTH, requesterAddressIn_SOUTH, readIn_SOUTH, 
        writeIn_SOUTH, dataIn_SOUTH, selectBit_EAST, destinationAddressIn_EAST, 
        requesterAddressIn_EAST, readIn_EAST, writeIn_EAST, dataIn_EAST, 
        selectBit_WEST, destinationAddressIn_WEST, requesterAddressIn_WEST, 
        readIn_WEST, writeIn_WEST, dataIn_WEST, readReady, 
        readRequesterAddress, cacheDataOut, destinationAddressOut, 
        requesterAddressOut, readOut, writeOut, dataOut );
  input [11:0] destinationAddressIn_NORTH;
  input [3:0] requesterAddressIn_NORTH;
  input [5:0] dataIn_NORTH;
  input [11:0] destinationAddressIn_SOUTH;
  input [3:0] requesterAddressIn_SOUTH;
  input [5:0] dataIn_SOUTH;
  input [11:0] destinationAddressIn_EAST;
  input [3:0] requesterAddressIn_EAST;
  input [5:0] dataIn_EAST;
  input [11:0] destinationAddressIn_WEST;
  input [3:0] requesterAddressIn_WEST;
  input [5:0] dataIn_WEST;
  input [3:0] readRequesterAddress;
  input [5:0] cacheDataOut;
  output [11:0] destinationAddressOut;
  output [3:0] requesterAddressOut;
  output [5:0] dataOut;
  input clk, reset, selectBit_NORTH, readIn_NORTH, writeIn_NORTH,
         selectBit_SOUTH, readIn_SOUTH, writeIn_SOUTH, selectBit_EAST,
         readIn_EAST, writeIn_EAST, selectBit_WEST, readIn_WEST, writeIn_WEST,
         readReady;
  output readOut, writeOut;
  wire   N373, N374, N375, \requesterAddressbuffer[0][3] ,
         \requesterAddressbuffer[0][2] , \requesterAddressbuffer[0][1] ,
         \requesterAddressbuffer[0][0] , \requesterAddressbuffer[1][3] ,
         \requesterAddressbuffer[1][2] , \requesterAddressbuffer[1][1] ,
         \requesterAddressbuffer[1][0] , \requesterAddressbuffer[2][3] ,
         \requesterAddressbuffer[2][2] , \requesterAddressbuffer[2][1] ,
         \requesterAddressbuffer[2][0] , \requesterAddressbuffer[3][3] ,
         \requesterAddressbuffer[3][2] , \requesterAddressbuffer[3][1] ,
         \requesterAddressbuffer[3][0] , \requesterAddressbuffer[4][3] ,
         \requesterAddressbuffer[4][2] , \requesterAddressbuffer[4][1] ,
         \requesterAddressbuffer[4][0] , \requesterAddressbuffer[5][3] ,
         \requesterAddressbuffer[5][2] , \requesterAddressbuffer[5][1] ,
         \requesterAddressbuffer[5][0] , \requesterAddressbuffer[6][3] ,
         \requesterAddressbuffer[6][2] , \requesterAddressbuffer[6][1] ,
         \requesterAddressbuffer[6][0] , \requesterAddressbuffer[7][3] ,
         \requesterAddressbuffer[7][2] , \requesterAddressbuffer[7][1] ,
         \requesterAddressbuffer[7][0] , \destinationAddressbuffer[0][11] ,
         \destinationAddressbuffer[0][10] , \destinationAddressbuffer[0][9] ,
         \destinationAddressbuffer[0][8] , \destinationAddressbuffer[0][7] ,
         \destinationAddressbuffer[0][6] , \destinationAddressbuffer[0][5] ,
         \destinationAddressbuffer[0][4] , \destinationAddressbuffer[0][3] ,
         \destinationAddressbuffer[0][2] , \destinationAddressbuffer[0][1] ,
         \destinationAddressbuffer[0][0] , \destinationAddressbuffer[1][11] ,
         \destinationAddressbuffer[1][10] , \destinationAddressbuffer[1][9] ,
         \destinationAddressbuffer[1][8] , \destinationAddressbuffer[1][7] ,
         \destinationAddressbuffer[1][6] , \destinationAddressbuffer[1][5] ,
         \destinationAddressbuffer[1][4] , \destinationAddressbuffer[1][3] ,
         \destinationAddressbuffer[1][2] , \destinationAddressbuffer[1][1] ,
         \destinationAddressbuffer[1][0] , \destinationAddressbuffer[2][11] ,
         \destinationAddressbuffer[2][10] , \destinationAddressbuffer[2][9] ,
         \destinationAddressbuffer[2][8] , \destinationAddressbuffer[2][7] ,
         \destinationAddressbuffer[2][6] , \destinationAddressbuffer[2][5] ,
         \destinationAddressbuffer[2][4] , \destinationAddressbuffer[2][3] ,
         \destinationAddressbuffer[2][2] , \destinationAddressbuffer[2][1] ,
         \destinationAddressbuffer[2][0] , \destinationAddressbuffer[3][11] ,
         \destinationAddressbuffer[3][10] , \destinationAddressbuffer[3][9] ,
         \destinationAddressbuffer[3][8] , \destinationAddressbuffer[3][7] ,
         \destinationAddressbuffer[3][6] , \destinationAddressbuffer[3][5] ,
         \destinationAddressbuffer[3][4] , \destinationAddressbuffer[3][3] ,
         \destinationAddressbuffer[3][2] , \destinationAddressbuffer[3][1] ,
         \destinationAddressbuffer[3][0] , \destinationAddressbuffer[4][11] ,
         \destinationAddressbuffer[4][10] , \destinationAddressbuffer[4][9] ,
         \destinationAddressbuffer[4][8] , \destinationAddressbuffer[4][7] ,
         \destinationAddressbuffer[4][6] , \destinationAddressbuffer[4][5] ,
         \destinationAddressbuffer[4][4] , \destinationAddressbuffer[4][3] ,
         \destinationAddressbuffer[4][2] , \destinationAddressbuffer[4][1] ,
         \destinationAddressbuffer[4][0] , \destinationAddressbuffer[5][11] ,
         \destinationAddressbuffer[5][10] , \destinationAddressbuffer[5][9] ,
         \destinationAddressbuffer[5][8] , \destinationAddressbuffer[5][7] ,
         \destinationAddressbuffer[5][6] , \destinationAddressbuffer[5][5] ,
         \destinationAddressbuffer[5][4] , \destinationAddressbuffer[5][3] ,
         \destinationAddressbuffer[5][2] , \destinationAddressbuffer[5][1] ,
         \destinationAddressbuffer[5][0] , \destinationAddressbuffer[6][11] ,
         \destinationAddressbuffer[6][10] , \destinationAddressbuffer[6][9] ,
         \destinationAddressbuffer[6][8] , \destinationAddressbuffer[6][7] ,
         \destinationAddressbuffer[6][6] , \destinationAddressbuffer[6][5] ,
         \destinationAddressbuffer[6][4] , \destinationAddressbuffer[6][3] ,
         \destinationAddressbuffer[6][2] , \destinationAddressbuffer[6][1] ,
         \destinationAddressbuffer[6][0] , \destinationAddressbuffer[7][11] ,
         \destinationAddressbuffer[7][10] , \destinationAddressbuffer[7][9] ,
         \destinationAddressbuffer[7][8] , \destinationAddressbuffer[7][7] ,
         \destinationAddressbuffer[7][6] , \destinationAddressbuffer[7][5] ,
         \destinationAddressbuffer[7][4] , \destinationAddressbuffer[7][3] ,
         \destinationAddressbuffer[7][2] , \destinationAddressbuffer[7][1] ,
         \destinationAddressbuffer[7][0] , \dataoutbuffer[7][5] ,
         \dataoutbuffer[7][4] , \dataoutbuffer[7][3] , \dataoutbuffer[7][2] ,
         \dataoutbuffer[7][1] , \dataoutbuffer[7][0] , \dataoutbuffer[6][5] ,
         \dataoutbuffer[6][4] , \dataoutbuffer[6][3] , \dataoutbuffer[6][2] ,
         \dataoutbuffer[6][1] , \dataoutbuffer[6][0] , \dataoutbuffer[5][5] ,
         \dataoutbuffer[5][4] , \dataoutbuffer[5][3] , \dataoutbuffer[5][2] ,
         \dataoutbuffer[5][1] , \dataoutbuffer[5][0] , \dataoutbuffer[4][5] ,
         \dataoutbuffer[4][4] , \dataoutbuffer[4][3] , \dataoutbuffer[4][2] ,
         \dataoutbuffer[4][1] , \dataoutbuffer[4][0] , \dataoutbuffer[3][5] ,
         \dataoutbuffer[3][4] , \dataoutbuffer[3][3] , \dataoutbuffer[3][2] ,
         \dataoutbuffer[3][1] , \dataoutbuffer[3][0] , \dataoutbuffer[2][5] ,
         \dataoutbuffer[2][4] , \dataoutbuffer[2][3] , \dataoutbuffer[2][2] ,
         \dataoutbuffer[2][1] , \dataoutbuffer[2][0] , \dataoutbuffer[1][5] ,
         \dataoutbuffer[1][4] , \dataoutbuffer[1][3] , \dataoutbuffer[1][2] ,
         \dataoutbuffer[1][1] , \dataoutbuffer[1][0] , \dataoutbuffer[0][5] ,
         \dataoutbuffer[0][4] , \dataoutbuffer[0][3] , \dataoutbuffer[0][2] ,
         \dataoutbuffer[0][1] , \dataoutbuffer[0][0] , empty_reg, N2624, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471;
  wire   [0:7] writeOutbuffer;
  wire   [0:7] readOutbuffer;
  wire   [2:0] read_reg;

  DFFNSRX1TS \readOutbuffer_reg[0]  ( .D(n1210), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[0]), .QN(n2471) );
  DFFNSRX1TS \readOutbuffer_reg[1]  ( .D(n1211), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[1]), .QN(n2470) );
  DFFNSRX1TS \readOutbuffer_reg[2]  ( .D(n1212), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[2]), .QN(n2469) );
  DFFNSRX1TS \readOutbuffer_reg[3]  ( .D(n1213), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[3]), .QN(n2468) );
  DFFNSRX1TS \readOutbuffer_reg[4]  ( .D(n1214), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[4]), .QN(n2467) );
  DFFNSRX1TS \readOutbuffer_reg[5]  ( .D(n1215), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[5]), .QN(n2466) );
  DFFNSRX1TS \readOutbuffer_reg[6]  ( .D(n1216), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[6]), .QN(n2465) );
  DFFNSRX1TS \readOutbuffer_reg[7]  ( .D(n1217), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[7]), .QN(n2464) );
  DFFNSRX1TS full_reg_reg ( .D(N2624), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(
        n2463) );
  DFFNSRX1TS \write_reg_reg[1]  ( .D(n1334), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(N374), .QN(n2462) );
  DFFNSRX1TS \read_reg_reg[1]  ( .D(n1330), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(read_reg[1]), .QN(n2461) );
  DFFNSRX1TS \read_reg_reg[0]  ( .D(n1336), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(read_reg[0]), .QN(n2460) );
  DFFNSRX1TS \write_reg_reg[2]  ( .D(n1333), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(N375), .QN(n2458) );
  DFFNSRX1TS \read_reg_reg[2]  ( .D(n1331), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(read_reg[2]), .QN(n2457) );
  DFFNSRX1TS \write_reg_reg[0]  ( .D(n1335), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(N373), .QN(n2456) );
  DFFNSRX1TS \requesterAddressbuffer_reg[2][0]  ( .D(n1285), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[2][1]  ( .D(n1284), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[2][2]  ( .D(n1283), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[2][3]  ( .D(n1282), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][0]  ( .D(n1149), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][1]  ( .D(n1148), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][2]  ( .D(n1147), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][3]  ( .D(n1146), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][0]  ( .D(n1273), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][1]  ( .D(n1272), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][2]  ( .D(n1271), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][3]  ( .D(n1270), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][4]  ( .D(n1269), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][5]  ( .D(n1268), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][5] ) );
  DFFNSRX1TS \writeOutbuffer_reg[7]  ( .D(n1225), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[7]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][4]  ( .D(n1205), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][5]  ( .D(n1204), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][6]  ( .D(n1203), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][7]  ( .D(n1202), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][8]  ( .D(n1201), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][9]  ( .D(n1200), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][10]  ( .D(n1199), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][11]  ( .D(n1198), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[6]  ( .D(n1224), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[6]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][4]  ( .D(n1193), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][5]  ( .D(n1192), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][6]  ( .D(n1191), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][7]  ( .D(n1190), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][8]  ( .D(n1189), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][9]  ( .D(n1188), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][10]  ( .D(n1187), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][11]  ( .D(n1186), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[3]  ( .D(n1221), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[3]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][4]  ( .D(n1157), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][5]  ( .D(n1156), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][6]  ( .D(n1155), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][7]  ( .D(n1154), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][8]  ( .D(n1153), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][9]  ( .D(n1152), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][10]  ( .D(n1151), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][11]  ( .D(n1150), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[2]  ( .D(n1220), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[2]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][4]  ( .D(n1145), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][5]  ( .D(n1144), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][6]  ( .D(n1143), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][7]  ( .D(n1142), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][8]  ( .D(n1141), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][9]  ( .D(n1140), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][10]  ( .D(n1139), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][11]  ( .D(n1138), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][11] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][0]  ( .D(n1231), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][1]  ( .D(n1230), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][2]  ( .D(n1229), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][3]  ( .D(n1228), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][4]  ( .D(n1227), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][5]  ( .D(n1226), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][0]  ( .D(n1237), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][1]  ( .D(n1236), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][2]  ( .D(n1235), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][3]  ( .D(n1234), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][4]  ( .D(n1233), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][5]  ( .D(n1232), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][5] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[5][0]  ( .D(n1297), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[5][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[5][1]  ( .D(n1296), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[5][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[5][2]  ( .D(n1295), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[5][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[5][3]  ( .D(n1294), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[5][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][0]  ( .D(n1185), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][1]  ( .D(n1184), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][2]  ( .D(n1183), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][3]  ( .D(n1182), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[4][0]  ( .D(n1293), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[4][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[4][1]  ( .D(n1292), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[4][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[4][2]  ( .D(n1291), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[4][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[4][3]  ( .D(n1290), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[4][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][0]  ( .D(n1173), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][1]  ( .D(n1172), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][2]  ( .D(n1171), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][3]  ( .D(n1170), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][0]  ( .D(n1255), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][1]  ( .D(n1254), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][2]  ( .D(n1253), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][3]  ( .D(n1252), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][4]  ( .D(n1251), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][5]  ( .D(n1250), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][0]  ( .D(n1261), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][1]  ( .D(n1260), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][2]  ( .D(n1259), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][3]  ( .D(n1258), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][4]  ( .D(n1257), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][5]  ( .D(n1256), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][5] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[1][0]  ( .D(n1281), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[1][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[1][1]  ( .D(n1280), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[1][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[1][2]  ( .D(n1279), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[1][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[1][3]  ( .D(n1278), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[1][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][0]  ( .D(n1137), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][1]  ( .D(n1136), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][2]  ( .D(n1135), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][3]  ( .D(n1134), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[0][0]  ( .D(n1277), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[0][1]  ( .D(n1276), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[0][2]  ( .D(n1275), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[0][3]  ( .D(n1274), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][0]  ( .D(n1125), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][1]  ( .D(n1124), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][2]  ( .D(n1123), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][3]  ( .D(n1122), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[7][0]  ( .D(n1305), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[7][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[7][1]  ( .D(n1304), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[7][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[7][2]  ( .D(n1303), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[7][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[7][3]  ( .D(n1302), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[7][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][0]  ( .D(n1209), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][1]  ( .D(n1208), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][2]  ( .D(n1207), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][3]  ( .D(n1206), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[6][0]  ( .D(n1301), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[6][1]  ( .D(n1300), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[6][2]  ( .D(n1299), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[6][3]  ( .D(n1298), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][0]  ( .D(n1197), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][1]  ( .D(n1196), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][2]  ( .D(n1195), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][3]  ( .D(n1194), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][0]  ( .D(n1243), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][1]  ( .D(n1242), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][2]  ( .D(n1241), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][3]  ( .D(n1240), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][4]  ( .D(n1239), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][5]  ( .D(n1238), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][0]  ( .D(n1249), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][1]  ( .D(n1248), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][2]  ( .D(n1247), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][3]  ( .D(n1246), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][4]  ( .D(n1245), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][5]  ( .D(n1244), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][5] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[3][0]  ( .D(n1289), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[3][1]  ( .D(n1288), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[3][2]  ( .D(n1287), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[3][3]  ( .D(n1286), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][0]  ( .D(n1161), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][1]  ( .D(n1160), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][2]  ( .D(n1159), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][3]  ( .D(n1158), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][0]  ( .D(n1267), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][1]  ( .D(n1266), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][2]  ( .D(n1265), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][3]  ( .D(n1264), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][4]  ( .D(n1263), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][5]  ( .D(n1262), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][5] ) );
  DFFNSRX1TS \writeOutbuffer_reg[5]  ( .D(n1223), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[5]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][4]  ( .D(n1181), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][5]  ( .D(n1180), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][6]  ( .D(n1179), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][7]  ( .D(n1178), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][8]  ( .D(n1177), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][9]  ( .D(n1176), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][10]  ( .D(n1175), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][11]  ( .D(n1174), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[4]  ( .D(n1222), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[4]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][4]  ( .D(n1169), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][5]  ( .D(n1168), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][6]  ( .D(n1167), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][7]  ( .D(n1166), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][8]  ( .D(n1165), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][9]  ( .D(n1164), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][10]  ( .D(n1163), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][11]  ( .D(n1162), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[1]  ( .D(n1219), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[1]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][4]  ( .D(n1133), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][5]  ( .D(n1132), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][6]  ( .D(n1131), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][7]  ( .D(n1130), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][8]  ( .D(n1129), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][9]  ( .D(n1128), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][10]  ( .D(n1127), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][11]  ( .D(n1126), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[0]  ( .D(n1218), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[0]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][4]  ( .D(n1121), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][5]  ( .D(n1120), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][6]  ( .D(n1119), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][7]  ( .D(n1118), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][8]  ( .D(n1117), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][9]  ( .D(n1116), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][10]  ( .D(n1115), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][11]  ( .D(n1114), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][11] ) );
  DFFNSRX1TS writeOut_reg ( .D(n1328), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        writeOut) );
  DFFNSRX1TS \destinationAddressOut_reg[4]  ( .D(n1319), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[4]) );
  DFFNSRX1TS \destinationAddressOut_reg[5]  ( .D(n1318), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[5]) );
  DFFNSRX1TS \destinationAddressOut_reg[6]  ( .D(n1317), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[6]) );
  DFFNSRX1TS \destinationAddressOut_reg[7]  ( .D(n1316), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[7]) );
  DFFNSRX1TS \destinationAddressOut_reg[8]  ( .D(n1315), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[8]) );
  DFFNSRX1TS \destinationAddressOut_reg[9]  ( .D(n1314), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[9]) );
  DFFNSRX1TS \destinationAddressOut_reg[10]  ( .D(n1313), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[10]) );
  DFFNSRX1TS \destinationAddressOut_reg[11]  ( .D(n1312), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[11]) );
  DFFNSRX1TS readOut_reg ( .D(n1329), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        readOut) );
  DFFNSRX1TS \requesterAddressOut_reg[0]  ( .D(n1327), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[0]) );
  DFFNSRX1TS \requesterAddressOut_reg[1]  ( .D(n1326), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[1]) );
  DFFNSRX1TS \requesterAddressOut_reg[2]  ( .D(n1325), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[2]) );
  DFFNSRX1TS \requesterAddressOut_reg[3]  ( .D(n1324), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[3]) );
  DFFNSRX1TS \destinationAddressOut_reg[0]  ( .D(n1323), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[0]) );
  DFFNSRX1TS \destinationAddressOut_reg[1]  ( .D(n1322), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[1]) );
  DFFNSRX1TS \destinationAddressOut_reg[2]  ( .D(n1321), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[2]) );
  DFFNSRX1TS \destinationAddressOut_reg[3]  ( .D(n1320), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[3]) );
  DFFNSRX1TS \dataOut_reg[0]  ( .D(n1311), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[0]) );
  DFFNSRX1TS \dataOut_reg[1]  ( .D(n1310), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[1]) );
  DFFNSRX1TS \dataOut_reg[2]  ( .D(n1309), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[2]) );
  DFFNSRX1TS \dataOut_reg[3]  ( .D(n1308), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[3]) );
  DFFNSRX1TS \dataOut_reg[4]  ( .D(n1307), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[4]) );
  DFFNSRX1TS \dataOut_reg[5]  ( .D(n1306), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[5]) );
  DFFNSRX2TS empty_reg_reg ( .D(n1332), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        empty_reg), .QN(n2459) );
  NOR2XLTS U1343 ( .A(n2456), .B(n1339), .Y(n1600) );
  NOR2XLTS U1344 ( .A(n1338), .B(n1340), .Y(n1698) );
  NOR2X2TS U1345 ( .A(n2271), .B(n1512), .Y(n1510) );
  NAND2BXLTS U1346 ( .AN(n1426), .B(n1344), .Y(n1504) );
  NAND2BXLTS U1347 ( .AN(n1532), .B(n1342), .Y(n1503) );
  NOR2X1TS U1348 ( .A(n1352), .B(n1341), .Y(n1598) );
  OAI21XLTS U1349 ( .A0(n1600), .A1(N374), .B0(n1353), .Y(n1597) );
  NOR2X2TS U1350 ( .A(n2459), .B(n1687), .Y(n1877) );
  NOR2X2TS U1351 ( .A(n2459), .B(n1688), .Y(n1682) );
  NOR2X2TS U1352 ( .A(read_reg[2]), .B(n1691), .Y(n1969) );
  NOR2X2TS U1353 ( .A(n1691), .B(n2457), .Y(n1971) );
  NAND2BXLTS U1354 ( .AN(n1456), .B(n1455), .Y(n1458) );
  NAND2BXLTS U1355 ( .AN(n1569), .B(n1568), .Y(n1570) );
  NAND2BXLTS U1356 ( .AN(n1537), .B(n1536), .Y(n1539) );
  NAND2BXLTS U1357 ( .AN(n1430), .B(n1429), .Y(n1431) );
  NOR2XLTS U1358 ( .A(n2232), .B(n2229), .Y(n1361) );
  NOR2XLTS U1359 ( .A(n2276), .B(n2273), .Y(n1508) );
  NAND2BXLTS U1360 ( .AN(n1604), .B(n1603), .Y(n1605) );
  NAND2BXLTS U1361 ( .AN(n1512), .B(n1508), .Y(n1511) );
  NAND2BXLTS U1362 ( .AN(n1362), .B(n1361), .Y(n1365) );
  NAND2BXLTS U1363 ( .AN(n1481), .B(n1480), .Y(n1483) );
  NOR2XLTS U1364 ( .A(n1452), .B(n1597), .Y(n1354) );
  NAND3XLTS U1365 ( .A(n1698), .B(empty_reg), .C(n1697), .Y(n1721) );
  NOR3XLTS U1366 ( .A(n1344), .B(n1346), .C(n1343), .Y(n1686) );
  NOR3XLTS U1367 ( .A(n1342), .B(n1346), .C(n1345), .Y(n1685) );
  CLKAND2X2TS U1368 ( .A(n1690), .B(n1978), .Y(n1707) );
  NOR2XLTS U1369 ( .A(n2292), .B(n1458), .Y(n1457) );
  NOR2XLTS U1370 ( .A(n2259), .B(n1570), .Y(n1571) );
  NOR2XLTS U1371 ( .A(n2237), .B(n1539), .Y(n1538) );
  NOR2XLTS U1372 ( .A(n2303), .B(n1431), .Y(n1432) );
  CLKBUFX2TS U1373 ( .A(n1482), .Y(n2416) );
  NOR2XLTS U1374 ( .A(n2281), .B(n1483), .Y(n1482) );
  XOR2XLTS U1375 ( .A(n1658), .B(n1657), .Y(n1670) );
  CLKAND2X2TS U1376 ( .A(n1655), .B(n1653), .Y(n1659) );
  NOR2XLTS U1377 ( .A(n1349), .B(n1634), .Y(n1671) );
  NAND4XLTS U1378 ( .A(n1596), .B(n1561), .C(n1532), .D(n1342), .Y(n2230) );
  NAND3XLTS U1379 ( .A(N374), .B(n1599), .C(n1598), .Y(n2225) );
  INVX2TS U1380 ( .A(n2229), .Y(n2227) );
  INVX2TS U1381 ( .A(n2243), .Y(n2241) );
  INVX2TS U1382 ( .A(n2240), .Y(n2238) );
  NAND3XLTS U1383 ( .A(n1599), .B(n1598), .C(n1597), .Y(n2247) );
  INVX2TS U1384 ( .A(n2254), .Y(n2252) );
  INVX2TS U1385 ( .A(n2251), .Y(n2249) );
  INVX2TS U1386 ( .A(n2265), .Y(n2263) );
  INVX2TS U1387 ( .A(n2262), .Y(n2260) );
  NAND2X1TS U1388 ( .A(n1354), .B(n1562), .Y(n2269) );
  INVX2TS U1389 ( .A(n2269), .Y(n2270) );
  INVX2TS U1390 ( .A(n2276), .Y(n2274) );
  INVX2TS U1391 ( .A(n2287), .Y(n2285) );
  INVX2TS U1392 ( .A(n2284), .Y(n2282) );
  INVX2TS U1393 ( .A(n2298), .Y(n2296) );
  INVX2TS U1394 ( .A(n2295), .Y(n2293) );
  INVX2TS U1395 ( .A(n2310), .Y(n2308) );
  INVX2TS U1396 ( .A(n2307), .Y(n2304) );
  ADDFX1TS U1397 ( .A(read_reg[1]), .B(n2462), .CI(n1639), .CO(n1635), .S(
        n1644) );
  NOR3XLTS U1398 ( .A(n1342), .B(n1344), .C(n1346), .Y(n1681) );
  XOR2XLTS U1399 ( .A(n1635), .B(n1636), .Y(n1650) );
  NOR2XLTS U1400 ( .A(n2243), .B(n2240), .Y(n1536) );
  NOR2XLTS U1401 ( .A(n2254), .B(n2251), .Y(n1603) );
  NOR2XLTS U1402 ( .A(n2265), .B(n2262), .Y(n1568) );
  NOR2XLTS U1403 ( .A(n2287), .B(n2284), .Y(n1480) );
  NOR2XLTS U1404 ( .A(n2298), .B(n2295), .Y(n1455) );
  ADDFX1TS U1405 ( .A(n1340), .B(n1338), .CI(n1344), .CO(n1641), .S(n1638) );
  NOR2XLTS U1406 ( .A(n2310), .B(n2307), .Y(n1429) );
  AO21XLTS U1407 ( .A0(n2456), .A1(n1339), .B0(n1600), .Y(n1352) );
  OAI21XLTS U1408 ( .A0(n1354), .A1(n1562), .B0(n2269), .Y(n1426) );
  NOR3BXLTS U1409 ( .AN(n1346), .B(n1342), .C(n1344), .Y(n1697) );
  NAND3XLTS U1410 ( .A(n1340), .B(n1681), .C(n1339), .Y(n1687) );
  NAND3XLTS U1411 ( .A(n1338), .B(n1681), .C(n1341), .Y(n1688) );
  ADDFX1TS U1412 ( .A(n1342), .B(n1346), .CI(n1638), .CO(n1640), .S(n1653) );
  AOI211XLTS U1413 ( .A0(n1650), .A1(n1649), .B0(n1648), .C0(n1647), .Y(n1651)
         );
  XOR2XLTS U1414 ( .A(N375), .B(n1356), .Y(n1532) );
  AOI31XLTS U1415 ( .A0(n1361), .A1(n1357), .A2(n2225), .B0(n1634), .Y(n1359)
         );
  AOI31XLTS U1416 ( .A0(n1603), .A1(n2247), .A2(n1601), .B0(n1634), .Y(n1602)
         );
  NAND3XLTS U1417 ( .A(n1600), .B(N375), .C(n2462), .Y(n1601) );
  AOI31XLTS U1418 ( .A0(n1508), .A1(n2269), .A2(n1507), .B0(n1634), .Y(n1509)
         );
  INVX2TS U1419 ( .A(n1561), .Y(n1595) );
  NOR2XLTS U1420 ( .A(n1598), .B(n1597), .Y(n1592) );
  ADDFX1TS U1421 ( .A(n1641), .B(N374), .CI(n1355), .CO(n1356), .S(n1596) );
  INVX2TS U1422 ( .A(n1562), .Y(n1599) );
  INVX2TS U1423 ( .A(n1597), .Y(n1564) );
  OAI21XLTS U1424 ( .A0(n1340), .A1(n1352), .B0(n1563), .Y(n1559) );
  ADDFX1TS U1425 ( .A(n1661), .B(N374), .CI(n1660), .CO(n1656), .S(n1669) );
  CLKAND2X2TS U1426 ( .A(n1655), .B(n1654), .Y(n1660) );
  NOR2XLTS U1427 ( .A(n1667), .B(n1349), .Y(n1672) );
  NAND4XLTS U1428 ( .A(N373), .B(N374), .C(N375), .D(n1346), .Y(n2233) );
  NOR2XLTS U1429 ( .A(n1505), .B(n1591), .Y(n2229) );
  NAND4XLTS U1430 ( .A(N374), .B(N375), .C(n1346), .D(n2456), .Y(n2244) );
  NOR3XLTS U1431 ( .A(n1560), .B(n1591), .C(n1559), .Y(n2240) );
  NOR3XLTS U1432 ( .A(n1596), .B(n1595), .C(n1594), .Y(n2254) );
  NAND4XLTS U1433 ( .A(N373), .B(N375), .C(n1346), .D(n2462), .Y(n2255) );
  NOR3XLTS U1434 ( .A(n1593), .B(n1592), .C(n1591), .Y(n2251) );
  NAND4XLTS U1435 ( .A(N375), .B(n1346), .C(n2456), .D(n2462), .Y(n2266) );
  NOR3XLTS U1436 ( .A(n1564), .B(n1563), .C(n1562), .Y(n2259) );
  NOR3BXLTS U1437 ( .AN(n1560), .B(n1591), .C(n1559), .Y(n2262) );
  NOR3XLTS U1438 ( .A(n1533), .B(n1595), .C(n1503), .Y(n2276) );
  NAND4XLTS U1439 ( .A(N374), .B(N373), .C(n1346), .D(n2458), .Y(n2277) );
  NOR2XLTS U1440 ( .A(n1505), .B(n1504), .Y(n2273) );
  INVX2TS U1441 ( .A(n2273), .Y(n2271) );
  NAND4XLTS U1442 ( .A(N374), .B(n1346), .C(n2456), .D(n2458), .Y(n2288) );
  NOR3XLTS U1443 ( .A(n1599), .B(n1563), .C(n1597), .Y(n2281) );
  NOR3XLTS U1444 ( .A(n1560), .B(n1559), .C(n1504), .Y(n2284) );
  NOR3XLTS U1445 ( .A(n1596), .B(n1595), .C(n1503), .Y(n2298) );
  NAND4XLTS U1446 ( .A(N373), .B(n1346), .C(n2458), .D(n2462), .Y(n2299) );
  NOR3XLTS U1447 ( .A(n1599), .B(n1564), .C(n1452), .Y(n2292) );
  NOR3XLTS U1448 ( .A(n1593), .B(n1592), .C(n1504), .Y(n2295) );
  NAND4XLTS U1449 ( .A(n1346), .B(n2456), .C(n2462), .D(n2458), .Y(n2311) );
  NOR3XLTS U1450 ( .A(n1599), .B(n1564), .C(n1563), .Y(n2303) );
  NOR3BXLTS U1451 ( .AN(n1560), .B(n1504), .C(n1559), .Y(n2307) );
  NAND4XLTS U1452 ( .A(n1984), .B(n1983), .C(n1982), .D(n1981), .Y(n1306) );
  NAND4XLTS U1453 ( .A(n1958), .B(n1957), .C(n1956), .D(n1955), .Y(n1307) );
  NAND4XLTS U1454 ( .A(n1944), .B(n1943), .C(n1942), .D(n1941), .Y(n1308) );
  NAND4XLTS U1455 ( .A(n1930), .B(n1929), .C(n1928), .D(n1927), .Y(n1309) );
  NAND4XLTS U1456 ( .A(n1915), .B(n1914), .C(n1913), .D(n1912), .Y(n1310) );
  NAND4XLTS U1457 ( .A(n1901), .B(n1900), .C(n1899), .D(n1898), .Y(n1311) );
  NAND4XLTS U1458 ( .A(n1816), .B(n1815), .C(n1814), .D(n1813), .Y(n1320) );
  NAND4XLTS U1459 ( .A(n1803), .B(n1802), .C(n1801), .D(n1800), .Y(n1321) );
  NAND4XLTS U1460 ( .A(n1790), .B(n1789), .C(n1788), .D(n1787), .Y(n1322) );
  NAND4XLTS U1461 ( .A(n1776), .B(n1775), .C(n1774), .D(n1773), .Y(n1323) );
  NAND4XLTS U1462 ( .A(n1763), .B(n1762), .C(n1761), .D(n1813), .Y(n1324) );
  NAND4XLTS U1463 ( .A(n1750), .B(n1749), .C(n1748), .D(n1800), .Y(n1325) );
  NAND4XLTS U1464 ( .A(n1737), .B(n1736), .C(n1735), .D(n1787), .Y(n1326) );
  NAND4XLTS U1465 ( .A(n1724), .B(n1723), .C(n1722), .D(n1773), .Y(n1327) );
  NAND4XLTS U1466 ( .A(n1701), .B(n1700), .C(n1699), .D(n1721), .Y(n1329) );
  NAND3XLTS U1467 ( .A(n1885), .B(n1884), .C(n1883), .Y(n1312) );
  NAND3XLTS U1468 ( .A(n1876), .B(n1875), .C(n1874), .Y(n1313) );
  NAND3XLTS U1469 ( .A(n1868), .B(n1867), .C(n1866), .Y(n1314) );
  NAND3XLTS U1470 ( .A(n1860), .B(n1859), .C(n1858), .Y(n1315) );
  NAND3XLTS U1471 ( .A(n1852), .B(n1851), .C(n1850), .Y(n1316) );
  NAND3XLTS U1472 ( .A(n1844), .B(n1843), .C(n1842), .Y(n1317) );
  NAND3XLTS U1473 ( .A(n1836), .B(n1835), .C(n1834), .Y(n1318) );
  NAND3XLTS U1474 ( .A(n1828), .B(n1827), .C(n1826), .Y(n1319) );
  NAND3XLTS U1475 ( .A(n1710), .B(n1709), .C(n1708), .Y(n1328) );
  OAI211XLTS U1476 ( .A0(n1451), .A1(n1617), .B0(n1434), .C0(n1433), .Y(n1114)
         );
  OAI211XLTS U1477 ( .A0(n1451), .A1(n1608), .B0(n1450), .C0(n1449), .Y(n1115)
         );
  OAI211XLTS U1478 ( .A0(n1451), .A1(n1611), .B0(n1438), .C0(n1437), .Y(n1116)
         );
  OAI211XLTS U1479 ( .A0(n1451), .A1(n1632), .B0(n1436), .C0(n1435), .Y(n1117)
         );
  OAI211XLTS U1480 ( .A0(n1451), .A1(n1614), .B0(n1440), .C0(n1439), .Y(n1118)
         );
  OAI211XLTS U1481 ( .A0(n1451), .A1(n1626), .B0(n1442), .C0(n1441), .Y(n1119)
         );
  OAI211XLTS U1482 ( .A0(n1451), .A1(n1629), .B0(n1444), .C0(n1443), .Y(n1120)
         );
  OAI211XLTS U1483 ( .A0(n1451), .A1(n1620), .B0(n1446), .C0(n1445), .Y(n1121)
         );
  OAI211XLTS U1484 ( .A0(n1451), .A1(n1623), .B0(n1448), .C0(n1447), .Y(n1218)
         );
  OAI211XLTS U1485 ( .A0(n1477), .A1(n1617), .B0(n1460), .C0(n1459), .Y(n1126)
         );
  OAI211XLTS U1486 ( .A0(n1477), .A1(n1608), .B0(n1472), .C0(n1471), .Y(n1127)
         );
  OAI211XLTS U1487 ( .A0(n1477), .A1(n1611), .B0(n1464), .C0(n1463), .Y(n1128)
         );
  OAI211XLTS U1488 ( .A0(n1477), .A1(n1632), .B0(n1462), .C0(n1461), .Y(n1129)
         );
  OAI211XLTS U1489 ( .A0(n1477), .A1(n1614), .B0(n1468), .C0(n1467), .Y(n1130)
         );
  OAI211XLTS U1490 ( .A0(n1477), .A1(n1626), .B0(n1470), .C0(n1469), .Y(n1131)
         );
  OAI211XLTS U1491 ( .A0(n1477), .A1(n1629), .B0(n1476), .C0(n1475), .Y(n1132)
         );
  OAI211XLTS U1492 ( .A0(n1477), .A1(n1620), .B0(n1474), .C0(n1473), .Y(n1133)
         );
  OAI211XLTS U1493 ( .A0(n1477), .A1(n1623), .B0(n1466), .C0(n1465), .Y(n1219)
         );
  OAI211XLTS U1494 ( .A0(n1590), .A1(n1617), .B0(n1575), .C0(n1574), .Y(n1162)
         );
  OAI211XLTS U1495 ( .A0(n1590), .A1(n1608), .B0(n1573), .C0(n1572), .Y(n1163)
         );
  OAI211XLTS U1496 ( .A0(n1590), .A1(n1611), .B0(n1579), .C0(n1578), .Y(n1164)
         );
  OAI211XLTS U1497 ( .A0(n1590), .A1(n1632), .B0(n1583), .C0(n1582), .Y(n1165)
         );
  OAI211XLTS U1498 ( .A0(n1590), .A1(n1614), .B0(n1587), .C0(n1586), .Y(n1166)
         );
  OAI211XLTS U1499 ( .A0(n1590), .A1(n1626), .B0(n1585), .C0(n1584), .Y(n1167)
         );
  OAI211XLTS U1500 ( .A0(n1590), .A1(n1629), .B0(n1589), .C0(n1588), .Y(n1168)
         );
  OAI211XLTS U1501 ( .A0(n1590), .A1(n1620), .B0(n1577), .C0(n1576), .Y(n1169)
         );
  OAI211XLTS U1502 ( .A0(n1590), .A1(n1623), .B0(n1581), .C0(n1580), .Y(n1222)
         );
  OAI211XLTS U1503 ( .A0(n1633), .A1(n1617), .B0(n1616), .C0(n1615), .Y(n1174)
         );
  OAI211XLTS U1504 ( .A0(n1633), .A1(n1608), .B0(n1607), .C0(n1606), .Y(n1175)
         );
  OAI211XLTS U1505 ( .A0(n1633), .A1(n1611), .B0(n1610), .C0(n1609), .Y(n1176)
         );
  OAI211XLTS U1506 ( .A0(n1633), .A1(n1632), .B0(n1631), .C0(n1630), .Y(n1177)
         );
  OAI211XLTS U1507 ( .A0(n1633), .A1(n1614), .B0(n1613), .C0(n1612), .Y(n1178)
         );
  OAI211XLTS U1508 ( .A0(n1633), .A1(n1626), .B0(n1625), .C0(n1624), .Y(n1179)
         );
  OAI211XLTS U1509 ( .A0(n1633), .A1(n1629), .B0(n1628), .C0(n1627), .Y(n1180)
         );
  OAI211XLTS U1510 ( .A0(n1633), .A1(n1620), .B0(n1619), .C0(n1618), .Y(n1181)
         );
  OAI211XLTS U1511 ( .A0(n1633), .A1(n1623), .B0(n1622), .C0(n1621), .Y(n1223)
         );
  NAND3XLTS U1512 ( .A(n2116), .B(n2115), .C(n2114), .Y(n1262) );
  NAND3XLTS U1513 ( .A(n2113), .B(n2112), .C(n2111), .Y(n1263) );
  NAND3XLTS U1514 ( .A(n2110), .B(n2109), .C(n2108), .Y(n1264) );
  NAND3XLTS U1515 ( .A(n2107), .B(n2106), .C(n2105), .Y(n1265) );
  NAND3XLTS U1516 ( .A(n2104), .B(n2103), .C(n2102), .Y(n1266) );
  NAND3XLTS U1517 ( .A(n2101), .B(n2100), .C(n2099), .Y(n1267) );
  NAND3XLTS U1518 ( .A(n2401), .B(n2400), .C(n2399), .Y(n1158) );
  NAND3XLTS U1519 ( .A(n2393), .B(n2392), .C(n2391), .Y(n1159) );
  NAND3XLTS U1520 ( .A(n2390), .B(n2389), .C(n2388), .Y(n1160) );
  NAND3XLTS U1521 ( .A(n2387), .B(n2386), .C(n2385), .Y(n1161) );
  NAND3XLTS U1522 ( .A(n2044), .B(n2043), .C(n2042), .Y(n1286) );
  NAND3XLTS U1523 ( .A(n2041), .B(n2040), .C(n2039), .Y(n1287) );
  NAND3XLTS U1524 ( .A(n2038), .B(n2037), .C(n2036), .Y(n1288) );
  NAND3XLTS U1525 ( .A(n2035), .B(n2034), .C(n2033), .Y(n1289) );
  NAND3XLTS U1526 ( .A(n2170), .B(n2169), .C(n2168), .Y(n1244) );
  NAND3XLTS U1527 ( .A(n2167), .B(n2166), .C(n2165), .Y(n1245) );
  NAND3XLTS U1528 ( .A(n2164), .B(n2163), .C(n2162), .Y(n1246) );
  NAND3XLTS U1529 ( .A(n2161), .B(n2160), .C(n2159), .Y(n1247) );
  NAND3XLTS U1530 ( .A(n2158), .B(n2157), .C(n2156), .Y(n1248) );
  NAND3XLTS U1531 ( .A(n2155), .B(n2154), .C(n2153), .Y(n1249) );
  NAND3XLTS U1532 ( .A(n2188), .B(n2187), .C(n2186), .Y(n1238) );
  NAND3XLTS U1533 ( .A(n2185), .B(n2184), .C(n2183), .Y(n1239) );
  NAND3XLTS U1534 ( .A(n2182), .B(n2181), .C(n2180), .Y(n1240) );
  NAND3XLTS U1535 ( .A(n2179), .B(n2178), .C(n2177), .Y(n1241) );
  NAND3XLTS U1536 ( .A(n2176), .B(n2175), .C(n2174), .Y(n1242) );
  NAND3XLTS U1537 ( .A(n2173), .B(n2172), .C(n2171), .Y(n1243) );
  NAND3XLTS U1538 ( .A(n2349), .B(n2348), .C(n2347), .Y(n1194) );
  NAND3XLTS U1539 ( .A(n2340), .B(n2339), .C(n2338), .Y(n1195) );
  NAND3XLTS U1540 ( .A(n2337), .B(n2336), .C(n2335), .Y(n1196) );
  NAND3XLTS U1541 ( .A(n2334), .B(n2333), .C(n2332), .Y(n1197) );
  NAND3XLTS U1542 ( .A(n2008), .B(n2007), .C(n2006), .Y(n1298) );
  NAND3XLTS U1543 ( .A(n2005), .B(n2004), .C(n2003), .Y(n1299) );
  NAND3XLTS U1544 ( .A(n2002), .B(n2001), .C(n2000), .Y(n1300) );
  NAND3XLTS U1545 ( .A(n1999), .B(n1998), .C(n1997), .Y(n1301) );
  NAND3XLTS U1546 ( .A(n2331), .B(n2330), .C(n2329), .Y(n1206) );
  NAND3XLTS U1547 ( .A(n2322), .B(n2321), .C(n2320), .Y(n1207) );
  NAND3XLTS U1548 ( .A(n2319), .B(n2318), .C(n2317), .Y(n1208) );
  NAND3XLTS U1549 ( .A(n2316), .B(n2315), .C(n2314), .Y(n1209) );
  NAND3XLTS U1550 ( .A(n1996), .B(n1995), .C(n1994), .Y(n1302) );
  NAND3XLTS U1551 ( .A(n1993), .B(n1992), .C(n1991), .Y(n1303) );
  NAND3XLTS U1552 ( .A(n1990), .B(n1989), .C(n1988), .Y(n1304) );
  NAND3XLTS U1553 ( .A(n1987), .B(n1986), .C(n1985), .Y(n1305) );
  NAND3XLTS U1554 ( .A(n2455), .B(n2454), .C(n2453), .Y(n1122) );
  NAND3XLTS U1555 ( .A(n2446), .B(n2445), .C(n2444), .Y(n1123) );
  NAND3XLTS U1556 ( .A(n2443), .B(n2442), .C(n2441), .Y(n1124) );
  NAND3XLTS U1557 ( .A(n2440), .B(n2439), .C(n2438), .Y(n1125) );
  NAND3XLTS U1558 ( .A(n2080), .B(n2079), .C(n2078), .Y(n1274) );
  NAND3XLTS U1559 ( .A(n2077), .B(n2076), .C(n2075), .Y(n1275) );
  NAND3XLTS U1560 ( .A(n2074), .B(n2073), .C(n2072), .Y(n1276) );
  NAND3XLTS U1561 ( .A(n2071), .B(n2070), .C(n2069), .Y(n1277) );
  NAND3XLTS U1562 ( .A(n2437), .B(n2436), .C(n2435), .Y(n1134) );
  NAND3XLTS U1563 ( .A(n2428), .B(n2427), .C(n2426), .Y(n1135) );
  NAND3XLTS U1564 ( .A(n2425), .B(n2424), .C(n2423), .Y(n1136) );
  NAND3XLTS U1565 ( .A(n2422), .B(n2421), .C(n2420), .Y(n1137) );
  NAND3XLTS U1566 ( .A(n2068), .B(n2067), .C(n2066), .Y(n1278) );
  NAND3XLTS U1567 ( .A(n2065), .B(n2064), .C(n2063), .Y(n1279) );
  NAND3XLTS U1568 ( .A(n2062), .B(n2061), .C(n2060), .Y(n1280) );
  NAND3XLTS U1569 ( .A(n2059), .B(n2058), .C(n2057), .Y(n1281) );
  NAND3XLTS U1570 ( .A(n2134), .B(n2133), .C(n2132), .Y(n1256) );
  NAND3XLTS U1571 ( .A(n2131), .B(n2130), .C(n2129), .Y(n1257) );
  NAND3XLTS U1572 ( .A(n2128), .B(n2127), .C(n2126), .Y(n1258) );
  NAND3XLTS U1573 ( .A(n2125), .B(n2124), .C(n2123), .Y(n1259) );
  NAND3XLTS U1574 ( .A(n2122), .B(n2121), .C(n2120), .Y(n1260) );
  NAND3XLTS U1575 ( .A(n2119), .B(n2118), .C(n2117), .Y(n1261) );
  NAND3XLTS U1576 ( .A(n2152), .B(n2151), .C(n2150), .Y(n1250) );
  NAND3XLTS U1577 ( .A(n2149), .B(n2148), .C(n2147), .Y(n1251) );
  NAND3XLTS U1578 ( .A(n2146), .B(n2145), .C(n2144), .Y(n1252) );
  NAND3XLTS U1579 ( .A(n2143), .B(n2142), .C(n2141), .Y(n1253) );
  NAND3XLTS U1580 ( .A(n2140), .B(n2139), .C(n2138), .Y(n1254) );
  NAND3XLTS U1581 ( .A(n2137), .B(n2136), .C(n2135), .Y(n1255) );
  NAND3XLTS U1582 ( .A(n2384), .B(n2383), .C(n2382), .Y(n1170) );
  NAND3XLTS U1583 ( .A(n2375), .B(n2374), .C(n2373), .Y(n1171) );
  NAND3XLTS U1584 ( .A(n2372), .B(n2371), .C(n2370), .Y(n1172) );
  NAND3XLTS U1585 ( .A(n2369), .B(n2368), .C(n2367), .Y(n1173) );
  NAND3XLTS U1586 ( .A(n2032), .B(n2031), .C(n2030), .Y(n1290) );
  NAND3XLTS U1587 ( .A(n2029), .B(n2028), .C(n2027), .Y(n1291) );
  NAND3XLTS U1588 ( .A(n2026), .B(n2025), .C(n2024), .Y(n1292) );
  NAND3XLTS U1589 ( .A(n2023), .B(n2022), .C(n2021), .Y(n1293) );
  NAND3XLTS U1590 ( .A(n2366), .B(n2365), .C(n2364), .Y(n1182) );
  NAND3XLTS U1591 ( .A(n2358), .B(n2357), .C(n2356), .Y(n1183) );
  NAND3XLTS U1592 ( .A(n2355), .B(n2354), .C(n2353), .Y(n1184) );
  NAND3XLTS U1593 ( .A(n2352), .B(n2351), .C(n2350), .Y(n1185) );
  NAND3XLTS U1594 ( .A(n2020), .B(n2019), .C(n2018), .Y(n1294) );
  NAND3XLTS U1595 ( .A(n2017), .B(n2016), .C(n2015), .Y(n1295) );
  NAND3XLTS U1596 ( .A(n2014), .B(n2013), .C(n2012), .Y(n1296) );
  NAND3XLTS U1597 ( .A(n2011), .B(n2010), .C(n2009), .Y(n1297) );
  NAND3XLTS U1598 ( .A(n2206), .B(n2205), .C(n2204), .Y(n1232) );
  NAND3XLTS U1599 ( .A(n2203), .B(n2202), .C(n2201), .Y(n1233) );
  NAND3XLTS U1600 ( .A(n2200), .B(n2199), .C(n2198), .Y(n1234) );
  NAND3XLTS U1601 ( .A(n2197), .B(n2196), .C(n2195), .Y(n1235) );
  NAND3XLTS U1602 ( .A(n2194), .B(n2193), .C(n2192), .Y(n1236) );
  NAND3XLTS U1603 ( .A(n2191), .B(n2190), .C(n2189), .Y(n1237) );
  NAND3XLTS U1604 ( .A(n2224), .B(n2223), .C(n2222), .Y(n1226) );
  NAND3XLTS U1605 ( .A(n2221), .B(n2220), .C(n2219), .Y(n1227) );
  NAND3XLTS U1606 ( .A(n2218), .B(n2217), .C(n2216), .Y(n1228) );
  NAND3XLTS U1607 ( .A(n2215), .B(n2214), .C(n2213), .Y(n1229) );
  NAND3XLTS U1608 ( .A(n2212), .B(n2211), .C(n2210), .Y(n1230) );
  NAND3XLTS U1609 ( .A(n2209), .B(n2208), .C(n2207), .Y(n1231) );
  OAI211XLTS U1610 ( .A0(n1502), .A1(n1617), .B0(n1487), .C0(n1486), .Y(n1138)
         );
  OAI211XLTS U1611 ( .A0(n1502), .A1(n1608), .B0(n1489), .C0(n1488), .Y(n1139)
         );
  OAI211XLTS U1612 ( .A0(n1502), .A1(n1611), .B0(n1491), .C0(n1490), .Y(n1140)
         );
  OAI211XLTS U1613 ( .A0(n1502), .A1(n1632), .B0(n1493), .C0(n1492), .Y(n1141)
         );
  OAI211XLTS U1614 ( .A0(n1502), .A1(n1614), .B0(n1495), .C0(n1494), .Y(n1142)
         );
  OAI211XLTS U1615 ( .A0(n1502), .A1(n1626), .B0(n1497), .C0(n1496), .Y(n1143)
         );
  OAI211XLTS U1616 ( .A0(n1502), .A1(n1629), .B0(n1485), .C0(n1484), .Y(n1144)
         );
  OAI211XLTS U1617 ( .A0(n1502), .A1(n1620), .B0(n1499), .C0(n1498), .Y(n1145)
         );
  OAI211XLTS U1618 ( .A0(n1502), .A1(n1623), .B0(n1501), .C0(n1500), .Y(n1220)
         );
  OAI211XLTS U1619 ( .A0(n1531), .A1(n1386), .B0(n1528), .C0(n1527), .Y(n1150)
         );
  OAI211XLTS U1620 ( .A0(n1531), .A1(n1379), .B0(n1526), .C0(n1525), .Y(n1151)
         );
  OAI211XLTS U1621 ( .A0(n1531), .A1(n1372), .B0(n1514), .C0(n1513), .Y(n1152)
         );
  OAI211XLTS U1622 ( .A0(n1531), .A1(n1400), .B0(n1516), .C0(n1515), .Y(n1153)
         );
  OAI211XLTS U1623 ( .A0(n1531), .A1(n1393), .B0(n1520), .C0(n1519), .Y(n1154)
         );
  OAI211XLTS U1624 ( .A0(n1531), .A1(n1364), .B0(n1518), .C0(n1517), .Y(n1155)
         );
  OAI211XLTS U1625 ( .A0(n1531), .A1(n1421), .B0(n1524), .C0(n1523), .Y(n1156)
         );
  OAI211XLTS U1626 ( .A0(n1531), .A1(n1414), .B0(n1530), .C0(n1529), .Y(n1157)
         );
  OAI211XLTS U1627 ( .A0(n1531), .A1(n1407), .B0(n1522), .C0(n1521), .Y(n1221)
         );
  OAI211XLTS U1628 ( .A0(n1558), .A1(n1617), .B0(n1557), .C0(n1556), .Y(n1186)
         );
  OAI211XLTS U1629 ( .A0(n1558), .A1(n1608), .B0(n1547), .C0(n1546), .Y(n1187)
         );
  OAI211XLTS U1630 ( .A0(n1558), .A1(n1611), .B0(n1543), .C0(n1542), .Y(n1188)
         );
  OAI211XLTS U1631 ( .A0(n1558), .A1(n1632), .B0(n1541), .C0(n1540), .Y(n1189)
         );
  OAI211XLTS U1632 ( .A0(n1558), .A1(n1614), .B0(n1545), .C0(n1544), .Y(n1190)
         );
  OAI211XLTS U1633 ( .A0(n1558), .A1(n1626), .B0(n1555), .C0(n1554), .Y(n1191)
         );
  OAI211XLTS U1634 ( .A0(n1558), .A1(n1629), .B0(n1551), .C0(n1550), .Y(n1192)
         );
  OAI211XLTS U1635 ( .A0(n1558), .A1(n1620), .B0(n1553), .C0(n1552), .Y(n1193)
         );
  OAI211XLTS U1636 ( .A0(n1558), .A1(n1623), .B0(n1549), .C0(n1548), .Y(n1224)
         );
  OAI211XLTS U1637 ( .A0(n1425), .A1(n1617), .B0(n1389), .C0(n1388), .Y(n1198)
         );
  OAI211XLTS U1638 ( .A0(n1425), .A1(n1608), .B0(n1382), .C0(n1381), .Y(n1199)
         );
  OAI211XLTS U1639 ( .A0(n1425), .A1(n1611), .B0(n1375), .C0(n1374), .Y(n1200)
         );
  OAI211XLTS U1640 ( .A0(n1425), .A1(n1632), .B0(n1403), .C0(n1402), .Y(n1201)
         );
  OAI211XLTS U1641 ( .A0(n1425), .A1(n1614), .B0(n1396), .C0(n1395), .Y(n1202)
         );
  OAI211XLTS U1642 ( .A0(n1425), .A1(n1626), .B0(n1368), .C0(n1367), .Y(n1203)
         );
  OAI211XLTS U1643 ( .A0(n1425), .A1(n1629), .B0(n1424), .C0(n1423), .Y(n1204)
         );
  OAI211XLTS U1644 ( .A0(n1425), .A1(n1620), .B0(n1417), .C0(n1416), .Y(n1205)
         );
  OAI211XLTS U1645 ( .A0(n1425), .A1(n1623), .B0(n1410), .C0(n1409), .Y(n1225)
         );
  NAND3XLTS U1646 ( .A(n2098), .B(n2097), .C(n2096), .Y(n1268) );
  NAND3XLTS U1647 ( .A(n2095), .B(n2094), .C(n2093), .Y(n1269) );
  NAND3XLTS U1648 ( .A(n2092), .B(n2091), .C(n2090), .Y(n1270) );
  NAND3XLTS U1649 ( .A(n2089), .B(n2088), .C(n2087), .Y(n1271) );
  NAND3XLTS U1650 ( .A(n2086), .B(n2085), .C(n2084), .Y(n1272) );
  NAND3XLTS U1651 ( .A(n2083), .B(n2082), .C(n2081), .Y(n1273) );
  NAND3XLTS U1652 ( .A(n2419), .B(n2418), .C(n2417), .Y(n1146) );
  NAND3XLTS U1653 ( .A(n2410), .B(n2409), .C(n2408), .Y(n1147) );
  NAND3XLTS U1654 ( .A(n2407), .B(n2406), .C(n2405), .Y(n1148) );
  NAND3XLTS U1655 ( .A(n2404), .B(n2403), .C(n2402), .Y(n1149) );
  NAND3XLTS U1656 ( .A(n2056), .B(n2055), .C(n2054), .Y(n1282) );
  NAND3XLTS U1657 ( .A(n2053), .B(n2052), .C(n2051), .Y(n1283) );
  NAND3XLTS U1658 ( .A(n2050), .B(n2049), .C(n2048), .Y(n1284) );
  NAND3XLTS U1659 ( .A(n2047), .B(n2046), .C(n2045), .Y(n1285) );
  AO22XLTS U1660 ( .A0(N373), .A1(n1672), .B0(n1671), .B1(n1668), .Y(n1335) );
  AO22XLTS U1661 ( .A0(N375), .A1(n1672), .B0(n1671), .B1(n1670), .Y(n1333) );
  AO22XLTS U1662 ( .A0(N374), .A1(n1672), .B0(n1671), .B1(n1669), .Y(n1334) );
  AOI211XLTS U1663 ( .A0(n1665), .A1(read_reg[2]), .B0(n1664), .C0(n1663), .Y(
        n1666) );
  XOR2XLTS U1664 ( .A(read_reg[0]), .B(n1668), .Y(n1664) );
  OAI21XLTS U1665 ( .A0(n1665), .A1(read_reg[2]), .B0(n1662), .Y(n1663) );
  NOR2X2TS U1666 ( .A(n1634), .B(n2255), .Y(n1337) );
  INVX2TS U1667 ( .A(n1338), .Y(n1339) );
  INVX2TS U1668 ( .A(n1340), .Y(n1341) );
  INVX2TS U1669 ( .A(n1342), .Y(n1343) );
  INVX2TS U1670 ( .A(n1344), .Y(n1345) );
  INVX2TS U1671 ( .A(n1349), .Y(n1350) );
  INVX2TS U1672 ( .A(n1371), .Y(n1372) );
  INVX2TS U1673 ( .A(n1399), .Y(n1400) );
  INVX2TS U1674 ( .A(n1363), .Y(n1364) );
  INVX2TS U1675 ( .A(n1392), .Y(n1393) );
  INVX2TS U1676 ( .A(n1406), .Y(n1407) );
  INVX2TS U1677 ( .A(n1420), .Y(n1421) );
  INVX2TS U1678 ( .A(n1378), .Y(n1379) );
  INVX2TS U1679 ( .A(n1385), .Y(n1386) );
  INVX2TS U1680 ( .A(n1413), .Y(n1414) );
  CLKBUFX2TS U1681 ( .A(selectBit_NORTH), .Y(n1338) );
  CLKBUFX2TS U1682 ( .A(selectBit_SOUTH), .Y(n1340) );
  CLKBUFX2TS U1683 ( .A(selectBit_WEST), .Y(n1342) );
  CLKBUFX2TS U1684 ( .A(selectBit_EAST), .Y(n1344) );
  CLKBUFX2TS U1685 ( .A(readReady), .Y(n1346) );
  NAND2X1TS U1686 ( .A(n1698), .B(n1681), .Y(n1690) );
  NAND2X2TS U1687 ( .A(n1690), .B(n2463), .Y(n1634) );
  INVX2TS U1688 ( .A(n1634), .Y(n1667) );
  NAND2X1TS U1689 ( .A(read_reg[0]), .B(read_reg[1]), .Y(n1691) );
  OAI21XLTS U1690 ( .A0(read_reg[0]), .A1(read_reg[1]), .B0(n1691), .Y(n1676)
         );
  AOI21X1TS U1691 ( .A0(n1691), .A1(n2457), .B0(n1971), .Y(n1673) );
  OAI22X1TS U1692 ( .A0(N374), .A1(n1676), .B0(n2458), .B1(n1673), .Y(n1347)
         );
  AOI221XLTS U1693 ( .A0(n1676), .A1(N374), .B0(n2458), .B1(n1673), .C0(n1347), 
        .Y(n1348) );
  NAND2X1TS U1694 ( .A(N373), .B(n2460), .Y(n1639) );
  OAI21XLTS U1695 ( .A0(N373), .A1(n2460), .B0(n1639), .Y(n1642) );
  AOI21X1TS U1696 ( .A0(n1348), .A1(n1642), .B0(empty_reg), .Y(n1351) );
  CLKBUFX2TS U1697 ( .A(reset), .Y(n1349) );
  OAI21XLTS U1698 ( .A0(n1667), .A1(n1351), .B0(n1350), .Y(n1332) );
  NAND2X1TS U1699 ( .A(n1600), .B(N374), .Y(n1353) );
  NAND2X1TS U1700 ( .A(n1340), .B(n1352), .Y(n1563) );
  NAND2X1TS U1701 ( .A(n1592), .B(n1559), .Y(n1505) );
  INVX2TS U1702 ( .A(n1598), .Y(n1452) );
  INVX2TS U1703 ( .A(n1353), .Y(n1506) );
  AOI22X1TS U1704 ( .A0(N375), .A1(n1353), .B0(n1506), .B1(n2458), .Y(n1562)
         );
  NAND2X1TS U1705 ( .A(n1344), .B(n1426), .Y(n1591) );
  ADDHXLTS U1706 ( .A(N373), .B(n1638), .CO(n1355), .S(n1561) );
  INVX2TS U1707 ( .A(n2230), .Y(n2232) );
  NAND2X1TS U1708 ( .A(N375), .B(n1506), .Y(n1357) );
  NAND2X1TS U1709 ( .A(n1359), .B(n2233), .Y(n1362) );
  NOR2X2TS U1710 ( .A(n2227), .B(n1362), .Y(n2325) );
  INVX2TS U1711 ( .A(n2325), .Y(n1425) );
  CLKBUFX2TS U1712 ( .A(destinationAddressIn_EAST[6]), .Y(n1358) );
  INVX2TS U1713 ( .A(n1358), .Y(n1626) );
  NOR2X2TS U1714 ( .A(n2233), .B(n1634), .Y(n2324) );
  OR2X1TS U1715 ( .A(n1359), .B(n2324), .Y(n2234) );
  INVX2TS U1716 ( .A(n2234), .Y(n2323) );
  NOR2X2TS U1717 ( .A(n2230), .B(n1362), .Y(n2326) );
  CLKBUFX2TS U1718 ( .A(destinationAddressIn_WEST[6]), .Y(n1360) );
  AOI22X1TS U1719 ( .A0(n2323), .A1(\destinationAddressbuffer[7][6] ), .B0(
        n2326), .B1(n1360), .Y(n1368) );
  NOR2X2TS U1720 ( .A(n2225), .B(n1365), .Y(n2328) );
  CLKBUFX2TS U1721 ( .A(destinationAddressIn_SOUTH[6]), .Y(n1363) );
  INVX2TS U1722 ( .A(n2225), .Y(n2226) );
  NOR2X2TS U1723 ( .A(n2226), .B(n1365), .Y(n2327) );
  CLKBUFX2TS U1724 ( .A(destinationAddressIn_NORTH[6]), .Y(n1366) );
  AOI22X1TS U1725 ( .A0(n2328), .A1(n1363), .B0(n2327), .B1(n1366), .Y(n1367)
         );
  CLKBUFX2TS U1726 ( .A(destinationAddressIn_EAST[9]), .Y(n1369) );
  INVX2TS U1727 ( .A(n1369), .Y(n1611) );
  CLKBUFX2TS U1728 ( .A(destinationAddressIn_WEST[9]), .Y(n1370) );
  AOI22X1TS U1729 ( .A0(n2323), .A1(\destinationAddressbuffer[7][9] ), .B0(
        n2326), .B1(n1370), .Y(n1375) );
  CLKBUFX2TS U1730 ( .A(destinationAddressIn_SOUTH[9]), .Y(n1371) );
  CLKBUFX2TS U1731 ( .A(destinationAddressIn_NORTH[9]), .Y(n1373) );
  AOI22X1TS U1732 ( .A0(n2328), .A1(n1371), .B0(n2327), .B1(n1373), .Y(n1374)
         );
  CLKBUFX2TS U1733 ( .A(destinationAddressIn_EAST[10]), .Y(n1376) );
  INVX2TS U1734 ( .A(n1376), .Y(n1608) );
  CLKBUFX2TS U1735 ( .A(destinationAddressIn_WEST[10]), .Y(n1377) );
  AOI22X1TS U1736 ( .A0(n2323), .A1(\destinationAddressbuffer[7][10] ), .B0(
        n2326), .B1(n1377), .Y(n1382) );
  CLKBUFX2TS U1737 ( .A(destinationAddressIn_SOUTH[10]), .Y(n1378) );
  CLKBUFX2TS U1738 ( .A(destinationAddressIn_NORTH[10]), .Y(n1380) );
  AOI22X1TS U1739 ( .A0(n2328), .A1(n1378), .B0(n2327), .B1(n1380), .Y(n1381)
         );
  CLKBUFX2TS U1740 ( .A(destinationAddressIn_EAST[11]), .Y(n1383) );
  INVX2TS U1741 ( .A(n1383), .Y(n1617) );
  CLKBUFX2TS U1742 ( .A(destinationAddressIn_WEST[11]), .Y(n1384) );
  AOI22X1TS U1743 ( .A0(n2323), .A1(\destinationAddressbuffer[7][11] ), .B0(
        n2326), .B1(n1384), .Y(n1389) );
  CLKBUFX2TS U1744 ( .A(destinationAddressIn_SOUTH[11]), .Y(n1385) );
  CLKBUFX2TS U1745 ( .A(destinationAddressIn_NORTH[11]), .Y(n1387) );
  AOI22X1TS U1746 ( .A0(n2328), .A1(n1385), .B0(n2327), .B1(n1387), .Y(n1388)
         );
  CLKBUFX2TS U1747 ( .A(destinationAddressIn_EAST[7]), .Y(n1390) );
  INVX2TS U1748 ( .A(n1390), .Y(n1614) );
  CLKBUFX2TS U1749 ( .A(destinationAddressIn_WEST[7]), .Y(n1391) );
  AOI22X1TS U1750 ( .A0(n2323), .A1(\destinationAddressbuffer[7][7] ), .B0(
        n2326), .B1(n1391), .Y(n1396) );
  CLKBUFX2TS U1751 ( .A(destinationAddressIn_SOUTH[7]), .Y(n1392) );
  CLKBUFX2TS U1752 ( .A(destinationAddressIn_NORTH[7]), .Y(n1394) );
  AOI22X1TS U1753 ( .A0(n2328), .A1(n1392), .B0(n2327), .B1(n1394), .Y(n1395)
         );
  CLKBUFX2TS U1754 ( .A(destinationAddressIn_EAST[8]), .Y(n1397) );
  INVX2TS U1755 ( .A(n1397), .Y(n1632) );
  CLKBUFX2TS U1756 ( .A(destinationAddressIn_WEST[8]), .Y(n1398) );
  AOI22X1TS U1757 ( .A0(n2323), .A1(\destinationAddressbuffer[7][8] ), .B0(
        n2326), .B1(n1398), .Y(n1403) );
  CLKBUFX2TS U1758 ( .A(destinationAddressIn_SOUTH[8]), .Y(n1399) );
  CLKBUFX2TS U1759 ( .A(destinationAddressIn_NORTH[8]), .Y(n1401) );
  AOI22X1TS U1760 ( .A0(n2328), .A1(n1399), .B0(n2327), .B1(n1401), .Y(n1402)
         );
  CLKBUFX2TS U1761 ( .A(writeIn_EAST), .Y(n1404) );
  INVX2TS U1762 ( .A(n1404), .Y(n1623) );
  CLKBUFX2TS U1763 ( .A(writeIn_WEST), .Y(n1405) );
  AOI22X1TS U1764 ( .A0(n2323), .A1(writeOutbuffer[7]), .B0(n2326), .B1(n1405), 
        .Y(n1410) );
  CLKBUFX2TS U1765 ( .A(writeIn_SOUTH), .Y(n1406) );
  CLKBUFX2TS U1766 ( .A(writeIn_NORTH), .Y(n1408) );
  AOI22X1TS U1767 ( .A0(n2328), .A1(n1406), .B0(n2327), .B1(n1408), .Y(n1409)
         );
  CLKBUFX2TS U1768 ( .A(destinationAddressIn_EAST[4]), .Y(n1411) );
  INVX2TS U1769 ( .A(n1411), .Y(n1620) );
  CLKBUFX2TS U1770 ( .A(destinationAddressIn_WEST[4]), .Y(n1412) );
  AOI22X1TS U1771 ( .A0(n2323), .A1(\destinationAddressbuffer[7][4] ), .B0(
        n2326), .B1(n1412), .Y(n1417) );
  CLKBUFX2TS U1772 ( .A(destinationAddressIn_SOUTH[4]), .Y(n1413) );
  CLKBUFX2TS U1773 ( .A(destinationAddressIn_NORTH[4]), .Y(n1415) );
  AOI22X1TS U1774 ( .A0(n2328), .A1(n1413), .B0(n2327), .B1(n1415), .Y(n1416)
         );
  CLKBUFX2TS U1775 ( .A(destinationAddressIn_EAST[5]), .Y(n1418) );
  INVX2TS U1776 ( .A(n1418), .Y(n1629) );
  CLKBUFX2TS U1777 ( .A(destinationAddressIn_WEST[5]), .Y(n1419) );
  AOI22X1TS U1778 ( .A0(n2323), .A1(\destinationAddressbuffer[7][5] ), .B0(
        n2326), .B1(n1419), .Y(n1424) );
  CLKBUFX2TS U1779 ( .A(destinationAddressIn_SOUTH[5]), .Y(n1420) );
  CLKBUFX2TS U1780 ( .A(destinationAddressIn_NORTH[5]), .Y(n1422) );
  AOI22X1TS U1781 ( .A0(n2328), .A1(n1420), .B0(n2327), .B1(n1422), .Y(n1423)
         );
  AOI21X1TS U1782 ( .A0(n1598), .A1(n1597), .B0(n1592), .Y(n1560) );
  NOR3XLTS U1783 ( .A(n1596), .B(n1561), .C(n1503), .Y(n2310) );
  NOR2XLTS U1784 ( .A(N373), .B(n1339), .Y(n1565) );
  AOI31XLTS U1785 ( .A0(n1565), .A1(n2462), .A2(n2458), .B0(n2303), .Y(n1427)
         );
  AOI21X1TS U1786 ( .A0(n1429), .A1(n1427), .B0(n1634), .Y(n1428) );
  NAND2X1TS U1787 ( .A(n1428), .B(n2311), .Y(n1430) );
  NOR2X2TS U1788 ( .A(n2304), .B(n1430), .Y(n2449) );
  INVX2TS U1789 ( .A(n2449), .Y(n1451) );
  NOR2X2TS U1790 ( .A(n1634), .B(n2311), .Y(n2448) );
  OR2X1TS U1791 ( .A(n1428), .B(n2448), .Y(n2312) );
  INVX2TS U1792 ( .A(n2312), .Y(n2447) );
  NOR2X2TS U1793 ( .A(n2308), .B(n1430), .Y(n2450) );
  AOI22X1TS U1794 ( .A0(n2447), .A1(\destinationAddressbuffer[0][11] ), .B0(
        n2450), .B1(n1384), .Y(n1434) );
  INVX2TS U1795 ( .A(n2303), .Y(n2302) );
  NOR2X2TS U1796 ( .A(n2302), .B(n1431), .Y(n2452) );
  CLKBUFX2TS U1797 ( .A(n1432), .Y(n2451) );
  AOI22X1TS U1798 ( .A0(n2452), .A1(n1385), .B0(n2451), .B1(n1387), .Y(n1433)
         );
  AOI22X1TS U1799 ( .A0(n2447), .A1(\destinationAddressbuffer[0][8] ), .B0(
        n2450), .B1(n1398), .Y(n1436) );
  AOI22X1TS U1800 ( .A0(n2452), .A1(n1399), .B0(n2451), .B1(n1401), .Y(n1435)
         );
  AOI22X1TS U1801 ( .A0(n2447), .A1(\destinationAddressbuffer[0][9] ), .B0(
        n2450), .B1(n1370), .Y(n1438) );
  AOI22X1TS U1802 ( .A0(n2452), .A1(n1371), .B0(n2451), .B1(n1373), .Y(n1437)
         );
  AOI22X1TS U1803 ( .A0(n2447), .A1(\destinationAddressbuffer[0][7] ), .B0(
        n2450), .B1(n1391), .Y(n1440) );
  AOI22X1TS U1804 ( .A0(n2452), .A1(n1392), .B0(n2451), .B1(n1394), .Y(n1439)
         );
  AOI22X1TS U1805 ( .A0(n2447), .A1(\destinationAddressbuffer[0][6] ), .B0(
        n2450), .B1(n1360), .Y(n1442) );
  AOI22X1TS U1806 ( .A0(n2452), .A1(n1363), .B0(n2451), .B1(n1366), .Y(n1441)
         );
  AOI22X1TS U1807 ( .A0(n2447), .A1(\destinationAddressbuffer[0][5] ), .B0(
        n2450), .B1(n1419), .Y(n1444) );
  AOI22X1TS U1808 ( .A0(n2452), .A1(n1420), .B0(n2451), .B1(n1422), .Y(n1443)
         );
  AOI22X1TS U1809 ( .A0(n2447), .A1(\destinationAddressbuffer[0][4] ), .B0(
        n2450), .B1(n1412), .Y(n1446) );
  AOI22X1TS U1810 ( .A0(n2452), .A1(n1413), .B0(n2451), .B1(n1415), .Y(n1445)
         );
  AOI22X1TS U1811 ( .A0(n2447), .A1(writeOutbuffer[0]), .B0(n2450), .B1(n1405), 
        .Y(n1448) );
  AOI22X1TS U1812 ( .A0(n2452), .A1(n1406), .B0(n2451), .B1(n1408), .Y(n1447)
         );
  AOI22X1TS U1813 ( .A0(n2447), .A1(\destinationAddressbuffer[0][10] ), .B0(
        n2450), .B1(n1377), .Y(n1450) );
  AOI22X1TS U1814 ( .A0(n2452), .A1(n1378), .B0(n2451), .B1(n1380), .Y(n1449)
         );
  INVX2TS U1815 ( .A(n1559), .Y(n1593) );
  AOI31XLTS U1816 ( .A0(n1600), .A1(n2462), .A2(n2458), .B0(n2292), .Y(n1453)
         );
  AOI21X1TS U1817 ( .A0(n1455), .A1(n1453), .B0(n1634), .Y(n1454) );
  NAND2X1TS U1818 ( .A(n1454), .B(n2299), .Y(n1456) );
  NOR2X2TS U1819 ( .A(n2293), .B(n1456), .Y(n2431) );
  INVX2TS U1820 ( .A(n2431), .Y(n1477) );
  NOR2X2TS U1821 ( .A(n1634), .B(n2299), .Y(n2430) );
  OR2X1TS U1822 ( .A(n1454), .B(n2430), .Y(n2300) );
  INVX2TS U1823 ( .A(n2300), .Y(n2429) );
  NOR2X2TS U1824 ( .A(n2296), .B(n1456), .Y(n2432) );
  AOI22X1TS U1825 ( .A0(n2429), .A1(\destinationAddressbuffer[1][11] ), .B0(
        n2432), .B1(n1384), .Y(n1460) );
  CLKBUFX2TS U1826 ( .A(n1457), .Y(n2434) );
  INVX2TS U1827 ( .A(n2292), .Y(n2291) );
  NOR2X2TS U1828 ( .A(n2291), .B(n1458), .Y(n2433) );
  AOI22X1TS U1829 ( .A0(n2434), .A1(n1387), .B0(n2433), .B1(n1385), .Y(n1459)
         );
  AOI22X1TS U1830 ( .A0(n2429), .A1(\destinationAddressbuffer[1][8] ), .B0(
        n2432), .B1(n1398), .Y(n1462) );
  AOI22X1TS U1831 ( .A0(n2434), .A1(n1401), .B0(n2433), .B1(n1399), .Y(n1461)
         );
  AOI22X1TS U1832 ( .A0(n2429), .A1(\destinationAddressbuffer[1][9] ), .B0(
        n2432), .B1(n1370), .Y(n1464) );
  AOI22X1TS U1833 ( .A0(n2434), .A1(n1373), .B0(n2433), .B1(n1371), .Y(n1463)
         );
  AOI22X1TS U1834 ( .A0(n2429), .A1(writeOutbuffer[1]), .B0(n2432), .B1(n1405), 
        .Y(n1466) );
  AOI22X1TS U1835 ( .A0(n2434), .A1(n1408), .B0(n2433), .B1(n1406), .Y(n1465)
         );
  AOI22X1TS U1836 ( .A0(n2429), .A1(\destinationAddressbuffer[1][7] ), .B0(
        n2432), .B1(n1391), .Y(n1468) );
  AOI22X1TS U1837 ( .A0(n2434), .A1(n1394), .B0(n2433), .B1(n1392), .Y(n1467)
         );
  AOI22X1TS U1838 ( .A0(n2429), .A1(\destinationAddressbuffer[1][6] ), .B0(
        n2432), .B1(n1360), .Y(n1470) );
  AOI22X1TS U1839 ( .A0(n2434), .A1(n1366), .B0(n2433), .B1(n1363), .Y(n1469)
         );
  AOI22X1TS U1840 ( .A0(n2429), .A1(\destinationAddressbuffer[1][10] ), .B0(
        n2432), .B1(n1377), .Y(n1472) );
  AOI22X1TS U1841 ( .A0(n2434), .A1(n1380), .B0(n2433), .B1(n1378), .Y(n1471)
         );
  AOI22X1TS U1842 ( .A0(n2429), .A1(\destinationAddressbuffer[1][4] ), .B0(
        n2432), .B1(n1412), .Y(n1474) );
  AOI22X1TS U1843 ( .A0(n2434), .A1(n1415), .B0(n2433), .B1(n1413), .Y(n1473)
         );
  AOI22X1TS U1844 ( .A0(n2429), .A1(\destinationAddressbuffer[1][5] ), .B0(
        n2432), .B1(n1419), .Y(n1476) );
  AOI22X1TS U1845 ( .A0(n2434), .A1(n1422), .B0(n2433), .B1(n1420), .Y(n1475)
         );
  INVX2TS U1846 ( .A(n1596), .Y(n1533) );
  NOR3XLTS U1847 ( .A(n1561), .B(n1533), .C(n1503), .Y(n2287) );
  AOI31XLTS U1848 ( .A0(N374), .A1(n1565), .A2(n2458), .B0(n2281), .Y(n1478)
         );
  AOI21X1TS U1849 ( .A0(n1480), .A1(n1478), .B0(n1634), .Y(n1479) );
  NAND2X1TS U1850 ( .A(n1479), .B(n2288), .Y(n1481) );
  NOR2X2TS U1851 ( .A(n2282), .B(n1481), .Y(n2413) );
  INVX2TS U1852 ( .A(n2413), .Y(n1502) );
  NOR2X2TS U1853 ( .A(n1634), .B(n2288), .Y(n2412) );
  OR2X1TS U1854 ( .A(n1479), .B(n2412), .Y(n2289) );
  INVX2TS U1855 ( .A(n2289), .Y(n2411) );
  NOR2X2TS U1856 ( .A(n2285), .B(n1481), .Y(n2414) );
  AOI22X1TS U1857 ( .A0(n2411), .A1(\destinationAddressbuffer[2][5] ), .B0(
        n2414), .B1(n1419), .Y(n1485) );
  INVX2TS U1858 ( .A(n2281), .Y(n2280) );
  NOR2X2TS U1859 ( .A(n2280), .B(n1483), .Y(n2415) );
  AOI22X1TS U1860 ( .A0(n2416), .A1(n1422), .B0(n2415), .B1(n1420), .Y(n1484)
         );
  AOI22X1TS U1861 ( .A0(n2411), .A1(\destinationAddressbuffer[2][11] ), .B0(
        n2414), .B1(n1384), .Y(n1487) );
  AOI22X1TS U1862 ( .A0(n2416), .A1(n1387), .B0(n2415), .B1(n1385), .Y(n1486)
         );
  AOI22X1TS U1863 ( .A0(n2411), .A1(\destinationAddressbuffer[2][10] ), .B0(
        n2414), .B1(n1377), .Y(n1489) );
  AOI22X1TS U1864 ( .A0(n2416), .A1(n1380), .B0(n2415), .B1(n1378), .Y(n1488)
         );
  AOI22X1TS U1865 ( .A0(n2411), .A1(\destinationAddressbuffer[2][9] ), .B0(
        n2414), .B1(n1370), .Y(n1491) );
  AOI22X1TS U1866 ( .A0(n2416), .A1(n1373), .B0(n2415), .B1(n1371), .Y(n1490)
         );
  AOI22X1TS U1867 ( .A0(n2411), .A1(\destinationAddressbuffer[2][8] ), .B0(
        n2414), .B1(n1398), .Y(n1493) );
  AOI22X1TS U1868 ( .A0(n2416), .A1(n1401), .B0(n2415), .B1(n1399), .Y(n1492)
         );
  AOI22X1TS U1869 ( .A0(n2411), .A1(\destinationAddressbuffer[2][7] ), .B0(
        n2414), .B1(n1391), .Y(n1495) );
  AOI22X1TS U1870 ( .A0(n2416), .A1(n1394), .B0(n2415), .B1(n1392), .Y(n1494)
         );
  AOI22X1TS U1871 ( .A0(n2411), .A1(\destinationAddressbuffer[2][6] ), .B0(
        n2414), .B1(n1360), .Y(n1497) );
  AOI22X1TS U1872 ( .A0(n2416), .A1(n1366), .B0(n2415), .B1(n1363), .Y(n1496)
         );
  AOI22X1TS U1873 ( .A0(n2411), .A1(\destinationAddressbuffer[2][4] ), .B0(
        n2414), .B1(n1412), .Y(n1499) );
  AOI22X1TS U1874 ( .A0(n2416), .A1(n1415), .B0(n2415), .B1(n1413), .Y(n1498)
         );
  AOI22X1TS U1875 ( .A0(n2411), .A1(writeOutbuffer[2]), .B0(n2414), .B1(n1405), 
        .Y(n1501) );
  AOI22X1TS U1876 ( .A0(n2416), .A1(n1408), .B0(n2415), .B1(n1406), .Y(n1500)
         );
  NAND2X1TS U1877 ( .A(n1506), .B(n2458), .Y(n1507) );
  NAND2X1TS U1878 ( .A(n1509), .B(n2277), .Y(n1512) );
  NOR2X2TS U1879 ( .A(n2269), .B(n1511), .Y(n2397) );
  INVX2TS U1880 ( .A(n2397), .Y(n1531) );
  NOR2X2TS U1881 ( .A(n1634), .B(n2277), .Y(n2395) );
  OR2X1TS U1882 ( .A(n1509), .B(n2395), .Y(n2278) );
  INVX2TS U1883 ( .A(n2278), .Y(n2394) );
  AOI22X1TS U1884 ( .A0(n2394), .A1(\destinationAddressbuffer[3][9] ), .B0(
        n1510), .B1(n1369), .Y(n1514) );
  NOR2X2TS U1885 ( .A(n2270), .B(n1511), .Y(n2398) );
  NOR2X2TS U1886 ( .A(n2274), .B(n1512), .Y(n2396) );
  AOI22X1TS U1887 ( .A0(n2398), .A1(n1373), .B0(n2396), .B1(n1370), .Y(n1513)
         );
  AOI22X1TS U1888 ( .A0(n2394), .A1(\destinationAddressbuffer[3][8] ), .B0(
        n1510), .B1(n1397), .Y(n1516) );
  AOI22X1TS U1889 ( .A0(n2398), .A1(n1401), .B0(n2396), .B1(n1398), .Y(n1515)
         );
  AOI22X1TS U1890 ( .A0(n2394), .A1(\destinationAddressbuffer[3][6] ), .B0(
        n1510), .B1(n1358), .Y(n1518) );
  AOI22X1TS U1891 ( .A0(n2398), .A1(n1366), .B0(n2396), .B1(n1360), .Y(n1517)
         );
  AOI22X1TS U1892 ( .A0(n2394), .A1(\destinationAddressbuffer[3][7] ), .B0(
        n1510), .B1(n1390), .Y(n1520) );
  AOI22X1TS U1893 ( .A0(n2398), .A1(n1394), .B0(n2396), .B1(n1391), .Y(n1519)
         );
  AOI22X1TS U1894 ( .A0(n2394), .A1(writeOutbuffer[3]), .B0(n1510), .B1(n1404), 
        .Y(n1522) );
  AOI22X1TS U1895 ( .A0(n2398), .A1(n1408), .B0(n2396), .B1(n1405), .Y(n1521)
         );
  AOI22X1TS U1896 ( .A0(n2394), .A1(\destinationAddressbuffer[3][5] ), .B0(
        n1510), .B1(n1418), .Y(n1524) );
  AOI22X1TS U1897 ( .A0(n2398), .A1(n1422), .B0(n2396), .B1(n1419), .Y(n1523)
         );
  AOI22X1TS U1898 ( .A0(n2394), .A1(\destinationAddressbuffer[3][10] ), .B0(
        n1510), .B1(n1376), .Y(n1526) );
  AOI22X1TS U1899 ( .A0(n2398), .A1(n1380), .B0(n2396), .B1(n1377), .Y(n1525)
         );
  AOI22X1TS U1900 ( .A0(n2394), .A1(\destinationAddressbuffer[3][11] ), .B0(
        n1510), .B1(n1383), .Y(n1528) );
  AOI22X1TS U1901 ( .A0(n2398), .A1(n1387), .B0(n2396), .B1(n1384), .Y(n1527)
         );
  AOI22X1TS U1902 ( .A0(n2394), .A1(\destinationAddressbuffer[3][4] ), .B0(
        n1510), .B1(n1411), .Y(n1530) );
  AOI22X1TS U1903 ( .A0(n2398), .A1(n1415), .B0(n2396), .B1(n1412), .Y(n1529)
         );
  NAND2X1TS U1904 ( .A(n1532), .B(n1342), .Y(n1594) );
  NOR3XLTS U1905 ( .A(n1561), .B(n1533), .C(n1594), .Y(n2243) );
  NOR3XLTS U1906 ( .A(n1562), .B(n1563), .C(n1597), .Y(n2237) );
  AOI31XLTS U1907 ( .A0(N375), .A1(N374), .A2(n1565), .B0(n2237), .Y(n1534) );
  AOI21X1TS U1908 ( .A0(n1536), .A1(n1534), .B0(n1634), .Y(n1535) );
  NAND2X1TS U1909 ( .A(n1535), .B(n2244), .Y(n1537) );
  NOR2X2TS U1910 ( .A(n2238), .B(n1537), .Y(n2343) );
  INVX2TS U1911 ( .A(n2343), .Y(n1558) );
  NOR2X2TS U1912 ( .A(n1634), .B(n2244), .Y(n2342) );
  OR2X1TS U1913 ( .A(n1535), .B(n2342), .Y(n2245) );
  INVX2TS U1914 ( .A(n2245), .Y(n2341) );
  NOR2X2TS U1915 ( .A(n2241), .B(n1537), .Y(n2344) );
  AOI22X1TS U1916 ( .A0(n2341), .A1(\destinationAddressbuffer[6][8] ), .B0(
        n2344), .B1(n1398), .Y(n1541) );
  CLKBUFX2TS U1917 ( .A(n1538), .Y(n2346) );
  INVX2TS U1918 ( .A(n2237), .Y(n2236) );
  NOR2X2TS U1919 ( .A(n2236), .B(n1539), .Y(n2345) );
  AOI22X1TS U1920 ( .A0(n2346), .A1(n1401), .B0(n2345), .B1(n1399), .Y(n1540)
         );
  AOI22X1TS U1921 ( .A0(n2341), .A1(\destinationAddressbuffer[6][9] ), .B0(
        n2344), .B1(n1370), .Y(n1543) );
  AOI22X1TS U1922 ( .A0(n2346), .A1(n1373), .B0(n2345), .B1(n1371), .Y(n1542)
         );
  AOI22X1TS U1923 ( .A0(n2341), .A1(\destinationAddressbuffer[6][7] ), .B0(
        n2344), .B1(n1391), .Y(n1545) );
  AOI22X1TS U1924 ( .A0(n2346), .A1(n1394), .B0(n2345), .B1(n1392), .Y(n1544)
         );
  AOI22X1TS U1925 ( .A0(n2341), .A1(\destinationAddressbuffer[6][10] ), .B0(
        n2344), .B1(n1377), .Y(n1547) );
  AOI22X1TS U1926 ( .A0(n2346), .A1(n1380), .B0(n2345), .B1(n1378), .Y(n1546)
         );
  AOI22X1TS U1927 ( .A0(n2341), .A1(writeOutbuffer[6]), .B0(n2344), .B1(n1405), 
        .Y(n1549) );
  AOI22X1TS U1928 ( .A0(n2346), .A1(n1408), .B0(n2345), .B1(n1406), .Y(n1548)
         );
  AOI22X1TS U1929 ( .A0(n2341), .A1(\destinationAddressbuffer[6][5] ), .B0(
        n2344), .B1(n1419), .Y(n1551) );
  AOI22X1TS U1930 ( .A0(n2346), .A1(n1422), .B0(n2345), .B1(n1420), .Y(n1550)
         );
  AOI22X1TS U1931 ( .A0(n2341), .A1(\destinationAddressbuffer[6][4] ), .B0(
        n2344), .B1(n1412), .Y(n1553) );
  AOI22X1TS U1932 ( .A0(n2346), .A1(n1415), .B0(n2345), .B1(n1413), .Y(n1552)
         );
  AOI22X1TS U1933 ( .A0(n2341), .A1(\destinationAddressbuffer[6][6] ), .B0(
        n2344), .B1(n1360), .Y(n1555) );
  AOI22X1TS U1934 ( .A0(n2346), .A1(n1366), .B0(n2345), .B1(n1363), .Y(n1554)
         );
  AOI22X1TS U1935 ( .A0(n2341), .A1(\destinationAddressbuffer[6][11] ), .B0(
        n2344), .B1(n1384), .Y(n1557) );
  AOI22X1TS U1936 ( .A0(n2346), .A1(n1387), .B0(n2345), .B1(n1385), .Y(n1556)
         );
  NOR3XLTS U1937 ( .A(n1596), .B(n1561), .C(n1594), .Y(n2265) );
  AOI31XLTS U1938 ( .A0(N375), .A1(n1565), .A2(n2462), .B0(n2259), .Y(n1566)
         );
  AOI21X1TS U1939 ( .A0(n1568), .A1(n1566), .B0(n1634), .Y(n1567) );
  NAND2X1TS U1940 ( .A(n1567), .B(n2266), .Y(n1569) );
  NOR2X2TS U1941 ( .A(n2260), .B(n1569), .Y(n2378) );
  INVX2TS U1942 ( .A(n2378), .Y(n1590) );
  NOR2X2TS U1943 ( .A(n1634), .B(n2266), .Y(n2377) );
  OR2X1TS U1944 ( .A(n1567), .B(n2377), .Y(n2267) );
  INVX2TS U1945 ( .A(n2267), .Y(n2376) );
  NOR2X2TS U1946 ( .A(n2263), .B(n1569), .Y(n2379) );
  AOI22X1TS U1947 ( .A0(n2376), .A1(\destinationAddressbuffer[4][10] ), .B0(
        n2379), .B1(n1377), .Y(n1573) );
  INVX2TS U1948 ( .A(n2259), .Y(n2258) );
  NOR2X2TS U1949 ( .A(n2258), .B(n1570), .Y(n2381) );
  CLKBUFX2TS U1950 ( .A(n1571), .Y(n2380) );
  AOI22X1TS U1951 ( .A0(n2381), .A1(n1378), .B0(n2380), .B1(n1380), .Y(n1572)
         );
  AOI22X1TS U1952 ( .A0(n2376), .A1(\destinationAddressbuffer[4][11] ), .B0(
        n2379), .B1(n1384), .Y(n1575) );
  AOI22X1TS U1953 ( .A0(n2381), .A1(n1385), .B0(n2380), .B1(n1387), .Y(n1574)
         );
  AOI22X1TS U1954 ( .A0(n2376), .A1(\destinationAddressbuffer[4][4] ), .B0(
        n2379), .B1(n1412), .Y(n1577) );
  AOI22X1TS U1955 ( .A0(n2381), .A1(n1413), .B0(n2380), .B1(n1415), .Y(n1576)
         );
  AOI22X1TS U1956 ( .A0(n2376), .A1(\destinationAddressbuffer[4][9] ), .B0(
        n2379), .B1(n1370), .Y(n1579) );
  AOI22X1TS U1957 ( .A0(n2381), .A1(n1371), .B0(n2380), .B1(n1373), .Y(n1578)
         );
  AOI22X1TS U1958 ( .A0(n2376), .A1(writeOutbuffer[4]), .B0(n2379), .B1(n1405), 
        .Y(n1581) );
  AOI22X1TS U1959 ( .A0(n2381), .A1(n1406), .B0(n2380), .B1(n1408), .Y(n1580)
         );
  AOI22X1TS U1960 ( .A0(n2376), .A1(\destinationAddressbuffer[4][8] ), .B0(
        n2379), .B1(n1398), .Y(n1583) );
  AOI22X1TS U1961 ( .A0(n2381), .A1(n1399), .B0(n2380), .B1(n1401), .Y(n1582)
         );
  AOI22X1TS U1962 ( .A0(n2376), .A1(\destinationAddressbuffer[4][6] ), .B0(
        n2379), .B1(n1360), .Y(n1585) );
  AOI22X1TS U1963 ( .A0(n2381), .A1(n1363), .B0(n2380), .B1(n1366), .Y(n1584)
         );
  AOI22X1TS U1964 ( .A0(n2376), .A1(\destinationAddressbuffer[4][7] ), .B0(
        n2379), .B1(n1391), .Y(n1587) );
  AOI22X1TS U1965 ( .A0(n2381), .A1(n1392), .B0(n2380), .B1(n1394), .Y(n1586)
         );
  AOI22X1TS U1966 ( .A0(n2376), .A1(\destinationAddressbuffer[4][5] ), .B0(
        n2379), .B1(n1419), .Y(n1589) );
  AOI22X1TS U1967 ( .A0(n2381), .A1(n1420), .B0(n2380), .B1(n1422), .Y(n1588)
         );
  NAND2X1TS U1968 ( .A(n1602), .B(n2255), .Y(n1604) );
  NOR2X2TS U1969 ( .A(n2249), .B(n1604), .Y(n2360) );
  INVX2TS U1970 ( .A(n2360), .Y(n1633) );
  OR2X1TS U1971 ( .A(n1602), .B(n1337), .Y(n2256) );
  INVX2TS U1972 ( .A(n2256), .Y(n2359) );
  NOR2X2TS U1973 ( .A(n2252), .B(n1604), .Y(n2361) );
  AOI22X1TS U1974 ( .A0(n2359), .A1(\destinationAddressbuffer[5][10] ), .B0(
        n2361), .B1(n1377), .Y(n1607) );
  INVX2TS U1975 ( .A(n2247), .Y(n2248) );
  NOR2X2TS U1976 ( .A(n2248), .B(n1605), .Y(n2363) );
  NOR2X2TS U1977 ( .A(n2247), .B(n1605), .Y(n2362) );
  AOI22X1TS U1978 ( .A0(n2363), .A1(n1380), .B0(n2362), .B1(n1378), .Y(n1606)
         );
  AOI22X1TS U1979 ( .A0(n2359), .A1(\destinationAddressbuffer[5][9] ), .B0(
        n2361), .B1(n1370), .Y(n1610) );
  AOI22X1TS U1980 ( .A0(n2363), .A1(n1373), .B0(n2362), .B1(n1371), .Y(n1609)
         );
  AOI22X1TS U1981 ( .A0(n2359), .A1(\destinationAddressbuffer[5][7] ), .B0(
        n2361), .B1(n1391), .Y(n1613) );
  AOI22X1TS U1982 ( .A0(n2363), .A1(n1394), .B0(n2362), .B1(n1392), .Y(n1612)
         );
  AOI22X1TS U1983 ( .A0(n2359), .A1(\destinationAddressbuffer[5][11] ), .B0(
        n2361), .B1(n1384), .Y(n1616) );
  AOI22X1TS U1984 ( .A0(n2363), .A1(n1387), .B0(n2362), .B1(n1385), .Y(n1615)
         );
  AOI22X1TS U1985 ( .A0(n2359), .A1(\destinationAddressbuffer[5][4] ), .B0(
        n2361), .B1(n1412), .Y(n1619) );
  AOI22X1TS U1986 ( .A0(n2363), .A1(n1415), .B0(n2362), .B1(n1413), .Y(n1618)
         );
  AOI22X1TS U1987 ( .A0(n2359), .A1(writeOutbuffer[5]), .B0(n2361), .B1(n1405), 
        .Y(n1622) );
  AOI22X1TS U1988 ( .A0(n2363), .A1(n1408), .B0(n2362), .B1(n1406), .Y(n1621)
         );
  AOI22X1TS U1989 ( .A0(n2359), .A1(\destinationAddressbuffer[5][6] ), .B0(
        n2361), .B1(n1360), .Y(n1625) );
  AOI22X1TS U1990 ( .A0(n2363), .A1(n1366), .B0(n2362), .B1(n1363), .Y(n1624)
         );
  AOI22X1TS U1991 ( .A0(n2359), .A1(\destinationAddressbuffer[5][5] ), .B0(
        n2361), .B1(n1419), .Y(n1628) );
  AOI22X1TS U1992 ( .A0(n2363), .A1(n1422), .B0(n2362), .B1(n1420), .Y(n1627)
         );
  AOI22X1TS U1993 ( .A0(n2359), .A1(\destinationAddressbuffer[5][8] ), .B0(
        n2361), .B1(n1398), .Y(n1631) );
  AOI22X1TS U1994 ( .A0(n2363), .A1(n1401), .B0(n2362), .B1(n1399), .Y(n1630)
         );
  NAND2X1TS U1995 ( .A(n1350), .B(empty_reg), .Y(n1677) );
  AOI22X1TS U1996 ( .A0(N375), .A1(n2457), .B0(read_reg[2]), .B1(n2458), .Y(
        n1636) );
  INVX2TS U1997 ( .A(n1652), .Y(n1649) );
  OAI21XLTS U1998 ( .A0(N374), .A1(n2461), .B0(n1636), .Y(n1637) );
  AOI21X1TS U1999 ( .A0(read_reg[0]), .A1(n2456), .B0(n1637), .Y(n1648) );
  ADDHXLTS U2000 ( .A(n1641), .B(n1640), .CO(n1652), .S(n1654) );
  INVX2TS U2001 ( .A(n1654), .Y(n1643) );
  AOI21X1TS U2002 ( .A0(n1644), .A1(n1643), .B0(n1642), .Y(n1646) );
  OAI22X1TS U2003 ( .A0(n1644), .A1(n1643), .B0(n1650), .B1(n1649), .Y(n1645)
         );
  AOI21X1TS U2004 ( .A0(n1653), .A1(n1646), .B0(n1645), .Y(n1647) );
  INVX2TS U2005 ( .A(n1651), .Y(n1655) );
  NAND2X1TS U2006 ( .A(n1655), .B(n1652), .Y(n1658) );
  XNOR2X1TS U2007 ( .A(N375), .B(n1656), .Y(n1657) );
  INVX2TS U2008 ( .A(n1670), .Y(n1665) );
  ADDHXLTS U2009 ( .A(N373), .B(n1659), .CO(n1661), .S(n1668) );
  XNOR2X1TS U2010 ( .A(read_reg[1]), .B(n1669), .Y(n1662) );
  OAI2BB2XLTS U2011 ( .B0(n2463), .B1(n1677), .A0N(n1671), .A1N(n1666), .Y(
        N2624) );
  NAND2X1TS U2012 ( .A(n1350), .B(n2459), .Y(n1675) );
  AOI22X1TS U2013 ( .A0(read_reg[0]), .A1(n1677), .B0(n1675), .B1(n2460), .Y(
        n1336) );
  INVX2TS U2014 ( .A(n1673), .Y(n1674) );
  OAI22X1TS U2015 ( .A0(n2457), .A1(n1677), .B0(n1674), .B1(n1675), .Y(n1331)
         );
  OAI22X1TS U2016 ( .A0(n2461), .A1(n1677), .B0(n1676), .B1(n1675), .Y(n1330)
         );
  CLKBUFX2TS U2017 ( .A(readIn_SOUTH), .Y(n1678) );
  CLKBUFX2TS U2018 ( .A(readIn_WEST), .Y(n1679) );
  NAND2X1TS U2019 ( .A(n1698), .B(empty_reg), .Y(n1684) );
  NOR4XLTS U2020 ( .A(n1346), .B(n1344), .C(n1343), .D(n1684), .Y(n1781) );
  CLKBUFX2TS U2021 ( .A(n1781), .Y(n1964) );
  AOI22X1TS U2022 ( .A0(n1678), .A1(n1877), .B0(n1679), .B1(n1964), .Y(n1701)
         );
  CLKBUFX2TS U2023 ( .A(readIn_NORTH), .Y(n1680) );
  CLKBUFX2TS U2024 ( .A(readIn_EAST), .Y(n1683) );
  NOR4XLTS U2025 ( .A(n1342), .B(n1346), .C(n1345), .D(n1684), .Y(n1918) );
  AOI22X1TS U2026 ( .A0(n1680), .A1(n1682), .B0(n1683), .B1(n1918), .Y(n1700)
         );
  OAI31X1TS U2027 ( .A0(n1686), .A1(n1697), .A2(n1685), .B0(n1698), .Y(n1689)
         );
  AND4X2TS U2028 ( .A(empty_reg), .B(n1689), .C(n1688), .D(n1687), .Y(n1978)
         );
  NOR3X1TS U2029 ( .A(read_reg[0]), .B(read_reg[2]), .C(n2461), .Y(n1965) );
  CLKBUFX2TS U2030 ( .A(n1965), .Y(n1890) );
  NOR3X1TS U2031 ( .A(read_reg[0]), .B(read_reg[1]), .C(read_reg[2]), .Y(n1817) );
  AOI22X1TS U2032 ( .A0(readOutbuffer[2]), .A1(n1890), .B0(readOutbuffer[0]), 
        .B1(n1817), .Y(n1695) );
  NOR3X1TS U2033 ( .A(read_reg[0]), .B(n2461), .C(n2457), .Y(n1967) );
  CLKBUFX2TS U2034 ( .A(n1967), .Y(n1891) );
  NOR3X1TS U2035 ( .A(read_reg[0]), .B(read_reg[1]), .C(n2457), .Y(n1818) );
  AOI22X1TS U2036 ( .A0(readOutbuffer[6]), .A1(n1891), .B0(readOutbuffer[4]), 
        .B1(n1818), .Y(n1694) );
  NOR3X1TS U2037 ( .A(read_reg[1]), .B(read_reg[2]), .C(n2460), .Y(n1819) );
  AOI22X1TS U2038 ( .A0(readOutbuffer[3]), .A1(n1969), .B0(readOutbuffer[1]), 
        .B1(n1819), .Y(n1693) );
  NOR3X1TS U2039 ( .A(read_reg[1]), .B(n2460), .C(n2457), .Y(n1820) );
  AOI22X1TS U2040 ( .A0(readOutbuffer[7]), .A1(n1971), .B0(readOutbuffer[5]), 
        .B1(n1820), .Y(n1692) );
  NAND4XLTS U2041 ( .A(n1695), .B(n1694), .C(n1693), .D(n1692), .Y(n1696) );
  AOI22X1TS U2042 ( .A0(readOut), .A1(n1707), .B0(n2459), .B1(n1696), .Y(n1699) );
  CLKBUFX2TS U2043 ( .A(n1918), .Y(n1961) );
  AOI22X1TS U2044 ( .A0(n1404), .A1(n1961), .B0(n1405), .B1(n1964), .Y(n1710)
         );
  AOI22X1TS U2045 ( .A0(n1408), .A1(n1682), .B0(n1406), .B1(n1877), .Y(n1709)
         );
  AOI22X1TS U2046 ( .A0(writeOutbuffer[2]), .A1(n1890), .B0(writeOutbuffer[0]), 
        .B1(n1817), .Y(n1705) );
  AOI22X1TS U2047 ( .A0(writeOutbuffer[6]), .A1(n1891), .B0(writeOutbuffer[4]), 
        .B1(n1818), .Y(n1704) );
  AOI22X1TS U2048 ( .A0(writeOutbuffer[3]), .A1(n1969), .B0(writeOutbuffer[1]), 
        .B1(n1819), .Y(n1703) );
  AOI22X1TS U2049 ( .A0(writeOutbuffer[7]), .A1(n1971), .B0(writeOutbuffer[5]), 
        .B1(n1820), .Y(n1702) );
  NAND4XLTS U2050 ( .A(n1705), .B(n1704), .C(n1703), .D(n1702), .Y(n1706) );
  AOI22X1TS U2051 ( .A0(writeOut), .A1(n1707), .B0(n2459), .B1(n1706), .Y(
        n1708) );
  CLKBUFX2TS U2052 ( .A(requesterAddressIn_NORTH[0]), .Y(n1711) );
  CLKBUFX2TS U2053 ( .A(requesterAddressIn_EAST[0]), .Y(n1712) );
  AOI22X1TS U2054 ( .A0(n1711), .A1(n1682), .B0(n1712), .B1(n1961), .Y(n1724)
         );
  CLKBUFX2TS U2055 ( .A(requesterAddressIn_SOUTH[0]), .Y(n1713) );
  CLKBUFX2TS U2056 ( .A(requesterAddressIn_WEST[0]), .Y(n1714) );
  AOI22X1TS U2057 ( .A0(n1713), .A1(n1877), .B0(n1714), .B1(n1964), .Y(n1723)
         );
  AOI22X1TS U2058 ( .A0(\requesterAddressbuffer[2][0] ), .A1(n1890), .B0(
        \requesterAddressbuffer[0][0] ), .B1(n1817), .Y(n1718) );
  AOI22X1TS U2059 ( .A0(\requesterAddressbuffer[6][0] ), .A1(n1891), .B0(
        \requesterAddressbuffer[4][0] ), .B1(n1818), .Y(n1717) );
  AOI22X1TS U2060 ( .A0(\requesterAddressbuffer[3][0] ), .A1(n1969), .B0(
        \requesterAddressbuffer[1][0] ), .B1(n1819), .Y(n1716) );
  AOI22X1TS U2061 ( .A0(\requesterAddressbuffer[7][0] ), .A1(n1971), .B0(
        \requesterAddressbuffer[5][0] ), .B1(n1820), .Y(n1715) );
  NAND4XLTS U2062 ( .A(n1718), .B(n1717), .C(n1716), .D(n1715), .Y(n1719) );
  AOI22X1TS U2063 ( .A0(requesterAddressOut[0]), .A1(n1978), .B0(n2459), .B1(
        n1719), .Y(n1722) );
  CLKBUFX2TS U2064 ( .A(readRequesterAddress[0]), .Y(n1720) );
  INVX2TS U2065 ( .A(n1721), .Y(n1980) );
  NAND2X1TS U2066 ( .A(n1720), .B(n1980), .Y(n1773) );
  CLKBUFX2TS U2067 ( .A(requesterAddressIn_NORTH[1]), .Y(n1725) );
  CLKBUFX2TS U2068 ( .A(requesterAddressIn_EAST[1]), .Y(n1726) );
  AOI22X1TS U2069 ( .A0(n1725), .A1(n1682), .B0(n1726), .B1(n1961), .Y(n1737)
         );
  CLKBUFX2TS U2070 ( .A(requesterAddressIn_SOUTH[1]), .Y(n1727) );
  CLKBUFX2TS U2071 ( .A(requesterAddressIn_WEST[1]), .Y(n1728) );
  AOI22X1TS U2072 ( .A0(n1727), .A1(n1877), .B0(n1728), .B1(n1781), .Y(n1736)
         );
  AOI22X1TS U2073 ( .A0(\requesterAddressbuffer[2][1] ), .A1(n1890), .B0(
        \requesterAddressbuffer[0][1] ), .B1(n1817), .Y(n1732) );
  AOI22X1TS U2074 ( .A0(\requesterAddressbuffer[6][1] ), .A1(n1891), .B0(
        \requesterAddressbuffer[4][1] ), .B1(n1818), .Y(n1731) );
  AOI22X1TS U2075 ( .A0(\requesterAddressbuffer[3][1] ), .A1(n1969), .B0(
        \requesterAddressbuffer[1][1] ), .B1(n1819), .Y(n1730) );
  AOI22X1TS U2076 ( .A0(\requesterAddressbuffer[7][1] ), .A1(n1971), .B0(
        \requesterAddressbuffer[5][1] ), .B1(n1820), .Y(n1729) );
  NAND4XLTS U2077 ( .A(n1732), .B(n1731), .C(n1730), .D(n1729), .Y(n1733) );
  AOI22X1TS U2078 ( .A0(requesterAddressOut[1]), .A1(n1978), .B0(n2459), .B1(
        n1733), .Y(n1735) );
  CLKBUFX2TS U2079 ( .A(readRequesterAddress[1]), .Y(n1734) );
  NAND2X1TS U2080 ( .A(n1734), .B(n1980), .Y(n1787) );
  CLKBUFX2TS U2081 ( .A(requesterAddressIn_NORTH[2]), .Y(n1738) );
  CLKBUFX2TS U2082 ( .A(requesterAddressIn_EAST[2]), .Y(n1739) );
  AOI22X1TS U2083 ( .A0(n1738), .A1(n1682), .B0(n1739), .B1(n1961), .Y(n1750)
         );
  CLKBUFX2TS U2084 ( .A(requesterAddressIn_SOUTH[2]), .Y(n1740) );
  CLKBUFX2TS U2085 ( .A(requesterAddressIn_WEST[2]), .Y(n1741) );
  AOI22X1TS U2086 ( .A0(n1740), .A1(n1877), .B0(n1741), .B1(n1964), .Y(n1749)
         );
  AOI22X1TS U2087 ( .A0(\requesterAddressbuffer[2][2] ), .A1(n1890), .B0(
        \requesterAddressbuffer[0][2] ), .B1(n1817), .Y(n1745) );
  AOI22X1TS U2088 ( .A0(\requesterAddressbuffer[6][2] ), .A1(n1891), .B0(
        \requesterAddressbuffer[4][2] ), .B1(n1818), .Y(n1744) );
  AOI22X1TS U2089 ( .A0(\requesterAddressbuffer[3][2] ), .A1(n1969), .B0(
        \requesterAddressbuffer[1][2] ), .B1(n1819), .Y(n1743) );
  AOI22X1TS U2090 ( .A0(\requesterAddressbuffer[7][2] ), .A1(n1971), .B0(
        \requesterAddressbuffer[5][2] ), .B1(n1820), .Y(n1742) );
  NAND4XLTS U2091 ( .A(n1745), .B(n1744), .C(n1743), .D(n1742), .Y(n1746) );
  AOI22X1TS U2092 ( .A0(requesterAddressOut[2]), .A1(n1978), .B0(n2459), .B1(
        n1746), .Y(n1748) );
  CLKBUFX2TS U2093 ( .A(readRequesterAddress[2]), .Y(n1747) );
  NAND2X1TS U2094 ( .A(n1747), .B(n1980), .Y(n1800) );
  CLKBUFX2TS U2095 ( .A(requesterAddressIn_NORTH[3]), .Y(n1751) );
  CLKBUFX2TS U2096 ( .A(requesterAddressIn_EAST[3]), .Y(n1752) );
  AOI22X1TS U2097 ( .A0(n1751), .A1(n1682), .B0(n1752), .B1(n1961), .Y(n1763)
         );
  CLKBUFX2TS U2098 ( .A(requesterAddressIn_SOUTH[3]), .Y(n1753) );
  CLKBUFX2TS U2099 ( .A(requesterAddressIn_WEST[3]), .Y(n1754) );
  AOI22X1TS U2100 ( .A0(n1753), .A1(n1877), .B0(n1754), .B1(n1781), .Y(n1762)
         );
  AOI22X1TS U2101 ( .A0(\requesterAddressbuffer[2][3] ), .A1(n1890), .B0(
        \requesterAddressbuffer[0][3] ), .B1(n1817), .Y(n1758) );
  AOI22X1TS U2102 ( .A0(\requesterAddressbuffer[6][3] ), .A1(n1891), .B0(
        \requesterAddressbuffer[4][3] ), .B1(n1818), .Y(n1757) );
  AOI22X1TS U2103 ( .A0(\requesterAddressbuffer[3][3] ), .A1(n1969), .B0(
        \requesterAddressbuffer[1][3] ), .B1(n1819), .Y(n1756) );
  AOI22X1TS U2104 ( .A0(\requesterAddressbuffer[7][3] ), .A1(n1971), .B0(
        \requesterAddressbuffer[5][3] ), .B1(n1820), .Y(n1755) );
  NAND4XLTS U2105 ( .A(n1758), .B(n1757), .C(n1756), .D(n1755), .Y(n1759) );
  AOI22X1TS U2106 ( .A0(requesterAddressOut[3]), .A1(n1978), .B0(n2459), .B1(
        n1759), .Y(n1761) );
  CLKBUFX2TS U2107 ( .A(readRequesterAddress[3]), .Y(n1760) );
  NAND2X1TS U2108 ( .A(n1760), .B(n1980), .Y(n1813) );
  CLKBUFX2TS U2109 ( .A(destinationAddressIn_NORTH[0]), .Y(n1764) );
  CLKBUFX2TS U2110 ( .A(destinationAddressIn_EAST[0]), .Y(n1765) );
  AOI22X1TS U2111 ( .A0(n1764), .A1(n1682), .B0(n1765), .B1(n1961), .Y(n1776)
         );
  CLKBUFX2TS U2112 ( .A(destinationAddressIn_SOUTH[0]), .Y(n1766) );
  CLKBUFX2TS U2113 ( .A(destinationAddressIn_WEST[0]), .Y(n1767) );
  AOI22X1TS U2114 ( .A0(n1766), .A1(n1877), .B0(n1767), .B1(n1964), .Y(n1775)
         );
  AOI22X1TS U2115 ( .A0(\destinationAddressbuffer[2][0] ), .A1(n1890), .B0(
        \destinationAddressbuffer[0][0] ), .B1(n1817), .Y(n1771) );
  AOI22X1TS U2116 ( .A0(\destinationAddressbuffer[6][0] ), .A1(n1891), .B0(
        \destinationAddressbuffer[4][0] ), .B1(n1818), .Y(n1770) );
  AOI22X1TS U2117 ( .A0(\destinationAddressbuffer[3][0] ), .A1(n1969), .B0(
        \destinationAddressbuffer[1][0] ), .B1(n1819), .Y(n1769) );
  AOI22X1TS U2118 ( .A0(\destinationAddressbuffer[7][0] ), .A1(n1971), .B0(
        \destinationAddressbuffer[5][0] ), .B1(n1820), .Y(n1768) );
  NAND4XLTS U2119 ( .A(n1771), .B(n1770), .C(n1769), .D(n1768), .Y(n1772) );
  AOI22X1TS U2120 ( .A0(destinationAddressOut[0]), .A1(n1978), .B0(n2459), 
        .B1(n1772), .Y(n1774) );
  CLKBUFX2TS U2121 ( .A(destinationAddressIn_NORTH[1]), .Y(n1777) );
  CLKBUFX2TS U2122 ( .A(destinationAddressIn_EAST[1]), .Y(n1778) );
  AOI22X1TS U2123 ( .A0(n1777), .A1(n1682), .B0(n1778), .B1(n1961), .Y(n1790)
         );
  CLKBUFX2TS U2124 ( .A(destinationAddressIn_SOUTH[1]), .Y(n1779) );
  CLKBUFX2TS U2125 ( .A(destinationAddressIn_WEST[1]), .Y(n1780) );
  AOI22X1TS U2126 ( .A0(n1779), .A1(n1877), .B0(n1780), .B1(n1781), .Y(n1789)
         );
  AOI22X1TS U2127 ( .A0(\destinationAddressbuffer[2][1] ), .A1(n1890), .B0(
        \destinationAddressbuffer[0][1] ), .B1(n1817), .Y(n1785) );
  AOI22X1TS U2128 ( .A0(\destinationAddressbuffer[6][1] ), .A1(n1891), .B0(
        \destinationAddressbuffer[4][1] ), .B1(n1818), .Y(n1784) );
  AOI22X1TS U2129 ( .A0(\destinationAddressbuffer[3][1] ), .A1(n1969), .B0(
        \destinationAddressbuffer[1][1] ), .B1(n1819), .Y(n1783) );
  AOI22X1TS U2130 ( .A0(\destinationAddressbuffer[7][1] ), .A1(n1971), .B0(
        \destinationAddressbuffer[5][1] ), .B1(n1820), .Y(n1782) );
  NAND4XLTS U2131 ( .A(n1785), .B(n1784), .C(n1783), .D(n1782), .Y(n1786) );
  AOI22X1TS U2132 ( .A0(destinationAddressOut[1]), .A1(n1978), .B0(n2459), 
        .B1(n1786), .Y(n1788) );
  CLKBUFX2TS U2133 ( .A(destinationAddressIn_NORTH[2]), .Y(n1791) );
  CLKBUFX2TS U2134 ( .A(destinationAddressIn_EAST[2]), .Y(n1792) );
  AOI22X1TS U2135 ( .A0(n1791), .A1(n1682), .B0(n1792), .B1(n1961), .Y(n1803)
         );
  CLKBUFX2TS U2136 ( .A(destinationAddressIn_SOUTH[2]), .Y(n1793) );
  CLKBUFX2TS U2137 ( .A(destinationAddressIn_WEST[2]), .Y(n1794) );
  AOI22X1TS U2138 ( .A0(n1793), .A1(n1877), .B0(n1794), .B1(n1964), .Y(n1802)
         );
  AOI22X1TS U2139 ( .A0(\destinationAddressbuffer[2][2] ), .A1(n1890), .B0(
        \destinationAddressbuffer[0][2] ), .B1(n1817), .Y(n1798) );
  AOI22X1TS U2140 ( .A0(\destinationAddressbuffer[6][2] ), .A1(n1891), .B0(
        \destinationAddressbuffer[4][2] ), .B1(n1818), .Y(n1797) );
  AOI22X1TS U2141 ( .A0(\destinationAddressbuffer[3][2] ), .A1(n1969), .B0(
        \destinationAddressbuffer[1][2] ), .B1(n1819), .Y(n1796) );
  AOI22X1TS U2142 ( .A0(\destinationAddressbuffer[7][2] ), .A1(n1971), .B0(
        \destinationAddressbuffer[5][2] ), .B1(n1820), .Y(n1795) );
  NAND4XLTS U2143 ( .A(n1798), .B(n1797), .C(n1796), .D(n1795), .Y(n1799) );
  AOI22X1TS U2144 ( .A0(destinationAddressOut[2]), .A1(n1978), .B0(n2459), 
        .B1(n1799), .Y(n1801) );
  CLKBUFX2TS U2145 ( .A(destinationAddressIn_NORTH[3]), .Y(n1804) );
  CLKBUFX2TS U2146 ( .A(destinationAddressIn_EAST[3]), .Y(n1805) );
  AOI22X1TS U2147 ( .A0(n1804), .A1(n1682), .B0(n1805), .B1(n1961), .Y(n1816)
         );
  CLKBUFX2TS U2148 ( .A(destinationAddressIn_SOUTH[3]), .Y(n1806) );
  CLKBUFX2TS U2149 ( .A(destinationAddressIn_WEST[3]), .Y(n1807) );
  AOI22X1TS U2150 ( .A0(n1806), .A1(n1877), .B0(n1807), .B1(n1964), .Y(n1815)
         );
  AOI22X1TS U2151 ( .A0(\destinationAddressbuffer[2][3] ), .A1(n1890), .B0(
        \destinationAddressbuffer[0][3] ), .B1(n1817), .Y(n1811) );
  AOI22X1TS U2152 ( .A0(\destinationAddressbuffer[6][3] ), .A1(n1891), .B0(
        \destinationAddressbuffer[4][3] ), .B1(n1818), .Y(n1810) );
  AOI22X1TS U2153 ( .A0(\destinationAddressbuffer[3][3] ), .A1(n1969), .B0(
        \destinationAddressbuffer[1][3] ), .B1(n1819), .Y(n1809) );
  AOI22X1TS U2154 ( .A0(\destinationAddressbuffer[7][3] ), .A1(n1971), .B0(
        \destinationAddressbuffer[5][3] ), .B1(n1820), .Y(n1808) );
  NAND4XLTS U2155 ( .A(n1811), .B(n1810), .C(n1809), .D(n1808), .Y(n1812) );
  AOI22X1TS U2156 ( .A0(destinationAddressOut[3]), .A1(n1978), .B0(n2459), 
        .B1(n1812), .Y(n1814) );
  AOI22X1TS U2157 ( .A0(n1411), .A1(n1961), .B0(n1412), .B1(n1964), .Y(n1828)
         );
  AOI22X1TS U2158 ( .A0(n1415), .A1(n1682), .B0(n1413), .B1(n1877), .Y(n1827)
         );
  CLKBUFX2TS U2159 ( .A(n1817), .Y(n1966) );
  AOI22X1TS U2160 ( .A0(\destinationAddressbuffer[2][4] ), .A1(n1890), .B0(
        \destinationAddressbuffer[0][4] ), .B1(n1966), .Y(n1824) );
  CLKBUFX2TS U2161 ( .A(n1818), .Y(n1968) );
  AOI22X1TS U2162 ( .A0(\destinationAddressbuffer[6][4] ), .A1(n1891), .B0(
        \destinationAddressbuffer[4][4] ), .B1(n1968), .Y(n1823) );
  CLKBUFX2TS U2163 ( .A(n1819), .Y(n1970) );
  AOI22X1TS U2164 ( .A0(\destinationAddressbuffer[3][4] ), .A1(n1969), .B0(
        \destinationAddressbuffer[1][4] ), .B1(n1970), .Y(n1822) );
  CLKBUFX2TS U2165 ( .A(n1820), .Y(n1972) );
  AOI22X1TS U2166 ( .A0(\destinationAddressbuffer[7][4] ), .A1(n1971), .B0(
        \destinationAddressbuffer[5][4] ), .B1(n1972), .Y(n1821) );
  NAND4XLTS U2167 ( .A(n1824), .B(n1823), .C(n1822), .D(n1821), .Y(n1825) );
  AOI22X1TS U2168 ( .A0(destinationAddressOut[4]), .A1(n1978), .B0(n2459), 
        .B1(n1825), .Y(n1826) );
  AOI22X1TS U2169 ( .A0(n1418), .A1(n1961), .B0(n1419), .B1(n1964), .Y(n1836)
         );
  AOI22X1TS U2170 ( .A0(n1422), .A1(n1682), .B0(n1420), .B1(n1877), .Y(n1835)
         );
  AOI22X1TS U2171 ( .A0(\destinationAddressbuffer[2][5] ), .A1(n1890), .B0(
        \destinationAddressbuffer[0][5] ), .B1(n1966), .Y(n1832) );
  AOI22X1TS U2172 ( .A0(\destinationAddressbuffer[6][5] ), .A1(n1891), .B0(
        \destinationAddressbuffer[4][5] ), .B1(n1968), .Y(n1831) );
  AOI22X1TS U2173 ( .A0(\destinationAddressbuffer[3][5] ), .A1(n1969), .B0(
        \destinationAddressbuffer[1][5] ), .B1(n1970), .Y(n1830) );
  AOI22X1TS U2174 ( .A0(\destinationAddressbuffer[7][5] ), .A1(n1971), .B0(
        \destinationAddressbuffer[5][5] ), .B1(n1972), .Y(n1829) );
  NAND4XLTS U2175 ( .A(n1832), .B(n1831), .C(n1830), .D(n1829), .Y(n1833) );
  AOI22X1TS U2176 ( .A0(destinationAddressOut[5]), .A1(n1978), .B0(n2459), 
        .B1(n1833), .Y(n1834) );
  AOI22X1TS U2177 ( .A0(n1358), .A1(n1961), .B0(n1360), .B1(n1964), .Y(n1844)
         );
  AOI22X1TS U2178 ( .A0(n1366), .A1(n1682), .B0(n1363), .B1(n1877), .Y(n1843)
         );
  AOI22X1TS U2179 ( .A0(\destinationAddressbuffer[2][6] ), .A1(n1965), .B0(
        \destinationAddressbuffer[0][6] ), .B1(n1966), .Y(n1840) );
  AOI22X1TS U2180 ( .A0(\destinationAddressbuffer[6][6] ), .A1(n1967), .B0(
        \destinationAddressbuffer[4][6] ), .B1(n1968), .Y(n1839) );
  AOI22X1TS U2181 ( .A0(\destinationAddressbuffer[3][6] ), .A1(n1969), .B0(
        \destinationAddressbuffer[1][6] ), .B1(n1970), .Y(n1838) );
  AOI22X1TS U2182 ( .A0(\destinationAddressbuffer[7][6] ), .A1(n1971), .B0(
        \destinationAddressbuffer[5][6] ), .B1(n1972), .Y(n1837) );
  NAND4XLTS U2183 ( .A(n1840), .B(n1839), .C(n1838), .D(n1837), .Y(n1841) );
  AOI22X1TS U2184 ( .A0(destinationAddressOut[6]), .A1(n1978), .B0(n2459), 
        .B1(n1841), .Y(n1842) );
  AOI22X1TS U2185 ( .A0(n1390), .A1(n1961), .B0(n1391), .B1(n1964), .Y(n1852)
         );
  AOI22X1TS U2186 ( .A0(n1394), .A1(n1682), .B0(n1392), .B1(n1877), .Y(n1851)
         );
  AOI22X1TS U2187 ( .A0(\destinationAddressbuffer[2][7] ), .A1(n1965), .B0(
        \destinationAddressbuffer[0][7] ), .B1(n1966), .Y(n1848) );
  AOI22X1TS U2188 ( .A0(\destinationAddressbuffer[6][7] ), .A1(n1967), .B0(
        \destinationAddressbuffer[4][7] ), .B1(n1968), .Y(n1847) );
  AOI22X1TS U2189 ( .A0(\destinationAddressbuffer[3][7] ), .A1(n1969), .B0(
        \destinationAddressbuffer[1][7] ), .B1(n1970), .Y(n1846) );
  AOI22X1TS U2190 ( .A0(\destinationAddressbuffer[7][7] ), .A1(n1971), .B0(
        \destinationAddressbuffer[5][7] ), .B1(n1972), .Y(n1845) );
  NAND4XLTS U2191 ( .A(n1848), .B(n1847), .C(n1846), .D(n1845), .Y(n1849) );
  AOI22X1TS U2192 ( .A0(destinationAddressOut[7]), .A1(n1978), .B0(n2459), 
        .B1(n1849), .Y(n1850) );
  AOI22X1TS U2193 ( .A0(n1397), .A1(n1961), .B0(n1398), .B1(n1964), .Y(n1860)
         );
  AOI22X1TS U2194 ( .A0(n1401), .A1(n1682), .B0(n1399), .B1(n1877), .Y(n1859)
         );
  AOI22X1TS U2195 ( .A0(\destinationAddressbuffer[2][8] ), .A1(n1965), .B0(
        \destinationAddressbuffer[0][8] ), .B1(n1966), .Y(n1856) );
  AOI22X1TS U2196 ( .A0(\destinationAddressbuffer[6][8] ), .A1(n1967), .B0(
        \destinationAddressbuffer[4][8] ), .B1(n1968), .Y(n1855) );
  AOI22X1TS U2197 ( .A0(\destinationAddressbuffer[3][8] ), .A1(n1969), .B0(
        \destinationAddressbuffer[1][8] ), .B1(n1970), .Y(n1854) );
  AOI22X1TS U2198 ( .A0(\destinationAddressbuffer[7][8] ), .A1(n1971), .B0(
        \destinationAddressbuffer[5][8] ), .B1(n1972), .Y(n1853) );
  NAND4XLTS U2199 ( .A(n1856), .B(n1855), .C(n1854), .D(n1853), .Y(n1857) );
  AOI22X1TS U2200 ( .A0(destinationAddressOut[8]), .A1(n1978), .B0(n2459), 
        .B1(n1857), .Y(n1858) );
  AOI22X1TS U2201 ( .A0(n1369), .A1(n1961), .B0(n1370), .B1(n1964), .Y(n1868)
         );
  AOI22X1TS U2202 ( .A0(n1373), .A1(n1682), .B0(n1371), .B1(n1877), .Y(n1867)
         );
  AOI22X1TS U2203 ( .A0(\destinationAddressbuffer[2][9] ), .A1(n1965), .B0(
        \destinationAddressbuffer[0][9] ), .B1(n1966), .Y(n1864) );
  AOI22X1TS U2204 ( .A0(\destinationAddressbuffer[6][9] ), .A1(n1967), .B0(
        \destinationAddressbuffer[4][9] ), .B1(n1968), .Y(n1863) );
  AOI22X1TS U2205 ( .A0(\destinationAddressbuffer[3][9] ), .A1(n1969), .B0(
        \destinationAddressbuffer[1][9] ), .B1(n1970), .Y(n1862) );
  AOI22X1TS U2206 ( .A0(\destinationAddressbuffer[7][9] ), .A1(n1971), .B0(
        \destinationAddressbuffer[5][9] ), .B1(n1972), .Y(n1861) );
  NAND4XLTS U2207 ( .A(n1864), .B(n1863), .C(n1862), .D(n1861), .Y(n1865) );
  AOI22X1TS U2208 ( .A0(destinationAddressOut[9]), .A1(n1978), .B0(n2459), 
        .B1(n1865), .Y(n1866) );
  AOI22X1TS U2209 ( .A0(n1376), .A1(n1961), .B0(n1377), .B1(n1964), .Y(n1876)
         );
  AOI22X1TS U2210 ( .A0(n1380), .A1(n1682), .B0(n1378), .B1(n1877), .Y(n1875)
         );
  AOI22X1TS U2211 ( .A0(\destinationAddressbuffer[2][10] ), .A1(n1890), .B0(
        \destinationAddressbuffer[0][10] ), .B1(n1966), .Y(n1872) );
  AOI22X1TS U2212 ( .A0(\destinationAddressbuffer[6][10] ), .A1(n1891), .B0(
        \destinationAddressbuffer[4][10] ), .B1(n1968), .Y(n1871) );
  AOI22X1TS U2213 ( .A0(\destinationAddressbuffer[3][10] ), .A1(n1969), .B0(
        \destinationAddressbuffer[1][10] ), .B1(n1970), .Y(n1870) );
  AOI22X1TS U2214 ( .A0(\destinationAddressbuffer[7][10] ), .A1(n1971), .B0(
        \destinationAddressbuffer[5][10] ), .B1(n1972), .Y(n1869) );
  NAND4XLTS U2215 ( .A(n1872), .B(n1871), .C(n1870), .D(n1869), .Y(n1873) );
  AOI22X1TS U2216 ( .A0(destinationAddressOut[10]), .A1(n1978), .B0(n2459), 
        .B1(n1873), .Y(n1874) );
  AOI22X1TS U2217 ( .A0(n1383), .A1(n1961), .B0(n1384), .B1(n1964), .Y(n1885)
         );
  AOI22X1TS U2218 ( .A0(n1387), .A1(n1682), .B0(n1385), .B1(n1877), .Y(n1884)
         );
  AOI22X1TS U2219 ( .A0(\destinationAddressbuffer[2][11] ), .A1(n1890), .B0(
        \destinationAddressbuffer[0][11] ), .B1(n1966), .Y(n1881) );
  AOI22X1TS U2220 ( .A0(\destinationAddressbuffer[6][11] ), .A1(n1891), .B0(
        \destinationAddressbuffer[4][11] ), .B1(n1968), .Y(n1880) );
  AOI22X1TS U2221 ( .A0(\destinationAddressbuffer[3][11] ), .A1(n1969), .B0(
        \destinationAddressbuffer[1][11] ), .B1(n1970), .Y(n1879) );
  AOI22X1TS U2222 ( .A0(\destinationAddressbuffer[7][11] ), .A1(n1971), .B0(
        \destinationAddressbuffer[5][11] ), .B1(n1972), .Y(n1878) );
  NAND4XLTS U2223 ( .A(n1881), .B(n1880), .C(n1879), .D(n1878), .Y(n1882) );
  AOI22X1TS U2224 ( .A0(destinationAddressOut[11]), .A1(n1978), .B0(n2459), 
        .B1(n1882), .Y(n1883) );
  CLKBUFX2TS U2225 ( .A(dataIn_NORTH[0]), .Y(n1886) );
  CLKBUFX2TS U2226 ( .A(dataIn_EAST[0]), .Y(n1887) );
  AOI22X1TS U2227 ( .A0(n1886), .A1(n1682), .B0(n1887), .B1(n1961), .Y(n1901)
         );
  CLKBUFX2TS U2228 ( .A(dataIn_SOUTH[0]), .Y(n1888) );
  CLKBUFX2TS U2229 ( .A(dataIn_WEST[0]), .Y(n1889) );
  AOI22X1TS U2230 ( .A0(n1888), .A1(n1877), .B0(n1889), .B1(n1964), .Y(n1900)
         );
  AOI22X1TS U2231 ( .A0(\dataoutbuffer[0][0] ), .A1(n1966), .B0(
        \dataoutbuffer[2][0] ), .B1(n1890), .Y(n1895) );
  AOI22X1TS U2232 ( .A0(\dataoutbuffer[4][0] ), .A1(n1968), .B0(
        \dataoutbuffer[6][0] ), .B1(n1891), .Y(n1894) );
  AOI22X1TS U2233 ( .A0(\dataoutbuffer[1][0] ), .A1(n1970), .B0(
        \dataoutbuffer[3][0] ), .B1(n1969), .Y(n1893) );
  AOI22X1TS U2234 ( .A0(\dataoutbuffer[5][0] ), .A1(n1972), .B0(
        \dataoutbuffer[7][0] ), .B1(n1971), .Y(n1892) );
  NAND4XLTS U2235 ( .A(n1895), .B(n1894), .C(n1893), .D(n1892), .Y(n1896) );
  AOI22X1TS U2236 ( .A0(dataOut[0]), .A1(n1978), .B0(n2459), .B1(n1896), .Y(
        n1899) );
  CLKBUFX2TS U2237 ( .A(cacheDataOut[0]), .Y(n1897) );
  NAND2X1TS U2238 ( .A(n1897), .B(n1980), .Y(n1898) );
  CLKBUFX2TS U2239 ( .A(dataIn_NORTH[1]), .Y(n1902) );
  CLKBUFX2TS U2240 ( .A(dataIn_EAST[1]), .Y(n1903) );
  AOI22X1TS U2241 ( .A0(n1902), .A1(n1682), .B0(n1903), .B1(n1918), .Y(n1915)
         );
  CLKBUFX2TS U2242 ( .A(dataIn_SOUTH[1]), .Y(n1904) );
  CLKBUFX2TS U2243 ( .A(dataIn_WEST[1]), .Y(n1905) );
  AOI22X1TS U2244 ( .A0(n1904), .A1(n1877), .B0(n1905), .B1(n1964), .Y(n1914)
         );
  AOI22X1TS U2245 ( .A0(\dataoutbuffer[0][1] ), .A1(n1966), .B0(
        \dataoutbuffer[2][1] ), .B1(n1965), .Y(n1909) );
  AOI22X1TS U2246 ( .A0(\dataoutbuffer[4][1] ), .A1(n1968), .B0(
        \dataoutbuffer[6][1] ), .B1(n1967), .Y(n1908) );
  AOI22X1TS U2247 ( .A0(\dataoutbuffer[1][1] ), .A1(n1970), .B0(
        \dataoutbuffer[3][1] ), .B1(n1969), .Y(n1907) );
  AOI22X1TS U2248 ( .A0(\dataoutbuffer[5][1] ), .A1(n1972), .B0(
        \dataoutbuffer[7][1] ), .B1(n1971), .Y(n1906) );
  NAND4XLTS U2249 ( .A(n1909), .B(n1908), .C(n1907), .D(n1906), .Y(n1910) );
  AOI22X1TS U2250 ( .A0(dataOut[1]), .A1(n1978), .B0(n2459), .B1(n1910), .Y(
        n1913) );
  CLKBUFX2TS U2251 ( .A(cacheDataOut[1]), .Y(n1911) );
  NAND2X1TS U2252 ( .A(n1911), .B(n1980), .Y(n1912) );
  CLKBUFX2TS U2253 ( .A(dataIn_NORTH[2]), .Y(n1916) );
  CLKBUFX2TS U2254 ( .A(dataIn_EAST[2]), .Y(n1917) );
  AOI22X1TS U2255 ( .A0(n1916), .A1(n1682), .B0(n1917), .B1(n1918), .Y(n1930)
         );
  CLKBUFX2TS U2256 ( .A(dataIn_SOUTH[2]), .Y(n1919) );
  CLKBUFX2TS U2257 ( .A(dataIn_WEST[2]), .Y(n1920) );
  AOI22X1TS U2258 ( .A0(n1919), .A1(n1877), .B0(n1920), .B1(n1964), .Y(n1929)
         );
  AOI22X1TS U2259 ( .A0(\dataoutbuffer[0][2] ), .A1(n1966), .B0(
        \dataoutbuffer[2][2] ), .B1(n1965), .Y(n1924) );
  AOI22X1TS U2260 ( .A0(\dataoutbuffer[4][2] ), .A1(n1968), .B0(
        \dataoutbuffer[6][2] ), .B1(n1967), .Y(n1923) );
  AOI22X1TS U2261 ( .A0(\dataoutbuffer[1][2] ), .A1(n1970), .B0(
        \dataoutbuffer[3][2] ), .B1(n1969), .Y(n1922) );
  AOI22X1TS U2262 ( .A0(\dataoutbuffer[5][2] ), .A1(n1972), .B0(
        \dataoutbuffer[7][2] ), .B1(n1971), .Y(n1921) );
  NAND4XLTS U2263 ( .A(n1924), .B(n1923), .C(n1922), .D(n1921), .Y(n1925) );
  AOI22X1TS U2264 ( .A0(dataOut[2]), .A1(n1978), .B0(n2459), .B1(n1925), .Y(
        n1928) );
  CLKBUFX2TS U2265 ( .A(cacheDataOut[2]), .Y(n1926) );
  NAND2X1TS U2266 ( .A(n1926), .B(n1980), .Y(n1927) );
  CLKBUFX2TS U2267 ( .A(dataIn_NORTH[3]), .Y(n1931) );
  CLKBUFX2TS U2268 ( .A(dataIn_EAST[3]), .Y(n1932) );
  AOI22X1TS U2269 ( .A0(n1931), .A1(n1682), .B0(n1932), .B1(n1961), .Y(n1944)
         );
  CLKBUFX2TS U2270 ( .A(dataIn_SOUTH[3]), .Y(n1933) );
  CLKBUFX2TS U2271 ( .A(dataIn_WEST[3]), .Y(n1934) );
  AOI22X1TS U2272 ( .A0(n1933), .A1(n1877), .B0(n1934), .B1(n1964), .Y(n1943)
         );
  AOI22X1TS U2273 ( .A0(\dataoutbuffer[0][3] ), .A1(n1966), .B0(
        \dataoutbuffer[2][3] ), .B1(n1965), .Y(n1938) );
  AOI22X1TS U2274 ( .A0(\dataoutbuffer[4][3] ), .A1(n1968), .B0(
        \dataoutbuffer[6][3] ), .B1(n1967), .Y(n1937) );
  AOI22X1TS U2275 ( .A0(\dataoutbuffer[1][3] ), .A1(n1970), .B0(
        \dataoutbuffer[3][3] ), .B1(n1969), .Y(n1936) );
  AOI22X1TS U2276 ( .A0(\dataoutbuffer[5][3] ), .A1(n1972), .B0(
        \dataoutbuffer[7][3] ), .B1(n1971), .Y(n1935) );
  NAND4XLTS U2277 ( .A(n1938), .B(n1937), .C(n1936), .D(n1935), .Y(n1939) );
  AOI22X1TS U2278 ( .A0(dataOut[3]), .A1(n1978), .B0(n2459), .B1(n1939), .Y(
        n1942) );
  CLKBUFX2TS U2279 ( .A(cacheDataOut[3]), .Y(n1940) );
  NAND2X1TS U2280 ( .A(n1940), .B(n1980), .Y(n1941) );
  CLKBUFX2TS U2281 ( .A(dataIn_NORTH[4]), .Y(n1945) );
  CLKBUFX2TS U2282 ( .A(dataIn_EAST[4]), .Y(n1946) );
  AOI22X1TS U2283 ( .A0(n1945), .A1(n1682), .B0(n1946), .B1(n1961), .Y(n1958)
         );
  CLKBUFX2TS U2284 ( .A(dataIn_SOUTH[4]), .Y(n1947) );
  CLKBUFX2TS U2285 ( .A(dataIn_WEST[4]), .Y(n1948) );
  AOI22X1TS U2286 ( .A0(n1947), .A1(n1877), .B0(n1948), .B1(n1964), .Y(n1957)
         );
  AOI22X1TS U2287 ( .A0(\dataoutbuffer[0][4] ), .A1(n1966), .B0(
        \dataoutbuffer[2][4] ), .B1(n1965), .Y(n1952) );
  AOI22X1TS U2288 ( .A0(\dataoutbuffer[4][4] ), .A1(n1968), .B0(
        \dataoutbuffer[6][4] ), .B1(n1967), .Y(n1951) );
  AOI22X1TS U2289 ( .A0(\dataoutbuffer[1][4] ), .A1(n1970), .B0(
        \dataoutbuffer[3][4] ), .B1(n1969), .Y(n1950) );
  AOI22X1TS U2290 ( .A0(\dataoutbuffer[5][4] ), .A1(n1972), .B0(
        \dataoutbuffer[7][4] ), .B1(n1971), .Y(n1949) );
  NAND4XLTS U2291 ( .A(n1952), .B(n1951), .C(n1950), .D(n1949), .Y(n1953) );
  AOI22X1TS U2292 ( .A0(dataOut[4]), .A1(n1978), .B0(n2459), .B1(n1953), .Y(
        n1956) );
  CLKBUFX2TS U2293 ( .A(cacheDataOut[4]), .Y(n1954) );
  NAND2X1TS U2294 ( .A(n1954), .B(n1980), .Y(n1955) );
  CLKBUFX2TS U2295 ( .A(dataIn_NORTH[5]), .Y(n1959) );
  CLKBUFX2TS U2296 ( .A(dataIn_EAST[5]), .Y(n1960) );
  AOI22X1TS U2297 ( .A0(n1959), .A1(n1682), .B0(n1960), .B1(n1961), .Y(n1984)
         );
  CLKBUFX2TS U2298 ( .A(dataIn_SOUTH[5]), .Y(n1962) );
  CLKBUFX2TS U2299 ( .A(dataIn_WEST[5]), .Y(n1963) );
  AOI22X1TS U2300 ( .A0(n1962), .A1(n1877), .B0(n1963), .B1(n1964), .Y(n1983)
         );
  AOI22X1TS U2301 ( .A0(\dataoutbuffer[0][5] ), .A1(n1966), .B0(
        \dataoutbuffer[2][5] ), .B1(n1965), .Y(n1976) );
  AOI22X1TS U2302 ( .A0(\dataoutbuffer[4][5] ), .A1(n1968), .B0(
        \dataoutbuffer[6][5] ), .B1(n1967), .Y(n1975) );
  AOI22X1TS U2303 ( .A0(\dataoutbuffer[1][5] ), .A1(n1970), .B0(
        \dataoutbuffer[3][5] ), .B1(n1969), .Y(n1974) );
  AOI22X1TS U2304 ( .A0(\dataoutbuffer[5][5] ), .A1(n1972), .B0(
        \dataoutbuffer[7][5] ), .B1(n1971), .Y(n1973) );
  NAND4XLTS U2305 ( .A(n1976), .B(n1975), .C(n1974), .D(n1973), .Y(n1977) );
  AOI22X1TS U2306 ( .A0(dataOut[5]), .A1(n1978), .B0(n2459), .B1(n1977), .Y(
        n1982) );
  CLKBUFX2TS U2307 ( .A(cacheDataOut[5]), .Y(n1979) );
  NAND2X1TS U2308 ( .A(n1979), .B(n1980), .Y(n1981) );
  AOI22X1TS U2309 ( .A0(n1720), .A1(n2324), .B0(n2323), .B1(
        \requesterAddressbuffer[7][0] ), .Y(n1987) );
  AOI22X1TS U2310 ( .A0(n2326), .A1(n1714), .B0(n2325), .B1(n1712), .Y(n1986)
         );
  AOI22X1TS U2311 ( .A0(n2328), .A1(n1713), .B0(n2327), .B1(n1711), .Y(n1985)
         );
  AOI22X1TS U2312 ( .A0(n2324), .A1(n1734), .B0(n2323), .B1(
        \requesterAddressbuffer[7][1] ), .Y(n1990) );
  AOI22X1TS U2313 ( .A0(n2326), .A1(n1728), .B0(n2325), .B1(n1726), .Y(n1989)
         );
  AOI22X1TS U2314 ( .A0(n2328), .A1(n1727), .B0(n2327), .B1(n1725), .Y(n1988)
         );
  AOI22X1TS U2315 ( .A0(n2324), .A1(n1747), .B0(n2323), .B1(
        \requesterAddressbuffer[7][2] ), .Y(n1993) );
  AOI22X1TS U2316 ( .A0(n2326), .A1(n1741), .B0(n2325), .B1(n1739), .Y(n1992)
         );
  AOI22X1TS U2317 ( .A0(n2328), .A1(n1740), .B0(n2327), .B1(n1738), .Y(n1991)
         );
  AOI22X1TS U2318 ( .A0(n2324), .A1(n1760), .B0(n2323), .B1(
        \requesterAddressbuffer[7][3] ), .Y(n1996) );
  AOI22X1TS U2319 ( .A0(n2326), .A1(n1754), .B0(n2325), .B1(n1752), .Y(n1995)
         );
  AOI22X1TS U2320 ( .A0(n2328), .A1(n1753), .B0(n2327), .B1(n1751), .Y(n1994)
         );
  AOI22X1TS U2321 ( .A0(n1720), .A1(n2342), .B0(n2341), .B1(
        \requesterAddressbuffer[6][0] ), .Y(n1999) );
  AOI22X1TS U2322 ( .A0(n1714), .A1(n2344), .B0(n1712), .B1(n2343), .Y(n1998)
         );
  AOI22X1TS U2323 ( .A0(n1713), .A1(n2345), .B0(n1711), .B1(n2346), .Y(n1997)
         );
  AOI22X1TS U2324 ( .A0(n1734), .A1(n2342), .B0(n2341), .B1(
        \requesterAddressbuffer[6][1] ), .Y(n2002) );
  AOI22X1TS U2325 ( .A0(n1728), .A1(n2344), .B0(n1726), .B1(n2343), .Y(n2001)
         );
  AOI22X1TS U2326 ( .A0(n1727), .A1(n2345), .B0(n1725), .B1(n2346), .Y(n2000)
         );
  AOI22X1TS U2327 ( .A0(n1747), .A1(n2342), .B0(n2341), .B1(
        \requesterAddressbuffer[6][2] ), .Y(n2005) );
  AOI22X1TS U2328 ( .A0(n1741), .A1(n2344), .B0(n1739), .B1(n2343), .Y(n2004)
         );
  AOI22X1TS U2329 ( .A0(n1740), .A1(n2345), .B0(n1738), .B1(n2346), .Y(n2003)
         );
  AOI22X1TS U2330 ( .A0(n1760), .A1(n2342), .B0(n2341), .B1(
        \requesterAddressbuffer[6][3] ), .Y(n2008) );
  AOI22X1TS U2331 ( .A0(n1754), .A1(n2344), .B0(n1752), .B1(n2343), .Y(n2007)
         );
  AOI22X1TS U2332 ( .A0(n1753), .A1(n2345), .B0(n1751), .B1(n2346), .Y(n2006)
         );
  AOI22X1TS U2333 ( .A0(n1720), .A1(n1337), .B0(n2359), .B1(
        \requesterAddressbuffer[5][0] ), .Y(n2011) );
  AOI22X1TS U2334 ( .A0(n1714), .A1(n2361), .B0(n1712), .B1(n2360), .Y(n2010)
         );
  AOI22X1TS U2335 ( .A0(n1713), .A1(n2362), .B0(n1711), .B1(n2363), .Y(n2009)
         );
  AOI22X1TS U2336 ( .A0(n1734), .A1(n1337), .B0(n2359), .B1(
        \requesterAddressbuffer[5][1] ), .Y(n2014) );
  AOI22X1TS U2337 ( .A0(n1728), .A1(n2361), .B0(n1726), .B1(n2360), .Y(n2013)
         );
  AOI22X1TS U2338 ( .A0(n1727), .A1(n2362), .B0(n1725), .B1(n2363), .Y(n2012)
         );
  AOI22X1TS U2339 ( .A0(n1747), .A1(n1337), .B0(n2359), .B1(
        \requesterAddressbuffer[5][2] ), .Y(n2017) );
  AOI22X1TS U2340 ( .A0(n1741), .A1(n2361), .B0(n1739), .B1(n2360), .Y(n2016)
         );
  AOI22X1TS U2341 ( .A0(n1740), .A1(n2362), .B0(n1738), .B1(n2363), .Y(n2015)
         );
  AOI22X1TS U2342 ( .A0(n1760), .A1(n1337), .B0(n2359), .B1(
        \requesterAddressbuffer[5][3] ), .Y(n2020) );
  AOI22X1TS U2343 ( .A0(n1754), .A1(n2361), .B0(n1752), .B1(n2360), .Y(n2019)
         );
  AOI22X1TS U2344 ( .A0(n1753), .A1(n2362), .B0(n1751), .B1(n2363), .Y(n2018)
         );
  AOI22X1TS U2345 ( .A0(n1720), .A1(n2377), .B0(n2376), .B1(
        \requesterAddressbuffer[4][0] ), .Y(n2023) );
  AOI22X1TS U2346 ( .A0(n1714), .A1(n2379), .B0(n1712), .B1(n2378), .Y(n2022)
         );
  AOI22X1TS U2347 ( .A0(n1713), .A1(n2381), .B0(n1711), .B1(n2380), .Y(n2021)
         );
  AOI22X1TS U2348 ( .A0(n1734), .A1(n2377), .B0(n2376), .B1(
        \requesterAddressbuffer[4][1] ), .Y(n2026) );
  AOI22X1TS U2349 ( .A0(n1728), .A1(n2379), .B0(n1726), .B1(n2378), .Y(n2025)
         );
  AOI22X1TS U2350 ( .A0(n1727), .A1(n2381), .B0(n1725), .B1(n2380), .Y(n2024)
         );
  AOI22X1TS U2351 ( .A0(n1747), .A1(n2377), .B0(n2376), .B1(
        \requesterAddressbuffer[4][2] ), .Y(n2029) );
  AOI22X1TS U2352 ( .A0(n1741), .A1(n2379), .B0(n1739), .B1(n2378), .Y(n2028)
         );
  AOI22X1TS U2353 ( .A0(n1740), .A1(n2381), .B0(n1738), .B1(n2380), .Y(n2027)
         );
  AOI22X1TS U2354 ( .A0(n1760), .A1(n2377), .B0(n2376), .B1(
        \requesterAddressbuffer[4][3] ), .Y(n2032) );
  AOI22X1TS U2355 ( .A0(n1754), .A1(n2379), .B0(n1752), .B1(n2378), .Y(n2031)
         );
  AOI22X1TS U2356 ( .A0(n1753), .A1(n2381), .B0(n1751), .B1(n2380), .Y(n2030)
         );
  AOI22X1TS U2357 ( .A0(n1720), .A1(n2395), .B0(n2394), .B1(
        \requesterAddressbuffer[3][0] ), .Y(n2035) );
  AOI22X1TS U2358 ( .A0(n1714), .A1(n2396), .B0(n1712), .B1(n1510), .Y(n2034)
         );
  AOI22X1TS U2359 ( .A0(n1713), .A1(n2397), .B0(n1711), .B1(n2398), .Y(n2033)
         );
  AOI22X1TS U2360 ( .A0(n1734), .A1(n2395), .B0(n2394), .B1(
        \requesterAddressbuffer[3][1] ), .Y(n2038) );
  AOI22X1TS U2361 ( .A0(n1728), .A1(n2396), .B0(n1726), .B1(n1510), .Y(n2037)
         );
  AOI22X1TS U2362 ( .A0(n1727), .A1(n2397), .B0(n1725), .B1(n2398), .Y(n2036)
         );
  AOI22X1TS U2363 ( .A0(n1747), .A1(n2395), .B0(n2394), .B1(
        \requesterAddressbuffer[3][2] ), .Y(n2041) );
  AOI22X1TS U2364 ( .A0(n1741), .A1(n2396), .B0(n1739), .B1(n1510), .Y(n2040)
         );
  AOI22X1TS U2365 ( .A0(n1740), .A1(n2397), .B0(n1738), .B1(n2398), .Y(n2039)
         );
  AOI22X1TS U2366 ( .A0(n1760), .A1(n2395), .B0(n2394), .B1(
        \requesterAddressbuffer[3][3] ), .Y(n2044) );
  AOI22X1TS U2367 ( .A0(n1754), .A1(n2396), .B0(n1752), .B1(n1510), .Y(n2043)
         );
  AOI22X1TS U2368 ( .A0(n1753), .A1(n2397), .B0(n1751), .B1(n2398), .Y(n2042)
         );
  AOI22X1TS U2369 ( .A0(n1720), .A1(n2412), .B0(n2411), .B1(
        \requesterAddressbuffer[2][0] ), .Y(n2047) );
  AOI22X1TS U2370 ( .A0(n1714), .A1(n2414), .B0(n1712), .B1(n2413), .Y(n2046)
         );
  AOI22X1TS U2371 ( .A0(n1713), .A1(n2415), .B0(n1711), .B1(n2416), .Y(n2045)
         );
  AOI22X1TS U2372 ( .A0(n1734), .A1(n2412), .B0(n2411), .B1(
        \requesterAddressbuffer[2][1] ), .Y(n2050) );
  AOI22X1TS U2373 ( .A0(n1728), .A1(n2414), .B0(n1726), .B1(n2413), .Y(n2049)
         );
  AOI22X1TS U2374 ( .A0(n1727), .A1(n2415), .B0(n1725), .B1(n2416), .Y(n2048)
         );
  AOI22X1TS U2375 ( .A0(n1747), .A1(n2412), .B0(n2411), .B1(
        \requesterAddressbuffer[2][2] ), .Y(n2053) );
  AOI22X1TS U2376 ( .A0(n1741), .A1(n2414), .B0(n1739), .B1(n2413), .Y(n2052)
         );
  AOI22X1TS U2377 ( .A0(n1740), .A1(n2415), .B0(n1738), .B1(n2416), .Y(n2051)
         );
  AOI22X1TS U2378 ( .A0(n1760), .A1(n2412), .B0(n2411), .B1(
        \requesterAddressbuffer[2][3] ), .Y(n2056) );
  AOI22X1TS U2379 ( .A0(n1754), .A1(n2414), .B0(n1752), .B1(n2413), .Y(n2055)
         );
  AOI22X1TS U2380 ( .A0(n1753), .A1(n2415), .B0(n1751), .B1(n2416), .Y(n2054)
         );
  AOI22X1TS U2381 ( .A0(n1720), .A1(n2430), .B0(n2429), .B1(
        \requesterAddressbuffer[1][0] ), .Y(n2059) );
  AOI22X1TS U2382 ( .A0(n1714), .A1(n2432), .B0(n1712), .B1(n2431), .Y(n2058)
         );
  AOI22X1TS U2383 ( .A0(n1713), .A1(n2433), .B0(n1711), .B1(n2434), .Y(n2057)
         );
  AOI22X1TS U2384 ( .A0(n1734), .A1(n2430), .B0(n2429), .B1(
        \requesterAddressbuffer[1][1] ), .Y(n2062) );
  AOI22X1TS U2385 ( .A0(n1728), .A1(n2432), .B0(n1726), .B1(n2431), .Y(n2061)
         );
  AOI22X1TS U2386 ( .A0(n1727), .A1(n2433), .B0(n1725), .B1(n2434), .Y(n2060)
         );
  AOI22X1TS U2387 ( .A0(n1747), .A1(n2430), .B0(n2429), .B1(
        \requesterAddressbuffer[1][2] ), .Y(n2065) );
  AOI22X1TS U2388 ( .A0(n1741), .A1(n2432), .B0(n1739), .B1(n2431), .Y(n2064)
         );
  AOI22X1TS U2389 ( .A0(n1740), .A1(n2433), .B0(n1738), .B1(n2434), .Y(n2063)
         );
  AOI22X1TS U2390 ( .A0(n1760), .A1(n2430), .B0(n2429), .B1(
        \requesterAddressbuffer[1][3] ), .Y(n2068) );
  AOI22X1TS U2391 ( .A0(n1754), .A1(n2432), .B0(n1752), .B1(n2431), .Y(n2067)
         );
  AOI22X1TS U2392 ( .A0(n1753), .A1(n2433), .B0(n1751), .B1(n2434), .Y(n2066)
         );
  AOI22X1TS U2393 ( .A0(n1720), .A1(n2448), .B0(n2447), .B1(
        \requesterAddressbuffer[0][0] ), .Y(n2071) );
  AOI22X1TS U2394 ( .A0(n1714), .A1(n2450), .B0(n1712), .B1(n2449), .Y(n2070)
         );
  AOI22X1TS U2395 ( .A0(n1713), .A1(n2452), .B0(n1711), .B1(n2451), .Y(n2069)
         );
  AOI22X1TS U2396 ( .A0(n1734), .A1(n2448), .B0(n2447), .B1(
        \requesterAddressbuffer[0][1] ), .Y(n2074) );
  AOI22X1TS U2397 ( .A0(n1728), .A1(n2450), .B0(n1726), .B1(n2449), .Y(n2073)
         );
  AOI22X1TS U2398 ( .A0(n1727), .A1(n2452), .B0(n1725), .B1(n2451), .Y(n2072)
         );
  AOI22X1TS U2399 ( .A0(n1747), .A1(n2448), .B0(n2447), .B1(
        \requesterAddressbuffer[0][2] ), .Y(n2077) );
  AOI22X1TS U2400 ( .A0(n1741), .A1(n2450), .B0(n1739), .B1(n2449), .Y(n2076)
         );
  AOI22X1TS U2401 ( .A0(n1740), .A1(n2452), .B0(n1738), .B1(n2451), .Y(n2075)
         );
  AOI22X1TS U2402 ( .A0(n1760), .A1(n2448), .B0(n2447), .B1(
        \requesterAddressbuffer[0][3] ), .Y(n2080) );
  AOI22X1TS U2403 ( .A0(n1754), .A1(n2450), .B0(n1752), .B1(n2449), .Y(n2079)
         );
  AOI22X1TS U2404 ( .A0(n1753), .A1(n2452), .B0(n1751), .B1(n2451), .Y(n2078)
         );
  AOI22X1TS U2405 ( .A0(n2448), .A1(n1897), .B0(n2447), .B1(
        \dataoutbuffer[0][0] ), .Y(n2083) );
  AOI22X1TS U2406 ( .A0(n2450), .A1(n1889), .B0(n2449), .B1(n1887), .Y(n2082)
         );
  AOI22X1TS U2407 ( .A0(n2452), .A1(n1888), .B0(n2451), .B1(n1886), .Y(n2081)
         );
  AOI22X1TS U2408 ( .A0(n2448), .A1(n1911), .B0(n2447), .B1(
        \dataoutbuffer[0][1] ), .Y(n2086) );
  AOI22X1TS U2409 ( .A0(n2450), .A1(n1905), .B0(n2449), .B1(n1903), .Y(n2085)
         );
  AOI22X1TS U2410 ( .A0(n2452), .A1(n1904), .B0(n2451), .B1(n1902), .Y(n2084)
         );
  AOI22X1TS U2411 ( .A0(n2448), .A1(n1926), .B0(n2447), .B1(
        \dataoutbuffer[0][2] ), .Y(n2089) );
  AOI22X1TS U2412 ( .A0(n2450), .A1(n1920), .B0(n2449), .B1(n1917), .Y(n2088)
         );
  AOI22X1TS U2413 ( .A0(n2452), .A1(n1919), .B0(n2451), .B1(n1916), .Y(n2087)
         );
  AOI22X1TS U2414 ( .A0(n2448), .A1(n1940), .B0(n2447), .B1(
        \dataoutbuffer[0][3] ), .Y(n2092) );
  AOI22X1TS U2415 ( .A0(n2450), .A1(n1934), .B0(n2449), .B1(n1932), .Y(n2091)
         );
  AOI22X1TS U2416 ( .A0(n2452), .A1(n1933), .B0(n2451), .B1(n1931), .Y(n2090)
         );
  AOI22X1TS U2417 ( .A0(n2448), .A1(n1954), .B0(n2447), .B1(
        \dataoutbuffer[0][4] ), .Y(n2095) );
  AOI22X1TS U2418 ( .A0(n2450), .A1(n1948), .B0(n2449), .B1(n1946), .Y(n2094)
         );
  AOI22X1TS U2419 ( .A0(n2452), .A1(n1947), .B0(n2451), .B1(n1945), .Y(n2093)
         );
  AOI22X1TS U2420 ( .A0(n2448), .A1(n1979), .B0(n2447), .B1(
        \dataoutbuffer[0][5] ), .Y(n2098) );
  AOI22X1TS U2421 ( .A0(n2450), .A1(n1963), .B0(n2449), .B1(n1960), .Y(n2097)
         );
  AOI22X1TS U2422 ( .A0(n2452), .A1(n1962), .B0(n2451), .B1(n1959), .Y(n2096)
         );
  AOI22X1TS U2423 ( .A0(n2430), .A1(n1897), .B0(n2429), .B1(
        \dataoutbuffer[1][0] ), .Y(n2101) );
  AOI22X1TS U2424 ( .A0(n2432), .A1(n1889), .B0(n2431), .B1(n1887), .Y(n2100)
         );
  AOI22X1TS U2425 ( .A0(n2434), .A1(n1886), .B0(n2433), .B1(n1888), .Y(n2099)
         );
  AOI22X1TS U2426 ( .A0(n2430), .A1(n1911), .B0(n2429), .B1(
        \dataoutbuffer[1][1] ), .Y(n2104) );
  AOI22X1TS U2427 ( .A0(n2432), .A1(n1905), .B0(n2431), .B1(n1903), .Y(n2103)
         );
  AOI22X1TS U2428 ( .A0(n2434), .A1(n1902), .B0(n2433), .B1(n1904), .Y(n2102)
         );
  AOI22X1TS U2429 ( .A0(n2430), .A1(n1926), .B0(n2429), .B1(
        \dataoutbuffer[1][2] ), .Y(n2107) );
  AOI22X1TS U2430 ( .A0(n2432), .A1(n1920), .B0(n2431), .B1(n1917), .Y(n2106)
         );
  AOI22X1TS U2431 ( .A0(n2434), .A1(n1916), .B0(n2433), .B1(n1919), .Y(n2105)
         );
  AOI22X1TS U2432 ( .A0(n2430), .A1(n1940), .B0(n2429), .B1(
        \dataoutbuffer[1][3] ), .Y(n2110) );
  AOI22X1TS U2433 ( .A0(n2432), .A1(n1934), .B0(n2431), .B1(n1932), .Y(n2109)
         );
  AOI22X1TS U2434 ( .A0(n2434), .A1(n1931), .B0(n2433), .B1(n1933), .Y(n2108)
         );
  AOI22X1TS U2435 ( .A0(n2430), .A1(n1954), .B0(n2429), .B1(
        \dataoutbuffer[1][4] ), .Y(n2113) );
  AOI22X1TS U2436 ( .A0(n2432), .A1(n1948), .B0(n2431), .B1(n1946), .Y(n2112)
         );
  AOI22X1TS U2437 ( .A0(n2434), .A1(n1945), .B0(n2433), .B1(n1947), .Y(n2111)
         );
  AOI22X1TS U2438 ( .A0(n2430), .A1(n1979), .B0(n2429), .B1(
        \dataoutbuffer[1][5] ), .Y(n2116) );
  AOI22X1TS U2439 ( .A0(n2432), .A1(n1963), .B0(n2431), .B1(n1960), .Y(n2115)
         );
  AOI22X1TS U2440 ( .A0(n2434), .A1(n1959), .B0(n2433), .B1(n1962), .Y(n2114)
         );
  AOI22X1TS U2441 ( .A0(n2412), .A1(n1897), .B0(n2411), .B1(
        \dataoutbuffer[2][0] ), .Y(n2119) );
  AOI22X1TS U2442 ( .A0(n2414), .A1(n1889), .B0(n2413), .B1(n1887), .Y(n2118)
         );
  AOI22X1TS U2443 ( .A0(n2416), .A1(n1886), .B0(n2415), .B1(n1888), .Y(n2117)
         );
  AOI22X1TS U2444 ( .A0(n2412), .A1(n1911), .B0(n2411), .B1(
        \dataoutbuffer[2][1] ), .Y(n2122) );
  AOI22X1TS U2445 ( .A0(n2414), .A1(n1905), .B0(n2413), .B1(n1903), .Y(n2121)
         );
  AOI22X1TS U2446 ( .A0(n2416), .A1(n1902), .B0(n2415), .B1(n1904), .Y(n2120)
         );
  AOI22X1TS U2447 ( .A0(n2412), .A1(n1926), .B0(n2411), .B1(
        \dataoutbuffer[2][2] ), .Y(n2125) );
  AOI22X1TS U2448 ( .A0(n2414), .A1(n1920), .B0(n2413), .B1(n1917), .Y(n2124)
         );
  AOI22X1TS U2449 ( .A0(n2416), .A1(n1916), .B0(n2415), .B1(n1919), .Y(n2123)
         );
  AOI22X1TS U2450 ( .A0(n2412), .A1(n1940), .B0(n2411), .B1(
        \dataoutbuffer[2][3] ), .Y(n2128) );
  AOI22X1TS U2451 ( .A0(n2414), .A1(n1934), .B0(n2413), .B1(n1932), .Y(n2127)
         );
  AOI22X1TS U2452 ( .A0(n2416), .A1(n1931), .B0(n2415), .B1(n1933), .Y(n2126)
         );
  AOI22X1TS U2453 ( .A0(n2412), .A1(n1954), .B0(n2411), .B1(
        \dataoutbuffer[2][4] ), .Y(n2131) );
  AOI22X1TS U2454 ( .A0(n2414), .A1(n1948), .B0(n2413), .B1(n1946), .Y(n2130)
         );
  AOI22X1TS U2455 ( .A0(n2416), .A1(n1945), .B0(n2415), .B1(n1947), .Y(n2129)
         );
  AOI22X1TS U2456 ( .A0(n2412), .A1(n1979), .B0(n2411), .B1(
        \dataoutbuffer[2][5] ), .Y(n2134) );
  AOI22X1TS U2457 ( .A0(n2414), .A1(n1963), .B0(n2413), .B1(n1960), .Y(n2133)
         );
  AOI22X1TS U2458 ( .A0(n2416), .A1(n1959), .B0(n2415), .B1(n1962), .Y(n2132)
         );
  AOI22X1TS U2459 ( .A0(n2395), .A1(n1897), .B0(n2394), .B1(
        \dataoutbuffer[3][0] ), .Y(n2137) );
  AOI22X1TS U2460 ( .A0(n2396), .A1(n1889), .B0(n1510), .B1(n1887), .Y(n2136)
         );
  AOI22X1TS U2461 ( .A0(n2398), .A1(n1886), .B0(n2397), .B1(n1888), .Y(n2135)
         );
  AOI22X1TS U2462 ( .A0(n2395), .A1(n1911), .B0(n2394), .B1(
        \dataoutbuffer[3][1] ), .Y(n2140) );
  AOI22X1TS U2463 ( .A0(n2396), .A1(n1905), .B0(n1510), .B1(n1903), .Y(n2139)
         );
  AOI22X1TS U2464 ( .A0(n2398), .A1(n1902), .B0(n2397), .B1(n1904), .Y(n2138)
         );
  AOI22X1TS U2465 ( .A0(n2395), .A1(n1926), .B0(n2394), .B1(
        \dataoutbuffer[3][2] ), .Y(n2143) );
  AOI22X1TS U2466 ( .A0(n2396), .A1(n1920), .B0(n1510), .B1(n1917), .Y(n2142)
         );
  AOI22X1TS U2467 ( .A0(n2398), .A1(n1916), .B0(n2397), .B1(n1919), .Y(n2141)
         );
  AOI22X1TS U2468 ( .A0(n2395), .A1(n1940), .B0(n2394), .B1(
        \dataoutbuffer[3][3] ), .Y(n2146) );
  AOI22X1TS U2469 ( .A0(n2396), .A1(n1934), .B0(n1510), .B1(n1932), .Y(n2145)
         );
  AOI22X1TS U2470 ( .A0(n2398), .A1(n1931), .B0(n2397), .B1(n1933), .Y(n2144)
         );
  AOI22X1TS U2471 ( .A0(n2395), .A1(n1954), .B0(n2394), .B1(
        \dataoutbuffer[3][4] ), .Y(n2149) );
  AOI22X1TS U2472 ( .A0(n2396), .A1(n1948), .B0(n1510), .B1(n1946), .Y(n2148)
         );
  AOI22X1TS U2473 ( .A0(n2398), .A1(n1945), .B0(n2397), .B1(n1947), .Y(n2147)
         );
  AOI22X1TS U2474 ( .A0(n2395), .A1(n1979), .B0(n2394), .B1(
        \dataoutbuffer[3][5] ), .Y(n2152) );
  AOI22X1TS U2475 ( .A0(n2396), .A1(n1963), .B0(n1510), .B1(n1960), .Y(n2151)
         );
  AOI22X1TS U2476 ( .A0(n2398), .A1(n1959), .B0(n2397), .B1(n1962), .Y(n2150)
         );
  AOI22X1TS U2477 ( .A0(n2377), .A1(n1897), .B0(n2376), .B1(
        \dataoutbuffer[4][0] ), .Y(n2155) );
  AOI22X1TS U2478 ( .A0(n2379), .A1(n1889), .B0(n2378), .B1(n1887), .Y(n2154)
         );
  AOI22X1TS U2479 ( .A0(n2381), .A1(n1888), .B0(n2380), .B1(n1886), .Y(n2153)
         );
  AOI22X1TS U2480 ( .A0(n2377), .A1(n1911), .B0(n2376), .B1(
        \dataoutbuffer[4][1] ), .Y(n2158) );
  AOI22X1TS U2481 ( .A0(n2379), .A1(n1905), .B0(n2378), .B1(n1903), .Y(n2157)
         );
  AOI22X1TS U2482 ( .A0(n2381), .A1(n1904), .B0(n2380), .B1(n1902), .Y(n2156)
         );
  AOI22X1TS U2483 ( .A0(n2377), .A1(n1926), .B0(n2376), .B1(
        \dataoutbuffer[4][2] ), .Y(n2161) );
  AOI22X1TS U2484 ( .A0(n2379), .A1(n1920), .B0(n2378), .B1(n1917), .Y(n2160)
         );
  AOI22X1TS U2485 ( .A0(n2381), .A1(n1919), .B0(n2380), .B1(n1916), .Y(n2159)
         );
  AOI22X1TS U2486 ( .A0(n2377), .A1(n1940), .B0(n2376), .B1(
        \dataoutbuffer[4][3] ), .Y(n2164) );
  AOI22X1TS U2487 ( .A0(n2379), .A1(n1934), .B0(n2378), .B1(n1932), .Y(n2163)
         );
  AOI22X1TS U2488 ( .A0(n2381), .A1(n1933), .B0(n2380), .B1(n1931), .Y(n2162)
         );
  AOI22X1TS U2489 ( .A0(n2377), .A1(n1954), .B0(n2376), .B1(
        \dataoutbuffer[4][4] ), .Y(n2167) );
  AOI22X1TS U2490 ( .A0(n2379), .A1(n1948), .B0(n2378), .B1(n1946), .Y(n2166)
         );
  AOI22X1TS U2491 ( .A0(n2381), .A1(n1947), .B0(n2380), .B1(n1945), .Y(n2165)
         );
  AOI22X1TS U2492 ( .A0(n2377), .A1(n1979), .B0(n2376), .B1(
        \dataoutbuffer[4][5] ), .Y(n2170) );
  AOI22X1TS U2493 ( .A0(n2379), .A1(n1963), .B0(n2378), .B1(n1960), .Y(n2169)
         );
  AOI22X1TS U2494 ( .A0(n2381), .A1(n1962), .B0(n2380), .B1(n1959), .Y(n2168)
         );
  AOI22X1TS U2495 ( .A0(n1337), .A1(n1897), .B0(n2359), .B1(
        \dataoutbuffer[5][0] ), .Y(n2173) );
  AOI22X1TS U2496 ( .A0(n2361), .A1(n1889), .B0(n2360), .B1(n1887), .Y(n2172)
         );
  AOI22X1TS U2497 ( .A0(n2363), .A1(n1886), .B0(n2362), .B1(n1888), .Y(n2171)
         );
  AOI22X1TS U2498 ( .A0(n1337), .A1(n1911), .B0(n2359), .B1(
        \dataoutbuffer[5][1] ), .Y(n2176) );
  AOI22X1TS U2499 ( .A0(n2361), .A1(n1905), .B0(n2360), .B1(n1903), .Y(n2175)
         );
  AOI22X1TS U2500 ( .A0(n2363), .A1(n1902), .B0(n2362), .B1(n1904), .Y(n2174)
         );
  AOI22X1TS U2501 ( .A0(n1337), .A1(n1926), .B0(n2359), .B1(
        \dataoutbuffer[5][2] ), .Y(n2179) );
  AOI22X1TS U2502 ( .A0(n2361), .A1(n1920), .B0(n2360), .B1(n1917), .Y(n2178)
         );
  AOI22X1TS U2503 ( .A0(n2363), .A1(n1916), .B0(n2362), .B1(n1919), .Y(n2177)
         );
  AOI22X1TS U2504 ( .A0(n1337), .A1(n1940), .B0(n2359), .B1(
        \dataoutbuffer[5][3] ), .Y(n2182) );
  AOI22X1TS U2505 ( .A0(n2361), .A1(n1934), .B0(n2360), .B1(n1932), .Y(n2181)
         );
  AOI22X1TS U2506 ( .A0(n2363), .A1(n1931), .B0(n2362), .B1(n1933), .Y(n2180)
         );
  AOI22X1TS U2507 ( .A0(n1337), .A1(n1954), .B0(n2359), .B1(
        \dataoutbuffer[5][4] ), .Y(n2185) );
  AOI22X1TS U2508 ( .A0(n2361), .A1(n1948), .B0(n2360), .B1(n1946), .Y(n2184)
         );
  AOI22X1TS U2509 ( .A0(n2363), .A1(n1945), .B0(n2362), .B1(n1947), .Y(n2183)
         );
  AOI22X1TS U2510 ( .A0(n1337), .A1(n1979), .B0(n2359), .B1(
        \dataoutbuffer[5][5] ), .Y(n2188) );
  AOI22X1TS U2511 ( .A0(n2361), .A1(n1963), .B0(n2360), .B1(n1960), .Y(n2187)
         );
  AOI22X1TS U2512 ( .A0(n2363), .A1(n1959), .B0(n2362), .B1(n1962), .Y(n2186)
         );
  AOI22X1TS U2513 ( .A0(n2342), .A1(n1897), .B0(n2341), .B1(
        \dataoutbuffer[6][0] ), .Y(n2191) );
  AOI22X1TS U2514 ( .A0(n2344), .A1(n1889), .B0(n2343), .B1(n1887), .Y(n2190)
         );
  AOI22X1TS U2515 ( .A0(n2346), .A1(n1886), .B0(n2345), .B1(n1888), .Y(n2189)
         );
  AOI22X1TS U2516 ( .A0(n2342), .A1(n1911), .B0(n2341), .B1(
        \dataoutbuffer[6][1] ), .Y(n2194) );
  AOI22X1TS U2517 ( .A0(n2344), .A1(n1905), .B0(n2343), .B1(n1903), .Y(n2193)
         );
  AOI22X1TS U2518 ( .A0(n2346), .A1(n1902), .B0(n2345), .B1(n1904), .Y(n2192)
         );
  AOI22X1TS U2519 ( .A0(n2342), .A1(n1926), .B0(n2341), .B1(
        \dataoutbuffer[6][2] ), .Y(n2197) );
  AOI22X1TS U2520 ( .A0(n2344), .A1(n1920), .B0(n2343), .B1(n1917), .Y(n2196)
         );
  AOI22X1TS U2521 ( .A0(n2346), .A1(n1916), .B0(n2345), .B1(n1919), .Y(n2195)
         );
  AOI22X1TS U2522 ( .A0(n2342), .A1(n1940), .B0(n2341), .B1(
        \dataoutbuffer[6][3] ), .Y(n2200) );
  AOI22X1TS U2523 ( .A0(n2344), .A1(n1934), .B0(n2343), .B1(n1932), .Y(n2199)
         );
  AOI22X1TS U2524 ( .A0(n2346), .A1(n1931), .B0(n2345), .B1(n1933), .Y(n2198)
         );
  AOI22X1TS U2525 ( .A0(n2342), .A1(n1954), .B0(n2341), .B1(
        \dataoutbuffer[6][4] ), .Y(n2203) );
  AOI22X1TS U2526 ( .A0(n2344), .A1(n1948), .B0(n2343), .B1(n1946), .Y(n2202)
         );
  AOI22X1TS U2527 ( .A0(n2346), .A1(n1945), .B0(n2345), .B1(n1947), .Y(n2201)
         );
  AOI22X1TS U2528 ( .A0(n2342), .A1(n1979), .B0(n2341), .B1(
        \dataoutbuffer[6][5] ), .Y(n2206) );
  AOI22X1TS U2529 ( .A0(n2344), .A1(n1963), .B0(n2343), .B1(n1960), .Y(n2205)
         );
  AOI22X1TS U2530 ( .A0(n2346), .A1(n1959), .B0(n2345), .B1(n1962), .Y(n2204)
         );
  AOI22X1TS U2531 ( .A0(n2324), .A1(n1897), .B0(n2323), .B1(
        \dataoutbuffer[7][0] ), .Y(n2209) );
  AOI22X1TS U2532 ( .A0(n2326), .A1(n1889), .B0(n2325), .B1(n1887), .Y(n2208)
         );
  AOI22X1TS U2533 ( .A0(n2328), .A1(n1888), .B0(n2327), .B1(n1886), .Y(n2207)
         );
  AOI22X1TS U2534 ( .A0(n2324), .A1(n1911), .B0(n2323), .B1(
        \dataoutbuffer[7][1] ), .Y(n2212) );
  AOI22X1TS U2535 ( .A0(n2326), .A1(n1905), .B0(n2325), .B1(n1903), .Y(n2211)
         );
  AOI22X1TS U2536 ( .A0(n2328), .A1(n1904), .B0(n2327), .B1(n1902), .Y(n2210)
         );
  AOI22X1TS U2537 ( .A0(n2324), .A1(n1926), .B0(n2323), .B1(
        \dataoutbuffer[7][2] ), .Y(n2215) );
  AOI22X1TS U2538 ( .A0(n2326), .A1(n1920), .B0(n2325), .B1(n1917), .Y(n2214)
         );
  AOI22X1TS U2539 ( .A0(n2328), .A1(n1919), .B0(n2327), .B1(n1916), .Y(n2213)
         );
  AOI22X1TS U2540 ( .A0(n2324), .A1(n1940), .B0(n2323), .B1(
        \dataoutbuffer[7][3] ), .Y(n2218) );
  AOI22X1TS U2541 ( .A0(n2326), .A1(n1934), .B0(n2325), .B1(n1932), .Y(n2217)
         );
  AOI22X1TS U2542 ( .A0(n2328), .A1(n1933), .B0(n2327), .B1(n1931), .Y(n2216)
         );
  AOI22X1TS U2543 ( .A0(n2324), .A1(n1954), .B0(n2323), .B1(
        \dataoutbuffer[7][4] ), .Y(n2221) );
  AOI22X1TS U2544 ( .A0(n2326), .A1(n1948), .B0(n2325), .B1(n1946), .Y(n2220)
         );
  AOI22X1TS U2545 ( .A0(n2328), .A1(n1947), .B0(n2327), .B1(n1945), .Y(n2219)
         );
  AOI22X1TS U2546 ( .A0(n2324), .A1(n1979), .B0(n2323), .B1(
        \dataoutbuffer[7][5] ), .Y(n2224) );
  AOI22X1TS U2547 ( .A0(n2326), .A1(n1963), .B0(n2325), .B1(n1960), .Y(n2223)
         );
  AOI22X1TS U2548 ( .A0(n2328), .A1(n1962), .B0(n2327), .B1(n1959), .Y(n2222)
         );
  INVX2TS U2549 ( .A(n1683), .Y(n2306) );
  AOI22X1TS U2550 ( .A0(n2226), .A1(n1678), .B0(n1680), .B1(n2225), .Y(n2228)
         );
  AOI22X1TS U2551 ( .A0(n2229), .A1(n2306), .B0(n2228), .B1(n2227), .Y(n2231)
         );
  AOI22X1TS U2552 ( .A0(n2232), .A1(n1679), .B0(n2231), .B1(n2230), .Y(n2235)
         );
  AOI32X1TS U2553 ( .A0(n2235), .A1(n2234), .A2(n2233), .B0(n2323), .B1(n2464), 
        .Y(n1217) );
  AOI22X1TS U2554 ( .A0(n2237), .A1(n1678), .B0(n1680), .B1(n2236), .Y(n2239)
         );
  AOI22X1TS U2555 ( .A0(n2240), .A1(n2306), .B0(n2239), .B1(n2238), .Y(n2242)
         );
  AOI22X1TS U2556 ( .A0(n2243), .A1(n1679), .B0(n2242), .B1(n2241), .Y(n2246)
         );
  AOI32X1TS U2557 ( .A0(n2246), .A1(n2245), .A2(n2244), .B0(n2341), .B1(n2465), 
        .Y(n1216) );
  AOI22X1TS U2558 ( .A0(n2248), .A1(n1678), .B0(n1680), .B1(n2247), .Y(n2250)
         );
  AOI22X1TS U2559 ( .A0(n2251), .A1(n2306), .B0(n2250), .B1(n2249), .Y(n2253)
         );
  AOI22X1TS U2560 ( .A0(n2254), .A1(n1679), .B0(n2253), .B1(n2252), .Y(n2257)
         );
  AOI32X1TS U2561 ( .A0(n2257), .A1(n2256), .A2(n2255), .B0(n2359), .B1(n2466), 
        .Y(n1215) );
  AOI22X1TS U2562 ( .A0(n2259), .A1(n1678), .B0(n1680), .B1(n2258), .Y(n2261)
         );
  AOI22X1TS U2563 ( .A0(n2262), .A1(n2306), .B0(n2261), .B1(n2260), .Y(n2264)
         );
  AOI22X1TS U2564 ( .A0(n2265), .A1(n1679), .B0(n2264), .B1(n2263), .Y(n2268)
         );
  AOI32X1TS U2565 ( .A0(n2268), .A1(n2267), .A2(n2266), .B0(n2376), .B1(n2467), 
        .Y(n1214) );
  AOI22X1TS U2566 ( .A0(n2270), .A1(n1678), .B0(n1680), .B1(n2269), .Y(n2272)
         );
  AOI22X1TS U2567 ( .A0(n2273), .A1(n2306), .B0(n2272), .B1(n2271), .Y(n2275)
         );
  AOI22X1TS U2568 ( .A0(n2276), .A1(n1679), .B0(n2275), .B1(n2274), .Y(n2279)
         );
  AOI32X1TS U2569 ( .A0(n2279), .A1(n2278), .A2(n2277), .B0(n2394), .B1(n2468), 
        .Y(n1213) );
  AOI22X1TS U2570 ( .A0(n2281), .A1(n1678), .B0(n1680), .B1(n2280), .Y(n2283)
         );
  AOI22X1TS U2571 ( .A0(n2284), .A1(n2306), .B0(n2283), .B1(n2282), .Y(n2286)
         );
  AOI22X1TS U2572 ( .A0(n2287), .A1(n1679), .B0(n2286), .B1(n2285), .Y(n2290)
         );
  AOI32X1TS U2573 ( .A0(n2290), .A1(n2289), .A2(n2288), .B0(n2411), .B1(n2469), 
        .Y(n1212) );
  AOI22X1TS U2574 ( .A0(n2292), .A1(n1678), .B0(n1680), .B1(n2291), .Y(n2294)
         );
  AOI22X1TS U2575 ( .A0(n2295), .A1(n2306), .B0(n2294), .B1(n2293), .Y(n2297)
         );
  AOI22X1TS U2576 ( .A0(n2298), .A1(n1679), .B0(n2297), .B1(n2296), .Y(n2301)
         );
  AOI32X1TS U2577 ( .A0(n2301), .A1(n2300), .A2(n2299), .B0(n2429), .B1(n2470), 
        .Y(n1211) );
  AOI22X1TS U2578 ( .A0(n2303), .A1(n1678), .B0(n1680), .B1(n2302), .Y(n2305)
         );
  AOI22X1TS U2579 ( .A0(n2307), .A1(n2306), .B0(n2305), .B1(n2304), .Y(n2309)
         );
  AOI22X1TS U2580 ( .A0(n2310), .A1(n1679), .B0(n2309), .B1(n2308), .Y(n2313)
         );
  AOI32X1TS U2581 ( .A0(n2313), .A1(n2312), .A2(n2311), .B0(n2447), .B1(n2471), 
        .Y(n1210) );
  AOI22X1TS U2582 ( .A0(n1720), .A1(n2324), .B0(n2323), .B1(
        \destinationAddressbuffer[7][0] ), .Y(n2316) );
  AOI22X1TS U2583 ( .A0(n2326), .A1(n1767), .B0(n2325), .B1(n1765), .Y(n2315)
         );
  AOI22X1TS U2584 ( .A0(n2328), .A1(n1766), .B0(n2327), .B1(n1764), .Y(n2314)
         );
  AOI22X1TS U2585 ( .A0(n2324), .A1(n1734), .B0(n2323), .B1(
        \destinationAddressbuffer[7][1] ), .Y(n2319) );
  AOI22X1TS U2586 ( .A0(n2326), .A1(n1780), .B0(n2325), .B1(n1778), .Y(n2318)
         );
  AOI22X1TS U2587 ( .A0(n2328), .A1(n1779), .B0(n2327), .B1(n1777), .Y(n2317)
         );
  AOI22X1TS U2588 ( .A0(n2324), .A1(n1747), .B0(n2323), .B1(
        \destinationAddressbuffer[7][2] ), .Y(n2322) );
  AOI22X1TS U2589 ( .A0(n2326), .A1(n1794), .B0(n2325), .B1(n1792), .Y(n2321)
         );
  AOI22X1TS U2590 ( .A0(n2328), .A1(n1793), .B0(n2327), .B1(n1791), .Y(n2320)
         );
  AOI22X1TS U2591 ( .A0(n2324), .A1(n1760), .B0(n2323), .B1(
        \destinationAddressbuffer[7][3] ), .Y(n2331) );
  AOI22X1TS U2592 ( .A0(n2326), .A1(n1807), .B0(n2325), .B1(n1805), .Y(n2330)
         );
  AOI22X1TS U2593 ( .A0(n2328), .A1(n1806), .B0(n2327), .B1(n1804), .Y(n2329)
         );
  AOI22X1TS U2594 ( .A0(n1720), .A1(n2342), .B0(n2341), .B1(
        \destinationAddressbuffer[6][0] ), .Y(n2334) );
  AOI22X1TS U2595 ( .A0(n2344), .A1(n1767), .B0(n2343), .B1(n1765), .Y(n2333)
         );
  AOI22X1TS U2596 ( .A0(n2346), .A1(n1764), .B0(n2345), .B1(n1766), .Y(n2332)
         );
  AOI22X1TS U2597 ( .A0(n1734), .A1(n2342), .B0(n2341), .B1(
        \destinationAddressbuffer[6][1] ), .Y(n2337) );
  AOI22X1TS U2598 ( .A0(n2344), .A1(n1780), .B0(n2343), .B1(n1778), .Y(n2336)
         );
  AOI22X1TS U2599 ( .A0(n2346), .A1(n1777), .B0(n2345), .B1(n1779), .Y(n2335)
         );
  AOI22X1TS U2600 ( .A0(n1747), .A1(n2342), .B0(n2341), .B1(
        \destinationAddressbuffer[6][2] ), .Y(n2340) );
  AOI22X1TS U2601 ( .A0(n2344), .A1(n1794), .B0(n2343), .B1(n1792), .Y(n2339)
         );
  AOI22X1TS U2602 ( .A0(n2346), .A1(n1791), .B0(n2345), .B1(n1793), .Y(n2338)
         );
  AOI22X1TS U2603 ( .A0(n1760), .A1(n2342), .B0(n2341), .B1(
        \destinationAddressbuffer[6][3] ), .Y(n2349) );
  AOI22X1TS U2604 ( .A0(n2344), .A1(n1807), .B0(n2343), .B1(n1805), .Y(n2348)
         );
  AOI22X1TS U2605 ( .A0(n2346), .A1(n1804), .B0(n2345), .B1(n1806), .Y(n2347)
         );
  AOI22X1TS U2606 ( .A0(n1720), .A1(n1337), .B0(n2359), .B1(
        \destinationAddressbuffer[5][0] ), .Y(n2352) );
  AOI22X1TS U2607 ( .A0(n2361), .A1(n1767), .B0(n2360), .B1(n1765), .Y(n2351)
         );
  AOI22X1TS U2608 ( .A0(n2363), .A1(n1764), .B0(n2362), .B1(n1766), .Y(n2350)
         );
  AOI22X1TS U2609 ( .A0(n1734), .A1(n1337), .B0(n2359), .B1(
        \destinationAddressbuffer[5][1] ), .Y(n2355) );
  AOI22X1TS U2610 ( .A0(n2361), .A1(n1780), .B0(n2360), .B1(n1778), .Y(n2354)
         );
  AOI22X1TS U2611 ( .A0(n2363), .A1(n1777), .B0(n2362), .B1(n1779), .Y(n2353)
         );
  AOI22X1TS U2612 ( .A0(n1747), .A1(n1337), .B0(n2359), .B1(
        \destinationAddressbuffer[5][2] ), .Y(n2358) );
  AOI22X1TS U2613 ( .A0(n2361), .A1(n1794), .B0(n2360), .B1(n1792), .Y(n2357)
         );
  AOI22X1TS U2614 ( .A0(n2363), .A1(n1791), .B0(n2362), .B1(n1793), .Y(n2356)
         );
  AOI22X1TS U2615 ( .A0(n1760), .A1(n1337), .B0(n2359), .B1(
        \destinationAddressbuffer[5][3] ), .Y(n2366) );
  AOI22X1TS U2616 ( .A0(n2361), .A1(n1807), .B0(n2360), .B1(n1805), .Y(n2365)
         );
  AOI22X1TS U2617 ( .A0(n2363), .A1(n1804), .B0(n2362), .B1(n1806), .Y(n2364)
         );
  AOI22X1TS U2618 ( .A0(n1720), .A1(n2377), .B0(n2376), .B1(
        \destinationAddressbuffer[4][0] ), .Y(n2369) );
  AOI22X1TS U2619 ( .A0(n2379), .A1(n1767), .B0(n2378), .B1(n1765), .Y(n2368)
         );
  AOI22X1TS U2620 ( .A0(n2381), .A1(n1766), .B0(n2380), .B1(n1764), .Y(n2367)
         );
  AOI22X1TS U2621 ( .A0(n1734), .A1(n2377), .B0(n2376), .B1(
        \destinationAddressbuffer[4][1] ), .Y(n2372) );
  AOI22X1TS U2622 ( .A0(n2379), .A1(n1780), .B0(n2378), .B1(n1778), .Y(n2371)
         );
  AOI22X1TS U2623 ( .A0(n2381), .A1(n1779), .B0(n2380), .B1(n1777), .Y(n2370)
         );
  AOI22X1TS U2624 ( .A0(n1747), .A1(n2377), .B0(n2376), .B1(
        \destinationAddressbuffer[4][2] ), .Y(n2375) );
  AOI22X1TS U2625 ( .A0(n2379), .A1(n1794), .B0(n2378), .B1(n1792), .Y(n2374)
         );
  AOI22X1TS U2626 ( .A0(n2381), .A1(n1793), .B0(n2380), .B1(n1791), .Y(n2373)
         );
  AOI22X1TS U2627 ( .A0(n1760), .A1(n2377), .B0(n2376), .B1(
        \destinationAddressbuffer[4][3] ), .Y(n2384) );
  AOI22X1TS U2628 ( .A0(n2379), .A1(n1807), .B0(n2378), .B1(n1805), .Y(n2383)
         );
  AOI22X1TS U2629 ( .A0(n2381), .A1(n1806), .B0(n2380), .B1(n1804), .Y(n2382)
         );
  AOI22X1TS U2630 ( .A0(n1720), .A1(n2395), .B0(n2394), .B1(
        \destinationAddressbuffer[3][0] ), .Y(n2387) );
  AOI22X1TS U2631 ( .A0(n2396), .A1(n1767), .B0(n1510), .B1(n1765), .Y(n2386)
         );
  AOI22X1TS U2632 ( .A0(n2398), .A1(n1764), .B0(n2397), .B1(n1766), .Y(n2385)
         );
  AOI22X1TS U2633 ( .A0(n1734), .A1(n2395), .B0(n2394), .B1(
        \destinationAddressbuffer[3][1] ), .Y(n2390) );
  AOI22X1TS U2634 ( .A0(n2396), .A1(n1780), .B0(n1510), .B1(n1778), .Y(n2389)
         );
  AOI22X1TS U2635 ( .A0(n2398), .A1(n1777), .B0(n2397), .B1(n1779), .Y(n2388)
         );
  AOI22X1TS U2636 ( .A0(n1747), .A1(n2395), .B0(n2394), .B1(
        \destinationAddressbuffer[3][2] ), .Y(n2393) );
  AOI22X1TS U2637 ( .A0(n2396), .A1(n1794), .B0(n1510), .B1(n1792), .Y(n2392)
         );
  AOI22X1TS U2638 ( .A0(n2398), .A1(n1791), .B0(n2397), .B1(n1793), .Y(n2391)
         );
  AOI22X1TS U2639 ( .A0(n1760), .A1(n2395), .B0(n2394), .B1(
        \destinationAddressbuffer[3][3] ), .Y(n2401) );
  AOI22X1TS U2640 ( .A0(n2396), .A1(n1807), .B0(n1510), .B1(n1805), .Y(n2400)
         );
  AOI22X1TS U2641 ( .A0(n2398), .A1(n1804), .B0(n2397), .B1(n1806), .Y(n2399)
         );
  AOI22X1TS U2642 ( .A0(n1720), .A1(n2412), .B0(n2411), .B1(
        \destinationAddressbuffer[2][0] ), .Y(n2404) );
  AOI22X1TS U2643 ( .A0(n2414), .A1(n1767), .B0(n2413), .B1(n1765), .Y(n2403)
         );
  AOI22X1TS U2644 ( .A0(n2416), .A1(n1764), .B0(n2415), .B1(n1766), .Y(n2402)
         );
  AOI22X1TS U2645 ( .A0(n1734), .A1(n2412), .B0(n2411), .B1(
        \destinationAddressbuffer[2][1] ), .Y(n2407) );
  AOI22X1TS U2646 ( .A0(n2414), .A1(n1780), .B0(n2413), .B1(n1778), .Y(n2406)
         );
  AOI22X1TS U2647 ( .A0(n2416), .A1(n1777), .B0(n2415), .B1(n1779), .Y(n2405)
         );
  AOI22X1TS U2648 ( .A0(n1747), .A1(n2412), .B0(n2411), .B1(
        \destinationAddressbuffer[2][2] ), .Y(n2410) );
  AOI22X1TS U2649 ( .A0(n2414), .A1(n1794), .B0(n2413), .B1(n1792), .Y(n2409)
         );
  AOI22X1TS U2650 ( .A0(n2416), .A1(n1791), .B0(n2415), .B1(n1793), .Y(n2408)
         );
  AOI22X1TS U2651 ( .A0(n1760), .A1(n2412), .B0(n2411), .B1(
        \destinationAddressbuffer[2][3] ), .Y(n2419) );
  AOI22X1TS U2652 ( .A0(n2414), .A1(n1807), .B0(n2413), .B1(n1805), .Y(n2418)
         );
  AOI22X1TS U2653 ( .A0(n2416), .A1(n1804), .B0(n2415), .B1(n1806), .Y(n2417)
         );
  AOI22X1TS U2654 ( .A0(n1720), .A1(n2430), .B0(n2429), .B1(
        \destinationAddressbuffer[1][0] ), .Y(n2422) );
  AOI22X1TS U2655 ( .A0(n2432), .A1(n1767), .B0(n2431), .B1(n1765), .Y(n2421)
         );
  AOI22X1TS U2656 ( .A0(n2434), .A1(n1764), .B0(n2433), .B1(n1766), .Y(n2420)
         );
  AOI22X1TS U2657 ( .A0(n1734), .A1(n2430), .B0(n2429), .B1(
        \destinationAddressbuffer[1][1] ), .Y(n2425) );
  AOI22X1TS U2658 ( .A0(n2432), .A1(n1780), .B0(n2431), .B1(n1778), .Y(n2424)
         );
  AOI22X1TS U2659 ( .A0(n2434), .A1(n1777), .B0(n2433), .B1(n1779), .Y(n2423)
         );
  AOI22X1TS U2660 ( .A0(n1747), .A1(n2430), .B0(n2429), .B1(
        \destinationAddressbuffer[1][2] ), .Y(n2428) );
  AOI22X1TS U2661 ( .A0(n2432), .A1(n1794), .B0(n2431), .B1(n1792), .Y(n2427)
         );
  AOI22X1TS U2662 ( .A0(n2434), .A1(n1791), .B0(n2433), .B1(n1793), .Y(n2426)
         );
  AOI22X1TS U2663 ( .A0(n1760), .A1(n2430), .B0(n2429), .B1(
        \destinationAddressbuffer[1][3] ), .Y(n2437) );
  AOI22X1TS U2664 ( .A0(n2432), .A1(n1807), .B0(n2431), .B1(n1805), .Y(n2436)
         );
  AOI22X1TS U2665 ( .A0(n2434), .A1(n1804), .B0(n2433), .B1(n1806), .Y(n2435)
         );
  AOI22X1TS U2666 ( .A0(n1720), .A1(n2448), .B0(n2447), .B1(
        \destinationAddressbuffer[0][0] ), .Y(n2440) );
  AOI22X1TS U2667 ( .A0(n2450), .A1(n1767), .B0(n2449), .B1(n1765), .Y(n2439)
         );
  AOI22X1TS U2668 ( .A0(n2452), .A1(n1766), .B0(n2451), .B1(n1764), .Y(n2438)
         );
  AOI22X1TS U2669 ( .A0(n1734), .A1(n2448), .B0(n2447), .B1(
        \destinationAddressbuffer[0][1] ), .Y(n2443) );
  AOI22X1TS U2670 ( .A0(n2450), .A1(n1780), .B0(n2449), .B1(n1778), .Y(n2442)
         );
  AOI22X1TS U2671 ( .A0(n2452), .A1(n1779), .B0(n2451), .B1(n1777), .Y(n2441)
         );
  AOI22X1TS U2672 ( .A0(n1747), .A1(n2448), .B0(n2447), .B1(
        \destinationAddressbuffer[0][2] ), .Y(n2446) );
  AOI22X1TS U2673 ( .A0(n2450), .A1(n1794), .B0(n2449), .B1(n1792), .Y(n2445)
         );
  AOI22X1TS U2674 ( .A0(n2452), .A1(n1793), .B0(n2451), .B1(n1791), .Y(n2444)
         );
  AOI22X1TS U2675 ( .A0(n1760), .A1(n2448), .B0(n2447), .B1(
        \destinationAddressbuffer[0][3] ), .Y(n2455) );
  AOI22X1TS U2676 ( .A0(n2450), .A1(n1807), .B0(n2449), .B1(n1805), .Y(n2454)
         );
  AOI22X1TS U2677 ( .A0(n2452), .A1(n1806), .B0(n2451), .B1(n1804), .Y(n2453)
         );
endmodule

