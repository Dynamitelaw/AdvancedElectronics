##
## LEF for PtnCells ;
## created by Encounter v14.23-s044_1 on Thu May 16 16:17:29 2019
##

VERSION 5.5 ;

NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO router
  CLASS BLOCK ;
  SIZE 666.0000 BY 612.0000 ;
  FOREIGN router 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 10.9000 0.6000 11.1000 ;
    END
  END clk
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MQ ;
        RECT 359.6000 0.0000 360.0000 1.2000 ;
    END
  END reset
  PIN localRouterAddress[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 26.9000 0.6000 27.1000 ;
    END
  END localRouterAddress[5]
  PIN localRouterAddress[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 24.9000 0.6000 25.1000 ;
    END
  END localRouterAddress[4]
  PIN localRouterAddress[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 22.9000 0.6000 23.1000 ;
    END
  END localRouterAddress[3]
  PIN localRouterAddress[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 20.9000 0.6000 21.1000 ;
    END
  END localRouterAddress[2]
  PIN localRouterAddress[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 18.9000 0.6000 19.1000 ;
    END
  END localRouterAddress[1]
  PIN localRouterAddress[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 16.9000 0.6000 17.1000 ;
    END
  END localRouterAddress[0]
  PIN destinationAddressIn_NORTH[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.4000 611.4000 31.6000 612.0000 ;
    END
  END destinationAddressIn_NORTH[13]
  PIN destinationAddressIn_NORTH[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.9000 611.4000 30.1000 612.0000 ;
    END
  END destinationAddressIn_NORTH[12]
  PIN destinationAddressIn_NORTH[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 28.4000 611.4000 28.6000 612.0000 ;
    END
  END destinationAddressIn_NORTH[11]
  PIN destinationAddressIn_NORTH[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 26.9000 611.4000 27.1000 612.0000 ;
    END
  END destinationAddressIn_NORTH[10]
  PIN destinationAddressIn_NORTH[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 25.4000 611.4000 25.6000 612.0000 ;
    END
  END destinationAddressIn_NORTH[9]
  PIN destinationAddressIn_NORTH[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 23.9000 611.4000 24.1000 612.0000 ;
    END
  END destinationAddressIn_NORTH[8]
  PIN destinationAddressIn_NORTH[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.4000 611.4000 22.6000 612.0000 ;
    END
  END destinationAddressIn_NORTH[7]
  PIN destinationAddressIn_NORTH[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20.9000 611.4000 21.1000 612.0000 ;
    END
  END destinationAddressIn_NORTH[6]
  PIN destinationAddressIn_NORTH[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19.4000 611.4000 19.6000 612.0000 ;
    END
  END destinationAddressIn_NORTH[5]
  PIN destinationAddressIn_NORTH[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17.9000 611.4000 18.1000 612.0000 ;
    END
  END destinationAddressIn_NORTH[4]
  PIN destinationAddressIn_NORTH[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16.4000 611.4000 16.6000 612.0000 ;
    END
  END destinationAddressIn_NORTH[3]
  PIN destinationAddressIn_NORTH[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14.9000 611.4000 15.1000 612.0000 ;
    END
  END destinationAddressIn_NORTH[2]
  PIN destinationAddressIn_NORTH[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13.4000 611.4000 13.6000 612.0000 ;
    END
  END destinationAddressIn_NORTH[1]
  PIN destinationAddressIn_NORTH[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11.9000 611.4000 12.1000 612.0000 ;
    END
  END destinationAddressIn_NORTH[0]
  PIN requesterAddressIn_NORTH[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 40.4000 611.4000 40.6000 612.0000 ;
    END
  END requesterAddressIn_NORTH[5]
  PIN requesterAddressIn_NORTH[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.9000 611.4000 39.1000 612.0000 ;
    END
  END requesterAddressIn_NORTH[4]
  PIN requesterAddressIn_NORTH[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 37.4000 611.4000 37.6000 612.0000 ;
    END
  END requesterAddressIn_NORTH[3]
  PIN requesterAddressIn_NORTH[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 35.9000 611.4000 36.1000 612.0000 ;
    END
  END requesterAddressIn_NORTH[2]
  PIN requesterAddressIn_NORTH[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.4000 611.4000 34.6000 612.0000 ;
    END
  END requesterAddressIn_NORTH[1]
  PIN requesterAddressIn_NORTH[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 32.9000 611.4000 33.1000 612.0000 ;
    END
  END requesterAddressIn_NORTH[0]
  PIN readIn_NORTH
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 41.9000 611.4000 42.1000 612.0000 ;
    END
  END readIn_NORTH
  PIN writeIn_NORTH
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 43.4000 611.4000 43.6000 612.0000 ;
    END
  END writeIn_NORTH
  PIN dataIn_NORTH[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 179.4000 611.4000 179.6000 612.0000 ;
    END
  END dataIn_NORTH[31]
  PIN dataIn_NORTH[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 177.9000 611.4000 178.1000 612.0000 ;
    END
  END dataIn_NORTH[30]
  PIN dataIn_NORTH[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 176.4000 611.4000 176.6000 612.0000 ;
    END
  END dataIn_NORTH[29]
  PIN dataIn_NORTH[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 174.9000 611.4000 175.1000 612.0000 ;
    END
  END dataIn_NORTH[28]
  PIN dataIn_NORTH[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 173.4000 611.4000 173.6000 612.0000 ;
    END
  END dataIn_NORTH[27]
  PIN dataIn_NORTH[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 171.9000 611.4000 172.1000 612.0000 ;
    END
  END dataIn_NORTH[26]
  PIN dataIn_NORTH[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 170.4000 611.4000 170.6000 612.0000 ;
    END
  END dataIn_NORTH[25]
  PIN dataIn_NORTH[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 168.9000 611.4000 169.1000 612.0000 ;
    END
  END dataIn_NORTH[24]
  PIN dataIn_NORTH[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 167.4000 611.4000 167.6000 612.0000 ;
    END
  END dataIn_NORTH[23]
  PIN dataIn_NORTH[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 165.9000 611.4000 166.1000 612.0000 ;
    END
  END dataIn_NORTH[22]
  PIN dataIn_NORTH[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 164.4000 611.4000 164.6000 612.0000 ;
    END
  END dataIn_NORTH[21]
  PIN dataIn_NORTH[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 162.9000 611.4000 163.1000 612.0000 ;
    END
  END dataIn_NORTH[20]
  PIN dataIn_NORTH[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 161.4000 611.4000 161.6000 612.0000 ;
    END
  END dataIn_NORTH[19]
  PIN dataIn_NORTH[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 159.9000 611.4000 160.1000 612.0000 ;
    END
  END dataIn_NORTH[18]
  PIN dataIn_NORTH[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 158.4000 611.4000 158.6000 612.0000 ;
    END
  END dataIn_NORTH[17]
  PIN dataIn_NORTH[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 156.9000 611.4000 157.1000 612.0000 ;
    END
  END dataIn_NORTH[16]
  PIN dataIn_NORTH[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 155.4000 611.4000 155.6000 612.0000 ;
    END
  END dataIn_NORTH[15]
  PIN dataIn_NORTH[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 153.9000 611.4000 154.1000 612.0000 ;
    END
  END dataIn_NORTH[14]
  PIN dataIn_NORTH[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 152.4000 611.4000 152.6000 612.0000 ;
    END
  END dataIn_NORTH[13]
  PIN dataIn_NORTH[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 150.9000 611.4000 151.1000 612.0000 ;
    END
  END dataIn_NORTH[12]
  PIN dataIn_NORTH[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 149.4000 611.4000 149.6000 612.0000 ;
    END
  END dataIn_NORTH[11]
  PIN dataIn_NORTH[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 147.9000 611.4000 148.1000 612.0000 ;
    END
  END dataIn_NORTH[10]
  PIN dataIn_NORTH[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 146.4000 611.4000 146.6000 612.0000 ;
    END
  END dataIn_NORTH[9]
  PIN dataIn_NORTH[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 144.9000 611.4000 145.1000 612.0000 ;
    END
  END dataIn_NORTH[8]
  PIN dataIn_NORTH[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 143.4000 611.4000 143.6000 612.0000 ;
    END
  END dataIn_NORTH[7]
  PIN dataIn_NORTH[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 141.9000 611.4000 142.1000 612.0000 ;
    END
  END dataIn_NORTH[6]
  PIN dataIn_NORTH[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 140.4000 611.4000 140.6000 612.0000 ;
    END
  END dataIn_NORTH[5]
  PIN dataIn_NORTH[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 138.9000 611.4000 139.1000 612.0000 ;
    END
  END dataIn_NORTH[4]
  PIN dataIn_NORTH[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 137.4000 611.4000 137.6000 612.0000 ;
    END
  END dataIn_NORTH[3]
  PIN dataIn_NORTH[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 135.9000 611.4000 136.1000 612.0000 ;
    END
  END dataIn_NORTH[2]
  PIN dataIn_NORTH[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 134.4000 611.4000 134.6000 612.0000 ;
    END
  END dataIn_NORTH[1]
  PIN dataIn_NORTH[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 132.9000 611.4000 133.1000 612.0000 ;
    END
  END dataIn_NORTH[0]
  PIN destinationAddressOut_NORTH[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 119.4000 611.4000 119.6000 612.0000 ;
    END
  END destinationAddressOut_NORTH[13]
  PIN destinationAddressOut_NORTH[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 117.9000 611.4000 118.1000 612.0000 ;
    END
  END destinationAddressOut_NORTH[12]
  PIN destinationAddressOut_NORTH[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 116.4000 611.4000 116.6000 612.0000 ;
    END
  END destinationAddressOut_NORTH[11]
  PIN destinationAddressOut_NORTH[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 114.9000 611.4000 115.1000 612.0000 ;
    END
  END destinationAddressOut_NORTH[10]
  PIN destinationAddressOut_NORTH[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 113.4000 611.4000 113.6000 612.0000 ;
    END
  END destinationAddressOut_NORTH[9]
  PIN destinationAddressOut_NORTH[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 111.9000 611.4000 112.1000 612.0000 ;
    END
  END destinationAddressOut_NORTH[8]
  PIN destinationAddressOut_NORTH[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 110.4000 611.4000 110.6000 612.0000 ;
    END
  END destinationAddressOut_NORTH[7]
  PIN destinationAddressOut_NORTH[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 108.9000 611.4000 109.1000 612.0000 ;
    END
  END destinationAddressOut_NORTH[6]
  PIN destinationAddressOut_NORTH[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 107.4000 611.4000 107.6000 612.0000 ;
    END
  END destinationAddressOut_NORTH[5]
  PIN destinationAddressOut_NORTH[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 105.9000 611.4000 106.1000 612.0000 ;
    END
  END destinationAddressOut_NORTH[4]
  PIN destinationAddressOut_NORTH[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 104.4000 611.4000 104.6000 612.0000 ;
    END
  END destinationAddressOut_NORTH[3]
  PIN destinationAddressOut_NORTH[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 102.9000 611.4000 103.1000 612.0000 ;
    END
  END destinationAddressOut_NORTH[2]
  PIN destinationAddressOut_NORTH[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 101.4000 611.4000 101.6000 612.0000 ;
    END
  END destinationAddressOut_NORTH[1]
  PIN destinationAddressOut_NORTH[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 99.9000 611.4000 100.1000 612.0000 ;
    END
  END destinationAddressOut_NORTH[0]
  PIN requesterAddressOut_NORTH[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 128.4000 611.4000 128.6000 612.0000 ;
    END
  END requesterAddressOut_NORTH[5]
  PIN requesterAddressOut_NORTH[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 126.9000 611.4000 127.1000 612.0000 ;
    END
  END requesterAddressOut_NORTH[4]
  PIN requesterAddressOut_NORTH[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 125.4000 611.4000 125.6000 612.0000 ;
    END
  END requesterAddressOut_NORTH[3]
  PIN requesterAddressOut_NORTH[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 123.9000 611.4000 124.1000 612.0000 ;
    END
  END requesterAddressOut_NORTH[2]
  PIN requesterAddressOut_NORTH[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 122.4000 611.4000 122.6000 612.0000 ;
    END
  END requesterAddressOut_NORTH[1]
  PIN requesterAddressOut_NORTH[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 120.9000 611.4000 121.1000 612.0000 ;
    END
  END requesterAddressOut_NORTH[0]
  PIN readOut_NORTH
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 129.9000 611.4000 130.1000 612.0000 ;
    END
  END readOut_NORTH
  PIN writeOut_NORTH
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 131.4000 611.4000 131.6000 612.0000 ;
    END
  END writeOut_NORTH
  PIN dataOut_NORTH[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 91.4000 611.4000 91.6000 612.0000 ;
    END
  END dataOut_NORTH[31]
  PIN dataOut_NORTH[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 89.9000 611.4000 90.1000 612.0000 ;
    END
  END dataOut_NORTH[30]
  PIN dataOut_NORTH[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 88.4000 611.4000 88.6000 612.0000 ;
    END
  END dataOut_NORTH[29]
  PIN dataOut_NORTH[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 86.9000 611.4000 87.1000 612.0000 ;
    END
  END dataOut_NORTH[28]
  PIN dataOut_NORTH[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 85.4000 611.4000 85.6000 612.0000 ;
    END
  END dataOut_NORTH[27]
  PIN dataOut_NORTH[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 83.9000 611.4000 84.1000 612.0000 ;
    END
  END dataOut_NORTH[26]
  PIN dataOut_NORTH[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 82.4000 611.4000 82.6000 612.0000 ;
    END
  END dataOut_NORTH[25]
  PIN dataOut_NORTH[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 80.9000 611.4000 81.1000 612.0000 ;
    END
  END dataOut_NORTH[24]
  PIN dataOut_NORTH[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 79.4000 611.4000 79.6000 612.0000 ;
    END
  END dataOut_NORTH[23]
  PIN dataOut_NORTH[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 77.9000 611.4000 78.1000 612.0000 ;
    END
  END dataOut_NORTH[22]
  PIN dataOut_NORTH[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 76.4000 611.4000 76.6000 612.0000 ;
    END
  END dataOut_NORTH[21]
  PIN dataOut_NORTH[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 74.9000 611.4000 75.1000 612.0000 ;
    END
  END dataOut_NORTH[20]
  PIN dataOut_NORTH[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 73.4000 611.4000 73.6000 612.0000 ;
    END
  END dataOut_NORTH[19]
  PIN dataOut_NORTH[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 71.9000 611.4000 72.1000 612.0000 ;
    END
  END dataOut_NORTH[18]
  PIN dataOut_NORTH[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 70.4000 611.4000 70.6000 612.0000 ;
    END
  END dataOut_NORTH[17]
  PIN dataOut_NORTH[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 68.9000 611.4000 69.1000 612.0000 ;
    END
  END dataOut_NORTH[16]
  PIN dataOut_NORTH[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 67.4000 611.4000 67.6000 612.0000 ;
    END
  END dataOut_NORTH[15]
  PIN dataOut_NORTH[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 65.9000 611.4000 66.1000 612.0000 ;
    END
  END dataOut_NORTH[14]
  PIN dataOut_NORTH[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 64.4000 611.4000 64.6000 612.0000 ;
    END
  END dataOut_NORTH[13]
  PIN dataOut_NORTH[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 62.9000 611.4000 63.1000 612.0000 ;
    END
  END dataOut_NORTH[12]
  PIN dataOut_NORTH[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 61.4000 611.4000 61.6000 612.0000 ;
    END
  END dataOut_NORTH[11]
  PIN dataOut_NORTH[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 59.9000 611.4000 60.1000 612.0000 ;
    END
  END dataOut_NORTH[10]
  PIN dataOut_NORTH[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 58.4000 611.4000 58.6000 612.0000 ;
    END
  END dataOut_NORTH[9]
  PIN dataOut_NORTH[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 56.9000 611.4000 57.1000 612.0000 ;
    END
  END dataOut_NORTH[8]
  PIN dataOut_NORTH[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 55.4000 611.4000 55.6000 612.0000 ;
    END
  END dataOut_NORTH[7]
  PIN dataOut_NORTH[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 53.9000 611.4000 54.1000 612.0000 ;
    END
  END dataOut_NORTH[6]
  PIN dataOut_NORTH[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 52.4000 611.4000 52.6000 612.0000 ;
    END
  END dataOut_NORTH[5]
  PIN dataOut_NORTH[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 50.9000 611.4000 51.1000 612.0000 ;
    END
  END dataOut_NORTH[4]
  PIN dataOut_NORTH[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 49.4000 611.4000 49.6000 612.0000 ;
    END
  END dataOut_NORTH[3]
  PIN dataOut_NORTH[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 47.9000 611.4000 48.1000 612.0000 ;
    END
  END dataOut_NORTH[2]
  PIN dataOut_NORTH[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.4000 611.4000 46.6000 612.0000 ;
    END
  END dataOut_NORTH[1]
  PIN dataOut_NORTH[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44.9000 611.4000 45.1000 612.0000 ;
    END
  END dataOut_NORTH[0]
  PIN destinationAddressIn_SOUTH[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.4000 0.0000 31.6000 0.6000 ;
    END
  END destinationAddressIn_SOUTH[13]
  PIN destinationAddressIn_SOUTH[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.9000 0.0000 30.1000 0.6000 ;
    END
  END destinationAddressIn_SOUTH[12]
  PIN destinationAddressIn_SOUTH[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 28.4000 0.0000 28.6000 0.6000 ;
    END
  END destinationAddressIn_SOUTH[11]
  PIN destinationAddressIn_SOUTH[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 26.9000 0.0000 27.1000 0.6000 ;
    END
  END destinationAddressIn_SOUTH[10]
  PIN destinationAddressIn_SOUTH[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 25.4000 0.0000 25.6000 0.6000 ;
    END
  END destinationAddressIn_SOUTH[9]
  PIN destinationAddressIn_SOUTH[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 23.9000 0.0000 24.1000 0.6000 ;
    END
  END destinationAddressIn_SOUTH[8]
  PIN destinationAddressIn_SOUTH[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.4000 0.0000 22.6000 0.6000 ;
    END
  END destinationAddressIn_SOUTH[7]
  PIN destinationAddressIn_SOUTH[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20.9000 0.0000 21.1000 0.6000 ;
    END
  END destinationAddressIn_SOUTH[6]
  PIN destinationAddressIn_SOUTH[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19.4000 0.0000 19.6000 0.6000 ;
    END
  END destinationAddressIn_SOUTH[5]
  PIN destinationAddressIn_SOUTH[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17.9000 0.0000 18.1000 0.6000 ;
    END
  END destinationAddressIn_SOUTH[4]
  PIN destinationAddressIn_SOUTH[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16.4000 0.0000 16.6000 0.6000 ;
    END
  END destinationAddressIn_SOUTH[3]
  PIN destinationAddressIn_SOUTH[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14.9000 0.0000 15.1000 0.6000 ;
    END
  END destinationAddressIn_SOUTH[2]
  PIN destinationAddressIn_SOUTH[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13.4000 0.0000 13.6000 0.6000 ;
    END
  END destinationAddressIn_SOUTH[1]
  PIN destinationAddressIn_SOUTH[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11.9000 0.0000 12.1000 0.6000 ;
    END
  END destinationAddressIn_SOUTH[0]
  PIN requesterAddressIn_SOUTH[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 40.4000 0.0000 40.6000 0.6000 ;
    END
  END requesterAddressIn_SOUTH[5]
  PIN requesterAddressIn_SOUTH[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.9000 0.0000 39.1000 0.6000 ;
    END
  END requesterAddressIn_SOUTH[4]
  PIN requesterAddressIn_SOUTH[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 37.4000 0.0000 37.6000 0.6000 ;
    END
  END requesterAddressIn_SOUTH[3]
  PIN requesterAddressIn_SOUTH[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 35.9000 0.0000 36.1000 0.6000 ;
    END
  END requesterAddressIn_SOUTH[2]
  PIN requesterAddressIn_SOUTH[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.4000 0.0000 34.6000 0.6000 ;
    END
  END requesterAddressIn_SOUTH[1]
  PIN requesterAddressIn_SOUTH[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 32.9000 0.0000 33.1000 0.6000 ;
    END
  END requesterAddressIn_SOUTH[0]
  PIN readIn_SOUTH
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 41.9000 0.0000 42.1000 0.6000 ;
    END
  END readIn_SOUTH
  PIN writeIn_SOUTH
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 43.4000 0.0000 43.6000 0.6000 ;
    END
  END writeIn_SOUTH
  PIN dataIn_SOUTH[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 91.4000 0.0000 91.6000 0.6000 ;
    END
  END dataIn_SOUTH[31]
  PIN dataIn_SOUTH[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 89.9000 0.0000 90.1000 0.6000 ;
    END
  END dataIn_SOUTH[30]
  PIN dataIn_SOUTH[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 88.4000 0.0000 88.6000 0.6000 ;
    END
  END dataIn_SOUTH[29]
  PIN dataIn_SOUTH[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 86.9000 0.0000 87.1000 0.6000 ;
    END
  END dataIn_SOUTH[28]
  PIN dataIn_SOUTH[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 85.4000 0.0000 85.6000 0.6000 ;
    END
  END dataIn_SOUTH[27]
  PIN dataIn_SOUTH[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 83.9000 0.0000 84.1000 0.6000 ;
    END
  END dataIn_SOUTH[26]
  PIN dataIn_SOUTH[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 82.4000 0.0000 82.6000 0.6000 ;
    END
  END dataIn_SOUTH[25]
  PIN dataIn_SOUTH[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 80.9000 0.0000 81.1000 0.6000 ;
    END
  END dataIn_SOUTH[24]
  PIN dataIn_SOUTH[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 79.4000 0.0000 79.6000 0.6000 ;
    END
  END dataIn_SOUTH[23]
  PIN dataIn_SOUTH[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 77.9000 0.0000 78.1000 0.6000 ;
    END
  END dataIn_SOUTH[22]
  PIN dataIn_SOUTH[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 76.4000 0.0000 76.6000 0.6000 ;
    END
  END dataIn_SOUTH[21]
  PIN dataIn_SOUTH[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 74.9000 0.0000 75.1000 0.6000 ;
    END
  END dataIn_SOUTH[20]
  PIN dataIn_SOUTH[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 73.4000 0.0000 73.6000 0.6000 ;
    END
  END dataIn_SOUTH[19]
  PIN dataIn_SOUTH[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 71.9000 0.0000 72.1000 0.6000 ;
    END
  END dataIn_SOUTH[18]
  PIN dataIn_SOUTH[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 70.4000 0.0000 70.6000 0.6000 ;
    END
  END dataIn_SOUTH[17]
  PIN dataIn_SOUTH[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 68.9000 0.0000 69.1000 0.6000 ;
    END
  END dataIn_SOUTH[16]
  PIN dataIn_SOUTH[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 67.4000 0.0000 67.6000 0.6000 ;
    END
  END dataIn_SOUTH[15]
  PIN dataIn_SOUTH[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 65.9000 0.0000 66.1000 0.6000 ;
    END
  END dataIn_SOUTH[14]
  PIN dataIn_SOUTH[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 64.4000 0.0000 64.6000 0.6000 ;
    END
  END dataIn_SOUTH[13]
  PIN dataIn_SOUTH[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 62.9000 0.0000 63.1000 0.6000 ;
    END
  END dataIn_SOUTH[12]
  PIN dataIn_SOUTH[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 61.4000 0.0000 61.6000 0.6000 ;
    END
  END dataIn_SOUTH[11]
  PIN dataIn_SOUTH[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 59.9000 0.0000 60.1000 0.6000 ;
    END
  END dataIn_SOUTH[10]
  PIN dataIn_SOUTH[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 58.4000 0.0000 58.6000 0.6000 ;
    END
  END dataIn_SOUTH[9]
  PIN dataIn_SOUTH[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 56.9000 0.0000 57.1000 0.6000 ;
    END
  END dataIn_SOUTH[8]
  PIN dataIn_SOUTH[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 55.4000 0.0000 55.6000 0.6000 ;
    END
  END dataIn_SOUTH[7]
  PIN dataIn_SOUTH[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 53.9000 0.0000 54.1000 0.6000 ;
    END
  END dataIn_SOUTH[6]
  PIN dataIn_SOUTH[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 52.4000 0.0000 52.6000 0.6000 ;
    END
  END dataIn_SOUTH[5]
  PIN dataIn_SOUTH[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 50.9000 0.0000 51.1000 0.6000 ;
    END
  END dataIn_SOUTH[4]
  PIN dataIn_SOUTH[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 49.4000 0.0000 49.6000 0.6000 ;
    END
  END dataIn_SOUTH[3]
  PIN dataIn_SOUTH[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 47.9000 0.0000 48.1000 0.6000 ;
    END
  END dataIn_SOUTH[2]
  PIN dataIn_SOUTH[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.4000 0.0000 46.6000 0.6000 ;
    END
  END dataIn_SOUTH[1]
  PIN dataIn_SOUTH[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44.9000 0.0000 45.1000 0.6000 ;
    END
  END dataIn_SOUTH[0]
  PIN destinationAddressOut_SOUTH[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 119.4000 0.0000 119.6000 0.6000 ;
    END
  END destinationAddressOut_SOUTH[13]
  PIN destinationAddressOut_SOUTH[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 117.9000 0.0000 118.1000 0.6000 ;
    END
  END destinationAddressOut_SOUTH[12]
  PIN destinationAddressOut_SOUTH[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 116.4000 0.0000 116.6000 0.6000 ;
    END
  END destinationAddressOut_SOUTH[11]
  PIN destinationAddressOut_SOUTH[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 114.9000 0.0000 115.1000 0.6000 ;
    END
  END destinationAddressOut_SOUTH[10]
  PIN destinationAddressOut_SOUTH[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 113.4000 0.0000 113.6000 0.6000 ;
    END
  END destinationAddressOut_SOUTH[9]
  PIN destinationAddressOut_SOUTH[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 111.9000 0.0000 112.1000 0.6000 ;
    END
  END destinationAddressOut_SOUTH[8]
  PIN destinationAddressOut_SOUTH[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 110.4000 0.0000 110.6000 0.6000 ;
    END
  END destinationAddressOut_SOUTH[7]
  PIN destinationAddressOut_SOUTH[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 108.9000 0.0000 109.1000 0.6000 ;
    END
  END destinationAddressOut_SOUTH[6]
  PIN destinationAddressOut_SOUTH[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 107.4000 0.0000 107.6000 0.6000 ;
    END
  END destinationAddressOut_SOUTH[5]
  PIN destinationAddressOut_SOUTH[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 105.9000 0.0000 106.1000 0.6000 ;
    END
  END destinationAddressOut_SOUTH[4]
  PIN destinationAddressOut_SOUTH[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 104.4000 0.0000 104.6000 0.6000 ;
    END
  END destinationAddressOut_SOUTH[3]
  PIN destinationAddressOut_SOUTH[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 102.9000 0.0000 103.1000 0.6000 ;
    END
  END destinationAddressOut_SOUTH[2]
  PIN destinationAddressOut_SOUTH[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 101.4000 0.0000 101.6000 0.6000 ;
    END
  END destinationAddressOut_SOUTH[1]
  PIN destinationAddressOut_SOUTH[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 99.9000 0.0000 100.1000 0.6000 ;
    END
  END destinationAddressOut_SOUTH[0]
  PIN requesterAddressOut_SOUTH[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 128.4000 0.0000 128.6000 0.6000 ;
    END
  END requesterAddressOut_SOUTH[5]
  PIN requesterAddressOut_SOUTH[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 126.9000 0.0000 127.1000 0.6000 ;
    END
  END requesterAddressOut_SOUTH[4]
  PIN requesterAddressOut_SOUTH[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 125.4000 0.0000 125.6000 0.6000 ;
    END
  END requesterAddressOut_SOUTH[3]
  PIN requesterAddressOut_SOUTH[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 123.9000 0.0000 124.1000 0.6000 ;
    END
  END requesterAddressOut_SOUTH[2]
  PIN requesterAddressOut_SOUTH[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 122.4000 0.0000 122.6000 0.6000 ;
    END
  END requesterAddressOut_SOUTH[1]
  PIN requesterAddressOut_SOUTH[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 120.9000 0.0000 121.1000 0.6000 ;
    END
  END requesterAddressOut_SOUTH[0]
  PIN readOut_SOUTH
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 129.9000 0.0000 130.1000 0.6000 ;
    END
  END readOut_SOUTH
  PIN writeOut_SOUTH
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 131.4000 0.0000 131.6000 0.6000 ;
    END
  END writeOut_SOUTH
  PIN dataOut_SOUTH[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 179.4000 0.0000 179.6000 0.6000 ;
    END
  END dataOut_SOUTH[31]
  PIN dataOut_SOUTH[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 177.9000 0.0000 178.1000 0.6000 ;
    END
  END dataOut_SOUTH[30]
  PIN dataOut_SOUTH[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 176.4000 0.0000 176.6000 0.6000 ;
    END
  END dataOut_SOUTH[29]
  PIN dataOut_SOUTH[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 174.9000 0.0000 175.1000 0.6000 ;
    END
  END dataOut_SOUTH[28]
  PIN dataOut_SOUTH[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 173.4000 0.0000 173.6000 0.6000 ;
    END
  END dataOut_SOUTH[27]
  PIN dataOut_SOUTH[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 171.9000 0.0000 172.1000 0.6000 ;
    END
  END dataOut_SOUTH[26]
  PIN dataOut_SOUTH[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 170.4000 0.0000 170.6000 0.6000 ;
    END
  END dataOut_SOUTH[25]
  PIN dataOut_SOUTH[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 168.9000 0.0000 169.1000 0.6000 ;
    END
  END dataOut_SOUTH[24]
  PIN dataOut_SOUTH[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 167.4000 0.0000 167.6000 0.6000 ;
    END
  END dataOut_SOUTH[23]
  PIN dataOut_SOUTH[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 165.9000 0.0000 166.1000 0.6000 ;
    END
  END dataOut_SOUTH[22]
  PIN dataOut_SOUTH[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 164.4000 0.0000 164.6000 0.6000 ;
    END
  END dataOut_SOUTH[21]
  PIN dataOut_SOUTH[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 162.9000 0.0000 163.1000 0.6000 ;
    END
  END dataOut_SOUTH[20]
  PIN dataOut_SOUTH[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 161.4000 0.0000 161.6000 0.6000 ;
    END
  END dataOut_SOUTH[19]
  PIN dataOut_SOUTH[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 159.9000 0.0000 160.1000 0.6000 ;
    END
  END dataOut_SOUTH[18]
  PIN dataOut_SOUTH[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 158.4000 0.0000 158.6000 0.6000 ;
    END
  END dataOut_SOUTH[17]
  PIN dataOut_SOUTH[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 156.9000 0.0000 157.1000 0.6000 ;
    END
  END dataOut_SOUTH[16]
  PIN dataOut_SOUTH[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 155.4000 0.0000 155.6000 0.6000 ;
    END
  END dataOut_SOUTH[15]
  PIN dataOut_SOUTH[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 153.9000 0.0000 154.1000 0.6000 ;
    END
  END dataOut_SOUTH[14]
  PIN dataOut_SOUTH[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 152.4000 0.0000 152.6000 0.6000 ;
    END
  END dataOut_SOUTH[13]
  PIN dataOut_SOUTH[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 150.9000 0.0000 151.1000 0.6000 ;
    END
  END dataOut_SOUTH[12]
  PIN dataOut_SOUTH[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 149.4000 0.0000 149.6000 0.6000 ;
    END
  END dataOut_SOUTH[11]
  PIN dataOut_SOUTH[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 147.9000 0.0000 148.1000 0.6000 ;
    END
  END dataOut_SOUTH[10]
  PIN dataOut_SOUTH[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 146.4000 0.0000 146.6000 0.6000 ;
    END
  END dataOut_SOUTH[9]
  PIN dataOut_SOUTH[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 144.9000 0.0000 145.1000 0.6000 ;
    END
  END dataOut_SOUTH[8]
  PIN dataOut_SOUTH[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 143.4000 0.0000 143.6000 0.6000 ;
    END
  END dataOut_SOUTH[7]
  PIN dataOut_SOUTH[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 141.9000 0.0000 142.1000 0.6000 ;
    END
  END dataOut_SOUTH[6]
  PIN dataOut_SOUTH[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 140.4000 0.0000 140.6000 0.6000 ;
    END
  END dataOut_SOUTH[5]
  PIN dataOut_SOUTH[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 138.9000 0.0000 139.1000 0.6000 ;
    END
  END dataOut_SOUTH[4]
  PIN dataOut_SOUTH[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 137.4000 0.0000 137.6000 0.6000 ;
    END
  END dataOut_SOUTH[3]
  PIN dataOut_SOUTH[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 135.9000 0.0000 136.1000 0.6000 ;
    END
  END dataOut_SOUTH[2]
  PIN dataOut_SOUTH[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 134.4000 0.0000 134.6000 0.6000 ;
    END
  END dataOut_SOUTH[1]
  PIN dataOut_SOUTH[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 132.9000 0.0000 133.1000 0.6000 ;
    END
  END dataOut_SOUTH[0]
  PIN destinationAddressIn_EAST[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 49.4000 666.0000 49.6000 ;
    END
  END destinationAddressIn_EAST[13]
  PIN destinationAddressIn_EAST[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 47.9000 666.0000 48.1000 ;
    END
  END destinationAddressIn_EAST[12]
  PIN destinationAddressIn_EAST[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 46.4000 666.0000 46.6000 ;
    END
  END destinationAddressIn_EAST[11]
  PIN destinationAddressIn_EAST[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 44.9000 666.0000 45.1000 ;
    END
  END destinationAddressIn_EAST[10]
  PIN destinationAddressIn_EAST[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 43.4000 666.0000 43.6000 ;
    END
  END destinationAddressIn_EAST[9]
  PIN destinationAddressIn_EAST[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 41.9000 666.0000 42.1000 ;
    END
  END destinationAddressIn_EAST[8]
  PIN destinationAddressIn_EAST[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 40.4000 666.0000 40.6000 ;
    END
  END destinationAddressIn_EAST[7]
  PIN destinationAddressIn_EAST[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 38.9000 666.0000 39.1000 ;
    END
  END destinationAddressIn_EAST[6]
  PIN destinationAddressIn_EAST[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 37.4000 666.0000 37.6000 ;
    END
  END destinationAddressIn_EAST[5]
  PIN destinationAddressIn_EAST[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 35.9000 666.0000 36.1000 ;
    END
  END destinationAddressIn_EAST[4]
  PIN destinationAddressIn_EAST[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 34.4000 666.0000 34.6000 ;
    END
  END destinationAddressIn_EAST[3]
  PIN destinationAddressIn_EAST[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 32.9000 666.0000 33.1000 ;
    END
  END destinationAddressIn_EAST[2]
  PIN destinationAddressIn_EAST[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 31.4000 666.0000 31.6000 ;
    END
  END destinationAddressIn_EAST[1]
  PIN destinationAddressIn_EAST[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 29.9000 666.0000 30.1000 ;
    END
  END destinationAddressIn_EAST[0]
  PIN requesterAddressIn_EAST[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 58.4000 666.0000 58.6000 ;
    END
  END requesterAddressIn_EAST[5]
  PIN requesterAddressIn_EAST[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 56.9000 666.0000 57.1000 ;
    END
  END requesterAddressIn_EAST[4]
  PIN requesterAddressIn_EAST[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 55.4000 666.0000 55.6000 ;
    END
  END requesterAddressIn_EAST[3]
  PIN requesterAddressIn_EAST[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 53.9000 666.0000 54.1000 ;
    END
  END requesterAddressIn_EAST[2]
  PIN requesterAddressIn_EAST[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 52.4000 666.0000 52.6000 ;
    END
  END requesterAddressIn_EAST[1]
  PIN requesterAddressIn_EAST[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 50.9000 666.0000 51.1000 ;
    END
  END requesterAddressIn_EAST[0]
  PIN readIn_EAST
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 59.9000 666.0000 60.1000 ;
    END
  END readIn_EAST
  PIN writeIn_EAST
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 61.4000 666.0000 61.6000 ;
    END
  END writeIn_EAST
  PIN dataIn_EAST[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 209.4000 666.0000 209.6000 ;
    END
  END dataIn_EAST[31]
  PIN dataIn_EAST[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 207.9000 666.0000 208.1000 ;
    END
  END dataIn_EAST[30]
  PIN dataIn_EAST[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 206.4000 666.0000 206.6000 ;
    END
  END dataIn_EAST[29]
  PIN dataIn_EAST[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 204.9000 666.0000 205.1000 ;
    END
  END dataIn_EAST[28]
  PIN dataIn_EAST[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 203.4000 666.0000 203.6000 ;
    END
  END dataIn_EAST[27]
  PIN dataIn_EAST[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 201.9000 666.0000 202.1000 ;
    END
  END dataIn_EAST[26]
  PIN dataIn_EAST[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 200.4000 666.0000 200.6000 ;
    END
  END dataIn_EAST[25]
  PIN dataIn_EAST[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 198.9000 666.0000 199.1000 ;
    END
  END dataIn_EAST[24]
  PIN dataIn_EAST[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 197.4000 666.0000 197.6000 ;
    END
  END dataIn_EAST[23]
  PIN dataIn_EAST[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 195.9000 666.0000 196.1000 ;
    END
  END dataIn_EAST[22]
  PIN dataIn_EAST[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 194.4000 666.0000 194.6000 ;
    END
  END dataIn_EAST[21]
  PIN dataIn_EAST[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 192.9000 666.0000 193.1000 ;
    END
  END dataIn_EAST[20]
  PIN dataIn_EAST[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 191.4000 666.0000 191.6000 ;
    END
  END dataIn_EAST[19]
  PIN dataIn_EAST[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 189.9000 666.0000 190.1000 ;
    END
  END dataIn_EAST[18]
  PIN dataIn_EAST[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 188.4000 666.0000 188.6000 ;
    END
  END dataIn_EAST[17]
  PIN dataIn_EAST[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 186.9000 666.0000 187.1000 ;
    END
  END dataIn_EAST[16]
  PIN dataIn_EAST[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 185.4000 666.0000 185.6000 ;
    END
  END dataIn_EAST[15]
  PIN dataIn_EAST[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 183.9000 666.0000 184.1000 ;
    END
  END dataIn_EAST[14]
  PIN dataIn_EAST[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 182.4000 666.0000 182.6000 ;
    END
  END dataIn_EAST[13]
  PIN dataIn_EAST[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 180.9000 666.0000 181.1000 ;
    END
  END dataIn_EAST[12]
  PIN dataIn_EAST[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 179.4000 666.0000 179.6000 ;
    END
  END dataIn_EAST[11]
  PIN dataIn_EAST[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 177.9000 666.0000 178.1000 ;
    END
  END dataIn_EAST[10]
  PIN dataIn_EAST[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 176.4000 666.0000 176.6000 ;
    END
  END dataIn_EAST[9]
  PIN dataIn_EAST[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 174.9000 666.0000 175.1000 ;
    END
  END dataIn_EAST[8]
  PIN dataIn_EAST[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 173.4000 666.0000 173.6000 ;
    END
  END dataIn_EAST[7]
  PIN dataIn_EAST[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 171.9000 666.0000 172.1000 ;
    END
  END dataIn_EAST[6]
  PIN dataIn_EAST[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 170.4000 666.0000 170.6000 ;
    END
  END dataIn_EAST[5]
  PIN dataIn_EAST[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 168.9000 666.0000 169.1000 ;
    END
  END dataIn_EAST[4]
  PIN dataIn_EAST[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 167.4000 666.0000 167.6000 ;
    END
  END dataIn_EAST[3]
  PIN dataIn_EAST[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 165.9000 666.0000 166.1000 ;
    END
  END dataIn_EAST[2]
  PIN dataIn_EAST[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 164.4000 666.0000 164.6000 ;
    END
  END dataIn_EAST[1]
  PIN dataIn_EAST[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 162.9000 666.0000 163.1000 ;
    END
  END dataIn_EAST[0]
  PIN destinationAddressOut_EAST[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 149.4000 666.0000 149.6000 ;
    END
  END destinationAddressOut_EAST[13]
  PIN destinationAddressOut_EAST[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 147.9000 666.0000 148.1000 ;
    END
  END destinationAddressOut_EAST[12]
  PIN destinationAddressOut_EAST[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 146.4000 666.0000 146.6000 ;
    END
  END destinationAddressOut_EAST[11]
  PIN destinationAddressOut_EAST[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 144.9000 666.0000 145.1000 ;
    END
  END destinationAddressOut_EAST[10]
  PIN destinationAddressOut_EAST[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 143.4000 666.0000 143.6000 ;
    END
  END destinationAddressOut_EAST[9]
  PIN destinationAddressOut_EAST[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 141.9000 666.0000 142.1000 ;
    END
  END destinationAddressOut_EAST[8]
  PIN destinationAddressOut_EAST[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 140.4000 666.0000 140.6000 ;
    END
  END destinationAddressOut_EAST[7]
  PIN destinationAddressOut_EAST[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 138.9000 666.0000 139.1000 ;
    END
  END destinationAddressOut_EAST[6]
  PIN destinationAddressOut_EAST[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 137.4000 666.0000 137.6000 ;
    END
  END destinationAddressOut_EAST[5]
  PIN destinationAddressOut_EAST[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 135.9000 666.0000 136.1000 ;
    END
  END destinationAddressOut_EAST[4]
  PIN destinationAddressOut_EAST[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 134.4000 666.0000 134.6000 ;
    END
  END destinationAddressOut_EAST[3]
  PIN destinationAddressOut_EAST[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 132.9000 666.0000 133.1000 ;
    END
  END destinationAddressOut_EAST[2]
  PIN destinationAddressOut_EAST[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 131.4000 666.0000 131.6000 ;
    END
  END destinationAddressOut_EAST[1]
  PIN destinationAddressOut_EAST[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 129.9000 666.0000 130.1000 ;
    END
  END destinationAddressOut_EAST[0]
  PIN requesterAddressOut_EAST[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 158.4000 666.0000 158.6000 ;
    END
  END requesterAddressOut_EAST[5]
  PIN requesterAddressOut_EAST[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 156.9000 666.0000 157.1000 ;
    END
  END requesterAddressOut_EAST[4]
  PIN requesterAddressOut_EAST[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 155.4000 666.0000 155.6000 ;
    END
  END requesterAddressOut_EAST[3]
  PIN requesterAddressOut_EAST[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 153.9000 666.0000 154.1000 ;
    END
  END requesterAddressOut_EAST[2]
  PIN requesterAddressOut_EAST[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 152.4000 666.0000 152.6000 ;
    END
  END requesterAddressOut_EAST[1]
  PIN requesterAddressOut_EAST[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 150.9000 666.0000 151.1000 ;
    END
  END requesterAddressOut_EAST[0]
  PIN readOut_EAST
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 159.9000 666.0000 160.1000 ;
    END
  END readOut_EAST
  PIN writeOut_EAST
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 161.4000 666.0000 161.6000 ;
    END
  END writeOut_EAST
  PIN dataOut_EAST[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 109.4000 666.0000 109.6000 ;
    END
  END dataOut_EAST[31]
  PIN dataOut_EAST[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 107.9000 666.0000 108.1000 ;
    END
  END dataOut_EAST[30]
  PIN dataOut_EAST[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 106.4000 666.0000 106.6000 ;
    END
  END dataOut_EAST[29]
  PIN dataOut_EAST[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 104.9000 666.0000 105.1000 ;
    END
  END dataOut_EAST[28]
  PIN dataOut_EAST[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 103.4000 666.0000 103.6000 ;
    END
  END dataOut_EAST[27]
  PIN dataOut_EAST[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 101.9000 666.0000 102.1000 ;
    END
  END dataOut_EAST[26]
  PIN dataOut_EAST[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 100.4000 666.0000 100.6000 ;
    END
  END dataOut_EAST[25]
  PIN dataOut_EAST[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 98.9000 666.0000 99.1000 ;
    END
  END dataOut_EAST[24]
  PIN dataOut_EAST[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 97.4000 666.0000 97.6000 ;
    END
  END dataOut_EAST[23]
  PIN dataOut_EAST[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 95.9000 666.0000 96.1000 ;
    END
  END dataOut_EAST[22]
  PIN dataOut_EAST[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 94.4000 666.0000 94.6000 ;
    END
  END dataOut_EAST[21]
  PIN dataOut_EAST[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 92.9000 666.0000 93.1000 ;
    END
  END dataOut_EAST[20]
  PIN dataOut_EAST[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 91.4000 666.0000 91.6000 ;
    END
  END dataOut_EAST[19]
  PIN dataOut_EAST[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 89.9000 666.0000 90.1000 ;
    END
  END dataOut_EAST[18]
  PIN dataOut_EAST[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 88.4000 666.0000 88.6000 ;
    END
  END dataOut_EAST[17]
  PIN dataOut_EAST[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 86.9000 666.0000 87.1000 ;
    END
  END dataOut_EAST[16]
  PIN dataOut_EAST[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 85.4000 666.0000 85.6000 ;
    END
  END dataOut_EAST[15]
  PIN dataOut_EAST[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 83.9000 666.0000 84.1000 ;
    END
  END dataOut_EAST[14]
  PIN dataOut_EAST[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 82.4000 666.0000 82.6000 ;
    END
  END dataOut_EAST[13]
  PIN dataOut_EAST[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 80.9000 666.0000 81.1000 ;
    END
  END dataOut_EAST[12]
  PIN dataOut_EAST[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 79.4000 666.0000 79.6000 ;
    END
  END dataOut_EAST[11]
  PIN dataOut_EAST[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 77.9000 666.0000 78.1000 ;
    END
  END dataOut_EAST[10]
  PIN dataOut_EAST[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 76.4000 666.0000 76.6000 ;
    END
  END dataOut_EAST[9]
  PIN dataOut_EAST[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 74.9000 666.0000 75.1000 ;
    END
  END dataOut_EAST[8]
  PIN dataOut_EAST[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 73.4000 666.0000 73.6000 ;
    END
  END dataOut_EAST[7]
  PIN dataOut_EAST[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 71.9000 666.0000 72.1000 ;
    END
  END dataOut_EAST[6]
  PIN dataOut_EAST[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 70.4000 666.0000 70.6000 ;
    END
  END dataOut_EAST[5]
  PIN dataOut_EAST[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 68.9000 666.0000 69.1000 ;
    END
  END dataOut_EAST[4]
  PIN dataOut_EAST[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 67.4000 666.0000 67.6000 ;
    END
  END dataOut_EAST[3]
  PIN dataOut_EAST[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 65.9000 666.0000 66.1000 ;
    END
  END dataOut_EAST[2]
  PIN dataOut_EAST[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 64.4000 666.0000 64.6000 ;
    END
  END dataOut_EAST[1]
  PIN dataOut_EAST[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 665.4000 62.9000 666.0000 63.1000 ;
    END
  END dataOut_EAST[0]
  PIN destinationAddressIn_WEST[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 53.4000 0.6000 53.6000 ;
    END
  END destinationAddressIn_WEST[13]
  PIN destinationAddressIn_WEST[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 51.9000 0.6000 52.1000 ;
    END
  END destinationAddressIn_WEST[12]
  PIN destinationAddressIn_WEST[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 50.4000 0.6000 50.6000 ;
    END
  END destinationAddressIn_WEST[11]
  PIN destinationAddressIn_WEST[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 48.9000 0.6000 49.1000 ;
    END
  END destinationAddressIn_WEST[10]
  PIN destinationAddressIn_WEST[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 47.4000 0.6000 47.6000 ;
    END
  END destinationAddressIn_WEST[9]
  PIN destinationAddressIn_WEST[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 45.9000 0.6000 46.1000 ;
    END
  END destinationAddressIn_WEST[8]
  PIN destinationAddressIn_WEST[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 44.4000 0.6000 44.6000 ;
    END
  END destinationAddressIn_WEST[7]
  PIN destinationAddressIn_WEST[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 42.9000 0.6000 43.1000 ;
    END
  END destinationAddressIn_WEST[6]
  PIN destinationAddressIn_WEST[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 41.4000 0.6000 41.6000 ;
    END
  END destinationAddressIn_WEST[5]
  PIN destinationAddressIn_WEST[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 39.9000 0.6000 40.1000 ;
    END
  END destinationAddressIn_WEST[4]
  PIN destinationAddressIn_WEST[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 38.4000 0.6000 38.6000 ;
    END
  END destinationAddressIn_WEST[3]
  PIN destinationAddressIn_WEST[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 36.9000 0.6000 37.1000 ;
    END
  END destinationAddressIn_WEST[2]
  PIN destinationAddressIn_WEST[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 35.4000 0.6000 35.6000 ;
    END
  END destinationAddressIn_WEST[1]
  PIN destinationAddressIn_WEST[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 33.9000 0.6000 34.1000 ;
    END
  END destinationAddressIn_WEST[0]
  PIN requesterAddressIn_WEST[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 62.4000 0.6000 62.6000 ;
    END
  END requesterAddressIn_WEST[5]
  PIN requesterAddressIn_WEST[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 60.9000 0.6000 61.1000 ;
    END
  END requesterAddressIn_WEST[4]
  PIN requesterAddressIn_WEST[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 59.4000 0.6000 59.6000 ;
    END
  END requesterAddressIn_WEST[3]
  PIN requesterAddressIn_WEST[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 57.9000 0.6000 58.1000 ;
    END
  END requesterAddressIn_WEST[2]
  PIN requesterAddressIn_WEST[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 56.4000 0.6000 56.6000 ;
    END
  END requesterAddressIn_WEST[1]
  PIN requesterAddressIn_WEST[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 54.9000 0.6000 55.1000 ;
    END
  END requesterAddressIn_WEST[0]
  PIN readIn_WEST
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 63.9000 0.6000 64.1000 ;
    END
  END readIn_WEST
  PIN writeIn_WEST
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 65.4000 0.6000 65.6000 ;
    END
  END writeIn_WEST
  PIN dataIn_WEST[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 113.4000 0.6000 113.6000 ;
    END
  END dataIn_WEST[31]
  PIN dataIn_WEST[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 111.9000 0.6000 112.1000 ;
    END
  END dataIn_WEST[30]
  PIN dataIn_WEST[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 110.4000 0.6000 110.6000 ;
    END
  END dataIn_WEST[29]
  PIN dataIn_WEST[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 108.9000 0.6000 109.1000 ;
    END
  END dataIn_WEST[28]
  PIN dataIn_WEST[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 107.4000 0.6000 107.6000 ;
    END
  END dataIn_WEST[27]
  PIN dataIn_WEST[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 105.9000 0.6000 106.1000 ;
    END
  END dataIn_WEST[26]
  PIN dataIn_WEST[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 104.4000 0.6000 104.6000 ;
    END
  END dataIn_WEST[25]
  PIN dataIn_WEST[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 102.9000 0.6000 103.1000 ;
    END
  END dataIn_WEST[24]
  PIN dataIn_WEST[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 101.4000 0.6000 101.6000 ;
    END
  END dataIn_WEST[23]
  PIN dataIn_WEST[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 99.9000 0.6000 100.1000 ;
    END
  END dataIn_WEST[22]
  PIN dataIn_WEST[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 98.4000 0.6000 98.6000 ;
    END
  END dataIn_WEST[21]
  PIN dataIn_WEST[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 96.9000 0.6000 97.1000 ;
    END
  END dataIn_WEST[20]
  PIN dataIn_WEST[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 95.4000 0.6000 95.6000 ;
    END
  END dataIn_WEST[19]
  PIN dataIn_WEST[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 93.9000 0.6000 94.1000 ;
    END
  END dataIn_WEST[18]
  PIN dataIn_WEST[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 92.4000 0.6000 92.6000 ;
    END
  END dataIn_WEST[17]
  PIN dataIn_WEST[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 90.9000 0.6000 91.1000 ;
    END
  END dataIn_WEST[16]
  PIN dataIn_WEST[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 89.4000 0.6000 89.6000 ;
    END
  END dataIn_WEST[15]
  PIN dataIn_WEST[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 87.9000 0.6000 88.1000 ;
    END
  END dataIn_WEST[14]
  PIN dataIn_WEST[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 86.4000 0.6000 86.6000 ;
    END
  END dataIn_WEST[13]
  PIN dataIn_WEST[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 84.9000 0.6000 85.1000 ;
    END
  END dataIn_WEST[12]
  PIN dataIn_WEST[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 83.4000 0.6000 83.6000 ;
    END
  END dataIn_WEST[11]
  PIN dataIn_WEST[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 81.9000 0.6000 82.1000 ;
    END
  END dataIn_WEST[10]
  PIN dataIn_WEST[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 80.4000 0.6000 80.6000 ;
    END
  END dataIn_WEST[9]
  PIN dataIn_WEST[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 78.9000 0.6000 79.1000 ;
    END
  END dataIn_WEST[8]
  PIN dataIn_WEST[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 77.4000 0.6000 77.6000 ;
    END
  END dataIn_WEST[7]
  PIN dataIn_WEST[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 75.9000 0.6000 76.1000 ;
    END
  END dataIn_WEST[6]
  PIN dataIn_WEST[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 74.4000 0.6000 74.6000 ;
    END
  END dataIn_WEST[5]
  PIN dataIn_WEST[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 72.9000 0.6000 73.1000 ;
    END
  END dataIn_WEST[4]
  PIN dataIn_WEST[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 71.4000 0.6000 71.6000 ;
    END
  END dataIn_WEST[3]
  PIN dataIn_WEST[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 69.9000 0.6000 70.1000 ;
    END
  END dataIn_WEST[2]
  PIN dataIn_WEST[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 68.4000 0.6000 68.6000 ;
    END
  END dataIn_WEST[1]
  PIN dataIn_WEST[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 66.9000 0.6000 67.1000 ;
    END
  END dataIn_WEST[0]
  PIN destinationAddressOut_WEST[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 130.4000 0.6000 130.6000 ;
    END
  END destinationAddressOut_WEST[13]
  PIN destinationAddressOut_WEST[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 128.9000 0.6000 129.1000 ;
    END
  END destinationAddressOut_WEST[12]
  PIN destinationAddressOut_WEST[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 127.4000 0.6000 127.6000 ;
    END
  END destinationAddressOut_WEST[11]
  PIN destinationAddressOut_WEST[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 125.9000 0.6000 126.1000 ;
    END
  END destinationAddressOut_WEST[10]
  PIN destinationAddressOut_WEST[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 124.4000 0.6000 124.6000 ;
    END
  END destinationAddressOut_WEST[9]
  PIN destinationAddressOut_WEST[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 122.9000 0.6000 123.1000 ;
    END
  END destinationAddressOut_WEST[8]
  PIN destinationAddressOut_WEST[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 121.4000 0.6000 121.6000 ;
    END
  END destinationAddressOut_WEST[7]
  PIN destinationAddressOut_WEST[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 119.9000 0.6000 120.1000 ;
    END
  END destinationAddressOut_WEST[6]
  PIN destinationAddressOut_WEST[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 118.4000 0.6000 118.6000 ;
    END
  END destinationAddressOut_WEST[5]
  PIN destinationAddressOut_WEST[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 116.9000 0.6000 117.1000 ;
    END
  END destinationAddressOut_WEST[4]
  PIN destinationAddressOut_WEST[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 115.4000 0.6000 115.6000 ;
    END
  END destinationAddressOut_WEST[3]
  PIN destinationAddressOut_WEST[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 113.9000 0.6000 114.1000 ;
    END
  END destinationAddressOut_WEST[2]
  PIN destinationAddressOut_WEST[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 112.4000 0.6000 112.6000 ;
    END
  END destinationAddressOut_WEST[1]
  PIN destinationAddressOut_WEST[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 110.9000 0.6000 111.1000 ;
    END
  END destinationAddressOut_WEST[0]
  PIN requesterAddressOut_WEST[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 139.4000 0.6000 139.6000 ;
    END
  END requesterAddressOut_WEST[5]
  PIN requesterAddressOut_WEST[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 137.9000 0.6000 138.1000 ;
    END
  END requesterAddressOut_WEST[4]
  PIN requesterAddressOut_WEST[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 136.4000 0.6000 136.6000 ;
    END
  END requesterAddressOut_WEST[3]
  PIN requesterAddressOut_WEST[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 134.9000 0.6000 135.1000 ;
    END
  END requesterAddressOut_WEST[2]
  PIN requesterAddressOut_WEST[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 133.4000 0.6000 133.6000 ;
    END
  END requesterAddressOut_WEST[1]
  PIN requesterAddressOut_WEST[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 131.9000 0.6000 132.1000 ;
    END
  END requesterAddressOut_WEST[0]
  PIN readOut_WEST
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 140.9000 0.6000 141.1000 ;
    END
  END readOut_WEST
  PIN writeOut_WEST
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 142.4000 0.6000 142.6000 ;
    END
  END writeOut_WEST
  PIN dataOut_WEST[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 190.4000 0.6000 190.6000 ;
    END
  END dataOut_WEST[31]
  PIN dataOut_WEST[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 188.9000 0.6000 189.1000 ;
    END
  END dataOut_WEST[30]
  PIN dataOut_WEST[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 187.4000 0.6000 187.6000 ;
    END
  END dataOut_WEST[29]
  PIN dataOut_WEST[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 185.9000 0.6000 186.1000 ;
    END
  END dataOut_WEST[28]
  PIN dataOut_WEST[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 184.4000 0.6000 184.6000 ;
    END
  END dataOut_WEST[27]
  PIN dataOut_WEST[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 182.9000 0.6000 183.1000 ;
    END
  END dataOut_WEST[26]
  PIN dataOut_WEST[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 181.4000 0.6000 181.6000 ;
    END
  END dataOut_WEST[25]
  PIN dataOut_WEST[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 179.9000 0.6000 180.1000 ;
    END
  END dataOut_WEST[24]
  PIN dataOut_WEST[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 178.4000 0.6000 178.6000 ;
    END
  END dataOut_WEST[23]
  PIN dataOut_WEST[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 176.9000 0.6000 177.1000 ;
    END
  END dataOut_WEST[22]
  PIN dataOut_WEST[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 175.4000 0.6000 175.6000 ;
    END
  END dataOut_WEST[21]
  PIN dataOut_WEST[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 173.9000 0.6000 174.1000 ;
    END
  END dataOut_WEST[20]
  PIN dataOut_WEST[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 172.4000 0.6000 172.6000 ;
    END
  END dataOut_WEST[19]
  PIN dataOut_WEST[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 170.9000 0.6000 171.1000 ;
    END
  END dataOut_WEST[18]
  PIN dataOut_WEST[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 169.4000 0.6000 169.6000 ;
    END
  END dataOut_WEST[17]
  PIN dataOut_WEST[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 167.9000 0.6000 168.1000 ;
    END
  END dataOut_WEST[16]
  PIN dataOut_WEST[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 166.4000 0.6000 166.6000 ;
    END
  END dataOut_WEST[15]
  PIN dataOut_WEST[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 164.9000 0.6000 165.1000 ;
    END
  END dataOut_WEST[14]
  PIN dataOut_WEST[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 163.4000 0.6000 163.6000 ;
    END
  END dataOut_WEST[13]
  PIN dataOut_WEST[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 161.9000 0.6000 162.1000 ;
    END
  END dataOut_WEST[12]
  PIN dataOut_WEST[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 160.4000 0.6000 160.6000 ;
    END
  END dataOut_WEST[11]
  PIN dataOut_WEST[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 158.9000 0.6000 159.1000 ;
    END
  END dataOut_WEST[10]
  PIN dataOut_WEST[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 157.4000 0.6000 157.6000 ;
    END
  END dataOut_WEST[9]
  PIN dataOut_WEST[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 155.9000 0.6000 156.1000 ;
    END
  END dataOut_WEST[8]
  PIN dataOut_WEST[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 154.4000 0.6000 154.6000 ;
    END
  END dataOut_WEST[7]
  PIN dataOut_WEST[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 152.9000 0.6000 153.1000 ;
    END
  END dataOut_WEST[6]
  PIN dataOut_WEST[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 151.4000 0.6000 151.6000 ;
    END
  END dataOut_WEST[5]
  PIN dataOut_WEST[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 149.9000 0.6000 150.1000 ;
    END
  END dataOut_WEST[4]
  PIN dataOut_WEST[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 148.4000 0.6000 148.6000 ;
    END
  END dataOut_WEST[3]
  PIN dataOut_WEST[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 146.9000 0.6000 147.1000 ;
    END
  END dataOut_WEST[2]
  PIN dataOut_WEST[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 145.4000 0.6000 145.6000 ;
    END
  END dataOut_WEST[1]
  PIN dataOut_WEST[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 143.9000 0.6000 144.1000 ;
    END
  END dataOut_WEST[0]
  PIN cacheDataIn_A[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 228.4000 0.0000 228.6000 0.6000 ;
    END
  END cacheDataIn_A[31]
  PIN cacheDataIn_A[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 226.9000 0.0000 227.1000 0.6000 ;
    END
  END cacheDataIn_A[30]
  PIN cacheDataIn_A[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 225.4000 0.0000 225.6000 0.6000 ;
    END
  END cacheDataIn_A[29]
  PIN cacheDataIn_A[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 223.9000 0.0000 224.1000 0.6000 ;
    END
  END cacheDataIn_A[28]
  PIN cacheDataIn_A[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 222.4000 0.0000 222.6000 0.6000 ;
    END
  END cacheDataIn_A[27]
  PIN cacheDataIn_A[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 220.9000 0.0000 221.1000 0.6000 ;
    END
  END cacheDataIn_A[26]
  PIN cacheDataIn_A[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 219.4000 0.0000 219.6000 0.6000 ;
    END
  END cacheDataIn_A[25]
  PIN cacheDataIn_A[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 217.9000 0.0000 218.1000 0.6000 ;
    END
  END cacheDataIn_A[24]
  PIN cacheDataIn_A[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 216.4000 0.0000 216.6000 0.6000 ;
    END
  END cacheDataIn_A[23]
  PIN cacheDataIn_A[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 214.9000 0.0000 215.1000 0.6000 ;
    END
  END cacheDataIn_A[22]
  PIN cacheDataIn_A[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 213.4000 0.0000 213.6000 0.6000 ;
    END
  END cacheDataIn_A[21]
  PIN cacheDataIn_A[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 211.9000 0.0000 212.1000 0.6000 ;
    END
  END cacheDataIn_A[20]
  PIN cacheDataIn_A[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 210.4000 0.0000 210.6000 0.6000 ;
    END
  END cacheDataIn_A[19]
  PIN cacheDataIn_A[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 208.9000 0.0000 209.1000 0.6000 ;
    END
  END cacheDataIn_A[18]
  PIN cacheDataIn_A[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 207.4000 0.0000 207.6000 0.6000 ;
    END
  END cacheDataIn_A[17]
  PIN cacheDataIn_A[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 205.9000 0.0000 206.1000 0.6000 ;
    END
  END cacheDataIn_A[16]
  PIN cacheDataIn_A[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 204.4000 0.0000 204.6000 0.6000 ;
    END
  END cacheDataIn_A[15]
  PIN cacheDataIn_A[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 202.9000 0.0000 203.1000 0.6000 ;
    END
  END cacheDataIn_A[14]
  PIN cacheDataIn_A[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 201.4000 0.0000 201.6000 0.6000 ;
    END
  END cacheDataIn_A[13]
  PIN cacheDataIn_A[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 199.9000 0.0000 200.1000 0.6000 ;
    END
  END cacheDataIn_A[12]
  PIN cacheDataIn_A[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 198.4000 0.0000 198.6000 0.6000 ;
    END
  END cacheDataIn_A[11]
  PIN cacheDataIn_A[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 196.9000 0.0000 197.1000 0.6000 ;
    END
  END cacheDataIn_A[10]
  PIN cacheDataIn_A[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 195.4000 0.0000 195.6000 0.6000 ;
    END
  END cacheDataIn_A[9]
  PIN cacheDataIn_A[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 193.9000 0.0000 194.1000 0.6000 ;
    END
  END cacheDataIn_A[8]
  PIN cacheDataIn_A[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 192.4000 0.0000 192.6000 0.6000 ;
    END
  END cacheDataIn_A[7]
  PIN cacheDataIn_A[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 190.9000 0.0000 191.1000 0.6000 ;
    END
  END cacheDataIn_A[6]
  PIN cacheDataIn_A[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 189.4000 0.0000 189.6000 0.6000 ;
    END
  END cacheDataIn_A[5]
  PIN cacheDataIn_A[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 187.9000 0.0000 188.1000 0.6000 ;
    END
  END cacheDataIn_A[4]
  PIN cacheDataIn_A[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 186.4000 0.0000 186.6000 0.6000 ;
    END
  END cacheDataIn_A[3]
  PIN cacheDataIn_A[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 184.9000 0.0000 185.1000 0.6000 ;
    END
  END cacheDataIn_A[2]
  PIN cacheDataIn_A[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 183.4000 0.0000 183.6000 0.6000 ;
    END
  END cacheDataIn_A[1]
  PIN cacheDataIn_A[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 181.9000 0.0000 182.1000 0.6000 ;
    END
  END cacheDataIn_A[0]
  PIN cacheAddressIn_A[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 240.4000 0.0000 240.6000 0.6000 ;
    END
  END cacheAddressIn_A[7]
  PIN cacheAddressIn_A[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 238.9000 0.0000 239.1000 0.6000 ;
    END
  END cacheAddressIn_A[6]
  PIN cacheAddressIn_A[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 237.4000 0.0000 237.6000 0.6000 ;
    END
  END cacheAddressIn_A[5]
  PIN cacheAddressIn_A[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 235.9000 0.0000 236.1000 0.6000 ;
    END
  END cacheAddressIn_A[4]
  PIN cacheAddressIn_A[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 234.4000 0.0000 234.6000 0.6000 ;
    END
  END cacheAddressIn_A[3]
  PIN cacheAddressIn_A[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 232.9000 0.0000 233.1000 0.6000 ;
    END
  END cacheAddressIn_A[2]
  PIN cacheAddressIn_A[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 231.4000 0.0000 231.6000 0.6000 ;
    END
  END cacheAddressIn_A[1]
  PIN cacheAddressIn_A[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 229.9000 0.0000 230.1000 0.6000 ;
    END
  END cacheAddressIn_A[0]
  PIN cacheDataOut_A[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 288.4000 0.0000 288.6000 0.6000 ;
    END
  END cacheDataOut_A[31]
  PIN cacheDataOut_A[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 286.9000 0.0000 287.1000 0.6000 ;
    END
  END cacheDataOut_A[30]
  PIN cacheDataOut_A[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 285.4000 0.0000 285.6000 0.6000 ;
    END
  END cacheDataOut_A[29]
  PIN cacheDataOut_A[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 283.9000 0.0000 284.1000 0.6000 ;
    END
  END cacheDataOut_A[28]
  PIN cacheDataOut_A[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 282.4000 0.0000 282.6000 0.6000 ;
    END
  END cacheDataOut_A[27]
  PIN cacheDataOut_A[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 280.9000 0.0000 281.1000 0.6000 ;
    END
  END cacheDataOut_A[26]
  PIN cacheDataOut_A[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 279.4000 0.0000 279.6000 0.6000 ;
    END
  END cacheDataOut_A[25]
  PIN cacheDataOut_A[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 277.9000 0.0000 278.1000 0.6000 ;
    END
  END cacheDataOut_A[24]
  PIN cacheDataOut_A[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 276.4000 0.0000 276.6000 0.6000 ;
    END
  END cacheDataOut_A[23]
  PIN cacheDataOut_A[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 274.9000 0.0000 275.1000 0.6000 ;
    END
  END cacheDataOut_A[22]
  PIN cacheDataOut_A[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 273.4000 0.0000 273.6000 0.6000 ;
    END
  END cacheDataOut_A[21]
  PIN cacheDataOut_A[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 271.9000 0.0000 272.1000 0.6000 ;
    END
  END cacheDataOut_A[20]
  PIN cacheDataOut_A[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 270.4000 0.0000 270.6000 0.6000 ;
    END
  END cacheDataOut_A[19]
  PIN cacheDataOut_A[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 268.9000 0.0000 269.1000 0.6000 ;
    END
  END cacheDataOut_A[18]
  PIN cacheDataOut_A[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 267.4000 0.0000 267.6000 0.6000 ;
    END
  END cacheDataOut_A[17]
  PIN cacheDataOut_A[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 265.9000 0.0000 266.1000 0.6000 ;
    END
  END cacheDataOut_A[16]
  PIN cacheDataOut_A[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 264.4000 0.0000 264.6000 0.6000 ;
    END
  END cacheDataOut_A[15]
  PIN cacheDataOut_A[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 262.9000 0.0000 263.1000 0.6000 ;
    END
  END cacheDataOut_A[14]
  PIN cacheDataOut_A[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 261.4000 0.0000 261.6000 0.6000 ;
    END
  END cacheDataOut_A[13]
  PIN cacheDataOut_A[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 259.9000 0.0000 260.1000 0.6000 ;
    END
  END cacheDataOut_A[12]
  PIN cacheDataOut_A[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 258.4000 0.0000 258.6000 0.6000 ;
    END
  END cacheDataOut_A[11]
  PIN cacheDataOut_A[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 256.9000 0.0000 257.1000 0.6000 ;
    END
  END cacheDataOut_A[10]
  PIN cacheDataOut_A[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 255.4000 0.0000 255.6000 0.6000 ;
    END
  END cacheDataOut_A[9]
  PIN cacheDataOut_A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 253.9000 0.0000 254.1000 0.6000 ;
    END
  END cacheDataOut_A[8]
  PIN cacheDataOut_A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 252.4000 0.0000 252.6000 0.6000 ;
    END
  END cacheDataOut_A[7]
  PIN cacheDataOut_A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 250.9000 0.0000 251.1000 0.6000 ;
    END
  END cacheDataOut_A[6]
  PIN cacheDataOut_A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 249.4000 0.0000 249.6000 0.6000 ;
    END
  END cacheDataOut_A[5]
  PIN cacheDataOut_A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 247.9000 0.0000 248.1000 0.6000 ;
    END
  END cacheDataOut_A[4]
  PIN cacheDataOut_A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 246.4000 0.0000 246.6000 0.6000 ;
    END
  END cacheDataOut_A[3]
  PIN cacheDataOut_A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 244.9000 0.0000 245.1000 0.6000 ;
    END
  END cacheDataOut_A[2]
  PIN cacheDataOut_A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 243.4000 0.0000 243.6000 0.6000 ;
    END
  END cacheDataOut_A[1]
  PIN cacheDataOut_A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 241.9000 0.0000 242.1000 0.6000 ;
    END
  END cacheDataOut_A[0]
  PIN memWrite_A
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 289.9000 0.0000 290.1000 0.6000 ;
    END
  END memWrite_A
  PIN portA_writtenTo
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 291.4000 0.0000 291.6000 0.6000 ;
    END
  END portA_writtenTo
  PIN cacheDataIn_B[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 341.4000 0.0000 341.6000 0.6000 ;
    END
  END cacheDataIn_B[31]
  PIN cacheDataIn_B[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 339.9000 0.0000 340.1000 0.6000 ;
    END
  END cacheDataIn_B[30]
  PIN cacheDataIn_B[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 338.4000 0.0000 338.6000 0.6000 ;
    END
  END cacheDataIn_B[29]
  PIN cacheDataIn_B[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 336.9000 0.0000 337.1000 0.6000 ;
    END
  END cacheDataIn_B[28]
  PIN cacheDataIn_B[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 335.4000 0.0000 335.6000 0.6000 ;
    END
  END cacheDataIn_B[27]
  PIN cacheDataIn_B[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 333.9000 0.0000 334.1000 0.6000 ;
    END
  END cacheDataIn_B[26]
  PIN cacheDataIn_B[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 332.4000 0.0000 332.6000 0.6000 ;
    END
  END cacheDataIn_B[25]
  PIN cacheDataIn_B[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 330.9000 0.0000 331.1000 0.6000 ;
    END
  END cacheDataIn_B[24]
  PIN cacheDataIn_B[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 329.4000 0.0000 329.6000 0.6000 ;
    END
  END cacheDataIn_B[23]
  PIN cacheDataIn_B[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 327.9000 0.0000 328.1000 0.6000 ;
    END
  END cacheDataIn_B[22]
  PIN cacheDataIn_B[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 326.4000 0.0000 326.6000 0.6000 ;
    END
  END cacheDataIn_B[21]
  PIN cacheDataIn_B[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 324.9000 0.0000 325.1000 0.6000 ;
    END
  END cacheDataIn_B[20]
  PIN cacheDataIn_B[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 323.4000 0.0000 323.6000 0.6000 ;
    END
  END cacheDataIn_B[19]
  PIN cacheDataIn_B[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 321.9000 0.0000 322.1000 0.6000 ;
    END
  END cacheDataIn_B[18]
  PIN cacheDataIn_B[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 320.4000 0.0000 320.6000 0.6000 ;
    END
  END cacheDataIn_B[17]
  PIN cacheDataIn_B[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 318.9000 0.0000 319.1000 0.6000 ;
    END
  END cacheDataIn_B[16]
  PIN cacheDataIn_B[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 317.4000 0.0000 317.6000 0.6000 ;
    END
  END cacheDataIn_B[15]
  PIN cacheDataIn_B[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 315.9000 0.0000 316.1000 0.6000 ;
    END
  END cacheDataIn_B[14]
  PIN cacheDataIn_B[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 314.4000 0.0000 314.6000 0.6000 ;
    END
  END cacheDataIn_B[13]
  PIN cacheDataIn_B[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 312.9000 0.0000 313.1000 0.6000 ;
    END
  END cacheDataIn_B[12]
  PIN cacheDataIn_B[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 311.4000 0.0000 311.6000 0.6000 ;
    END
  END cacheDataIn_B[11]
  PIN cacheDataIn_B[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 309.9000 0.0000 310.1000 0.6000 ;
    END
  END cacheDataIn_B[10]
  PIN cacheDataIn_B[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 308.4000 0.0000 308.6000 0.6000 ;
    END
  END cacheDataIn_B[9]
  PIN cacheDataIn_B[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 306.9000 0.0000 307.1000 0.6000 ;
    END
  END cacheDataIn_B[8]
  PIN cacheDataIn_B[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 305.4000 0.0000 305.6000 0.6000 ;
    END
  END cacheDataIn_B[7]
  PIN cacheDataIn_B[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 303.9000 0.0000 304.1000 0.6000 ;
    END
  END cacheDataIn_B[6]
  PIN cacheDataIn_B[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 302.4000 0.0000 302.6000 0.6000 ;
    END
  END cacheDataIn_B[5]
  PIN cacheDataIn_B[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 300.9000 0.0000 301.1000 0.6000 ;
    END
  END cacheDataIn_B[4]
  PIN cacheDataIn_B[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 299.4000 0.0000 299.6000 0.6000 ;
    END
  END cacheDataIn_B[3]
  PIN cacheDataIn_B[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 297.9000 0.0000 298.1000 0.6000 ;
    END
  END cacheDataIn_B[2]
  PIN cacheDataIn_B[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 296.4000 0.0000 296.6000 0.6000 ;
    END
  END cacheDataIn_B[1]
  PIN cacheDataIn_B[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 294.9000 0.0000 295.1000 0.6000 ;
    END
  END cacheDataIn_B[0]
  PIN cacheAddressIn_B[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 353.4000 0.0000 353.6000 0.6000 ;
    END
  END cacheAddressIn_B[7]
  PIN cacheAddressIn_B[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 351.9000 0.0000 352.1000 0.6000 ;
    END
  END cacheAddressIn_B[6]
  PIN cacheAddressIn_B[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 350.4000 0.0000 350.6000 0.6000 ;
    END
  END cacheAddressIn_B[5]
  PIN cacheAddressIn_B[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 348.9000 0.0000 349.1000 0.6000 ;
    END
  END cacheAddressIn_B[4]
  PIN cacheAddressIn_B[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 347.4000 0.0000 347.6000 0.6000 ;
    END
  END cacheAddressIn_B[3]
  PIN cacheAddressIn_B[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 345.9000 0.0000 346.1000 0.6000 ;
    END
  END cacheAddressIn_B[2]
  PIN cacheAddressIn_B[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 344.4000 0.0000 344.6000 0.6000 ;
    END
  END cacheAddressIn_B[1]
  PIN cacheAddressIn_B[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 342.9000 0.0000 343.1000 0.6000 ;
    END
  END cacheAddressIn_B[0]
  PIN cacheDataOut_B[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 401.4000 0.0000 401.6000 0.6000 ;
    END
  END cacheDataOut_B[31]
  PIN cacheDataOut_B[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 399.9000 0.0000 400.1000 0.6000 ;
    END
  END cacheDataOut_B[30]
  PIN cacheDataOut_B[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 398.4000 0.0000 398.6000 0.6000 ;
    END
  END cacheDataOut_B[29]
  PIN cacheDataOut_B[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 396.9000 0.0000 397.1000 0.6000 ;
    END
  END cacheDataOut_B[28]
  PIN cacheDataOut_B[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 395.4000 0.0000 395.6000 0.6000 ;
    END
  END cacheDataOut_B[27]
  PIN cacheDataOut_B[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 393.9000 0.0000 394.1000 0.6000 ;
    END
  END cacheDataOut_B[26]
  PIN cacheDataOut_B[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 392.4000 0.0000 392.6000 0.6000 ;
    END
  END cacheDataOut_B[25]
  PIN cacheDataOut_B[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 390.9000 0.0000 391.1000 0.6000 ;
    END
  END cacheDataOut_B[24]
  PIN cacheDataOut_B[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 389.4000 0.0000 389.6000 0.6000 ;
    END
  END cacheDataOut_B[23]
  PIN cacheDataOut_B[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 387.9000 0.0000 388.1000 0.6000 ;
    END
  END cacheDataOut_B[22]
  PIN cacheDataOut_B[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 386.4000 0.0000 386.6000 0.6000 ;
    END
  END cacheDataOut_B[21]
  PIN cacheDataOut_B[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 384.9000 0.0000 385.1000 0.6000 ;
    END
  END cacheDataOut_B[20]
  PIN cacheDataOut_B[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 383.4000 0.0000 383.6000 0.6000 ;
    END
  END cacheDataOut_B[19]
  PIN cacheDataOut_B[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 381.9000 0.0000 382.1000 0.6000 ;
    END
  END cacheDataOut_B[18]
  PIN cacheDataOut_B[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 380.4000 0.0000 380.6000 0.6000 ;
    END
  END cacheDataOut_B[17]
  PIN cacheDataOut_B[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 378.9000 0.0000 379.1000 0.6000 ;
    END
  END cacheDataOut_B[16]
  PIN cacheDataOut_B[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 377.4000 0.0000 377.6000 0.6000 ;
    END
  END cacheDataOut_B[15]
  PIN cacheDataOut_B[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 375.9000 0.0000 376.1000 0.6000 ;
    END
  END cacheDataOut_B[14]
  PIN cacheDataOut_B[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 374.4000 0.0000 374.6000 0.6000 ;
    END
  END cacheDataOut_B[13]
  PIN cacheDataOut_B[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 372.9000 0.0000 373.1000 0.6000 ;
    END
  END cacheDataOut_B[12]
  PIN cacheDataOut_B[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 371.4000 0.0000 371.6000 0.6000 ;
    END
  END cacheDataOut_B[11]
  PIN cacheDataOut_B[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 369.9000 0.0000 370.1000 0.6000 ;
    END
  END cacheDataOut_B[10]
  PIN cacheDataOut_B[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 368.4000 0.0000 368.6000 0.6000 ;
    END
  END cacheDataOut_B[9]
  PIN cacheDataOut_B[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 366.9000 0.0000 367.1000 0.6000 ;
    END
  END cacheDataOut_B[8]
  PIN cacheDataOut_B[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 365.4000 0.0000 365.6000 0.6000 ;
    END
  END cacheDataOut_B[7]
  PIN cacheDataOut_B[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 363.9000 0.0000 364.1000 0.6000 ;
    END
  END cacheDataOut_B[6]
  PIN cacheDataOut_B[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 362.4000 0.0000 362.6000 0.6000 ;
    END
  END cacheDataOut_B[5]
  PIN cacheDataOut_B[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 360.9000 0.0000 361.1000 0.6000 ;
    END
  END cacheDataOut_B[4]
  PIN cacheDataOut_B[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 359.4000 0.0000 359.6000 0.6000 ;
    END
  END cacheDataOut_B[3]
  PIN cacheDataOut_B[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 357.9000 0.0000 358.1000 0.6000 ;
    END
  END cacheDataOut_B[2]
  PIN cacheDataOut_B[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 356.4000 0.0000 356.6000 0.6000 ;
    END
  END cacheDataOut_B[1]
  PIN cacheDataOut_B[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 354.9000 0.0000 355.1000 0.6000 ;
    END
  END cacheDataOut_B[0]
  PIN memWrite_B
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 402.9000 0.0000 403.1000 0.6000 ;
    END
  END memWrite_B
  PIN portB_writtenTo
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 404.4000 0.0000 404.6000 0.6000 ;
    END
  END portB_writtenTo
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 666.0000 612.0000 ;
    LAYER M2 ;
      RECT 181.5200 609.4800 666.0000 612.0000 ;
      RECT 93.5200 609.4800 97.9800 612.0000 ;
      RECT 0.0000 609.4800 9.9800 612.0000 ;
      RECT 0.0000 211.5200 666.0000 609.4800 ;
      RECT 0.0000 192.5200 663.4800 211.5200 ;
      RECT 2.5200 127.9800 663.4800 192.5200 ;
      RECT 2.5200 111.5200 666.0000 127.9800 ;
      RECT 2.5200 31.9800 663.4800 111.5200 ;
      RECT 0.0000 29.0200 663.4800 31.9800 ;
      RECT 2.5200 27.9800 663.4800 29.0200 ;
      RECT 2.5200 14.9800 666.0000 27.9800 ;
      RECT 0.0000 2.5200 666.0000 14.9800 ;
      RECT 406.5200 0.0000 666.0000 2.5200 ;
      RECT 93.5200 0.0000 97.9800 2.5200 ;
      RECT 0.0000 0.0000 9.9800 2.5200 ;
    LAYER M3 ;
      RECT 0.0000 13.0200 666.0000 612.0000 ;
      RECT 2.5200 8.9800 666.0000 13.0200 ;
      RECT 0.0000 0.0000 666.0000 8.9800 ;
    LAYER MQ ;
      RECT 0.0000 3.1200 666.0000 612.0000 ;
      RECT 361.9200 0.0000 666.0000 3.1200 ;
      RECT 0.0000 0.0000 357.6800 3.1200 ;
  END
END router

END LIBRARY
