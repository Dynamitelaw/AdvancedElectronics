
module cacheAccessArbiter ( clk, reset, cacheAddressIn_NORTH, 
        requesterAddressIn_NORTH, memRead_NORTH, memWrite_NORTH, dataIn_NORTH, 
        readReady_NORTH, requesterAddressOut_NORTH, cacheDataOut_NORTH, 
        cacheAddressIn_SOUTH, requesterAddressIn_SOUTH, memRead_SOUTH, 
        memWrite_SOUTH, dataIn_SOUTH, readReady_SOUTH, 
        requesterAddressOut_SOUTH, cacheDataOut_SOUTH, cacheAddressIn_EAST, 
        requesterAddressIn_EAST, memRead_EAST, memWrite_EAST, dataIn_EAST, 
        readReady_EAST, requesterAddressOut_EAST, cacheDataOut_EAST, 
        cacheAddressIn_WEST, requesterAddressIn_WEST, memRead_WEST, 
        memWrite_WEST, dataIn_WEST, readReady_WEST, requesterAddressOut_WEST, 
        cacheDataOut_WEST, cacheDataIn_A, cacheAddressIn_A, cacheDataOut_A, 
        memWrite_A, cacheDataIn_B, cacheAddressIn_B, cacheDataOut_B, 
        memWrite_B );
  input [7:0] cacheAddressIn_NORTH;
  input [3:0] requesterAddressIn_NORTH;
  input [5:0] dataIn_NORTH;
  output [3:0] requesterAddressOut_NORTH;
  output [5:0] cacheDataOut_NORTH;
  input [7:0] cacheAddressIn_SOUTH;
  input [3:0] requesterAddressIn_SOUTH;
  input [5:0] dataIn_SOUTH;
  output [3:0] requesterAddressOut_SOUTH;
  output [5:0] cacheDataOut_SOUTH;
  input [7:0] cacheAddressIn_EAST;
  input [3:0] requesterAddressIn_EAST;
  input [5:0] dataIn_EAST;
  output [3:0] requesterAddressOut_EAST;
  output [5:0] cacheDataOut_EAST;
  input [7:0] cacheAddressIn_WEST;
  input [3:0] requesterAddressIn_WEST;
  input [5:0] dataIn_WEST;
  output [3:0] requesterAddressOut_WEST;
  output [5:0] cacheDataOut_WEST;
  output [5:0] cacheDataIn_A;
  output [7:0] cacheAddressIn_A;
  input [5:0] cacheDataOut_A;
  output [5:0] cacheDataIn_B;
  output [7:0] cacheAddressIn_B;
  input [5:0] cacheDataOut_B;
  input clk, reset, memRead_NORTH, memWrite_NORTH, memRead_SOUTH,
         memWrite_SOUTH, memRead_EAST, memWrite_EAST, memRead_WEST,
         memWrite_WEST;
  output readReady_NORTH, readReady_SOUTH, readReady_EAST, readReady_WEST,
         memWrite_A, memWrite_B;
  wire   N882, N883, N884, \dataToWriteBuffer[6][5] ,
         \dataToWriteBuffer[6][4] , \dataToWriteBuffer[6][3] ,
         \dataToWriteBuffer[6][2] , \dataToWriteBuffer[6][1] ,
         \dataToWriteBuffer[6][0] , \dataToWriteBuffer[5][5] ,
         \dataToWriteBuffer[5][4] , \dataToWriteBuffer[5][3] ,
         \dataToWriteBuffer[5][2] , \dataToWriteBuffer[5][1] ,
         \dataToWriteBuffer[5][0] , \dataToWriteBuffer[4][5] ,
         \dataToWriteBuffer[4][4] , \dataToWriteBuffer[4][3] ,
         \dataToWriteBuffer[4][2] , \dataToWriteBuffer[4][1] ,
         \dataToWriteBuffer[4][0] , \dataToWriteBuffer[3][5] ,
         \dataToWriteBuffer[3][4] , \dataToWriteBuffer[3][3] ,
         \dataToWriteBuffer[3][2] , \dataToWriteBuffer[3][1] ,
         \dataToWriteBuffer[3][0] , \dataToWriteBuffer[2][5] ,
         \dataToWriteBuffer[2][4] , \dataToWriteBuffer[2][3] ,
         \dataToWriteBuffer[2][2] , \dataToWriteBuffer[2][1] ,
         \dataToWriteBuffer[2][0] , \dataToWriteBuffer[1][5] ,
         \dataToWriteBuffer[1][4] , \dataToWriteBuffer[1][3] ,
         \dataToWriteBuffer[1][2] , \dataToWriteBuffer[1][1] ,
         \dataToWriteBuffer[1][0] , \dataToWriteBuffer[0][5] ,
         \dataToWriteBuffer[0][4] , \dataToWriteBuffer[0][3] ,
         \dataToWriteBuffer[0][2] , \dataToWriteBuffer[0][1] ,
         \dataToWriteBuffer[0][0] , \addressToWriteBuffer[6][7] ,
         \addressToWriteBuffer[6][6] , \addressToWriteBuffer[6][5] ,
         \addressToWriteBuffer[6][4] , \addressToWriteBuffer[6][3] ,
         \addressToWriteBuffer[6][2] , \addressToWriteBuffer[6][1] ,
         \addressToWriteBuffer[6][0] , \addressToWriteBuffer[5][7] ,
         \addressToWriteBuffer[5][6] , \addressToWriteBuffer[5][5] ,
         \addressToWriteBuffer[5][4] , \addressToWriteBuffer[5][3] ,
         \addressToWriteBuffer[5][2] , \addressToWriteBuffer[5][1] ,
         \addressToWriteBuffer[5][0] , \addressToWriteBuffer[4][7] ,
         \addressToWriteBuffer[4][6] , \addressToWriteBuffer[4][5] ,
         \addressToWriteBuffer[4][4] , \addressToWriteBuffer[4][3] ,
         \addressToWriteBuffer[4][2] , \addressToWriteBuffer[4][1] ,
         \addressToWriteBuffer[4][0] , \addressToWriteBuffer[3][7] ,
         \addressToWriteBuffer[3][6] , \addressToWriteBuffer[3][5] ,
         \addressToWriteBuffer[3][4] , \addressToWriteBuffer[3][3] ,
         \addressToWriteBuffer[3][2] , \addressToWriteBuffer[3][1] ,
         \addressToWriteBuffer[3][0] , \addressToWriteBuffer[2][7] ,
         \addressToWriteBuffer[2][6] , \addressToWriteBuffer[2][5] ,
         \addressToWriteBuffer[2][4] , \addressToWriteBuffer[2][3] ,
         \addressToWriteBuffer[2][2] , \addressToWriteBuffer[2][1] ,
         \addressToWriteBuffer[2][0] , \addressToWriteBuffer[1][7] ,
         \addressToWriteBuffer[1][6] , \addressToWriteBuffer[1][5] ,
         \addressToWriteBuffer[1][4] , \addressToWriteBuffer[1][3] ,
         \addressToWriteBuffer[1][2] , \addressToWriteBuffer[1][1] ,
         \addressToWriteBuffer[1][0] , \addressToWriteBuffer[0][7] ,
         \addressToWriteBuffer[0][6] , \addressToWriteBuffer[0][5] ,
         \addressToWriteBuffer[0][4] , \addressToWriteBuffer[0][3] ,
         \addressToWriteBuffer[0][2] , \addressToWriteBuffer[0][1] ,
         \addressToWriteBuffer[0][0] , \requesterAddressBuffer[1][3] ,
         \requesterAddressBuffer[1][2] , \requesterAddressBuffer[1][1] ,
         \requesterAddressBuffer[1][0] , \requesterAddressBuffer[0][3] ,
         \requesterAddressBuffer[0][2] , \requesterAddressBuffer[0][1] ,
         \requesterAddressBuffer[0][0] , \requesterPortBuffer[5][1] ,
         \requesterPortBuffer[5][0] , \requesterPortBuffer[4][1] ,
         \requesterPortBuffer[4][0] , \requesterPortBuffer[3][1] ,
         \requesterPortBuffer[3][0] , \requesterPortBuffer[2][1] ,
         \requesterPortBuffer[2][0] , \requesterPortBuffer[1][1] ,
         \requesterPortBuffer[1][0] , \requesterPortBuffer[0][1] ,
         \requesterPortBuffer[0][0] , \prevRequesterPort_B[0] , prevMemRead_B,
         prevMemRead_A, N5457, N5465, N5473, N5481, n1155, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1214, n1215, n1216, n1217, n1218, n1219, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1272,
         n1273, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808;
  wire   [7:0] isWrite;
  wire   [3:0] prevRequesterAddress_B;
  wire   [1:0] prevRequesterPort_A;
  wire   [3:0] prevRequesterAddress_A;

  EDFFX1TS \readReady_Concatenated_reg[3]  ( .D(N5481), .E(n297), .CK(clk), 
        .Q(readReady_WEST) );
  EDFFX1TS \readReady_Concatenated_reg[2]  ( .D(N5473), .E(n808), .CK(clk), 
        .Q(readReady_EAST) );
  EDFFX1TS \readReady_Concatenated_reg[1]  ( .D(N5465), .E(n442), .CK(clk), 
        .Q(readReady_SOUTH) );
  EDFFX1TS \readReady_Concatenated_reg[0]  ( .D(N5457), .E(n297), .CK(clk), 
        .Q(readReady_NORTH) );
  DFFNSRX1TS \requesterAddressBuffer_reg[1][3]  ( .D(n1347), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressBuffer[1][3] ) );
  DFFNSRX1TS \requesterAddressBuffer_reg[1][2]  ( .D(n1348), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressBuffer[1][2] ) );
  DFFNSRX1TS \requesterAddressBuffer_reg[1][1]  ( .D(n1349), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressBuffer[1][1] ) );
  DFFNSRX1TS \requesterAddressBuffer_reg[1][0]  ( .D(n1350), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressBuffer[1][0] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[0][5]  ( .D(n1262), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[0][5] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[0][4]  ( .D(n1263), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[0][4] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[0][3]  ( .D(n1264), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[0][3] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[0][2]  ( .D(n1265), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[0][2] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[0][1]  ( .D(n1266), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[0][1] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[0][0]  ( .D(n1267), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[0][0] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[0][7]  ( .D(n1339), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[0][7] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[0][6]  ( .D(n1340), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[0][6] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[0][5]  ( .D(n1341), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[0][5] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[0][4]  ( .D(n1342), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[0][4] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[0][3]  ( .D(n1343), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[0][3] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[0][2]  ( .D(n1344), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[0][2] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[0][1]  ( .D(n1345), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[0][1] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[0][0]  ( .D(n1346), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[0][0] ) );
  DFFNSRX1TS \requesterPortBuffer_reg[0][1]  ( .D(n1282), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[0][1] ) );
  DFFNSRX1TS \requesterPortBuffer_reg[0][0]  ( .D(n1363), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[0][0] ) );
  DFFNSRX1TS \requesterAddressBuffer_reg[0][3]  ( .D(n1351), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressBuffer[0][3] ) );
  DFFNSRX1TS \requesterAddressBuffer_reg[0][2]  ( .D(n1352), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressBuffer[0][2] ) );
  DFFNSRX1TS \requesterAddressBuffer_reg[0][1]  ( .D(n1353), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressBuffer[0][1] ) );
  DFFNSRX1TS \requesterAddressBuffer_reg[0][0]  ( .D(n1354), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressBuffer[0][0] ) );
  DFFNSRX1TS \requesterPortBuffer_reg[4][1]  ( .D(n799), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[4][1] ) );
  DFFNSRX1TS \requesterPortBuffer_reg[4][0]  ( .D(n798), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[4][0] ) );
  DFFNSRX1TS \requesterPortBuffer_reg[1][1]  ( .D(n1280), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[1][1] ) );
  DFFNSRX1TS \requesterPortBuffer_reg[1][0]  ( .D(n1281), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[1][0] ) );
  DFFNSRX1TS \isWrite_reg[3]  ( .D(n1216), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(isWrite[3]) );
  DFFNSRX1TS \isWrite_reg[4]  ( .D(n1215), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(isWrite[4]) );
  DFFNSRX1TS \dataToWriteBuffer_reg[4][5]  ( .D(n1238), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[4][5] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[4][4]  ( .D(n1239), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[4][4] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[4][3]  ( .D(n1240), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[4][3] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[4][2]  ( .D(n1241), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[4][2] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[4][1]  ( .D(n1242), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[4][1] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[4][0]  ( .D(n1243), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[4][0] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[4][7]  ( .D(n1307), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[4][7] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[4][6]  ( .D(n1308), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[4][6] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[4][5]  ( .D(n1309), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[4][5] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[4][4]  ( .D(n1310), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[4][4] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[4][3]  ( .D(n1311), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[4][3] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[4][2]  ( .D(n1312), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[4][2] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[4][1]  ( .D(n1313), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[4][1] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[4][0]  ( .D(n1314), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[4][0] ) );
  DFFNSRX1TS \isWrite_reg[2]  ( .D(n1217), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(isWrite[2]) );
  DFFNSRX1TS \dataToWriteBuffer_reg[1][5]  ( .D(n1256), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[1][5] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[1][4]  ( .D(n1257), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[1][4] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[1][3]  ( .D(n1258), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[1][3] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[1][2]  ( .D(n1259), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[1][2] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[1][1]  ( .D(n1260), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[1][1] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[1][0]  ( .D(n1261), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[1][0] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[1][7]  ( .D(n1331), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[1][7] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[1][6]  ( .D(n1332), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[1][6] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[1][5]  ( .D(n1333), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[1][5] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[1][4]  ( .D(n1334), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[1][4] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[1][3]  ( .D(n1335), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[1][3] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[1][2]  ( .D(n1336), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[1][2] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[1][1]  ( .D(n1337), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[1][1] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[1][0]  ( .D(n1338), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[1][0] ) );
  DFFNSRX1TS \requesterPortBuffer_reg[3][0]  ( .D(n1277), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[3][0] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[3][5]  ( .D(n1244), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[3][5] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[3][4]  ( .D(n1245), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[3][4] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[3][3]  ( .D(n1246), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[3][3] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[3][2]  ( .D(n1247), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[3][2] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[3][1]  ( .D(n1248), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[3][1] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[3][0]  ( .D(n1249), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[3][0] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[3][7]  ( .D(n1315), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[3][7] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[3][6]  ( .D(n1316), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[3][6] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[3][5]  ( .D(n1317), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[3][5] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[3][4]  ( .D(n1318), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[3][4] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[3][3]  ( .D(n1319), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[3][3] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[3][2]  ( .D(n1320), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[3][2] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[3][1]  ( .D(n1321), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[3][1] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[3][0]  ( .D(n1322), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[3][0] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[2][5]  ( .D(n1250), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[2][5] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[2][4]  ( .D(n1251), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[2][4] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[2][3]  ( .D(n1252), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[2][3] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[2][2]  ( .D(n1253), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[2][2] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[2][1]  ( .D(n1254), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[2][1] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[2][0]  ( .D(n1255), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[2][0] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[2][7]  ( .D(n1323), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[2][7] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[2][6]  ( .D(n1324), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[2][6] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[2][5]  ( .D(n1325), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[2][5] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[2][4]  ( .D(n1326), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[2][4] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[2][3]  ( .D(n1327), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[2][3] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[2][2]  ( .D(n1328), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[2][2] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[2][1]  ( .D(n1329), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[2][1] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[2][0]  ( .D(n1330), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[2][0] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[5][5]  ( .D(n1232), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[5][5] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[5][4]  ( .D(n1233), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[5][4] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[5][3]  ( .D(n1234), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[5][3] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[5][2]  ( .D(n1235), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[5][2] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[5][1]  ( .D(n1236), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[5][1] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[5][0]  ( .D(n1237), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[5][0] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[5][7]  ( .D(n1299), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[5][7] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[5][6]  ( .D(n1300), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[5][6] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[5][5]  ( .D(n1301), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[5][5] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[5][4]  ( .D(n1302), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[5][4] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[5][3]  ( .D(n1303), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[5][3] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[5][2]  ( .D(n1304), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[5][2] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[5][1]  ( .D(n1305), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[5][1] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[5][0]  ( .D(n1306), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[5][0] ) );
  DFFNSRX1TS \requesterPortBuffer_reg[3][1]  ( .D(n1276), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[3][1] ) );
  DFFNSRX1TS \requesterPortBuffer_reg[2][1]  ( .D(n1278), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[2][1] ) );
  DFFNSRX1TS \requesterPortBuffer_reg[2][0]  ( .D(n1279), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[2][0] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[6][5]  ( .D(n1226), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[6][5] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[6][4]  ( .D(n1227), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[6][4] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[6][3]  ( .D(n1228), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[6][3] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[6][2]  ( .D(n1229), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[6][2] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[6][1]  ( .D(n1230), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[6][1] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[6][0]  ( .D(n1231), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[6][0] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[6][7]  ( .D(n1291), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[6][7] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[6][6]  ( .D(n1292), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[6][6] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[6][5]  ( .D(n1293), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[6][5] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[6][4]  ( .D(n1294), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[6][4] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[6][3]  ( .D(n1295), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[6][3] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[6][2]  ( .D(n1296), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[6][2] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[6][1]  ( .D(n1297), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[6][1] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[6][0]  ( .D(n1298), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[6][0] ) );
  DFFNSRX1TS \isWrite_reg[0]  ( .D(n1219), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(isWrite[0]) );
  DFFNSRX1TS \requesterPortBuffer_reg[5][1]  ( .D(n1272), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[5][1] ) );
  DFFNSRX1TS \requesterPortBuffer_reg[5][0]  ( .D(n1273), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[5][0] ) );
  DFFNSRX1TS \nextEmptyBuffer_reg[0]  ( .D(n1211), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(N882) );
  DFFNSRX1TS prevMemRead_B_reg ( .D(n1204), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(prevMemRead_B) );
  DFFNSRX1TS prevMemRead_A_reg ( .D(n1203), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(prevMemRead_A) );
  DFFNSRX1TS \prevRequesterAddress_A_reg[3]  ( .D(n1205), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_A[3]), .QN(n5) );
  DFFNSRX1TS \prevRequesterAddress_A_reg[2]  ( .D(n1206), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_A[2]), .QN(n6) );
  DFFNSRX1TS \prevRequesterAddress_A_reg[1]  ( .D(n1207), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_A[1]), .QN(n7) );
  DFFNSRX1TS \prevRequesterAddress_A_reg[0]  ( .D(n1208), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_A[0]), .QN(n8) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[3][3]  ( .D(n1171), .CK(clk), 
        .Q(requesterAddressOut_WEST[3]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[3][2]  ( .D(n1170), .CK(clk), 
        .Q(requesterAddressOut_WEST[2]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[3][1]  ( .D(n1169), .CK(clk), 
        .Q(requesterAddressOut_WEST[1]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[2][3]  ( .D(n1167), .CK(clk), 
        .Q(requesterAddressOut_EAST[3]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[2][2]  ( .D(n1166), .CK(clk), 
        .Q(requesterAddressOut_EAST[2]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[2][1]  ( .D(n1165), .CK(clk), 
        .Q(requesterAddressOut_EAST[1]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[1][3]  ( .D(n1163), .CK(clk), 
        .Q(requesterAddressOut_SOUTH[3]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[1][2]  ( .D(n1162), .CK(clk), 
        .Q(requesterAddressOut_SOUTH[2]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[1][1]  ( .D(n1161), .CK(clk), 
        .Q(requesterAddressOut_SOUTH[1]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[3][0]  ( .D(n1168), .CK(clk), 
        .Q(requesterAddressOut_WEST[0]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[2][0]  ( .D(n1164), .CK(clk), 
        .Q(requesterAddressOut_EAST[0]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[1][0]  ( .D(n1160), .CK(clk), 
        .Q(requesterAddressOut_SOUTH[0]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[0][3]  ( .D(n1159), .CK(clk), 
        .Q(requesterAddressOut_NORTH[3]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[0][2]  ( .D(n1158), .CK(clk), 
        .Q(requesterAddressOut_NORTH[2]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[0][1]  ( .D(n1157), .CK(clk), 
        .Q(requesterAddressOut_NORTH[1]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[0][0]  ( .D(n1155), .CK(clk), 
        .Q(requesterAddressOut_NORTH[0]) );
  DFFNSRX1TS memWrite_A_reg ( .D(n1181), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        memWrite_A) );
  DFFNSRX1TS \cacheDataIn_A_reg[5]  ( .D(n1196), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[5]) );
  DFFNSRX1TS \cacheDataIn_A_reg[4]  ( .D(n1197), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[4]) );
  DFFNSRX1TS \cacheDataIn_A_reg[3]  ( .D(n1198), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[3]) );
  DFFNSRX1TS \cacheDataIn_A_reg[2]  ( .D(n1199), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[2]) );
  DFFNSRX1TS \cacheDataIn_A_reg[1]  ( .D(n1200), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[1]) );
  DFFNSRX1TS \cacheDataIn_A_reg[0]  ( .D(n1201), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[0]) );
  DFFNSRX1TS \cacheAddressIn_B_reg[7]  ( .D(n1195), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_B[7]) );
  DFFNSRX1TS \cacheAddressIn_B_reg[6]  ( .D(n1194), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_B[6]) );
  DFFNSRX1TS \cacheAddressIn_B_reg[5]  ( .D(n1193), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_B[5]) );
  DFFNSRX1TS \cacheAddressIn_B_reg[4]  ( .D(n1192), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_B[4]) );
  DFFNSRX1TS \cacheAddressIn_B_reg[3]  ( .D(n1191), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_B[3]) );
  DFFNSRX1TS \cacheAddressIn_B_reg[2]  ( .D(n1190), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_B[2]) );
  DFFNSRX1TS \cacheAddressIn_B_reg[1]  ( .D(n1189), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_B[1]) );
  DFFNSRX1TS \cacheAddressIn_B_reg[0]  ( .D(n1188), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_B[0]) );
  DFFNSRX1TS \cacheDataIn_B_reg[5]  ( .D(n1187), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[5]) );
  DFFNSRX1TS \cacheDataIn_B_reg[4]  ( .D(n1186), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[4]) );
  DFFNSRX1TS \cacheDataIn_B_reg[3]  ( .D(n1185), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[3]) );
  DFFNSRX1TS \cacheDataIn_B_reg[2]  ( .D(n1184), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[2]) );
  DFFNSRX1TS \cacheDataIn_B_reg[1]  ( .D(n1183), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[1]) );
  DFFNSRX1TS \cacheDataIn_B_reg[0]  ( .D(n1182), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[0]) );
  DFFNSRX1TS \cacheAddressIn_A_reg[7]  ( .D(n1180), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_A[7]) );
  DFFNSRX1TS \cacheAddressIn_A_reg[6]  ( .D(n1179), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_A[6]) );
  DFFNSRX1TS \cacheAddressIn_A_reg[5]  ( .D(n1178), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_A[5]) );
  DFFNSRX1TS \cacheAddressIn_A_reg[4]  ( .D(n1177), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_A[4]) );
  DFFNSRX1TS \cacheAddressIn_A_reg[3]  ( .D(n1176), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_A[3]) );
  DFFNSRX1TS \cacheAddressIn_A_reg[2]  ( .D(n1175), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_A[2]) );
  DFFNSRX1TS \cacheAddressIn_A_reg[1]  ( .D(n1174), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_A[1]) );
  DFFNSRX1TS \cacheAddressIn_A_reg[0]  ( .D(n1173), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_A[0]) );
  DFFNSRX1TS \prevRequesterPort_A_reg[0]  ( .D(n1356), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterPort_A[0]), .QN(n795) );
  DFFNSRX1TS \nextEmptyBuffer_reg[2]  ( .D(n1209), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(N884), .QN(n804) );
  DFFNSRX1TS \isWrite_reg[5]  ( .D(n1214), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(isWrite[5]), .QN(n806) );
  DFFNSRX1TS memWrite_B_reg ( .D(n1202), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        memWrite_B), .QN(n807) );
  DFFNSRX1TS \prevRequesterPort_B_reg[1]  ( .D(n1357), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n793), .QN(n792) );
  DFFNSRX1TS \prevRequesterPort_B_reg[0]  ( .D(n1358), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\prevRequesterPort_B[0] ), .QN(n794) );
  DFFNSRX1TS \prevRequesterAddress_B_reg[3]  ( .D(n1359), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_B[3]), .QN(n800) );
  DFFNSRX1TS \prevRequesterAddress_B_reg[2]  ( .D(n1360), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_B[2]), .QN(n801) );
  DFFNSRX1TS \prevRequesterAddress_B_reg[1]  ( .D(n1361), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_B[1]), .QN(n802) );
  DFFNSRX1TS \prevRequesterAddress_B_reg[0]  ( .D(n1362), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_B[0]), .QN(n803) );
  DFFNSRX1TS \nextEmptyBuffer_reg[1]  ( .D(n1210), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(N883), .QN(n796) );
  DFFNSRX1TS \isWrite_reg[1]  ( .D(n1218), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(isWrite[1]), .QN(n805) );
  DFFNSRX1TS \prevRequesterPort_A_reg[1]  ( .D(n1355), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterPort_A[1]), .QN(n797) );
  CLKBUFX2TS U3 ( .A(n660), .Y(n692) );
  CLKBUFX2TS U4 ( .A(n38), .Y(n441) );
  OAI21XLTS U5 ( .A0(n421), .A1(n204), .B0(n456), .Y(n58) );
  CLKBUFX2TS U6 ( .A(n25), .Y(n77) );
  OAI21XLTS U7 ( .A0(n26), .A1(n202), .B0(n196), .Y(n27) );
  NOR2XLTS U8 ( .A(n654), .B(n397), .Y(n39) );
  NOR2XLTS U9 ( .A(n464), .B(n425), .Y(n64) );
  INVX2TS U10 ( .A(n196), .Y(n134) );
  NOR2XLTS U11 ( .A(N882), .B(n581), .Y(n17) );
  NOR3XLTS U12 ( .A(n420), .B(n602), .C(n31), .Y(n642) );
  INVX2TS U13 ( .A(n685), .Y(n770) );
  INVX2TS U14 ( .A(memWrite_NORTH), .Y(n643) );
  INVX2TS U15 ( .A(n424), .Y(n522) );
  NOR2XLTS U16 ( .A(n654), .B(n87), .Y(n88) );
  NOR2XLTS U17 ( .A(n80), .B(n203), .Y(n59) );
  INVX2TS U18 ( .A(n45), .Y(n370) );
  INVX2TS U19 ( .A(n55), .Y(n403) );
  INVX2TS U20 ( .A(n55), .Y(n382) );
  INVX2TS U21 ( .A(n45), .Y(n225) );
  NOR2XLTS U22 ( .A(prevRequesterPort_A[0]), .B(n797), .Y(n418) );
  NAND2X1TS U23 ( .A(n26), .B(n202), .Y(n196) );
  NOR2XLTS U24 ( .A(memRead_EAST), .B(memWrite_EAST), .Y(n25) );
  NOR4XLTS U25 ( .A(n464), .B(n470), .C(n463), .D(n462), .Y(n465) );
  INVX2TS U26 ( .A(n42), .Y(n749) );
  CLKBUFX2TS U27 ( .A(n444), .Y(n447) );
  AO21XLTS U28 ( .A0(n560), .A1(dataIn_NORTH[1]), .B0(n535), .Y(n1236) );
  AO21XLTS U29 ( .A0(n551), .A1(dataIn_NORTH[3]), .B0(n550), .Y(n1234) );
  AO21XLTS U30 ( .A0(n551), .A1(dataIn_NORTH[0]), .B0(n530), .Y(n1237) );
  AO21XLTS U31 ( .A0(n560), .A1(dataIn_NORTH[4]), .B0(n559), .Y(n1233) );
  AO21XLTS U32 ( .A0(cacheAddressIn_NORTH[0]), .A1(n495), .B0(n474), .Y(n1306)
         );
  AO21XLTS U33 ( .A0(n551), .A1(cacheAddressIn_NORTH[5]), .B0(n500), .Y(n1301)
         );
  AO21XLTS U34 ( .A0(n495), .A1(cacheAddressIn_NORTH[4]), .B0(n494), .Y(n1302)
         );
  AO21XLTS U35 ( .A0(n495), .A1(cacheAddressIn_NORTH[3]), .B0(n490), .Y(n1303)
         );
  AO21XLTS U36 ( .A0(n560), .A1(cacheAddressIn_NORTH[2]), .B0(n482), .Y(n1304)
         );
  AO21XLTS U37 ( .A0(n551), .A1(cacheAddressIn_NORTH[1]), .B0(n478), .Y(n1305)
         );
  AO21XLTS U38 ( .A0(n560), .A1(cacheAddressIn_NORTH[6]), .B0(n505), .Y(n1300)
         );
  OAI211XLTS U39 ( .A0(n568), .A1(n504), .B0(n503), .C0(n502), .Y(n505) );
  OAI211XLTS U40 ( .A0(n568), .A1(n477), .B0(n476), .C0(n475), .Y(n478) );
  OAI211XLTS U41 ( .A0(n558), .A1(n481), .B0(n480), .C0(n479), .Y(n482) );
  OAI211XLTS U42 ( .A0(n549), .A1(n489), .B0(n488), .C0(n487), .Y(n490) );
  OAI211XLTS U43 ( .A0(n467), .A1(n499), .B0(n498), .C0(n497), .Y(n500) );
  OAI211XLTS U44 ( .A0(n558), .A1(n557), .B0(n556), .C0(n555), .Y(n559) );
  OAI211XLTS U45 ( .A0(n549), .A1(n548), .B0(n547), .C0(n546), .Y(n550) );
  OAI211XLTS U46 ( .A0(n558), .A1(n534), .B0(n533), .C0(n532), .Y(n535) );
  OAI211XLTS U47 ( .A0(n568), .A1(n529), .B0(n528), .C0(n527), .Y(n530) );
  OAI211XLTS U48 ( .A0(n549), .A1(n493), .B0(n492), .C0(n491), .Y(n494) );
  OAI211XLTS U49 ( .A0(n473), .A1(n467), .B0(n472), .C0(n471), .Y(n474) );
  NAND2BXLTS U50 ( .AN(n461), .B(n469), .Y(n462) );
  NOR3BX1TS U51 ( .AN(n460), .B(n463), .C(n470), .Y(n461) );
  NOR4BX1TS U52 ( .AN(n87), .B(n770), .C(n83), .D(n85), .Y(n84) );
  NAND2BX1TS U53 ( .AN(n466), .B(n469), .Y(n467) );
  NAND2X1TS U54 ( .A(n466), .B(n468), .Y(n463) );
  CLKBUFX2TS U55 ( .A(n732), .Y(n707) );
  CLKBUFX2TS U56 ( .A(n194), .Y(n347) );
  INVX1TS U57 ( .A(n55), .Y(n390) );
  NAND3X1TS U58 ( .A(n587), .B(n513), .C(n58), .Y(n55) );
  NAND3X1TS U59 ( .A(n762), .B(n33), .C(n642), .Y(n619) );
  OAI21X1TS U60 ( .A0(n602), .A1(n198), .B0(n316), .Y(n608) );
  NAND3BX1TS U61 ( .AN(n609), .B(n459), .C(n78), .Y(n513) );
  CLKBUFX2TS U62 ( .A(n601), .Y(n606) );
  INVX2TS U63 ( .A(n4), .Y(n26) );
  OR2X2TS U64 ( .A(n24), .B(n641), .Y(n4) );
  NOR2X1TS U65 ( .A(n747), .B(n440), .Y(n41) );
  INVX1TS U66 ( .A(n3), .Y(n420) );
  CLKAND2X2TS U67 ( .A(n464), .B(N882), .Y(n16) );
  OR2X2TS U68 ( .A(memRead_WEST), .B(n591), .Y(n136) );
  CLKBUFX2TS U69 ( .A(n417), .Y(n769) );
  CLKBUFX2TS U70 ( .A(n418), .Y(n759) );
  INVX1TS U71 ( .A(n424), .Y(n21) );
  NOR2X1TS U72 ( .A(memRead_SOUTH), .B(memWrite_SOUTH), .Y(n424) );
  INVX1TS U73 ( .A(memWrite_SOUTH), .Y(n645) );
  AOI211XLTS U74 ( .A0(n199), .A1(n422), .B0(n642), .C0(n421), .Y(n621) );
  NOR2X1TS U75 ( .A(n23), .B(n522), .Y(n641) );
  AOI211XLTS U76 ( .A0(n19), .A1(n18), .B0(n454), .C0(n453), .Y(n470) );
  NOR2XLTS U77 ( .A(n82), .B(n81), .Y(n459) );
  OAI21XLTS U78 ( .A0(N883), .A1(n22), .B0(N884), .Y(n78) );
  AOI211XLTS U79 ( .A0(n794), .A1(n792), .B0(n770), .C0(n415), .Y(n310) );
  NAND3XLTS U80 ( .A(n592), .B(n524), .C(n303), .Y(n589) );
  INVX2TS U81 ( .A(cacheAddressIn_EAST[5]), .Y(n373) );
  INVX2TS U82 ( .A(cacheAddressIn_EAST[6]), .Y(n377) );
  OAI211XLTS U83 ( .A0(n365), .A1(n360), .B0(n364), .C0(n363), .Y(n1362) );
  OAI211XLTS U84 ( .A0(n351), .A1(n360), .B0(n350), .C0(n349), .Y(n1361) );
  OAI211XLTS U85 ( .A0(n361), .A1(n360), .B0(n359), .C0(n358), .Y(n1360) );
  OAI211XLTS U86 ( .A0(n356), .A1(n360), .B0(n355), .C0(n354), .Y(n1359) );
  OAI21XLTS U87 ( .A0(n425), .A1(n319), .B0(n318), .Y(n1279) );
  OAI211XLTS U88 ( .A0(n344), .A1(n504), .B0(n331), .C0(n330), .Y(n1324) );
  OAI211XLTS U89 ( .A0(n336), .A1(n540), .B0(n324), .C0(n323), .Y(n1253) );
  OAI211XLTS U90 ( .A0(n60), .A1(n548), .B0(n333), .C0(n332), .Y(n1252) );
  NAND3XLTS U91 ( .A(N884), .B(N883), .C(n522), .Y(n453) );
  OAI21XLTS U92 ( .A0(n352), .A1(n37), .B0(n600), .Y(n36) );
  AOI2BB2XLTS U93 ( .B0(n201), .B1(n299), .A0N(n28), .A1N(n201), .Y(n81) );
  NOR2XLTS U94 ( .A(n77), .B(n78), .Y(n458) );
  NAND3XLTS U95 ( .A(n80), .B(n79), .C(n455), .Y(n87) );
  NOR2XLTS U96 ( .A(n302), .B(n203), .Y(n646) );
  CLKAND2X2TS U97 ( .A(n85), .B(n685), .Y(n86) );
  INVX2TS U98 ( .A(cacheAddressIn_EAST[4]), .Y(n142) );
  INVX2TS U99 ( .A(cacheAddressIn_EAST[7]), .Y(n148) );
  NAND2BXLTS U100 ( .AN(n574), .B(n440), .Y(n449) );
  OAI21XLTS U101 ( .A0(n618), .A1(n617), .B0(n615), .Y(n616) );
  AOI211XLTS U102 ( .A0(n606), .A1(n613), .B0(n612), .C0(n611), .Y(n618) );
  NAND3BXLTS U103 ( .AN(n692), .B(n426), .C(n619), .Y(n1356) );
  NAND3BXLTS U104 ( .AN(n715), .B(n429), .C(n619), .Y(n1355) );
  OAI21XLTS U105 ( .A0(n576), .A1(n38), .B0(n575), .Y(n577) );
  OAI21XLTS U106 ( .A0(n601), .A1(n605), .B0(n615), .Y(n604) );
  OAI32X1TS U107 ( .A0(memRead_EAST), .A1(memRead_SOUTH), .A2(n643), .B0(n645), 
        .B1(memRead_EAST), .Y(n594) );
  NAND3XLTS U108 ( .A(n744), .B(n743), .C(n742), .Y(n1173) );
  NAND3XLTS U109 ( .A(n736), .B(n735), .C(n734), .Y(n1174) );
  NAND3XLTS U110 ( .A(n728), .B(n727), .C(n726), .Y(n1175) );
  NAND3XLTS U111 ( .A(n721), .B(n720), .C(n719), .Y(n1176) );
  NAND3XLTS U112 ( .A(n713), .B(n712), .C(n711), .Y(n1177) );
  NAND3XLTS U113 ( .A(n706), .B(n705), .C(n704), .Y(n1178) );
  NAND3XLTS U114 ( .A(n700), .B(n699), .C(n698), .Y(n1179) );
  NAND3XLTS U115 ( .A(n695), .B(n694), .C(n693), .Y(n1180) );
  NAND3XLTS U116 ( .A(n658), .B(n657), .C(n656), .Y(n1201) );
  NAND3XLTS U117 ( .A(n663), .B(n662), .C(n661), .Y(n1200) );
  NAND3XLTS U118 ( .A(n667), .B(n666), .C(n665), .Y(n1199) );
  NAND3XLTS U119 ( .A(n674), .B(n673), .C(n672), .Y(n1198) );
  NAND3XLTS U120 ( .A(n679), .B(n678), .C(n677), .Y(n1197) );
  NAND3XLTS U121 ( .A(n684), .B(n683), .C(n682), .Y(n1196) );
  OAI21XLTS U122 ( .A0(n803), .A1(n313), .B0(n308), .Y(n1155) );
  OAI21XLTS U123 ( .A0(n802), .A1(n313), .B0(n312), .Y(n1157) );
  OAI21XLTS U124 ( .A0(n801), .A1(n313), .B0(n307), .Y(n1158) );
  OAI21XLTS U125 ( .A0(n800), .A1(n313), .B0(n309), .Y(n1159) );
  NAND3XLTS U126 ( .A(n625), .B(n624), .C(n623), .Y(n1208) );
  NAND3XLTS U127 ( .A(n628), .B(n627), .C(n626), .Y(n1207) );
  NAND3XLTS U128 ( .A(n632), .B(n631), .C(n630), .Y(n1206) );
  NAND3XLTS U129 ( .A(n639), .B(n638), .C(n637), .Y(n1205) );
  NAND3XLTS U130 ( .A(n589), .B(n526), .C(n525), .Y(n1273) );
  AO21XLTS U131 ( .A0(n465), .A1(cacheAddressIn_NORTH[7]), .B0(n510), .Y(n1299) );
  OAI211XLTS U132 ( .A0(n549), .A1(n509), .B0(n508), .C0(n507), .Y(n510) );
  AO21XLTS U133 ( .A0(n465), .A1(dataIn_NORTH[2]), .B0(n541), .Y(n1235) );
  OAI211XLTS U134 ( .A0(n558), .A1(n540), .B0(n539), .C0(n538), .Y(n541) );
  AO21XLTS U135 ( .A0(n465), .A1(dataIn_NORTH[5]), .B0(n569), .Y(n1232) );
  OAI211XLTS U136 ( .A0(n568), .A1(n567), .B0(n566), .C0(n565), .Y(n569) );
  OAI211XLTS U137 ( .A0(n341), .A1(n473), .B0(n327), .C0(n326), .Y(n1330) );
  OAI211XLTS U138 ( .A0(n341), .A1(n493), .B0(n340), .C0(n339), .Y(n1326) );
  OAI211XLTS U139 ( .A0(n60), .A1(n509), .B0(n321), .C0(n320), .Y(n1323) );
  OAI211XLTS U140 ( .A0(n344), .A1(n534), .B0(n343), .C0(n342), .Y(n1254) );
  OAI211XLTS U141 ( .A0(n336), .A1(n567), .B0(n335), .C0(n334), .Y(n1250) );
  OAI211XLTS U142 ( .A0(n389), .A1(n388), .B0(n387), .C0(n386), .Y(n1337) );
  OAI211XLTS U143 ( .A0(n369), .A1(n388), .B0(n368), .C0(n367), .Y(n1335) );
  OAI211XLTS U144 ( .A0(n373), .A1(n395), .B0(n372), .C0(n371), .Y(n1333) );
  OAI211XLTS U145 ( .A0(n377), .A1(n401), .B0(n376), .C0(n375), .Y(n1332) );
  OAI211XLTS U146 ( .A0(n381), .A1(n409), .B0(n380), .C0(n379), .Y(n1261) );
  OAI211XLTS U147 ( .A0(n410), .A1(n409), .B0(n408), .C0(n407), .Y(n1259) );
  OAI211XLTS U148 ( .A0(n402), .A1(n401), .B0(n400), .C0(n399), .Y(n1258) );
  OAI211XLTS U149 ( .A0(n396), .A1(n395), .B0(n394), .C0(n393), .Y(n1257) );
  AO21XLTS U150 ( .A0(n516), .A1(\requesterPortBuffer[1][0] ), .B0(n512), .Y(
        n1281) );
  AO21XLTS U151 ( .A0(n516), .A1(\requesterPortBuffer[1][1] ), .B0(n515), .Y(
        n1280) );
  AOI31XLTS U152 ( .A0(n514), .A1(n513), .A2(n441), .B0(n447), .Y(n515) );
  AO22XLTS U153 ( .A0(n775), .A1(prevMemRead_A), .B0(n769), .B1(prevMemRead_B), 
        .Y(N5465) );
  AO22XLTS U154 ( .A0(n759), .A1(prevMemRead_A), .B0(n764), .B1(prevMemRead_B), 
        .Y(N5473) );
  NOR2XLTS U155 ( .A(n28), .B(n27), .Y(n29) );
  OA21XLTS U156 ( .A0(n77), .A1(n641), .B0(n219), .Y(n3) );
  NOR2BX1TS U157 ( .AN(n39), .B(n441), .Y(n40) );
  AND2X2TS U158 ( .A(n443), .B(n653), .Y(n9) );
  NOR3BX1TS U159 ( .AN(n641), .B(n25), .C(n427), .Y(n428) );
  INVX2TS U160 ( .A(n219), .Y(n22) );
  OAI211XLTS U161 ( .A0(n581), .A1(n608), .B0(n808), .C0(n440), .Y(n194) );
  NOR2BX1TS U162 ( .AN(n621), .B(n620), .Y(n622) );
  NOR2X1TS U163 ( .A(memRead_NORTH), .B(memWrite_NORTH), .Y(n19) );
  OR3X1TS U164 ( .A(n792), .B(n794), .C(n746), .Y(n10) );
  OR2X1TS U165 ( .A(n795), .B(n797), .Y(n11) );
  NOR3XLTS U166 ( .A(n416), .B(n775), .C(n794), .Y(n417) );
  OAI21XLTS U167 ( .A0(N882), .A1(n33), .B0(n314), .Y(n18) );
  INVX2TS U168 ( .A(n600), .Y(n601) );
  NAND2X1TS U169 ( .A(n796), .B(n804), .Y(n14) );
  INVX2TS U170 ( .A(n804), .Y(n12) );
  NOR2XLTS U171 ( .A(prevRequesterPort_A[1]), .B(n795), .Y(n13) );
  INVX2TS U185 ( .A(dataIn_EAST[1]), .Y(n152) );
  INVX2TS U186 ( .A(n14), .Y(n137) );
  INVX2TS U187 ( .A(n137), .Y(n15) );
  INVX2TS U188 ( .A(n15), .Y(n464) );
  INVX2TS U189 ( .A(n16), .Y(n314) );
  NAND2X1TS U190 ( .A(n796), .B(n314), .Y(n600) );
  INVX2TS U191 ( .A(n137), .Y(n581) );
  INVX2TS U192 ( .A(n17), .Y(n423) );
  INVX2TS U193 ( .A(n423), .Y(n33) );
  INVX2TS U194 ( .A(n18), .Y(n35) );
  INVX2TS U195 ( .A(n35), .Y(n28) );
  INVX2TS U196 ( .A(n19), .Y(n20) );
  INVX2TS U197 ( .A(n20), .Y(n199) );
  INVX2TS U198 ( .A(n199), .Y(n23) );
  NAND2X1TS U199 ( .A(n23), .B(n21), .Y(n219) );
  INVX2TS U200 ( .A(n22), .Y(n34) );
  INVX2TS U201 ( .A(n34), .Y(n24) );
  INVX2TS U202 ( .A(n77), .Y(n202) );
  INVX2TS U203 ( .A(n27), .Y(n31) );
  INVX2TS U204 ( .A(n34), .Y(n352) );
  NAND2X1TS U205 ( .A(n352), .B(n202), .Y(n609) );
  OAI22X1TS U206 ( .A0(n29), .A1(n420), .B0(n609), .B1(n28), .Y(n30) );
  XOR2X1TS U207 ( .A(n600), .B(n30), .Y(n317) );
  INVX2TS U208 ( .A(n31), .Y(n198) );
  XNOR2X1TS U209 ( .A(n198), .B(n28), .Y(n79) );
  NOR2X1TS U210 ( .A(n317), .B(n79), .Y(n457) );
  INVX2TS U211 ( .A(memWrite_WEST), .Y(n576) );
  INVX2TS U212 ( .A(n576), .Y(n591) );
  INVX2TS U213 ( .A(n136), .Y(n610) );
  INVX2TS U214 ( .A(n136), .Y(n197) );
  INVX2TS U215 ( .A(n197), .Y(n456) );
  INVX2TS U216 ( .A(n423), .Y(n687) );
  INVX2TS U217 ( .A(n687), .Y(n32) );
  INVX2TS U218 ( .A(n32), .Y(n315) );
  INVX2TS U219 ( .A(n315), .Y(n421) );
  AOI21X1TS U220 ( .A0(n457), .A1(n456), .B0(n421), .Y(n574) );
  INVX2TS U221 ( .A(reset), .Y(n297) );
  CLKBUFX2TS U222 ( .A(n297), .Y(n42) );
  CLKBUFX2TS U223 ( .A(n42), .Y(n469) );
  INVX2TS U224 ( .A(n469), .Y(n654) );
  CLKBUFX2TS U225 ( .A(n297), .Y(n306) );
  CLKBUFX2TS U226 ( .A(n306), .Y(n442) );
  NAND2X1TS U227 ( .A(n442), .B(n33), .Y(n203) );
  INVX2TS U228 ( .A(n203), .Y(n413) );
  CLKBUFX2TS U229 ( .A(n413), .Y(n269) );
  CLKBUFX2TS U230 ( .A(n269), .Y(n241) );
  CLKBUFX2TS U231 ( .A(n241), .Y(n243) );
  CLKBUFX2TS U232 ( .A(n243), .Y(n587) );
  INVX2TS U233 ( .A(n4), .Y(n201) );
  INVX2TS U234 ( .A(n35), .Y(n299) );
  NOR2BX1TS U235 ( .AN(n201), .B(n299), .Y(n37) );
  OAI31X1TS U236 ( .A0(n24), .A1(n600), .A2(n37), .B0(n36), .Y(n82) );
  INVX2TS U237 ( .A(n3), .Y(n204) );
  INVX2TS U238 ( .A(n55), .Y(n397) );
  CLKAND2X2TS U239 ( .A(n574), .B(n39), .Y(n50) );
  INVX2TS U240 ( .A(n50), .Y(n401) );
  INVX2TS U241 ( .A(dataIn_WEST[1]), .Y(n534) );
  INVX2TS U242 ( .A(n534), .Y(n659) );
  NAND2X1TS U243 ( .A(n457), .B(n315), .Y(n38) );
  INVX2TS U244 ( .A(n40), .Y(n366) );
  AOI22X1TS U245 ( .A0(n659), .A1(n40), .B0(n382), .B1(
        \dataToWriteBuffer[1][1] ), .Y(n44) );
  CLKBUFX2TS U246 ( .A(n42), .Y(n685) );
  INVX2TS U247 ( .A(n685), .Y(n747) );
  INVX2TS U248 ( .A(n16), .Y(n440) );
  INVX2TS U249 ( .A(n41), .Y(n45) );
  INVX2TS U250 ( .A(n45), .Y(n406) );
  CLKBUFX2TS U251 ( .A(n42), .Y(n443) );
  INVX2TS U252 ( .A(n443), .Y(n425) );
  CLKBUFX2TS U253 ( .A(n64), .Y(n245) );
  CLKBUFX2TS U254 ( .A(n245), .Y(n398) );
  AOI22X1TS U255 ( .A0(n406), .A1(\dataToWriteBuffer[2][1] ), .B0(n398), .B1(
        \dataToWriteBuffer[3][1] ), .Y(n43) );
  OAI211XLTS U256 ( .A0(n152), .A1(n401), .B0(n44), .C0(n43), .Y(n1260) );
  INVX2TS U257 ( .A(cacheAddressIn_EAST[0]), .Y(n168) );
  INVX2TS U258 ( .A(n50), .Y(n409) );
  INVX2TS U259 ( .A(cacheAddressIn_WEST[0]), .Y(n473) );
  INVX2TS U260 ( .A(n473), .Y(n739) );
  INVX2TS U261 ( .A(n366), .Y(n404) );
  AOI22X1TS U262 ( .A0(n739), .A1(n404), .B0(n390), .B1(
        \addressToWriteBuffer[1][0] ), .Y(n47) );
  INVX2TS U263 ( .A(n45), .Y(n61) );
  CLKBUFX2TS U264 ( .A(n61), .Y(n271) );
  CLKBUFX2TS U265 ( .A(n271), .Y(n573) );
  CLKBUFX2TS U266 ( .A(n64), .Y(n145) );
  CLKBUFX2TS U267 ( .A(n145), .Y(n436) );
  CLKBUFX2TS U268 ( .A(n436), .Y(n253) );
  CLKBUFX2TS U269 ( .A(n253), .Y(n70) );
  CLKBUFX2TS U270 ( .A(n70), .Y(n337) );
  AOI22X1TS U271 ( .A0(n573), .A1(\addressToWriteBuffer[2][0] ), .B0(n337), 
        .B1(\addressToWriteBuffer[3][0] ), .Y(n46) );
  OAI211XLTS U272 ( .A0(n168), .A1(n409), .B0(n47), .C0(n46), .Y(n1338) );
  INVX2TS U273 ( .A(dataIn_EAST[5]), .Y(n173) );
  INVX2TS U274 ( .A(n50), .Y(n388) );
  INVX2TS U275 ( .A(dataIn_WEST[5]), .Y(n567) );
  INVX2TS U276 ( .A(n567), .Y(n680) );
  INVX2TS U277 ( .A(n366), .Y(n391) );
  AOI22X1TS U278 ( .A0(n680), .A1(n391), .B0(n382), .B1(
        \dataToWriteBuffer[1][5] ), .Y(n49) );
  CLKBUFX2TS U279 ( .A(n70), .Y(n405) );
  AOI22X1TS U280 ( .A0(n41), .A1(\dataToWriteBuffer[2][5] ), .B0(n405), .B1(
        \dataToWriteBuffer[3][5] ), .Y(n48) );
  OAI211XLTS U281 ( .A0(n173), .A1(n388), .B0(n49), .C0(n48), .Y(n1256) );
  INVX2TS U282 ( .A(n50), .Y(n395) );
  INVX2TS U283 ( .A(cacheAddressIn_WEST[7]), .Y(n509) );
  INVX2TS U284 ( .A(n509), .Y(n691) );
  AOI22X1TS U285 ( .A0(n691), .A1(n404), .B0(n397), .B1(
        \addressToWriteBuffer[1][7] ), .Y(n52) );
  CLKBUFX2TS U286 ( .A(n64), .Y(n346) );
  CLKBUFX2TS U287 ( .A(n346), .Y(n384) );
  AOI22X1TS U288 ( .A0(n41), .A1(\addressToWriteBuffer[2][7] ), .B0(n384), 
        .B1(\addressToWriteBuffer[3][7] ), .Y(n51) );
  OAI211XLTS U289 ( .A0(n148), .A1(n395), .B0(n52), .C0(n51), .Y(n1331) );
  INVX2TS U290 ( .A(cacheAddressIn_WEST[4]), .Y(n493) );
  INVX2TS U291 ( .A(n493), .Y(n709) );
  AOI22X1TS U292 ( .A0(n709), .A1(n391), .B0(n390), .B1(
        \addressToWriteBuffer[1][4] ), .Y(n54) );
  CLKBUFX2TS U293 ( .A(n70), .Y(n374) );
  AOI22X1TS U294 ( .A0(n370), .A1(\addressToWriteBuffer[2][4] ), .B0(n374), 
        .B1(\addressToWriteBuffer[3][4] ), .Y(n53) );
  OAI211XLTS U295 ( .A0(n142), .A1(n401), .B0(n54), .C0(n53), .Y(n1334) );
  INVX2TS U296 ( .A(cacheAddressIn_EAST[2]), .Y(n161) );
  INVX2TS U297 ( .A(cacheAddressIn_WEST[2]), .Y(n481) );
  INVX2TS U298 ( .A(n481), .Y(n724) );
  AOI22X1TS U299 ( .A0(n724), .A1(n40), .B0(n403), .B1(
        \addressToWriteBuffer[1][2] ), .Y(n57) );
  CLKBUFX2TS U300 ( .A(n61), .Y(n385) );
  AOI22X1TS U301 ( .A0(n385), .A1(\addressToWriteBuffer[2][2] ), .B0(n384), 
        .B1(\addressToWriteBuffer[3][2] ), .Y(n56) );
  OAI211XLTS U302 ( .A0(n161), .A1(n409), .B0(n57), .C0(n56), .Y(n1336) );
  NOR2BX1TS U303 ( .AN(n317), .B(n58), .Y(n80) );
  INVX2TS U304 ( .A(n59), .Y(n325) );
  INVX2TS U305 ( .A(n325), .Y(n517) );
  NAND3BX1TS U306 ( .AN(n517), .B(n315), .C(n443), .Y(n60) );
  INVX2TS U307 ( .A(n60), .Y(n69) );
  INVX2TS U308 ( .A(n69), .Y(n341) );
  INVX2TS U309 ( .A(dataIn_WEST[0]), .Y(n529) );
  CLKBUFX2TS U310 ( .A(n61), .Y(n545) );
  CLKBUFX2TS U311 ( .A(n545), .Y(n437) );
  AOI22X1TS U312 ( .A0(\dataToWriteBuffer[3][0] ), .A1(n437), .B0(n405), .B1(
        \dataToWriteBuffer[4][0] ), .Y(n63) );
  INVX2TS U313 ( .A(n325), .Y(n322) );
  NAND2X1TS U314 ( .A(\dataToWriteBuffer[2][0] ), .B(n322), .Y(n62) );
  OAI211XLTS U315 ( .A0(n341), .A1(n529), .B0(n63), .C0(n62), .Y(n1255) );
  INVX2TS U316 ( .A(n69), .Y(n344) );
  CLKBUFX2TS U317 ( .A(n545), .Y(n275) );
  CLKBUFX2TS U318 ( .A(n275), .Y(n328) );
  CLKBUFX2TS U319 ( .A(n64), .Y(n518) );
  AOI22X1TS U320 ( .A0(\addressToWriteBuffer[3][2] ), .A1(n328), .B0(n518), 
        .B1(\addressToWriteBuffer[4][2] ), .Y(n66) );
  INVX2TS U321 ( .A(n325), .Y(n329) );
  NAND2X1TS U322 ( .A(\addressToWriteBuffer[2][2] ), .B(n329), .Y(n65) );
  OAI211XLTS U323 ( .A0(n344), .A1(n481), .B0(n66), .C0(n65), .Y(n1328) );
  INVX2TS U324 ( .A(cacheAddressIn_WEST[3]), .Y(n489) );
  CLKBUFX2TS U325 ( .A(n275), .Y(n519) );
  AOI22X1TS U326 ( .A0(\addressToWriteBuffer[3][3] ), .A1(n519), .B0(n337), 
        .B1(\addressToWriteBuffer[4][3] ), .Y(n68) );
  NAND2X1TS U327 ( .A(\addressToWriteBuffer[2][3] ), .B(n517), .Y(n67) );
  OAI211XLTS U328 ( .A0(n336), .A1(n489), .B0(n68), .C0(n67), .Y(n1327) );
  INVX2TS U329 ( .A(n69), .Y(n336) );
  INVX2TS U330 ( .A(cacheAddressIn_WEST[1]), .Y(n477) );
  CLKBUFX2TS U331 ( .A(n70), .Y(n378) );
  AOI22X1TS U332 ( .A0(\addressToWriteBuffer[3][1] ), .A1(n519), .B0(n378), 
        .B1(\addressToWriteBuffer[4][1] ), .Y(n72) );
  NAND2X1TS U333 ( .A(\addressToWriteBuffer[2][1] ), .B(n582), .Y(n71) );
  OAI211XLTS U334 ( .A0(n336), .A1(n477), .B0(n72), .C0(n71), .Y(n1329) );
  INVX2TS U335 ( .A(cacheAddressIn_WEST[5]), .Y(n499) );
  AOI22X1TS U336 ( .A0(\addressToWriteBuffer[3][5] ), .A1(n519), .B0(n337), 
        .B1(\addressToWriteBuffer[4][5] ), .Y(n74) );
  NAND2X1TS U337 ( .A(\addressToWriteBuffer[2][5] ), .B(n329), .Y(n73) );
  OAI211XLTS U338 ( .A0(n341), .A1(n499), .B0(n74), .C0(n73), .Y(n1325) );
  INVX2TS U339 ( .A(dataIn_WEST[4]), .Y(n557) );
  CLKBUFX2TS U340 ( .A(n275), .Y(n506) );
  CLKBUFX2TS U341 ( .A(n506), .Y(n338) );
  CLKBUFX2TS U342 ( .A(n346), .Y(n392) );
  AOI22X1TS U343 ( .A0(\dataToWriteBuffer[3][4] ), .A1(n338), .B0(n392), .B1(
        \dataToWriteBuffer[4][4] ), .Y(n76) );
  NAND2X1TS U344 ( .A(\dataToWriteBuffer[2][4] ), .B(n322), .Y(n75) );
  OAI211XLTS U345 ( .A0(n344), .A1(n557), .B0(n76), .C0(n75), .Y(n1251) );
  CLKBUFX2TS U346 ( .A(n306), .Y(n762) );
  AND4X1TS U347 ( .A(n458), .B(n82), .C(n81), .D(n762), .Y(n95) );
  INVX2TS U348 ( .A(n95), .Y(n127) );
  INVX2TS U349 ( .A(n204), .Y(n316) );
  AOI21X1TS U350 ( .A0(n316), .A1(n796), .B0(n804), .Y(n455) );
  AND3X1TS U351 ( .A(n458), .B(n82), .C(n81), .Y(n83) );
  NOR2XLTS U352 ( .A(n19), .B(n299), .Y(n454) );
  NOR2BX1TS U353 ( .AN(n454), .B(n453), .Y(n85) );
  INVX2TS U354 ( .A(n84), .Y(n102) );
  INVX2TS U355 ( .A(n102), .Y(n123) );
  INVX2TS U356 ( .A(n86), .Y(n107) );
  AOI22X1TS U357 ( .A0(\dataToWriteBuffer[6][1] ), .A1(n123), .B0(
        dataIn_SOUTH[1]), .B1(n128), .Y(n90) );
  INVX2TS U358 ( .A(n88), .Y(n108) );
  INVX2TS U359 ( .A(n108), .Y(n118) );
  NAND2X1TS U360 ( .A(n659), .B(n118), .Y(n89) );
  OAI211XLTS U361 ( .A0(n127), .A1(n152), .B0(n90), .C0(n89), .Y(n1230) );
  INVX2TS U362 ( .A(n95), .Y(n133) );
  INVX2TS U363 ( .A(cacheAddressIn_EAST[1]), .Y(n389) );
  INVX2TS U364 ( .A(n107), .Y(n114) );
  AOI22X1TS U365 ( .A0(\addressToWriteBuffer[6][1] ), .A1(n123), .B0(
        cacheAddressIn_SOUTH[1]), .B1(n114), .Y(n92) );
  INVX2TS U366 ( .A(n477), .Y(n733) );
  INVX2TS U367 ( .A(n108), .Y(n130) );
  NAND2X1TS U368 ( .A(n733), .B(n130), .Y(n91) );
  OAI211XLTS U369 ( .A0(n133), .A1(n389), .B0(n92), .C0(n91), .Y(n1297) );
  INVX2TS U370 ( .A(n95), .Y(n117) );
  INVX2TS U371 ( .A(n102), .Y(n111) );
  AOI22X1TS U372 ( .A0(\addressToWriteBuffer[6][0] ), .A1(n111), .B0(
        cacheAddressIn_SOUTH[0]), .B1(n114), .Y(n94) );
  NAND2X1TS U373 ( .A(n739), .B(n130), .Y(n93) );
  OAI211XLTS U374 ( .A0(n117), .A1(n168), .B0(n94), .C0(n93), .Y(n1298) );
  INVX2TS U375 ( .A(n95), .Y(n121) );
  INVX2TS U376 ( .A(dataIn_EAST[4]), .Y(n396) );
  INVX2TS U377 ( .A(n107), .Y(n128) );
  AOI22X1TS U378 ( .A0(\dataToWriteBuffer[6][4] ), .A1(n111), .B0(
        dataIn_SOUTH[4]), .B1(n128), .Y(n97) );
  INVX2TS U379 ( .A(n557), .Y(n676) );
  NAND2X1TS U380 ( .A(n676), .B(n118), .Y(n96) );
  OAI211XLTS U381 ( .A0(n121), .A1(n396), .B0(n97), .C0(n96), .Y(n1227) );
  AOI22X1TS U382 ( .A0(\addressToWriteBuffer[6][4] ), .A1(n111), .B0(
        cacheAddressIn_SOUTH[4]), .B1(n114), .Y(n99) );
  INVX2TS U383 ( .A(n108), .Y(n124) );
  NAND2X1TS U384 ( .A(n709), .B(n124), .Y(n98) );
  OAI211XLTS U385 ( .A0(n127), .A1(n142), .B0(n99), .C0(n98), .Y(n1294) );
  INVX2TS U386 ( .A(n102), .Y(n129) );
  AOI22X1TS U387 ( .A0(\addressToWriteBuffer[6][7] ), .A1(n129), .B0(
        cacheAddressIn_SOUTH[7]), .B1(n86), .Y(n101) );
  NAND2X1TS U388 ( .A(n691), .B(n124), .Y(n100) );
  OAI211XLTS U389 ( .A0(n133), .A1(n148), .B0(n101), .C0(n100), .Y(n1291) );
  AOI22X1TS U390 ( .A0(\addressToWriteBuffer[6][2] ), .A1(n129), .B0(
        cacheAddressIn_SOUTH[2]), .B1(n86), .Y(n104) );
  NAND2X1TS U391 ( .A(n724), .B(n130), .Y(n103) );
  OAI211XLTS U392 ( .A0(n117), .A1(n161), .B0(n104), .C0(n103), .Y(n1296) );
  INVX2TS U393 ( .A(dataIn_EAST[2]), .Y(n410) );
  AOI22X1TS U394 ( .A0(\dataToWriteBuffer[6][2] ), .A1(n84), .B0(
        dataIn_SOUTH[2]), .B1(n128), .Y(n106) );
  INVX2TS U395 ( .A(dataIn_WEST[2]), .Y(n540) );
  INVX2TS U396 ( .A(n540), .Y(n664) );
  NAND2X1TS U397 ( .A(n664), .B(n124), .Y(n105) );
  OAI211XLTS U398 ( .A0(n121), .A1(n410), .B0(n106), .C0(n105), .Y(n1229) );
  INVX2TS U399 ( .A(dataIn_EAST[3]), .Y(n402) );
  INVX2TS U400 ( .A(n107), .Y(n122) );
  AOI22X1TS U401 ( .A0(\dataToWriteBuffer[6][3] ), .A1(n129), .B0(
        dataIn_SOUTH[3]), .B1(n122), .Y(n110) );
  INVX2TS U402 ( .A(dataIn_WEST[3]), .Y(n548) );
  INVX2TS U403 ( .A(n548), .Y(n670) );
  NAND2X1TS U404 ( .A(n670), .B(n118), .Y(n109) );
  OAI211XLTS U405 ( .A0(n127), .A1(n402), .B0(n110), .C0(n109), .Y(n1228) );
  INVX2TS U406 ( .A(dataIn_EAST[0]), .Y(n381) );
  AOI22X1TS U407 ( .A0(\dataToWriteBuffer[6][0] ), .A1(n111), .B0(
        dataIn_SOUTH[0]), .B1(n122), .Y(n113) );
  INVX2TS U408 ( .A(n529), .Y(n655) );
  NAND2X1TS U409 ( .A(n655), .B(n88), .Y(n112) );
  OAI211XLTS U410 ( .A0(n133), .A1(n381), .B0(n113), .C0(n112), .Y(n1231) );
  AOI22X1TS U411 ( .A0(\addressToWriteBuffer[6][5] ), .A1(n123), .B0(
        cacheAddressIn_SOUTH[5]), .B1(n114), .Y(n116) );
  INVX2TS U412 ( .A(n499), .Y(n702) );
  NAND2X1TS U413 ( .A(n702), .B(n88), .Y(n115) );
  OAI211XLTS U414 ( .A0(n117), .A1(n373), .B0(n116), .C0(n115), .Y(n1293) );
  AOI22X1TS U415 ( .A0(\addressToWriteBuffer[6][6] ), .A1(n84), .B0(
        cacheAddressIn_SOUTH[6]), .B1(n122), .Y(n120) );
  INVX2TS U416 ( .A(cacheAddressIn_WEST[6]), .Y(n504) );
  INVX2TS U417 ( .A(n504), .Y(n697) );
  NAND2X1TS U418 ( .A(n697), .B(n118), .Y(n119) );
  OAI211XLTS U419 ( .A0(n121), .A1(n377), .B0(n120), .C0(n119), .Y(n1292) );
  AOI22X1TS U420 ( .A0(\dataToWriteBuffer[6][5] ), .A1(n123), .B0(
        dataIn_SOUTH[5]), .B1(n122), .Y(n126) );
  NAND2X1TS U421 ( .A(n680), .B(n124), .Y(n125) );
  OAI211XLTS U422 ( .A0(n127), .A1(n173), .B0(n126), .C0(n125), .Y(n1226) );
  INVX2TS U423 ( .A(cacheAddressIn_EAST[3]), .Y(n369) );
  AOI22X1TS U424 ( .A0(\addressToWriteBuffer[6][3] ), .A1(n129), .B0(
        cacheAddressIn_SOUTH[3]), .B1(n128), .Y(n132) );
  INVX2TS U425 ( .A(n489), .Y(n717) );
  NAND2X1TS U426 ( .A(n717), .B(n130), .Y(n131) );
  OAI211XLTS U427 ( .A0(n133), .A1(n369), .B0(n132), .C0(n131), .Y(n1295) );
  INVX2TS U428 ( .A(n196), .Y(n135) );
  CLKBUFX2TS U429 ( .A(n269), .Y(n430) );
  CLKBUFX2TS U430 ( .A(n430), .Y(n282) );
  CLKBUFX2TS U431 ( .A(n282), .Y(n411) );
  CLKAND2X2TS U432 ( .A(n135), .B(n411), .Y(n149) );
  INVX2TS U433 ( .A(n149), .Y(n187) );
  OR2X1TS U434 ( .A(n219), .B(n203), .Y(n162) );
  INVX2TS U435 ( .A(n162), .Y(n183) );
  CLKBUFX2TS U436 ( .A(n145), .Y(n220) );
  CLKBUFX2TS U437 ( .A(n220), .Y(n158) );
  AOI22X1TS U438 ( .A0(cacheAddressIn_SOUTH[4]), .A1(n183), .B0(
        \addressToWriteBuffer[1][4] ), .B1(n158), .Y(n141) );
  INVX2TS U439 ( .A(n136), .Y(n602) );
  NOR3XLTS U440 ( .A(n204), .B(n198), .C(n602), .Y(n200) );
  NAND2X1TS U441 ( .A(n411), .B(n200), .Y(n217) );
  CLKBUFX2TS U442 ( .A(n217), .Y(n155) );
  INVX2TS U443 ( .A(n155), .Y(n170) );
  AOI21X1TS U444 ( .A0(n687), .A1(n608), .B0(n15), .Y(n138) );
  NAND2X1TS U445 ( .A(n442), .B(n138), .Y(n649) );
  INVX2TS U446 ( .A(n649), .Y(n139) );
  INVX2TS U447 ( .A(n139), .Y(n163) );
  INVX2TS U448 ( .A(n163), .Y(n189) );
  AOI22X1TS U449 ( .A0(n709), .A1(n170), .B0(n189), .B1(cacheAddressIn_B[4]), 
        .Y(n140) );
  OAI211XLTS U450 ( .A0(n142), .A1(n187), .B0(n141), .C0(n140), .Y(n1192) );
  INVX2TS U451 ( .A(n149), .Y(n192) );
  INVX2TS U452 ( .A(n162), .Y(n174) );
  AOI22X1TS U453 ( .A0(cacheAddressIn_SOUTH[6]), .A1(n174), .B0(
        \addressToWriteBuffer[1][6] ), .B1(n158), .Y(n144) );
  INVX2TS U454 ( .A(n155), .Y(n362) );
  INVX2TS U455 ( .A(n217), .Y(n353) );
  AOI22X1TS U456 ( .A0(n697), .A1(n353), .B0(n189), .B1(cacheAddressIn_B[6]), 
        .Y(n143) );
  OAI211XLTS U457 ( .A0(n377), .A1(n192), .B0(n144), .C0(n143), .Y(n1194) );
  INVX2TS U458 ( .A(n149), .Y(n177) );
  INVX2TS U459 ( .A(n162), .Y(n169) );
  CLKBUFX2TS U460 ( .A(n145), .Y(n178) );
  AOI22X1TS U461 ( .A0(cacheAddressIn_SOUTH[7]), .A1(n169), .B0(
        \addressToWriteBuffer[1][7] ), .B1(n178), .Y(n147) );
  AOI22X1TS U462 ( .A0(n691), .A1(n362), .B0(n189), .B1(cacheAddressIn_B[7]), 
        .Y(n146) );
  OAI211XLTS U463 ( .A0(n148), .A1(n177), .B0(n147), .C0(n146), .Y(n1195) );
  INVX2TS U464 ( .A(n149), .Y(n182) );
  AOI22X1TS U465 ( .A0(dataIn_SOUTH[1]), .A1(n169), .B0(
        \dataToWriteBuffer[1][1] ), .B1(n158), .Y(n151) );
  INVX2TS U466 ( .A(n155), .Y(n348) );
  INVX2TS U467 ( .A(n163), .Y(n179) );
  AOI22X1TS U468 ( .A0(n659), .A1(n348), .B0(n179), .B1(cacheDataIn_B[1]), .Y(
        n150) );
  OAI211XLTS U469 ( .A0(n152), .A1(n182), .B0(n151), .C0(n150), .Y(n1183) );
  CLKBUFX2TS U470 ( .A(n220), .Y(n303) );
  AOI22X1TS U471 ( .A0(dataIn_SOUTH[0]), .A1(n174), .B0(
        \dataToWriteBuffer[1][0] ), .B1(n303), .Y(n154) );
  INVX2TS U472 ( .A(n163), .Y(n184) );
  AOI22X1TS U473 ( .A0(n655), .A1(n357), .B0(n184), .B1(cacheDataIn_B[0]), .Y(
        n153) );
  OAI211XLTS U474 ( .A0(n381), .A1(n187), .B0(n154), .C0(n153), .Y(n1182) );
  CLKBUFX2TS U475 ( .A(n220), .Y(n570) );
  AOI22X1TS U476 ( .A0(cacheAddressIn_SOUTH[3]), .A1(n169), .B0(
        \addressToWriteBuffer[1][3] ), .B1(n570), .Y(n157) );
  INVX2TS U477 ( .A(n155), .Y(n357) );
  AOI22X1TS U478 ( .A0(n717), .A1(n357), .B0(n179), .B1(cacheAddressIn_B[3]), 
        .Y(n156) );
  OAI211XLTS U479 ( .A0(n369), .A1(n192), .B0(n157), .C0(n156), .Y(n1191) );
  AOI22X1TS U480 ( .A0(cacheAddressIn_SOUTH[2]), .A1(n174), .B0(
        \addressToWriteBuffer[1][2] ), .B1(n158), .Y(n160) );
  AOI22X1TS U481 ( .A0(n724), .A1(n353), .B0(n184), .B1(cacheAddressIn_B[2]), 
        .Y(n159) );
  OAI211XLTS U482 ( .A0(n161), .A1(n177), .B0(n160), .C0(n159), .Y(n1190) );
  INVX2TS U483 ( .A(n162), .Y(n188) );
  AOI22X1TS U484 ( .A0(cacheAddressIn_SOUTH[1]), .A1(n188), .B0(
        \addressToWriteBuffer[1][1] ), .B1(n178), .Y(n165) );
  AOI22X1TS U485 ( .A0(n733), .A1(n170), .B0(n139), .B1(cacheAddressIn_B[1]), 
        .Y(n164) );
  OAI211XLTS U486 ( .A0(n389), .A1(n182), .B0(n165), .C0(n164), .Y(n1189) );
  AOI22X1TS U487 ( .A0(cacheAddressIn_SOUTH[0]), .A1(n183), .B0(
        \addressToWriteBuffer[1][0] ), .B1(n570), .Y(n167) );
  AOI22X1TS U488 ( .A0(n739), .A1(n348), .B0(n179), .B1(cacheAddressIn_B[0]), 
        .Y(n166) );
  OAI211XLTS U489 ( .A0(n168), .A1(n187), .B0(n167), .C0(n166), .Y(n1188) );
  AOI22X1TS U490 ( .A0(dataIn_SOUTH[5]), .A1(n169), .B0(
        \dataToWriteBuffer[1][5] ), .B1(n178), .Y(n172) );
  AOI22X1TS U491 ( .A0(n680), .A1(n170), .B0(n184), .B1(cacheDataIn_B[5]), .Y(
        n171) );
  OAI211XLTS U492 ( .A0(n173), .A1(n192), .B0(n172), .C0(n171), .Y(n1187) );
  AOI22X1TS U493 ( .A0(dataIn_SOUTH[4]), .A1(n174), .B0(
        \dataToWriteBuffer[1][4] ), .B1(n398), .Y(n176) );
  AOI22X1TS U494 ( .A0(n676), .A1(n170), .B0(n139), .B1(cacheDataIn_B[4]), .Y(
        n175) );
  OAI211XLTS U495 ( .A0(n396), .A1(n177), .B0(n176), .C0(n175), .Y(n1186) );
  AOI22X1TS U496 ( .A0(dataIn_SOUTH[3]), .A1(n188), .B0(
        \dataToWriteBuffer[1][3] ), .B1(n178), .Y(n181) );
  AOI22X1TS U497 ( .A0(n670), .A1(n348), .B0(n179), .B1(cacheDataIn_B[3]), .Y(
        n180) );
  OAI211XLTS U498 ( .A0(n402), .A1(n182), .B0(n181), .C0(n180), .Y(n1185) );
  AOI22X1TS U499 ( .A0(dataIn_SOUTH[2]), .A1(n183), .B0(
        \dataToWriteBuffer[1][2] ), .B1(n398), .Y(n186) );
  AOI22X1TS U500 ( .A0(n664), .A1(n362), .B0(n184), .B1(cacheDataIn_B[2]), .Y(
        n185) );
  OAI211XLTS U501 ( .A0(n410), .A1(n187), .B0(n186), .C0(n185), .Y(n1184) );
  AOI22X1TS U502 ( .A0(cacheAddressIn_SOUTH[5]), .A1(n188), .B0(
        \addressToWriteBuffer[1][5] ), .B1(n570), .Y(n191) );
  AOI22X1TS U503 ( .A0(n702), .A1(n357), .B0(n189), .B1(cacheAddressIn_B[5]), 
        .Y(n190) );
  OAI211XLTS U504 ( .A0(n373), .A1(n192), .B0(n191), .C0(n190), .Y(n1193) );
  CLKBUFX2TS U505 ( .A(n282), .Y(n571) );
  INVX2TS U506 ( .A(n571), .Y(n193) );
  INVX2TS U507 ( .A(n193), .Y(n345) );
  CLKBUFX2TS U508 ( .A(n346), .Y(n523) );
  CLKBUFX2TS U509 ( .A(n306), .Y(n808) );
  AOI22X1TS U510 ( .A0(\requesterPortBuffer[1][1] ), .A1(n523), .B0(n793), 
        .B1(n194), .Y(n195) );
  OAI211XLTS U511 ( .A0(n193), .A1(n196), .B0(n195), .C0(n217), .Y(n1357) );
  INVX2TS U512 ( .A(n197), .Y(n592) );
  AOI22X1TS U513 ( .A0(n610), .A1(n31), .B0(n198), .B1(n592), .Y(n300) );
  AOI222XLTS U514 ( .A0(n20), .A1(memWrite_SOUTH), .B0(memWrite_EAST), .B1(
        n201), .C0(memWrite_WEST), .C1(n200), .Y(n648) );
  NOR4XLTS U515 ( .A(n592), .B(n202), .C(n20), .D(n522), .Y(n302) );
  OAI211XLTS U516 ( .A0(n204), .A1(n300), .B0(n648), .C0(n646), .Y(n205) );
  INVX2TS U517 ( .A(n205), .Y(n1204) );
  CLKBUFX2TS U518 ( .A(n245), .Y(n256) );
  CLKBUFX2TS U519 ( .A(n241), .Y(n246) );
  CLKBUFX2TS U520 ( .A(n246), .Y(n212) );
  AOI222XLTS U521 ( .A0(\addressToWriteBuffer[6][1] ), .A1(n256), .B0(
        \addressToWriteBuffer[5][1] ), .B1(n225), .C0(n212), .C1(
        \addressToWriteBuffer[4][1] ), .Y(n206) );
  INVX2TS U522 ( .A(n206), .Y(n1313) );
  CLKBUFX2TS U523 ( .A(n385), .Y(n260) );
  CLKBUFX2TS U524 ( .A(n260), .Y(n214) );
  AOI222XLTS U525 ( .A0(\addressToWriteBuffer[6][7] ), .A1(n256), .B0(
        \addressToWriteBuffer[5][7] ), .B1(n214), .C0(n212), .C1(
        \addressToWriteBuffer[4][7] ), .Y(n207) );
  INVX2TS U526 ( .A(n207), .Y(n1307) );
  CLKBUFX2TS U527 ( .A(n436), .Y(n228) );
  CLKBUFX2TS U528 ( .A(n228), .Y(n279) );
  CLKBUFX2TS U529 ( .A(n246), .Y(n255) );
  AOI222XLTS U530 ( .A0(\addressToWriteBuffer[6][6] ), .A1(n279), .B0(
        \addressToWriteBuffer[5][6] ), .B1(n214), .C0(n255), .C1(
        \addressToWriteBuffer[4][6] ), .Y(n208) );
  INVX2TS U531 ( .A(n208), .Y(n1308) );
  AOI222XLTS U532 ( .A0(\addressToWriteBuffer[6][4] ), .A1(n256), .B0(
        \addressToWriteBuffer[5][4] ), .B1(n214), .C0(n255), .C1(
        \addressToWriteBuffer[4][4] ), .Y(n209) );
  INVX2TS U533 ( .A(n209), .Y(n1310) );
  CLKBUFX2TS U534 ( .A(n228), .Y(n276) );
  CLKBUFX2TS U535 ( .A(n276), .Y(n215) );
  CLKBUFX2TS U536 ( .A(n260), .Y(n258) );
  CLKBUFX2TS U537 ( .A(n243), .Y(n239) );
  AOI222XLTS U538 ( .A0(\addressToWriteBuffer[6][3] ), .A1(n215), .B0(
        \addressToWriteBuffer[5][3] ), .B1(n258), .C0(n239), .C1(
        \addressToWriteBuffer[4][3] ), .Y(n210) );
  INVX2TS U539 ( .A(n210), .Y(n1311) );
  AOI222XLTS U540 ( .A0(\addressToWriteBuffer[6][2] ), .A1(n215), .B0(
        \addressToWriteBuffer[5][2] ), .B1(n258), .C0(n212), .C1(
        \addressToWriteBuffer[4][2] ), .Y(n211) );
  INVX2TS U541 ( .A(n211), .Y(n1312) );
  AOI222XLTS U542 ( .A0(\addressToWriteBuffer[6][0] ), .A1(n215), .B0(
        \addressToWriteBuffer[5][0] ), .B1(n258), .C0(n212), .C1(
        \addressToWriteBuffer[4][0] ), .Y(n213) );
  INVX2TS U543 ( .A(n213), .Y(n1314) );
  AOI222XLTS U544 ( .A0(\addressToWriteBuffer[6][5] ), .A1(n215), .B0(
        \addressToWriteBuffer[5][5] ), .B1(n214), .C0(n239), .C1(
        \addressToWriteBuffer[4][5] ), .Y(n216) );
  INVX2TS U545 ( .A(n216), .Y(n1309) );
  AOI22X1TS U546 ( .A0(\requesterPortBuffer[1][0] ), .A1(n523), .B0(
        \prevRequesterPort_B[0] ), .B1(n194), .Y(n218) );
  OAI211XLTS U547 ( .A0(n193), .A1(n219), .B0(n218), .C0(n217), .Y(n1358) );
  CLKBUFX2TS U548 ( .A(n220), .Y(n288) );
  AOI222XLTS U549 ( .A0(\dataToWriteBuffer[6][3] ), .A1(n288), .B0(
        \dataToWriteBuffer[5][3] ), .B1(n225), .C0(n241), .C1(
        \dataToWriteBuffer[4][3] ), .Y(n221) );
  INVX2TS U550 ( .A(n221), .Y(n1240) );
  CLKBUFX2TS U551 ( .A(n430), .Y(n230) );
  CLKBUFX2TS U552 ( .A(n436), .Y(n433) );
  CLKBUFX2TS U553 ( .A(n433), .Y(n236) );
  AOI222XLTS U554 ( .A0(n230), .A1(\addressToWriteBuffer[0][2] ), .B0(
        \addressToWriteBuffer[2][2] ), .B1(n236), .C0(
        \addressToWriteBuffer[1][2] ), .C1(n271), .Y(n222) );
  INVX2TS U555 ( .A(n222), .Y(n1344) );
  CLKBUFX2TS U556 ( .A(n433), .Y(n439) );
  AOI222XLTS U557 ( .A0(n230), .A1(\addressToWriteBuffer[0][0] ), .B0(
        \addressToWriteBuffer[2][0] ), .B1(n439), .C0(
        \addressToWriteBuffer[1][0] ), .C1(n271), .Y(n223) );
  INVX2TS U558 ( .A(n223), .Y(n1346) );
  CLKBUFX2TS U559 ( .A(n245), .Y(n285) );
  AOI222XLTS U560 ( .A0(\dataToWriteBuffer[6][1] ), .A1(n285), .B0(
        \dataToWriteBuffer[5][1] ), .B1(n225), .C0(n239), .C1(
        \dataToWriteBuffer[4][1] ), .Y(n224) );
  INVX2TS U561 ( .A(n224), .Y(n1242) );
  AOI222XLTS U562 ( .A0(\dataToWriteBuffer[6][2] ), .A1(n285), .B0(
        \dataToWriteBuffer[5][2] ), .B1(n225), .C0(n587), .C1(
        \dataToWriteBuffer[4][2] ), .Y(n226) );
  INVX2TS U563 ( .A(n226), .Y(n1241) );
  CLKBUFX2TS U564 ( .A(n228), .Y(n265) );
  CLKBUFX2TS U565 ( .A(n573), .Y(n234) );
  AOI222XLTS U566 ( .A0(n243), .A1(\dataToWriteBuffer[0][3] ), .B0(
        \dataToWriteBuffer[2][3] ), .B1(n265), .C0(\dataToWriteBuffer[1][3] ), 
        .C1(n234), .Y(n227) );
  INVX2TS U567 ( .A(n227), .Y(n1264) );
  CLKBUFX2TS U568 ( .A(n228), .Y(n262) );
  AOI222XLTS U569 ( .A0(n230), .A1(\addressToWriteBuffer[0][7] ), .B0(
        \addressToWriteBuffer[2][7] ), .B1(n262), .C0(
        \addressToWriteBuffer[1][7] ), .C1(n234), .Y(n229) );
  INVX2TS U570 ( .A(n229), .Y(n1339) );
  CLKBUFX2TS U571 ( .A(n573), .Y(n273) );
  AOI222XLTS U572 ( .A0(n230), .A1(\addressToWriteBuffer[0][3] ), .B0(
        \addressToWriteBuffer[2][3] ), .B1(n236), .C0(
        \addressToWriteBuffer[1][3] ), .C1(n273), .Y(n231) );
  INVX2TS U573 ( .A(n231), .Y(n1343) );
  AOI222XLTS U574 ( .A0(n246), .A1(\requesterPortBuffer[0][1] ), .B0(
        \requesterPortBuffer[2][1] ), .B1(n262), .C0(
        \requesterPortBuffer[1][1] ), .C1(n234), .Y(n232) );
  INVX2TS U575 ( .A(n232), .Y(n1282) );
  CLKBUFX2TS U576 ( .A(n430), .Y(n266) );
  AOI222XLTS U577 ( .A0(n266), .A1(\addressToWriteBuffer[0][6] ), .B0(
        \addressToWriteBuffer[2][6] ), .B1(n262), .C0(
        \addressToWriteBuffer[1][6] ), .C1(n273), .Y(n233) );
  INVX2TS U578 ( .A(n233), .Y(n1340) );
  AOI222XLTS U579 ( .A0(n266), .A1(\addressToWriteBuffer[0][4] ), .B0(
        \addressToWriteBuffer[2][4] ), .B1(n236), .C0(
        \addressToWriteBuffer[1][4] ), .C1(n234), .Y(n235) );
  INVX2TS U580 ( .A(n235), .Y(n1342) );
  AOI222XLTS U581 ( .A0(n266), .A1(\addressToWriteBuffer[0][5] ), .B0(
        \addressToWriteBuffer[2][5] ), .B1(n236), .C0(
        \addressToWriteBuffer[1][5] ), .C1(n273), .Y(n237) );
  INVX2TS U582 ( .A(n237), .Y(n1341) );
  CLKBUFX2TS U583 ( .A(n269), .Y(n263) );
  CLKBUFX2TS U584 ( .A(n385), .Y(n251) );
  CLKBUFX2TS U585 ( .A(n251), .Y(n412) );
  AOI222XLTS U586 ( .A0(n263), .A1(\requesterPortBuffer[3][1] ), .B0(n412), 
        .B1(\requesterPortBuffer[4][1] ), .C0(n276), .C1(
        \requesterPortBuffer[5][1] ), .Y(n238) );
  INVX2TS U587 ( .A(n238), .Y(n1276) );
  CLKBUFX2TS U588 ( .A(n260), .Y(n287) );
  AOI222XLTS U589 ( .A0(\dataToWriteBuffer[6][0] ), .A1(n288), .B0(
        \dataToWriteBuffer[5][0] ), .B1(n287), .C0(n239), .C1(
        \dataToWriteBuffer[4][0] ), .Y(n240) );
  INVX2TS U590 ( .A(n240), .Y(n1243) );
  AOI222XLTS U591 ( .A0(\dataToWriteBuffer[6][4] ), .A1(n285), .B0(
        \dataToWriteBuffer[5][4] ), .B1(n287), .C0(n241), .C1(
        \dataToWriteBuffer[4][4] ), .Y(n242) );
  INVX2TS U592 ( .A(n242), .Y(n1239) );
  AOI222XLTS U593 ( .A0(\dataToWriteBuffer[6][5] ), .A1(n303), .B0(
        \dataToWriteBuffer[5][5] ), .B1(n287), .C0(n243), .C1(
        \dataToWriteBuffer[4][5] ), .Y(n244) );
  INVX2TS U594 ( .A(n244), .Y(n1238) );
  CLKBUFX2TS U595 ( .A(n245), .Y(n295) );
  CLKBUFX2TS U596 ( .A(n246), .Y(n252) );
  AOI222XLTS U597 ( .A0(\addressToWriteBuffer[5][5] ), .A1(n295), .B0(n252), 
        .B1(\addressToWriteBuffer[3][5] ), .C0(n412), .C1(
        \addressToWriteBuffer[4][5] ), .Y(n247) );
  INVX2TS U598 ( .A(n247), .Y(n1317) );
  CLKBUFX2TS U599 ( .A(n251), .Y(n284) );
  AOI222XLTS U600 ( .A0(\addressToWriteBuffer[5][7] ), .A1(n253), .B0(n252), 
        .B1(\addressToWriteBuffer[3][7] ), .C0(n284), .C1(
        \addressToWriteBuffer[4][7] ), .Y(n248) );
  INVX2TS U601 ( .A(n248), .Y(n1315) );
  CLKBUFX2TS U602 ( .A(n251), .Y(n293) );
  AOI222XLTS U603 ( .A0(\addressToWriteBuffer[5][1] ), .A1(n279), .B0(n252), 
        .B1(\addressToWriteBuffer[3][1] ), .C0(n293), .C1(
        \addressToWriteBuffer[4][1] ), .Y(n249) );
  INVX2TS U604 ( .A(n249), .Y(n1321) );
  AOI222XLTS U605 ( .A0(\addressToWriteBuffer[5][0] ), .A1(n253), .B0(n255), 
        .B1(\addressToWriteBuffer[3][0] ), .C0(n284), .C1(
        \addressToWriteBuffer[4][0] ), .Y(n250) );
  INVX2TS U606 ( .A(n250), .Y(n1322) );
  CLKBUFX2TS U607 ( .A(n251), .Y(n290) );
  AOI222XLTS U608 ( .A0(\addressToWriteBuffer[5][3] ), .A1(n253), .B0(n252), 
        .B1(\addressToWriteBuffer[3][3] ), .C0(n290), .C1(
        \addressToWriteBuffer[4][3] ), .Y(n254) );
  INVX2TS U609 ( .A(n254), .Y(n1319) );
  AOI222XLTS U610 ( .A0(\addressToWriteBuffer[5][4] ), .A1(n256), .B0(n255), 
        .B1(\addressToWriteBuffer[3][4] ), .C0(n293), .C1(
        \addressToWriteBuffer[4][4] ), .Y(n257) );
  INVX2TS U611 ( .A(n257), .Y(n1318) );
  AOI222XLTS U612 ( .A0(n263), .A1(\dataToWriteBuffer[0][4] ), .B0(
        \dataToWriteBuffer[2][4] ), .B1(n265), .C0(\dataToWriteBuffer[1][4] ), 
        .C1(n258), .Y(n259) );
  INVX2TS U613 ( .A(n259), .Y(n1263) );
  CLKBUFX2TS U614 ( .A(n260), .Y(n268) );
  AOI222XLTS U615 ( .A0(n263), .A1(\dataToWriteBuffer[0][0] ), .B0(
        \dataToWriteBuffer[2][0] ), .B1(n265), .C0(\dataToWriteBuffer[1][0] ), 
        .C1(n268), .Y(n261) );
  INVX2TS U616 ( .A(n261), .Y(n1267) );
  AOI222XLTS U617 ( .A0(n263), .A1(\dataToWriteBuffer[0][2] ), .B0(
        \dataToWriteBuffer[2][2] ), .B1(n262), .C0(\dataToWriteBuffer[1][2] ), 
        .C1(n268), .Y(n264) );
  INVX2TS U618 ( .A(n264), .Y(n1265) );
  AOI222XLTS U619 ( .A0(n266), .A1(\dataToWriteBuffer[0][1] ), .B0(
        \dataToWriteBuffer[2][1] ), .B1(n265), .C0(\dataToWriteBuffer[1][1] ), 
        .C1(n268), .Y(n267) );
  INVX2TS U620 ( .A(n267), .Y(n1266) );
  AOI222XLTS U621 ( .A0(n269), .A1(\dataToWriteBuffer[0][5] ), .B0(
        \dataToWriteBuffer[2][5] ), .B1(n276), .C0(\dataToWriteBuffer[1][5] ), 
        .C1(n268), .Y(n270) );
  INVX2TS U622 ( .A(n270), .Y(n1262) );
  AOI222XLTS U623 ( .A0(n571), .A1(\addressToWriteBuffer[0][1] ), .B0(
        \addressToWriteBuffer[2][1] ), .B1(n439), .C0(
        \addressToWriteBuffer[1][1] ), .C1(n271), .Y(n272) );
  INVX2TS U624 ( .A(n272), .Y(n1345) );
  AOI222XLTS U625 ( .A0(n571), .A1(\requesterPortBuffer[0][0] ), .B0(
        \requesterPortBuffer[2][0] ), .B1(n439), .C0(
        \requesterPortBuffer[1][0] ), .C1(n273), .Y(n274) );
  INVX2TS U626 ( .A(n274), .Y(n1363) );
  CLKBUFX2TS U627 ( .A(n275), .Y(n434) );
  AOI222XLTS U628 ( .A0(n411), .A1(\requesterPortBuffer[3][0] ), .B0(n434), 
        .B1(\requesterPortBuffer[4][0] ), .C0(n276), .C1(
        \requesterPortBuffer[5][0] ), .Y(n277) );
  INVX2TS U629 ( .A(n277), .Y(n1277) );
  CLKBUFX2TS U630 ( .A(n282), .Y(n291) );
  AOI222XLTS U631 ( .A0(\addressToWriteBuffer[5][6] ), .A1(n279), .B0(n291), 
        .B1(\addressToWriteBuffer[3][6] ), .C0(n290), .C1(
        \addressToWriteBuffer[4][6] ), .Y(n278) );
  INVX2TS U632 ( .A(n278), .Y(n1316) );
  AOI222XLTS U633 ( .A0(\addressToWriteBuffer[5][2] ), .A1(n279), .B0(n291), 
        .B1(\addressToWriteBuffer[3][2] ), .C0(n293), .C1(
        \addressToWriteBuffer[4][2] ), .Y(n280) );
  INVX2TS U634 ( .A(n280), .Y(n1320) );
  AOI222XLTS U635 ( .A0(\dataToWriteBuffer[5][3] ), .A1(n295), .B0(n291), .B1(
        \dataToWriteBuffer[3][3] ), .C0(n290), .C1(\dataToWriteBuffer[4][3] ), 
        .Y(n281) );
  INVX2TS U636 ( .A(n281), .Y(n1246) );
  CLKBUFX2TS U637 ( .A(n282), .Y(n294) );
  AOI222XLTS U638 ( .A0(\dataToWriteBuffer[5][2] ), .A1(n288), .B0(n294), .B1(
        \dataToWriteBuffer[3][2] ), .C0(n284), .C1(\dataToWriteBuffer[4][2] ), 
        .Y(n283) );
  INVX2TS U639 ( .A(n283), .Y(n1247) );
  AOI222XLTS U640 ( .A0(\dataToWriteBuffer[5][0] ), .A1(n285), .B0(n294), .B1(
        \dataToWriteBuffer[3][0] ), .C0(n284), .C1(\dataToWriteBuffer[4][0] ), 
        .Y(n286) );
  INVX2TS U641 ( .A(n286), .Y(n1249) );
  AOI222XLTS U642 ( .A0(\dataToWriteBuffer[5][4] ), .A1(n288), .B0(n294), .B1(
        \dataToWriteBuffer[3][4] ), .C0(n287), .C1(\dataToWriteBuffer[4][4] ), 
        .Y(n289) );
  INVX2TS U643 ( .A(n289), .Y(n1245) );
  AOI222XLTS U644 ( .A0(\dataToWriteBuffer[5][1] ), .A1(n295), .B0(n291), .B1(
        \dataToWriteBuffer[3][1] ), .C0(n290), .C1(\dataToWriteBuffer[4][1] ), 
        .Y(n292) );
  INVX2TS U645 ( .A(n292), .Y(n1248) );
  AOI222XLTS U646 ( .A0(\dataToWriteBuffer[5][5] ), .A1(n295), .B0(n294), .B1(
        \dataToWriteBuffer[3][5] ), .C0(n293), .C1(\dataToWriteBuffer[4][5] ), 
        .Y(n296) );
  INVX2TS U647 ( .A(n296), .Y(n1244) );
  NOR2XLTS U648 ( .A(n300), .B(n18), .Y(n607) );
  AOI21X1TS U649 ( .A0(n687), .A1(n302), .B0(n425), .Y(n615) );
  INVX2TS U650 ( .A(n615), .Y(n298) );
  AOI211XLTS U651 ( .A0(n300), .A1(n299), .B0(n607), .C0(n298), .Y(n1211) );
  NAND3XLTS U652 ( .A(N883), .B(n12), .C(N882), .Y(n301) );
  INVX2TS U653 ( .A(n301), .Y(n524) );
  NAND2X1TS U654 ( .A(n524), .B(n303), .Y(n305) );
  OAI211XLTS U655 ( .A0(n302), .A1(n301), .B0(n440), .C0(n762), .Y(n598) );
  INVX2TS U656 ( .A(n598), .Y(n596) );
  NAND2X1TS U657 ( .A(n596), .B(\requesterPortBuffer[5][1] ), .Y(n304) );
  OAI211XLTS U658 ( .A0(n25), .A1(n305), .B0(n304), .C0(n589), .Y(n1272) );
  NOR2XLTS U659 ( .A(prevRequesterPort_A[0]), .B(prevRequesterPort_A[1]), .Y(
        n415) );
  NOR3XLTS U660 ( .A(\prevRequesterPort_B[0] ), .B(n793), .C(n415), .Y(n414)
         );
  CLKBUFX2TS U661 ( .A(n306), .Y(n640) );
  NAND2X1TS U662 ( .A(n414), .B(n640), .Y(n313) );
  INVX2TS U663 ( .A(n6), .Y(n750) );
  NOR2BX1TS U664 ( .AN(n415), .B(n749), .Y(n311) );
  AOI22X1TS U665 ( .A0(n750), .A1(n311), .B0(n310), .B1(
        requesterAddressOut_NORTH[2]), .Y(n307) );
  INVX2TS U666 ( .A(n8), .Y(n756) );
  AOI22X1TS U667 ( .A0(n756), .A1(n311), .B0(n310), .B1(
        requesterAddressOut_NORTH[0]), .Y(n308) );
  INVX2TS U668 ( .A(n5), .Y(n745) );
  AOI22X1TS U669 ( .A0(n745), .A1(n311), .B0(n310), .B1(
        requesterAddressOut_NORTH[3]), .Y(n309) );
  INVX2TS U670 ( .A(n7), .Y(n752) );
  AOI22X1TS U671 ( .A0(n752), .A1(n311), .B0(n310), .B1(
        requesterAddressOut_NORTH[1]), .Y(n312) );
  INVX2TS U672 ( .A(n314), .Y(n586) );
  NOR4BXLTS U673 ( .AN(n317), .B(n421), .C(n610), .D(n316), .Y(n580) );
  AOI21X1TS U674 ( .A0(\requesterPortBuffer[3][0] ), .A1(n586), .B0(n580), .Y(
        n319) );
  AOI22X1TS U675 ( .A0(\requesterPortBuffer[2][0] ), .A1(n329), .B0(n518), 
        .B1(\requesterPortBuffer[4][0] ), .Y(n318) );
  AOI22X1TS U676 ( .A0(\addressToWriteBuffer[3][7] ), .A1(n328), .B0(n374), 
        .B1(\addressToWriteBuffer[4][7] ), .Y(n321) );
  NAND2X1TS U677 ( .A(\addressToWriteBuffer[2][7] ), .B(n517), .Y(n320) );
  AOI22X1TS U678 ( .A0(\dataToWriteBuffer[3][2] ), .A1(n338), .B0(n405), .B1(
        \dataToWriteBuffer[4][2] ), .Y(n324) );
  NAND2X1TS U679 ( .A(\dataToWriteBuffer[2][2] ), .B(n322), .Y(n323) );
  AOI22X1TS U680 ( .A0(\addressToWriteBuffer[3][0] ), .A1(n328), .B0(n384), 
        .B1(\addressToWriteBuffer[4][0] ), .Y(n327) );
  INVX2TS U681 ( .A(n325), .Y(n582) );
  NAND2X1TS U682 ( .A(\addressToWriteBuffer[2][0] ), .B(n582), .Y(n326) );
  AOI22X1TS U683 ( .A0(\addressToWriteBuffer[3][6] ), .A1(n328), .B0(n392), 
        .B1(\addressToWriteBuffer[4][6] ), .Y(n331) );
  NAND2X1TS U684 ( .A(\addressToWriteBuffer[2][6] ), .B(n329), .Y(n330) );
  AOI22X1TS U685 ( .A0(\dataToWriteBuffer[3][3] ), .A1(n437), .B0(n392), .B1(
        \dataToWriteBuffer[4][3] ), .Y(n333) );
  NAND2X1TS U686 ( .A(\dataToWriteBuffer[2][3] ), .B(n322), .Y(n332) );
  AOI22X1TS U687 ( .A0(\dataToWriteBuffer[3][5] ), .A1(n338), .B0(n518), .B1(
        \dataToWriteBuffer[4][5] ), .Y(n335) );
  NAND2X1TS U688 ( .A(\dataToWriteBuffer[2][5] ), .B(n582), .Y(n334) );
  AOI22X1TS U689 ( .A0(\addressToWriteBuffer[3][4] ), .A1(n338), .B0(n337), 
        .B1(\addressToWriteBuffer[4][4] ), .Y(n340) );
  NAND2X1TS U690 ( .A(\addressToWriteBuffer[2][4] ), .B(n59), .Y(n339) );
  AOI22X1TS U691 ( .A0(\dataToWriteBuffer[3][1] ), .A1(n437), .B0(n374), .B1(
        \dataToWriteBuffer[4][1] ), .Y(n343) );
  NAND2X1TS U692 ( .A(\dataToWriteBuffer[2][1] ), .B(n59), .Y(n342) );
  AOI22X1TS U693 ( .A0(n352), .A1(requesterAddressIn_SOUTH[1]), .B0(n135), 
        .B1(requesterAddressIn_EAST[1]), .Y(n351) );
  INVX2TS U694 ( .A(n345), .Y(n360) );
  CLKBUFX2TS U695 ( .A(n346), .Y(n593) );
  AOI22X1TS U696 ( .A0(\requesterAddressBuffer[1][1] ), .A1(n593), .B0(
        prevRequesterAddress_B[1]), .B1(n347), .Y(n350) );
  NAND2X1TS U697 ( .A(requesterAddressIn_WEST[1]), .B(n348), .Y(n349) );
  AOI22X1TS U698 ( .A0(n352), .A1(requesterAddressIn_SOUTH[3]), .B0(n135), 
        .B1(requesterAddressIn_EAST[3]), .Y(n356) );
  AOI22X1TS U699 ( .A0(\requesterAddressBuffer[1][3] ), .A1(n593), .B0(
        prevRequesterAddress_B[3]), .B1(n347), .Y(n355) );
  NAND2X1TS U700 ( .A(requesterAddressIn_WEST[3]), .B(n353), .Y(n354) );
  AOI22X1TS U701 ( .A0(n22), .A1(requesterAddressIn_SOUTH[2]), .B0(n135), .B1(
        requesterAddressIn_EAST[2]), .Y(n361) );
  AOI22X1TS U702 ( .A0(\requesterAddressBuffer[1][2] ), .A1(n523), .B0(
        prevRequesterAddress_B[2]), .B1(n347), .Y(n359) );
  NAND2X1TS U703 ( .A(requesterAddressIn_WEST[2]), .B(n357), .Y(n358) );
  AOI22X1TS U704 ( .A0(n22), .A1(requesterAddressIn_SOUTH[0]), .B0(n134), .B1(
        requesterAddressIn_EAST[0]), .Y(n365) );
  AOI22X1TS U705 ( .A0(\requesterAddressBuffer[1][0] ), .A1(n593), .B0(
        prevRequesterAddress_B[0]), .B1(n347), .Y(n364) );
  NAND2X1TS U706 ( .A(requesterAddressIn_WEST[0]), .B(n362), .Y(n363) );
  INVX2TS U707 ( .A(n366), .Y(n383) );
  AOI22X1TS U708 ( .A0(n717), .A1(n383), .B0(n397), .B1(
        \addressToWriteBuffer[1][3] ), .Y(n368) );
  AOI22X1TS U709 ( .A0(n370), .A1(\addressToWriteBuffer[2][3] ), .B0(n378), 
        .B1(\addressToWriteBuffer[3][3] ), .Y(n367) );
  AOI22X1TS U710 ( .A0(n702), .A1(n383), .B0(n382), .B1(
        \addressToWriteBuffer[1][5] ), .Y(n372) );
  AOI22X1TS U711 ( .A0(n370), .A1(\addressToWriteBuffer[2][5] ), .B0(n378), 
        .B1(\addressToWriteBuffer[3][5] ), .Y(n371) );
  AOI22X1TS U712 ( .A0(n697), .A1(n383), .B0(n403), .B1(
        \addressToWriteBuffer[1][6] ), .Y(n376) );
  AOI22X1TS U713 ( .A0(n406), .A1(\addressToWriteBuffer[2][6] ), .B0(n374), 
        .B1(\addressToWriteBuffer[3][6] ), .Y(n375) );
  AOI22X1TS U714 ( .A0(n655), .A1(n391), .B0(n390), .B1(
        \dataToWriteBuffer[1][0] ), .Y(n380) );
  AOI22X1TS U715 ( .A0(n61), .A1(\dataToWriteBuffer[2][0] ), .B0(n378), .B1(
        \dataToWriteBuffer[3][0] ), .Y(n379) );
  AOI22X1TS U716 ( .A0(n733), .A1(n383), .B0(n382), .B1(
        \addressToWriteBuffer[1][1] ), .Y(n387) );
  AOI22X1TS U717 ( .A0(n385), .A1(\addressToWriteBuffer[2][1] ), .B0(n384), 
        .B1(\addressToWriteBuffer[3][1] ), .Y(n386) );
  AOI22X1TS U718 ( .A0(n676), .A1(n391), .B0(n390), .B1(
        \dataToWriteBuffer[1][4] ), .Y(n394) );
  AOI22X1TS U719 ( .A0(n406), .A1(\dataToWriteBuffer[2][4] ), .B0(n392), .B1(
        \dataToWriteBuffer[3][4] ), .Y(n393) );
  AOI22X1TS U720 ( .A0(n670), .A1(n404), .B0(n397), .B1(
        \dataToWriteBuffer[1][3] ), .Y(n400) );
  AOI22X1TS U721 ( .A0(n41), .A1(\dataToWriteBuffer[2][3] ), .B0(n398), .B1(
        \dataToWriteBuffer[3][3] ), .Y(n399) );
  AOI22X1TS U722 ( .A0(n664), .A1(n404), .B0(n403), .B1(
        \dataToWriteBuffer[1][2] ), .Y(n408) );
  AOI22X1TS U723 ( .A0(n406), .A1(\dataToWriteBuffer[2][2] ), .B0(n405), .B1(
        \dataToWriteBuffer[3][2] ), .Y(n407) );
  AO22XLTS U724 ( .A0(n411), .A1(\requesterPortBuffer[4][0] ), .B0(n412), .B1(
        \requesterPortBuffer[5][0] ), .Y(n798) );
  AO22XLTS U725 ( .A0(n413), .A1(\requesterPortBuffer[4][1] ), .B0(n412), .B1(
        \requesterPortBuffer[5][1] ), .Y(n799) );
  AO22XLTS U726 ( .A0(n415), .A1(prevMemRead_A), .B0(n414), .B1(prevMemRead_B), 
        .Y(N5457) );
  NOR2XLTS U727 ( .A(prevRequesterPort_A[1]), .B(n795), .Y(n775) );
  INVX2TS U728 ( .A(n792), .Y(n416) );
  NOR3XLTS U729 ( .A(\prevRequesterPort_B[0] ), .B(n759), .C(n792), .Y(n764)
         );
  INVX2TS U730 ( .A(n11), .Y(n746) );
  INVX2TS U731 ( .A(n10), .Y(n419) );
  AO22XLTS U732 ( .A0(n746), .A1(prevMemRead_A), .B0(n419), .B1(prevMemRead_B), 
        .Y(N5481) );
  NAND2X1TS U733 ( .A(n77), .B(n424), .Y(n422) );
  NAND2X1TS U734 ( .A(n19), .B(n621), .Y(n653) );
  INVX2TS U735 ( .A(n9), .Y(n620) );
  NAND2BX1TS U736 ( .AN(n620), .B(n33), .Y(n427) );
  OR3X1TS U737 ( .A(n424), .B(n20), .C(n427), .Y(n671) );
  INVX2TS U738 ( .A(n671), .Y(n660) );
  NOR2XLTS U739 ( .A(n17), .B(n425), .Y(n629) );
  CLKBUFX2TS U740 ( .A(n629), .Y(n635) );
  AOI22X1TS U741 ( .A0(\requesterPortBuffer[0][0] ), .A1(n635), .B0(
        prevRequesterPort_A[0]), .B1(n620), .Y(n426) );
  INVX2TS U742 ( .A(n428), .Y(n634) );
  INVX2TS U743 ( .A(n634), .Y(n715) );
  AOI22X1TS U744 ( .A0(\requesterPortBuffer[0][1] ), .A1(n635), .B0(
        prevRequesterPort_A[1]), .B1(n620), .Y(n429) );
  AOI22X1TS U745 ( .A0(n345), .A1(\requesterAddressBuffer[0][0] ), .B0(
        requesterAddressIn_SOUTH[0]), .B1(n434), .Y(n431) );
  OAI2BB1X1TS U746 ( .A0N(requesterAddressIn_EAST[0]), .A1N(n433), .B0(n431), 
        .Y(n1354) );
  AOI22X1TS U747 ( .A0(n345), .A1(\requesterAddressBuffer[0][1] ), .B0(
        requesterAddressIn_SOUTH[1]), .B1(n434), .Y(n432) );
  OAI2BB1X1TS U748 ( .A0N(requesterAddressIn_EAST[1]), .A1N(n433), .B0(n432), 
        .Y(n1353) );
  AOI22X1TS U749 ( .A0(n430), .A1(\requesterAddressBuffer[0][2] ), .B0(
        requesterAddressIn_SOUTH[2]), .B1(n434), .Y(n435) );
  OAI2BB1X1TS U750 ( .A0N(requesterAddressIn_EAST[2]), .A1N(n436), .B0(n435), 
        .Y(n1352) );
  AOI22X1TS U751 ( .A0(n413), .A1(\requesterAddressBuffer[0][3] ), .B0(
        requesterAddressIn_SOUTH[3]), .B1(n437), .Y(n438) );
  OAI2BB1X1TS U752 ( .A0N(requesterAddressIn_EAST[3]), .A1N(n439), .B0(n438), 
        .Y(n1351) );
  NAND2X1TS U753 ( .A(n464), .B(n441), .Y(n450) );
  AOI22X1TS U754 ( .A0(requesterAddressIn_EAST[0]), .A1(n449), .B0(
        requesterAddressIn_WEST[0]), .B1(n450), .Y(n445) );
  NAND3X1TS U755 ( .A(n574), .B(n442), .C(n513), .Y(n578) );
  NAND2X1TS U756 ( .A(n443), .B(n578), .Y(n444) );
  INVX2TS U757 ( .A(n578), .Y(n516) );
  OAI2BB2XLTS U758 ( .B0(n445), .B1(n444), .A0N(n516), .A1N(
        \requesterAddressBuffer[1][0] ), .Y(n1350) );
  AOI22X1TS U759 ( .A0(requesterAddressIn_WEST[1]), .A1(n450), .B0(
        requesterAddressIn_EAST[1]), .B1(n449), .Y(n446) );
  OAI2BB2XLTS U760 ( .B0(n446), .B1(n444), .A0N(n516), .A1N(
        \requesterAddressBuffer[1][1] ), .Y(n1349) );
  AOI22X1TS U761 ( .A0(requesterAddressIn_WEST[2]), .A1(n450), .B0(
        requesterAddressIn_EAST[2]), .B1(n449), .Y(n448) );
  INVX2TS U762 ( .A(n578), .Y(n451) );
  OAI2BB2XLTS U763 ( .B0(n448), .B1(n447), .A0N(n451), .A1N(
        \requesterAddressBuffer[1][2] ), .Y(n1348) );
  AOI22X1TS U764 ( .A0(requesterAddressIn_WEST[3]), .A1(n450), .B0(
        requesterAddressIn_EAST[3]), .B1(n449), .Y(n452) );
  OAI2BB2XLTS U765 ( .B0(n452), .B1(n447), .A0N(n451), .A1N(
        \requesterAddressBuffer[1][3] ), .Y(n1347) );
  NAND3X1TS U766 ( .A(n457), .B(n456), .C(n455), .Y(n466) );
  NAND2X1TS U767 ( .A(n459), .B(n458), .Y(n468) );
  INVX2TS U768 ( .A(n314), .Y(n584) );
  AOI211XLTS U769 ( .A0(n524), .A1(n23), .B0(n584), .C0(n747), .Y(n460) );
  INVX2TS U770 ( .A(n461), .Y(n485) );
  INVX2TS U771 ( .A(n465), .Y(n483) );
  INVX2TS U772 ( .A(n483), .Y(n495) );
  INVX2TS U773 ( .A(n467), .Y(n484) );
  OR2X1TS U774 ( .A(n747), .B(n468), .Y(n496) );
  INVX2TS U775 ( .A(n496), .Y(n542) );
  AOI22X1TS U776 ( .A0(n461), .A1(\addressToWriteBuffer[5][0] ), .B0(
        cacheAddressIn_EAST[0]), .B1(n542), .Y(n472) );
  CLKBUFX2TS U777 ( .A(n545), .Y(n531) );
  CLKBUFX2TS U778 ( .A(n531), .Y(n564) );
  NAND2X1TS U779 ( .A(n470), .B(n469), .Y(n486) );
  INVX2TS U780 ( .A(n486), .Y(n554) );
  AOI22X1TS U781 ( .A0(n564), .A1(\addressToWriteBuffer[6][0] ), .B0(
        cacheAddressIn_SOUTH[0]), .B1(n554), .Y(n471) );
  INVX2TS U782 ( .A(n483), .Y(n551) );
  INVX2TS U783 ( .A(n484), .Y(n568) );
  INVX2TS U784 ( .A(n485), .Y(n543) );
  INVX2TS U785 ( .A(n496), .Y(n536) );
  AOI22X1TS U786 ( .A0(n543), .A1(\addressToWriteBuffer[5][1] ), .B0(n536), 
        .B1(cacheAddressIn_EAST[1]), .Y(n476) );
  INVX2TS U787 ( .A(n486), .Y(n563) );
  AOI22X1TS U788 ( .A0(n506), .A1(\addressToWriteBuffer[6][1] ), .B0(n563), 
        .B1(cacheAddressIn_SOUTH[1]), .Y(n475) );
  INVX2TS U789 ( .A(n483), .Y(n560) );
  INVX2TS U790 ( .A(n484), .Y(n558) );
  INVX2TS U791 ( .A(n485), .Y(n553) );
  AOI22X1TS U792 ( .A0(n553), .A1(\addressToWriteBuffer[5][2] ), .B0(n542), 
        .B1(cacheAddressIn_EAST[2]), .Y(n480) );
  CLKBUFX2TS U793 ( .A(n531), .Y(n501) );
  INVX2TS U794 ( .A(n486), .Y(n537) );
  AOI22X1TS U795 ( .A0(n501), .A1(\addressToWriteBuffer[6][2] ), .B0(n537), 
        .B1(cacheAddressIn_SOUTH[2]), .Y(n479) );
  INVX2TS U796 ( .A(n484), .Y(n549) );
  INVX2TS U797 ( .A(n485), .Y(n562) );
  INVX2TS U798 ( .A(n496), .Y(n552) );
  AOI22X1TS U799 ( .A0(n562), .A1(\addressToWriteBuffer[5][3] ), .B0(n552), 
        .B1(cacheAddressIn_EAST[3]), .Y(n488) );
  INVX2TS U800 ( .A(n486), .Y(n544) );
  AOI22X1TS U801 ( .A0(n506), .A1(\addressToWriteBuffer[6][3] ), .B0(n544), 
        .B1(cacheAddressIn_SOUTH[3]), .Y(n487) );
  AOI22X1TS U802 ( .A0(n461), .A1(\addressToWriteBuffer[5][4] ), .B0(n552), 
        .B1(cacheAddressIn_EAST[4]), .Y(n492) );
  AOI22X1TS U803 ( .A0(n501), .A1(\addressToWriteBuffer[6][4] ), .B0(n554), 
        .B1(cacheAddressIn_SOUTH[4]), .Y(n491) );
  INVX2TS U804 ( .A(n496), .Y(n561) );
  AOI22X1TS U805 ( .A0(n543), .A1(\addressToWriteBuffer[5][5] ), .B0(n561), 
        .B1(cacheAddressIn_EAST[5]), .Y(n498) );
  AOI22X1TS U806 ( .A0(n501), .A1(\addressToWriteBuffer[6][5] ), .B0(n563), 
        .B1(cacheAddressIn_SOUTH[5]), .Y(n497) );
  AOI22X1TS U807 ( .A0(n553), .A1(\addressToWriteBuffer[5][6] ), .B0(n536), 
        .B1(cacheAddressIn_EAST[6]), .Y(n503) );
  AOI22X1TS U808 ( .A0(n501), .A1(\addressToWriteBuffer[6][6] ), .B0(n537), 
        .B1(cacheAddressIn_SOUTH[6]), .Y(n502) );
  AOI22X1TS U809 ( .A0(n562), .A1(\addressToWriteBuffer[5][7] ), .B0(n542), 
        .B1(cacheAddressIn_EAST[7]), .Y(n508) );
  AOI22X1TS U810 ( .A0(n506), .A1(\addressToWriteBuffer[6][7] ), .B0(n544), 
        .B1(cacheAddressIn_SOUTH[7]), .Y(n507) );
  AOI22X1TS U811 ( .A0(\requesterPortBuffer[2][0] ), .A1(n586), .B0(
        \requesterPortBuffer[3][0] ), .B1(n15), .Y(n511) );
  AOI21X1TS U812 ( .A0(n511), .A1(n38), .B0(n447), .Y(n512) );
  AOI22X1TS U813 ( .A0(\requesterPortBuffer[2][1] ), .A1(n584), .B0(
        \requesterPortBuffer[3][1] ), .B1(n15), .Y(n514) );
  AOI22X1TS U814 ( .A0(n517), .A1(\requesterPortBuffer[2][1] ), .B0(n580), 
        .B1(n640), .Y(n521) );
  AOI22X1TS U815 ( .A0(\requesterPortBuffer[3][1] ), .A1(n519), .B0(n518), 
        .B1(\requesterPortBuffer[4][1] ), .Y(n520) );
  NAND2X1TS U816 ( .A(n521), .B(n520), .Y(n1278) );
  NAND2X1TS U817 ( .A(n596), .B(\requesterPortBuffer[5][0] ), .Y(n526) );
  NAND4XLTS U818 ( .A(n25), .B(n524), .C(n523), .D(n522), .Y(n525) );
  AOI22X1TS U819 ( .A0(n543), .A1(\dataToWriteBuffer[5][0] ), .B0(n552), .B1(
        dataIn_EAST[0]), .Y(n528) );
  AOI22X1TS U820 ( .A0(n531), .A1(\dataToWriteBuffer[6][0] ), .B0(n554), .B1(
        dataIn_SOUTH[0]), .Y(n527) );
  AOI22X1TS U821 ( .A0(n553), .A1(\dataToWriteBuffer[5][1] ), .B0(n561), .B1(
        dataIn_EAST[1]), .Y(n533) );
  AOI22X1TS U822 ( .A0(n531), .A1(\dataToWriteBuffer[6][1] ), .B0(n563), .B1(
        dataIn_SOUTH[1]), .Y(n532) );
  AOI22X1TS U823 ( .A0(n562), .A1(\dataToWriteBuffer[5][2] ), .B0(n536), .B1(
        dataIn_EAST[2]), .Y(n539) );
  AOI22X1TS U824 ( .A0(n564), .A1(\dataToWriteBuffer[6][2] ), .B0(n537), .B1(
        dataIn_SOUTH[2]), .Y(n538) );
  AOI22X1TS U825 ( .A0(n543), .A1(\dataToWriteBuffer[5][3] ), .B0(n542), .B1(
        dataIn_EAST[3]), .Y(n547) );
  AOI22X1TS U826 ( .A0(n545), .A1(\dataToWriteBuffer[6][3] ), .B0(n544), .B1(
        dataIn_SOUTH[3]), .Y(n546) );
  AOI22X1TS U827 ( .A0(n553), .A1(\dataToWriteBuffer[5][4] ), .B0(n552), .B1(
        dataIn_EAST[4]), .Y(n556) );
  AOI22X1TS U828 ( .A0(n564), .A1(\dataToWriteBuffer[6][4] ), .B0(n554), .B1(
        dataIn_SOUTH[4]), .Y(n555) );
  AOI22X1TS U829 ( .A0(n562), .A1(\dataToWriteBuffer[5][5] ), .B0(n561), .B1(
        dataIn_EAST[5]), .Y(n566) );
  AOI22X1TS U830 ( .A0(n564), .A1(\dataToWriteBuffer[6][5] ), .B0(n563), .B1(
        dataIn_SOUTH[5]), .Y(n565) );
  AOI22X1TS U831 ( .A0(n571), .A1(isWrite[0]), .B0(isWrite[2]), .B1(n570), .Y(
        n572) );
  OAI2BB1X1TS U832 ( .A0N(isWrite[1]), .A1N(n573), .B0(n572), .Y(n1219) );
  CLKBUFX2TS U833 ( .A(memWrite_EAST), .Y(n595) );
  AOI22X1TS U834 ( .A0(n574), .A1(n595), .B0(isWrite[3]), .B1(n581), .Y(n575)
         );
  AOI21X1TS U835 ( .A0(n584), .A1(isWrite[2]), .B0(n577), .Y(n579) );
  OAI22X1TS U836 ( .A0(n579), .A1(n444), .B0(n578), .B1(n805), .Y(n1218) );
  INVX2TS U837 ( .A(n640), .Y(n774) );
  AOI222XLTS U838 ( .A0(n581), .A1(isWrite[4]), .B0(isWrite[3]), .B1(n586), 
        .C0(memWrite_WEST), .C1(n580), .Y(n583) );
  OAI2BB2XLTS U839 ( .B0(n774), .B1(n583), .A0N(n582), .A1N(isWrite[2]), .Y(
        n1217) );
  AOI22X1TS U840 ( .A0(isWrite[4]), .A1(n584), .B0(isWrite[5]), .B1(n14), .Y(
        n585) );
  OAI2BB2XLTS U841 ( .B0(n749), .B1(n585), .A0N(isWrite[3]), .A1N(n587), .Y(
        n1216) );
  NAND2X1TS U842 ( .A(isWrite[5]), .B(n586), .Y(n588) );
  OAI2BB2XLTS U843 ( .B0(n749), .B1(n588), .A0N(isWrite[4]), .A1N(n587), .Y(
        n1215) );
  INVX2TS U844 ( .A(n589), .Y(n590) );
  NAND2X1TS U845 ( .A(n591), .B(n590), .Y(n599) );
  OAI211XLTS U846 ( .A0(n595), .A1(n594), .B0(n593), .C0(n197), .Y(n597) );
  AOI32X1TS U847 ( .A0(n599), .A1(n598), .A2(n597), .B0(n596), .B1(n806), .Y(
        n1214) );
  CLKBUFX2TS U848 ( .A(n608), .Y(n613) );
  OAI21XLTS U849 ( .A0(n602), .A1(n609), .B0(n613), .Y(n603) );
  XNOR2X1TS U850 ( .A(n607), .B(n603), .Y(n605) );
  AOI21X1TS U851 ( .A0(n601), .A1(n605), .B0(n604), .Y(n1210) );
  OA21XLTS U852 ( .A0(n608), .A1(n606), .B0(n607), .Y(n612) );
  NOR2XLTS U853 ( .A(n610), .B(n609), .Y(n611) );
  NAND2X1TS U854 ( .A(N884), .B(n796), .Y(n614) );
  OAI21XLTS U855 ( .A0(N884), .A1(n606), .B0(n614), .Y(n617) );
  AOI21X1TS U856 ( .A0(n618), .A1(n617), .B0(n616), .Y(n1209) );
  CLKBUFX2TS U857 ( .A(n619), .Y(n675) );
  INVX2TS U858 ( .A(n675), .Y(n732) );
  INVX2TS U859 ( .A(n9), .Y(n633) );
  AOI22X1TS U860 ( .A0(requesterAddressIn_WEST[0]), .A1(n732), .B0(n756), .B1(
        n633), .Y(n625) );
  INVX2TS U861 ( .A(n634), .Y(n731) );
  AOI22X1TS U862 ( .A0(requesterAddressIn_EAST[0]), .A1(n731), .B0(n629), .B1(
        \requesterAddressBuffer[0][0] ), .Y(n624) );
  INVX2TS U863 ( .A(n622), .Y(n636) );
  INVX2TS U864 ( .A(n636), .Y(n718) );
  AOI22X1TS U865 ( .A0(n692), .A1(requesterAddressIn_SOUTH[0]), .B0(n718), 
        .B1(requesterAddressIn_NORTH[0]), .Y(n623) );
  INVX2TS U866 ( .A(n675), .Y(n701) );
  AOI22X1TS U867 ( .A0(requesterAddressIn_WEST[1]), .A1(n701), .B0(n752), .B1(
        n633), .Y(n628) );
  INVX2TS U868 ( .A(n634), .Y(n708) );
  AOI22X1TS U869 ( .A0(requesterAddressIn_EAST[1]), .A1(n708), .B0(n629), .B1(
        \requesterAddressBuffer[0][1] ), .Y(n627) );
  INVX2TS U870 ( .A(n671), .Y(n710) );
  INVX2TS U871 ( .A(n636), .Y(n741) );
  AOI22X1TS U872 ( .A0(n710), .A1(requesterAddressIn_SOUTH[1]), .B0(n741), 
        .B1(requesterAddressIn_NORTH[1]), .Y(n626) );
  INVX2TS U873 ( .A(n675), .Y(n723) );
  AOI22X1TS U874 ( .A0(requesterAddressIn_WEST[2]), .A1(n723), .B0(n750), .B1(
        n633), .Y(n632) );
  AOI22X1TS U875 ( .A0(requesterAddressIn_EAST[2]), .A1(n428), .B0(n629), .B1(
        \requesterAddressBuffer[0][2] ), .Y(n631) );
  INVX2TS U876 ( .A(n671), .Y(n740) );
  INVX2TS U877 ( .A(n636), .Y(n703) );
  AOI22X1TS U878 ( .A0(n740), .A1(requesterAddressIn_SOUTH[2]), .B0(n703), 
        .B1(requesterAddressIn_NORTH[2]), .Y(n630) );
  AOI22X1TS U879 ( .A0(requesterAddressIn_WEST[3]), .A1(n707), .B0(n745), .B1(
        n633), .Y(n639) );
  INVX2TS U880 ( .A(n634), .Y(n696) );
  AOI22X1TS U881 ( .A0(requesterAddressIn_EAST[3]), .A1(n696), .B0(n635), .B1(
        \requesterAddressBuffer[0][3] ), .Y(n638) );
  INVX2TS U882 ( .A(n636), .Y(n725) );
  AOI22X1TS U883 ( .A0(n660), .A1(requesterAddressIn_SOUTH[3]), .B0(n725), 
        .B1(requesterAddressIn_NORTH[3]), .Y(n637) );
  NAND2X1TS U884 ( .A(n32), .B(n640), .Y(n651) );
  AOI22X1TS U885 ( .A0(memWrite_WEST), .A1(n642), .B0(memWrite_EAST), .B1(n641), .Y(n644) );
  OAI211XLTS U886 ( .A0(memRead_NORTH), .A1(n645), .B0(n644), .C0(n643), .Y(
        n686) );
  INVX2TS U887 ( .A(n646), .Y(n647) );
  OAI22X1TS U888 ( .A0(isWrite[0]), .A1(n651), .B0(n686), .B1(n647), .Y(n1203)
         );
  AOI22X1TS U889 ( .A0(n17), .A1(n648), .B0(n805), .B1(n32), .Y(n650) );
  AOI32X1TS U890 ( .A0(n650), .A1(n649), .A2(n808), .B0(n139), .B1(n807), .Y(
        n1202) );
  INVX2TS U891 ( .A(n651), .Y(n652) );
  INVX2TS U892 ( .A(n652), .Y(n690) );
  INVX2TS U893 ( .A(n690), .Y(n669) );
  OR2X1TS U894 ( .A(n654), .B(n653), .Y(n668) );
  INVX2TS U895 ( .A(n668), .Y(n729) );
  AOI22X1TS U896 ( .A0(n669), .A1(\dataToWriteBuffer[0][0] ), .B0(n729), .B1(
        cacheDataIn_A[0]), .Y(n658) );
  AOI22X1TS U897 ( .A0(n655), .A1(n723), .B0(dataIn_EAST[0]), .B1(n696), .Y(
        n657) );
  AOI22X1TS U898 ( .A0(dataIn_NORTH[0]), .A1(n718), .B0(dataIn_SOUTH[0]), .B1(
        n660), .Y(n656) );
  INVX2TS U899 ( .A(n668), .Y(n737) );
  AOI22X1TS U900 ( .A0(n669), .A1(\dataToWriteBuffer[0][1] ), .B0(n737), .B1(
        cacheDataIn_A[1]), .Y(n663) );
  AOI22X1TS U901 ( .A0(n659), .A1(n707), .B0(dataIn_EAST[1]), .B1(n715), .Y(
        n662) );
  AOI22X1TS U902 ( .A0(dataIn_NORTH[1]), .A1(n703), .B0(dataIn_SOUTH[1]), .B1(
        n660), .Y(n661) );
  INVX2TS U903 ( .A(n668), .Y(n714) );
  AOI22X1TS U904 ( .A0(n669), .A1(\dataToWriteBuffer[0][2] ), .B0(n714), .B1(
        cacheDataIn_A[2]), .Y(n667) );
  AOI22X1TS U905 ( .A0(n664), .A1(n732), .B0(dataIn_EAST[2]), .B1(n708), .Y(
        n666) );
  AOI22X1TS U906 ( .A0(dataIn_NORTH[2]), .A1(n718), .B0(dataIn_SOUTH[2]), .B1(
        n692), .Y(n665) );
  INVX2TS U907 ( .A(n668), .Y(n722) );
  AOI22X1TS U908 ( .A0(n669), .A1(\dataToWriteBuffer[0][3] ), .B0(n722), .B1(
        cacheDataIn_A[3]), .Y(n674) );
  AOI22X1TS U909 ( .A0(n670), .A1(n701), .B0(dataIn_EAST[3]), .B1(n731), .Y(
        n673) );
  INVX2TS U910 ( .A(n671), .Y(n681) );
  AOI22X1TS U911 ( .A0(dataIn_NORTH[3]), .A1(n703), .B0(dataIn_SOUTH[3]), .B1(
        n681), .Y(n672) );
  INVX2TS U912 ( .A(n690), .Y(n738) );
  AOI22X1TS U913 ( .A0(n738), .A1(\dataToWriteBuffer[0][4] ), .B0(n729), .B1(
        cacheDataIn_A[4]), .Y(n679) );
  INVX2TS U914 ( .A(n675), .Y(n716) );
  AOI22X1TS U915 ( .A0(n676), .A1(n716), .B0(dataIn_EAST[4]), .B1(n696), .Y(
        n678) );
  AOI22X1TS U916 ( .A0(dataIn_NORTH[4]), .A1(n725), .B0(dataIn_SOUTH[4]), .B1(
        n681), .Y(n677) );
  AOI22X1TS U917 ( .A0(n730), .A1(\dataToWriteBuffer[0][5] ), .B0(n737), .B1(
        cacheDataIn_A[5]), .Y(n684) );
  AOI22X1TS U918 ( .A0(n680), .A1(n707), .B0(dataIn_EAST[5]), .B1(n731), .Y(
        n683) );
  AOI22X1TS U919 ( .A0(dataIn_NORTH[5]), .A1(n741), .B0(dataIn_SOUTH[5]), .B1(
        n681), .Y(n682) );
  OAI221XLTS U920 ( .A0(n687), .A1(isWrite[0]), .B0(n32), .B1(n686), .C0(n685), 
        .Y(n688) );
  INVX2TS U921 ( .A(n688), .Y(n689) );
  OAI2BB2XLTS U922 ( .B0(n722), .B1(n689), .A0N(n714), .A1N(memWrite_A), .Y(
        n1181) );
  INVX2TS U923 ( .A(n690), .Y(n730) );
  AOI22X1TS U924 ( .A0(n730), .A1(\addressToWriteBuffer[0][7] ), .B0(n714), 
        .B1(cacheAddressIn_A[7]), .Y(n695) );
  AOI22X1TS U925 ( .A0(n691), .A1(n701), .B0(cacheAddressIn_EAST[7]), .B1(n715), .Y(n694) );
  AOI22X1TS U926 ( .A0(cacheAddressIn_NORTH[7]), .A1(n741), .B0(
        cacheAddressIn_SOUTH[7]), .B1(n681), .Y(n693) );
  AOI22X1TS U927 ( .A0(n738), .A1(\addressToWriteBuffer[0][6] ), .B0(n722), 
        .B1(cacheAddressIn_A[6]), .Y(n700) );
  AOI22X1TS U928 ( .A0(n697), .A1(n716), .B0(cacheAddressIn_EAST[6]), .B1(n696), .Y(n699) );
  AOI22X1TS U929 ( .A0(cacheAddressIn_NORTH[6]), .A1(n725), .B0(
        cacheAddressIn_SOUTH[6]), .B1(n710), .Y(n698) );
  AOI22X1TS U930 ( .A0(n652), .A1(\addressToWriteBuffer[0][5] ), .B0(n729), 
        .B1(cacheAddressIn_A[5]), .Y(n706) );
  AOI22X1TS U931 ( .A0(n702), .A1(n701), .B0(cacheAddressIn_EAST[5]), .B1(n708), .Y(n705) );
  AOI22X1TS U932 ( .A0(cacheAddressIn_NORTH[5]), .A1(n703), .B0(
        cacheAddressIn_SOUTH[5]), .B1(n710), .Y(n704) );
  AOI22X1TS U933 ( .A0(n730), .A1(\addressToWriteBuffer[0][4] ), .B0(n737), 
        .B1(cacheAddressIn_A[4]), .Y(n713) );
  AOI22X1TS U934 ( .A0(n709), .A1(n716), .B0(cacheAddressIn_EAST[4]), .B1(n708), .Y(n712) );
  AOI22X1TS U935 ( .A0(cacheAddressIn_NORTH[4]), .A1(n622), .B0(
        cacheAddressIn_SOUTH[4]), .B1(n710), .Y(n711) );
  AOI22X1TS U936 ( .A0(n738), .A1(\addressToWriteBuffer[0][3] ), .B0(n714), 
        .B1(cacheAddressIn_A[3]), .Y(n721) );
  AOI22X1TS U937 ( .A0(n717), .A1(n716), .B0(cacheAddressIn_EAST[3]), .B1(n715), .Y(n720) );
  AOI22X1TS U938 ( .A0(cacheAddressIn_NORTH[3]), .A1(n718), .B0(
        cacheAddressIn_SOUTH[3]), .B1(n692), .Y(n719) );
  AOI22X1TS U939 ( .A0(n652), .A1(\addressToWriteBuffer[0][2] ), .B0(n722), 
        .B1(cacheAddressIn_A[2]), .Y(n728) );
  AOI22X1TS U940 ( .A0(n724), .A1(n723), .B0(cacheAddressIn_EAST[2]), .B1(n428), .Y(n727) );
  AOI22X1TS U941 ( .A0(cacheAddressIn_NORTH[2]), .A1(n725), .B0(
        cacheAddressIn_SOUTH[2]), .B1(n740), .Y(n726) );
  AOI22X1TS U942 ( .A0(n730), .A1(\addressToWriteBuffer[0][1] ), .B0(n729), 
        .B1(cacheAddressIn_A[1]), .Y(n736) );
  AOI22X1TS U943 ( .A0(n733), .A1(n732), .B0(cacheAddressIn_EAST[1]), .B1(n731), .Y(n735) );
  AOI22X1TS U944 ( .A0(cacheAddressIn_NORTH[1]), .A1(n622), .B0(
        cacheAddressIn_SOUTH[1]), .B1(n740), .Y(n734) );
  AOI22X1TS U945 ( .A0(n738), .A1(\addressToWriteBuffer[0][0] ), .B0(n737), 
        .B1(cacheAddressIn_A[0]), .Y(n744) );
  AOI22X1TS U946 ( .A0(n739), .A1(n723), .B0(cacheAddressIn_EAST[0]), .B1(n428), .Y(n743) );
  AOI22X1TS U947 ( .A0(cacheAddressIn_NORTH[0]), .A1(n741), .B0(
        cacheAddressIn_SOUTH[0]), .B1(n740), .Y(n742) );
  INVX2TS U948 ( .A(n11), .Y(n755) );
  INVX2TS U949 ( .A(n10), .Y(n754) );
  AOI22X1TS U950 ( .A0(n745), .A1(n755), .B0(prevRequesterAddress_B[3]), .B1(
        n754), .Y(n748) );
  AOI211XLTS U951 ( .A0(\prevRequesterPort_B[0] ), .A1(n793), .B0(n747), .C0(
        n746), .Y(n757) );
  OAI2BB2XLTS U952 ( .B0(n749), .B1(n748), .A0N(requesterAddressOut_WEST[3]), 
        .A1N(n757), .Y(n1171) );
  INVX2TS U953 ( .A(n808), .Y(n761) );
  AOI22X1TS U954 ( .A0(n750), .A1(n755), .B0(prevRequesterAddress_B[2]), .B1(
        n754), .Y(n751) );
  OAI2BB2XLTS U955 ( .B0(n761), .B1(n751), .A0N(requesterAddressOut_WEST[2]), 
        .A1N(n757), .Y(n1170) );
  AOI22X1TS U956 ( .A0(n752), .A1(n755), .B0(prevRequesterAddress_B[1]), .B1(
        n754), .Y(n753) );
  OAI2BB2XLTS U957 ( .B0(n761), .B1(n753), .A0N(requesterAddressOut_WEST[1]), 
        .A1N(n757), .Y(n1169) );
  AOI22X1TS U958 ( .A0(n756), .A1(n755), .B0(prevRequesterAddress_B[0]), .B1(
        n754), .Y(n758) );
  OAI2BB2XLTS U959 ( .B0(n761), .B1(n758), .A0N(requesterAddressOut_WEST[0]), 
        .A1N(n757), .Y(n1168) );
  AOI22X1TS U960 ( .A0(n745), .A1(n759), .B0(prevRequesterAddress_B[3]), .B1(
        n764), .Y(n760) );
  AOI211XLTS U961 ( .A0(n793), .A1(n794), .B0(n770), .C0(n759), .Y(n767) );
  OAI2BB2XLTS U962 ( .B0(n761), .B1(n760), .A0N(requesterAddressOut_EAST[3]), 
        .A1N(n767), .Y(n1167) );
  INVX2TS U963 ( .A(n762), .Y(n778) );
  AOI22X1TS U964 ( .A0(n750), .A1(n418), .B0(prevRequesterAddress_B[2]), .B1(
        n764), .Y(n763) );
  OAI2BB2XLTS U965 ( .B0(n778), .B1(n763), .A0N(requesterAddressOut_EAST[2]), 
        .A1N(n767), .Y(n1166) );
  CLKBUFX2TS U966 ( .A(n764), .Y(n766) );
  AOI22X1TS U967 ( .A0(prevRequesterAddress_A[1]), .A1(n418), .B0(
        prevRequesterAddress_B[1]), .B1(n766), .Y(n765) );
  OAI2BB2XLTS U968 ( .B0(n778), .B1(n765), .A0N(requesterAddressOut_EAST[1]), 
        .A1N(n767), .Y(n1165) );
  AOI22X1TS U969 ( .A0(prevRequesterAddress_A[0]), .A1(n418), .B0(
        prevRequesterAddress_B[0]), .B1(n766), .Y(n768) );
  OAI2BB2XLTS U970 ( .B0(n778), .B1(n768), .A0N(requesterAddressOut_EAST[0]), 
        .A1N(n767), .Y(n1164) );
  AOI22X1TS U971 ( .A0(prevRequesterAddress_A[3]), .A1(n13), .B0(
        prevRequesterAddress_B[3]), .B1(n769), .Y(n771) );
  NOR3XLTS U972 ( .A(n770), .B(n775), .C(n769), .Y(n776) );
  OAI2BB2XLTS U973 ( .B0(n774), .B1(n771), .A0N(requesterAddressOut_SOUTH[3]), 
        .A1N(n776), .Y(n1163) );
  AOI22X1TS U974 ( .A0(prevRequesterAddress_A[2]), .A1(n13), .B0(
        prevRequesterAddress_B[2]), .B1(n769), .Y(n772) );
  OAI2BB2XLTS U975 ( .B0(n774), .B1(n772), .A0N(requesterAddressOut_SOUTH[2]), 
        .A1N(n776), .Y(n1162) );
  AOI22X1TS U976 ( .A0(n752), .A1(n13), .B0(prevRequesterAddress_B[1]), .B1(
        n417), .Y(n773) );
  OAI2BB2XLTS U977 ( .B0(n774), .B1(n773), .A0N(requesterAddressOut_SOUTH[1]), 
        .A1N(n776), .Y(n1161) );
  AOI22X1TS U978 ( .A0(n756), .A1(n13), .B0(prevRequesterAddress_B[0]), .B1(
        n417), .Y(n777) );
  OAI2BB2XLTS U979 ( .B0(n778), .B1(n777), .A0N(requesterAddressOut_SOUTH[0]), 
        .A1N(n776), .Y(n1160) );
endmodule


module outputPortArbiter_0 ( clk, reset, selectBit_NORTH, 
        destinationAddressIn_NORTH, requesterAddressIn_NORTH, readIn_NORTH, 
        writeIn_NORTH, dataIn_NORTH, selectBit_SOUTH, 
        destinationAddressIn_SOUTH, requesterAddressIn_SOUTH, readIn_SOUTH, 
        writeIn_SOUTH, dataIn_SOUTH, selectBit_EAST, destinationAddressIn_EAST, 
        requesterAddressIn_EAST, readIn_EAST, writeIn_EAST, dataIn_EAST, 
        selectBit_WEST, destinationAddressIn_WEST, requesterAddressIn_WEST, 
        readIn_WEST, writeIn_WEST, dataIn_WEST, readReady, 
        readRequesterAddress, cacheDataOut, destinationAddressOut, 
        requesterAddressOut, readOut, writeOut, dataOut );
  input [11:0] destinationAddressIn_NORTH;
  input [3:0] requesterAddressIn_NORTH;
  input [5:0] dataIn_NORTH;
  input [11:0] destinationAddressIn_SOUTH;
  input [3:0] requesterAddressIn_SOUTH;
  input [5:0] dataIn_SOUTH;
  input [11:0] destinationAddressIn_EAST;
  input [3:0] requesterAddressIn_EAST;
  input [5:0] dataIn_EAST;
  input [11:0] destinationAddressIn_WEST;
  input [3:0] requesterAddressIn_WEST;
  input [5:0] dataIn_WEST;
  input [3:0] readRequesterAddress;
  input [5:0] cacheDataOut;
  output [11:0] destinationAddressOut;
  output [3:0] requesterAddressOut;
  output [5:0] dataOut;
  input clk, reset, selectBit_NORTH, readIn_NORTH, writeIn_NORTH,
         selectBit_SOUTH, readIn_SOUTH, writeIn_SOUTH, selectBit_EAST,
         readIn_EAST, writeIn_EAST, selectBit_WEST, readIn_WEST, writeIn_WEST,
         readReady;
  output readOut, writeOut;
  wire   \requesterAddressbuffer[0][3] , \requesterAddressbuffer[0][2] ,
         \requesterAddressbuffer[0][1] , \requesterAddressbuffer[0][0] ,
         \requesterAddressbuffer[1][3] , \requesterAddressbuffer[1][2] ,
         \requesterAddressbuffer[1][1] , \requesterAddressbuffer[1][0] ,
         \requesterAddressbuffer[2][3] , \requesterAddressbuffer[2][2] ,
         \requesterAddressbuffer[2][1] , \requesterAddressbuffer[2][0] ,
         \requesterAddressbuffer[3][3] , \requesterAddressbuffer[3][2] ,
         \requesterAddressbuffer[3][1] , \requesterAddressbuffer[3][0] ,
         \requesterAddressbuffer[4][3] , \requesterAddressbuffer[4][2] ,
         \requesterAddressbuffer[4][1] , \requesterAddressbuffer[4][0] ,
         \requesterAddressbuffer[5][3] , \requesterAddressbuffer[5][2] ,
         \requesterAddressbuffer[5][1] , \requesterAddressbuffer[5][0] ,
         \requesterAddressbuffer[6][3] , \requesterAddressbuffer[6][2] ,
         \requesterAddressbuffer[6][1] , \requesterAddressbuffer[6][0] ,
         \requesterAddressbuffer[7][3] , \requesterAddressbuffer[7][2] ,
         \requesterAddressbuffer[7][1] , \requesterAddressbuffer[7][0] ,
         \destinationAddressbuffer[0][11] , \destinationAddressbuffer[0][10] ,
         \destinationAddressbuffer[0][9] , \destinationAddressbuffer[0][8] ,
         \destinationAddressbuffer[0][7] , \destinationAddressbuffer[0][6] ,
         \destinationAddressbuffer[0][5] , \destinationAddressbuffer[0][4] ,
         \destinationAddressbuffer[0][3] , \destinationAddressbuffer[0][2] ,
         \destinationAddressbuffer[0][1] , \destinationAddressbuffer[0][0] ,
         \destinationAddressbuffer[1][11] , \destinationAddressbuffer[1][10] ,
         \destinationAddressbuffer[1][9] , \destinationAddressbuffer[1][8] ,
         \destinationAddressbuffer[1][7] , \destinationAddressbuffer[1][6] ,
         \destinationAddressbuffer[1][5] , \destinationAddressbuffer[1][4] ,
         \destinationAddressbuffer[1][3] , \destinationAddressbuffer[1][2] ,
         \destinationAddressbuffer[1][1] , \destinationAddressbuffer[1][0] ,
         \destinationAddressbuffer[2][11] , \destinationAddressbuffer[2][10] ,
         \destinationAddressbuffer[2][9] , \destinationAddressbuffer[2][8] ,
         \destinationAddressbuffer[2][7] , \destinationAddressbuffer[2][6] ,
         \destinationAddressbuffer[2][5] , \destinationAddressbuffer[2][4] ,
         \destinationAddressbuffer[2][3] , \destinationAddressbuffer[2][2] ,
         \destinationAddressbuffer[2][1] , \destinationAddressbuffer[2][0] ,
         \destinationAddressbuffer[3][11] , \destinationAddressbuffer[3][10] ,
         \destinationAddressbuffer[3][9] , \destinationAddressbuffer[3][8] ,
         \destinationAddressbuffer[3][7] , \destinationAddressbuffer[3][6] ,
         \destinationAddressbuffer[3][5] , \destinationAddressbuffer[3][4] ,
         \destinationAddressbuffer[3][3] , \destinationAddressbuffer[3][2] ,
         \destinationAddressbuffer[3][1] , \destinationAddressbuffer[3][0] ,
         \destinationAddressbuffer[4][11] , \destinationAddressbuffer[4][10] ,
         \destinationAddressbuffer[4][9] , \destinationAddressbuffer[4][8] ,
         \destinationAddressbuffer[4][7] , \destinationAddressbuffer[4][6] ,
         \destinationAddressbuffer[4][5] , \destinationAddressbuffer[4][4] ,
         \destinationAddressbuffer[4][3] , \destinationAddressbuffer[4][2] ,
         \destinationAddressbuffer[4][1] , \destinationAddressbuffer[4][0] ,
         \destinationAddressbuffer[5][11] , \destinationAddressbuffer[5][10] ,
         \destinationAddressbuffer[5][9] , \destinationAddressbuffer[5][8] ,
         \destinationAddressbuffer[5][7] , \destinationAddressbuffer[5][6] ,
         \destinationAddressbuffer[5][5] , \destinationAddressbuffer[5][4] ,
         \destinationAddressbuffer[5][3] , \destinationAddressbuffer[5][2] ,
         \destinationAddressbuffer[5][1] , \destinationAddressbuffer[5][0] ,
         \destinationAddressbuffer[6][11] , \destinationAddressbuffer[6][10] ,
         \destinationAddressbuffer[6][9] , \destinationAddressbuffer[6][8] ,
         \destinationAddressbuffer[6][7] , \destinationAddressbuffer[6][6] ,
         \destinationAddressbuffer[6][5] , \destinationAddressbuffer[6][4] ,
         \destinationAddressbuffer[6][3] , \destinationAddressbuffer[6][2] ,
         \destinationAddressbuffer[6][1] , \destinationAddressbuffer[6][0] ,
         \destinationAddressbuffer[7][11] , \destinationAddressbuffer[7][10] ,
         \destinationAddressbuffer[7][9] , \destinationAddressbuffer[7][8] ,
         \destinationAddressbuffer[7][7] , \destinationAddressbuffer[7][6] ,
         \destinationAddressbuffer[7][5] , \destinationAddressbuffer[7][4] ,
         \destinationAddressbuffer[7][3] , \destinationAddressbuffer[7][2] ,
         \destinationAddressbuffer[7][1] , \destinationAddressbuffer[7][0] ,
         \dataoutbuffer[7][5] , \dataoutbuffer[7][4] , \dataoutbuffer[7][3] ,
         \dataoutbuffer[7][2] , \dataoutbuffer[7][1] , \dataoutbuffer[7][0] ,
         \dataoutbuffer[6][5] , \dataoutbuffer[6][4] , \dataoutbuffer[6][3] ,
         \dataoutbuffer[6][2] , \dataoutbuffer[6][1] , \dataoutbuffer[6][0] ,
         \dataoutbuffer[5][5] , \dataoutbuffer[5][4] , \dataoutbuffer[5][3] ,
         \dataoutbuffer[5][2] , \dataoutbuffer[5][1] , \dataoutbuffer[5][0] ,
         \dataoutbuffer[4][5] , \dataoutbuffer[4][4] , \dataoutbuffer[4][3] ,
         \dataoutbuffer[4][2] , \dataoutbuffer[4][1] , \dataoutbuffer[4][0] ,
         \dataoutbuffer[3][5] , \dataoutbuffer[3][4] , \dataoutbuffer[3][3] ,
         \dataoutbuffer[3][2] , \dataoutbuffer[3][1] , \dataoutbuffer[3][0] ,
         \dataoutbuffer[2][5] , \dataoutbuffer[2][4] , \dataoutbuffer[2][3] ,
         \dataoutbuffer[2][2] , \dataoutbuffer[2][1] , \dataoutbuffer[2][0] ,
         \dataoutbuffer[1][5] , \dataoutbuffer[1][4] , \dataoutbuffer[1][3] ,
         \dataoutbuffer[1][2] , \dataoutbuffer[1][1] , \dataoutbuffer[1][0] ,
         \dataoutbuffer[0][5] , \dataoutbuffer[0][4] , \dataoutbuffer[0][3] ,
         \dataoutbuffer[0][2] , \dataoutbuffer[0][1] , \dataoutbuffer[0][0] ,
         N2624, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1904, n1905, n1906, n1907,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926;
  wire   [0:7] writeOutbuffer;
  wire   [0:7] readOutbuffer;

  DFFNSRX1TS full_reg_reg ( .D(N2624), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(
        n1918) );
  DFFNSRX1TS \dataoutbuffer_reg[0][0]  ( .D(n1273), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][1]  ( .D(n1272), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][2]  ( .D(n1271), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][3]  ( .D(n1270), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][4]  ( .D(n1269), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][5]  ( .D(n1268), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][5] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[2][0]  ( .D(n1285), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[2][1]  ( .D(n1284), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[2][2]  ( .D(n1283), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[2][3]  ( .D(n1282), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][0]  ( .D(n1149), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][1]  ( .D(n1148), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][2]  ( .D(n1147), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][3]  ( .D(n1146), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][3] ) );
  DFFNSRX1TS \writeOutbuffer_reg[7]  ( .D(n1225), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[7]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][4]  ( .D(n1205), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][5]  ( .D(n1204), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][6]  ( .D(n1203), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][7]  ( .D(n1202), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][8]  ( .D(n1201), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][9]  ( .D(n1200), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][11]  ( .D(n1198), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[6]  ( .D(n1224), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[6]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][4]  ( .D(n1193), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][5]  ( .D(n1192), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][6]  ( .D(n1191), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][7]  ( .D(n1190), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][8]  ( .D(n1189), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][9]  ( .D(n1188), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][10]  ( .D(n1187), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][11]  ( .D(n1186), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[3]  ( .D(n1221), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[3]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][4]  ( .D(n1157), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][5]  ( .D(n1156), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][6]  ( .D(n1155), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][7]  ( .D(n1154), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][8]  ( .D(n1153), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][9]  ( .D(n1152), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][10]  ( .D(n1151), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][11]  ( .D(n1150), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[2]  ( .D(n1220), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[2]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][4]  ( .D(n1145), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][5]  ( .D(n1144), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][6]  ( .D(n1143), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][7]  ( .D(n1142), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][8]  ( .D(n1141), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][9]  ( .D(n1140), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][10]  ( .D(n1139), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][11]  ( .D(n1138), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][11] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][0]  ( .D(n1231), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][1]  ( .D(n1230), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][2]  ( .D(n1229), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][3]  ( .D(n1228), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][4]  ( .D(n1227), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][5]  ( .D(n1226), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][0]  ( .D(n1237), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][1]  ( .D(n1236), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][2]  ( .D(n1235), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][3]  ( .D(n1234), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][4]  ( .D(n1233), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][5]  ( .D(n1232), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][0]  ( .D(n1255), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][1]  ( .D(n1254), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][2]  ( .D(n1253), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][3]  ( .D(n1252), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][4]  ( .D(n1251), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][5]  ( .D(n1250), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][0]  ( .D(n1261), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][1]  ( .D(n1260), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][2]  ( .D(n1259), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][3]  ( .D(n1258), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][4]  ( .D(n1257), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][5]  ( .D(n1256), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][5] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[5][0]  ( .D(n1297), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[5][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[5][1]  ( .D(n1296), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[5][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[5][2]  ( .D(n1295), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[5][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[5][3]  ( .D(n1294), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[5][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][0]  ( .D(n1185), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][1]  ( .D(n1184), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][2]  ( .D(n1183), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][3]  ( .D(n1182), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[4][0]  ( .D(n1293), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[4][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[4][1]  ( .D(n1292), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[4][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[4][2]  ( .D(n1291), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[4][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[4][3]  ( .D(n1290), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[4][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][0]  ( .D(n1173), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][1]  ( .D(n1172), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][2]  ( .D(n1171), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][3]  ( .D(n1170), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[1][0]  ( .D(n1281), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[1][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[1][1]  ( .D(n1280), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[1][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[1][2]  ( .D(n1279), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[1][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[1][3]  ( .D(n1278), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[1][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][0]  ( .D(n1137), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][1]  ( .D(n1136), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][2]  ( .D(n1135), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][3]  ( .D(n1134), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[0][0]  ( .D(n1277), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[0][1]  ( .D(n1276), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[0][2]  ( .D(n1275), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[0][3]  ( .D(n1274), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][0]  ( .D(n1125), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][1]  ( .D(n1124), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][2]  ( .D(n1123), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][3]  ( .D(n1122), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][0]  ( .D(n1243), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][1]  ( .D(n1242), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][2]  ( .D(n1241), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][3]  ( .D(n1240), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][4]  ( .D(n1239), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][5]  ( .D(n1238), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][0]  ( .D(n1249), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][1]  ( .D(n1248), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][2]  ( .D(n1247), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][3]  ( .D(n1246), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][4]  ( .D(n1245), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][5]  ( .D(n1244), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][0]  ( .D(n1267), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][1]  ( .D(n1266), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][2]  ( .D(n1265), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][3]  ( .D(n1264), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][4]  ( .D(n1263), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][5]  ( .D(n1262), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][5] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[7][0]  ( .D(n1305), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[7][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[7][1]  ( .D(n1304), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[7][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[7][2]  ( .D(n1303), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[7][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[7][3]  ( .D(n1302), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[7][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][0]  ( .D(n1209), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][1]  ( .D(n1208), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][2]  ( .D(n1207), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][3]  ( .D(n1206), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[6][0]  ( .D(n1301), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[6][1]  ( .D(n1300), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[6][2]  ( .D(n1299), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[6][3]  ( .D(n1298), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][0]  ( .D(n1197), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][1]  ( .D(n1196), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][2]  ( .D(n1195), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][3]  ( .D(n1194), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[3][0]  ( .D(n1289), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[3][1]  ( .D(n1288), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[3][2]  ( .D(n1287), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[3][3]  ( .D(n1286), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][0]  ( .D(n1161), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][1]  ( .D(n1160), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][2]  ( .D(n1159), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][3]  ( .D(n1158), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][3] ) );
  DFFNSRX1TS \writeOutbuffer_reg[5]  ( .D(n1223), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[5]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][4]  ( .D(n1181), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][5]  ( .D(n1180), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][6]  ( .D(n1179), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][7]  ( .D(n1178), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][8]  ( .D(n1177), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][9]  ( .D(n1176), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][10]  ( .D(n1175), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][11]  ( .D(n1174), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[4]  ( .D(n1222), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[4]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][4]  ( .D(n1169), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][5]  ( .D(n1168), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][6]  ( .D(n1167), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][7]  ( .D(n1166), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][8]  ( .D(n1165), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][9]  ( .D(n1164), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][10]  ( .D(n1163), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][11]  ( .D(n1162), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[1]  ( .D(n1219), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[1]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][4]  ( .D(n1133), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][5]  ( .D(n1132), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][6]  ( .D(n1131), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][7]  ( .D(n1130), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][8]  ( .D(n1129), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][9]  ( .D(n1128), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][10]  ( .D(n1127), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][11]  ( .D(n1126), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[0]  ( .D(n1218), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[0]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][4]  ( .D(n1121), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][5]  ( .D(n1120), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][6]  ( .D(n1119), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][7]  ( .D(n1118), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][8]  ( .D(n1117), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][9]  ( .D(n1116), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][10]  ( .D(n1115), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][11]  ( .D(n1114), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][11] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][10]  ( .D(n1199), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][10] ) );
  DFFNSRX1TS writeOut_reg ( .D(n1328), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        writeOut) );
  DFFNSRX1TS \destinationAddressOut_reg[4]  ( .D(n1319), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[4]) );
  DFFNSRX1TS \destinationAddressOut_reg[5]  ( .D(n1318), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[5]) );
  DFFNSRX1TS \destinationAddressOut_reg[6]  ( .D(n1317), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[6]) );
  DFFNSRX1TS \destinationAddressOut_reg[7]  ( .D(n1316), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[7]) );
  DFFNSRX1TS \destinationAddressOut_reg[8]  ( .D(n1315), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[8]) );
  DFFNSRX1TS \destinationAddressOut_reg[9]  ( .D(n1314), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[9]) );
  DFFNSRX1TS \destinationAddressOut_reg[10]  ( .D(n1313), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[10]) );
  DFFNSRX1TS \destinationAddressOut_reg[11]  ( .D(n1312), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[11]) );
  DFFNSRX1TS readOut_reg ( .D(n1329), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        readOut) );
  DFFNSRX1TS \requesterAddressOut_reg[0]  ( .D(n1327), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[0]) );
  DFFNSRX1TS \requesterAddressOut_reg[1]  ( .D(n1326), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[1]) );
  DFFNSRX1TS \requesterAddressOut_reg[2]  ( .D(n1325), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[2]) );
  DFFNSRX1TS \requesterAddressOut_reg[3]  ( .D(n1324), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[3]) );
  DFFNSRX1TS \destinationAddressOut_reg[0]  ( .D(n1323), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[0]) );
  DFFNSRX1TS \destinationAddressOut_reg[1]  ( .D(n1322), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[1]) );
  DFFNSRX1TS \destinationAddressOut_reg[2]  ( .D(n1321), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[2]) );
  DFFNSRX1TS \destinationAddressOut_reg[3]  ( .D(n1320), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[3]) );
  DFFNSRX1TS \dataOut_reg[0]  ( .D(n1311), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[0]) );
  DFFNSRX1TS \dataOut_reg[1]  ( .D(n1310), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[1]) );
  DFFNSRX1TS \dataOut_reg[2]  ( .D(n1309), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[2]) );
  DFFNSRX1TS \dataOut_reg[3]  ( .D(n1308), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[3]) );
  DFFNSRX1TS \dataOut_reg[4]  ( .D(n1307), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[4]) );
  DFFNSRX1TS \dataOut_reg[5]  ( .D(n1306), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[5]) );
  DFFNSRX1TS \read_reg_reg[1]  ( .D(n1330), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1911), .QN(n1910) );
  DFFNSRX1TS \write_reg_reg[0]  ( .D(n1335), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1909), .QN(n1913) );
  DFFNSRX1TS \write_reg_reg[2]  ( .D(n1333), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1914), .QN(n1915) );
  DFFNSRX1TS \read_reg_reg[0]  ( .D(n1336), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1904), .QN(n1917) );
  DFFNSRX1TS \read_reg_reg[2]  ( .D(n1331), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1907), .QN(n1908) );
  DFFNSRX1TS empty_reg_reg ( .D(n1332), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        n1906), .QN(n1905) );
  DFFNSRX1TS \readOutbuffer_reg[7]  ( .D(n1217), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[7]), .QN(n1919) );
  DFFNSRX1TS \readOutbuffer_reg[4]  ( .D(n1214), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[4]), .QN(n1922) );
  DFFNSRX1TS \readOutbuffer_reg[6]  ( .D(n1216), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[6]), .QN(n1920) );
  DFFNSRX1TS \readOutbuffer_reg[5]  ( .D(n1215), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[5]), .QN(n1921) );
  DFFNSRX1TS \readOutbuffer_reg[3]  ( .D(n1213), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[3]), .QN(n1923) );
  DFFNSRX1TS \readOutbuffer_reg[2]  ( .D(n1212), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[2]), .QN(n1924) );
  DFFNSRX1TS \readOutbuffer_reg[0]  ( .D(n1210), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[0]), .QN(n1926) );
  DFFNSRX1TS \readOutbuffer_reg[1]  ( .D(n1211), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[1]), .QN(n1925) );
  DFFNSRX1TS \write_reg_reg[1]  ( .D(n1334), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1912), .QN(n1916) );
  CMPR32X2TS U3 ( .A(n474), .B(n485), .C(n473), .CO(n468), .S(n492) );
  NAND2BX1TS U4 ( .AN(n122), .B(selectBit_WEST), .Y(n379) );
  CMPR32X2TS U5 ( .A(n453), .B(n482), .C(n16), .CO(n17), .S(n14) );
  CMPR32X2TS U6 ( .A(n529), .B(n451), .C(n454), .CO(n443), .S(n456) );
  CLKBUFX2TS U7 ( .A(n20), .Y(n80) );
  ADDHXLTS U8 ( .A(n440), .B(n449), .CO(n16), .S(n15) );
  CLKBUFX2TS U9 ( .A(n18), .Y(n19) );
  AO21X2TS U10 ( .A0(n448), .A1(n503), .B0(n19), .Y(n21) );
  INVX2TS U11 ( .A(n8), .Y(n222) );
  OAI31X1TS U12 ( .A0(n515), .A1(n514), .A2(n536), .B0(n537), .Y(n517) );
  OR2X1TS U13 ( .A(n21), .B(n505), .Y(n9) );
  NOR2XLTS U14 ( .A(n1589), .B(n1586), .Y(n129) );
  NOR2XLTS U15 ( .A(n124), .B(n381), .Y(n1586) );
  NOR3XLTS U16 ( .A(n382), .B(n270), .C(n181), .Y(n1555) );
  CLKBUFX2TS U17 ( .A(n14), .Y(n78) );
  NAND2X1TS U18 ( .A(n537), .B(n519), .Y(n507) );
  NOR2XLTS U19 ( .A(n838), .B(n516), .Y(n542) );
  NOR2XLTS U20 ( .A(n838), .B(n518), .Y(n687) );
  INVX2TS U21 ( .A(n1567), .Y(n1565) );
  INVX2TS U22 ( .A(n141), .Y(n951) );
  INVX2TS U23 ( .A(n1545), .Y(n1543) );
  INVX2TS U24 ( .A(n1625), .Y(n1622) );
  INVX2TS U25 ( .A(n1614), .Y(n1611) );
  NOR3XLTS U26 ( .A(n15), .B(n180), .C(n379), .Y(n1600) );
  INVX2TS U27 ( .A(n1558), .Y(n1556) );
  AOI31XLTS U28 ( .A0(n33), .A1(n28), .A2(n1541), .B0(n81), .Y(n31) );
  NOR2XLTS U29 ( .A(n1607), .B(n323), .Y(n321) );
  NOR2XLTS U30 ( .A(n1542), .B(n36), .Y(n40) );
  NOR3XLTS U31 ( .A(n1614), .B(n1608), .C(n320), .Y(n315) );
  CLKBUFX2TS U32 ( .A(n1084), .Y(n1079) );
  NOR2XLTS U33 ( .A(n1564), .B(n229), .Y(n228) );
  NOR2XLTS U34 ( .A(n480), .B(n1590), .Y(n132) );
  NOR2XLTS U35 ( .A(n81), .B(n1559), .Y(n84) );
  NOR3XLTS U36 ( .A(n1600), .B(n1594), .C(n188), .Y(n183) );
  NOR2XLTS U37 ( .A(n1551), .B(n89), .Y(n90) );
  NOR3XLTS U38 ( .A(n1548), .B(n1543), .C(n34), .Y(n29) );
  NOR2XLTS U39 ( .A(n480), .B(n1601), .Y(n184) );
  NOR2XLTS U40 ( .A(n1592), .B(n189), .Y(n190) );
  NOR3XLTS U41 ( .A(n1629), .B(n1622), .C(n394), .Y(n389) );
  NOR3XLTS U42 ( .A(n1570), .B(n1565), .C(n227), .Y(n1) );
  OAI211XLTS U43 ( .A0(n221), .A1(n236), .B0(n200), .C0(n199), .Y(n1140) );
  NOR2X1TS U44 ( .A(n1593), .B(n189), .Y(n198) );
  NOR2X1TS U45 ( .A(n24), .B(n134), .Y(n130) );
  NAND2BX1TS U46 ( .AN(n320), .B(n319), .Y(n323) );
  NAND2BX1TS U47 ( .AN(n278), .B(n277), .Y(n279) );
  NAND2BX1TS U48 ( .AN(n136), .B(n129), .Y(n134) );
  NOR2X1TS U49 ( .A(n1587), .B(n136), .Y(n137) );
  NAND2BXLTS U50 ( .AN(n87), .B(n86), .Y(n89) );
  AOI31X1TS U51 ( .A0(n226), .A1(n1561), .A2(n224), .B0(n390), .Y(n225) );
  AOI31X1TS U52 ( .A0(n129), .A1(n24), .A2(n127), .B0(n390), .Y(n133) );
  NOR2X1TS U53 ( .A(n1548), .B(n1545), .Y(n33) );
  NOR2X1TS U54 ( .A(n1581), .B(n1577), .Y(n277) );
  INVX1TS U55 ( .A(n1610), .Y(n1608) );
  INVX1TS U56 ( .A(n1597), .Y(n1594) );
  NOR2X1TS U57 ( .A(n124), .B(n270), .Y(n1545) );
  NOR3X1TS U58 ( .A(n383), .B(n80), .C(n272), .Y(n1574) );
  NOR3X1TS U59 ( .A(n384), .B(n383), .C(n80), .Y(n1621) );
  OAI21X1TS U60 ( .A0(selectBit_SOUTH), .A1(n21), .B0(n80), .Y(n380) );
  NOR3X1TS U61 ( .A(n272), .B(n80), .C(n222), .Y(n1552) );
  NAND3X1TS U62 ( .A(n384), .B(n223), .C(n222), .Y(n1561) );
  NOR3X1TS U63 ( .A(n26), .B(n383), .C(n9), .Y(n1607) );
  AND2X2TS U64 ( .A(n25), .B(n79), .Y(n23) );
  NAND3X1TS U65 ( .A(n493), .B(n384), .C(n223), .Y(n1541) );
  INVX1TS U66 ( .A(n1589), .Y(n1587) );
  NOR3X1TS U67 ( .A(n384), .B(n20), .C(n222), .Y(n1593) );
  INVX1TS U68 ( .A(n1600), .Y(n1598) );
  NOR2X1TS U69 ( .A(n223), .B(n271), .Y(n311) );
  NOR2X1TS U70 ( .A(n9), .B(n271), .Y(n25) );
  INVX1TS U71 ( .A(n271), .Y(n383) );
  INVX1TS U72 ( .A(n1581), .Y(n1578) );
  INVX1TS U73 ( .A(n1629), .Y(n1626) );
  INVX1TS U74 ( .A(n8), .Y(n271) );
  NOR3X1TS U75 ( .A(n14), .B(n77), .C(n379), .Y(n1614) );
  INVX1TS U76 ( .A(n79), .Y(n26) );
  NOR3X1TS U77 ( .A(n78), .B(n121), .C(n269), .Y(n1581) );
  NOR3X1TS U78 ( .A(n78), .B(n15), .C(n379), .Y(n1629) );
  INVX1TS U79 ( .A(n22), .Y(n125) );
  NOR2X1TS U80 ( .A(selectBit_NORTH), .B(n504), .Y(n537) );
  CLKBUFX2TS U81 ( .A(n53), .Y(n295) );
  NOR2X1TS U82 ( .A(n448), .B(n503), .Y(n18) );
  CLKBUFX2TS U83 ( .A(readIn_EAST), .Y(n1540) );
  INVX1TS U84 ( .A(n1915), .Y(n497) );
  NOR3BX1TS U85 ( .AN(n382), .B(n270), .C(n380), .Y(n1577) );
  CLKINVX1TS U86 ( .A(n1570), .Y(n1568) );
  INVX2TS U87 ( .A(n464), .Y(n461) );
  XOR2X1TS U88 ( .A(n471), .B(n470), .Y(n494) );
  INVX2TS U89 ( .A(n322), .Y(n344) );
  INVX2TS U90 ( .A(n228), .Y(n254) );
  NAND2X1TS U91 ( .A(n133), .B(n1590), .Y(n136) );
  NAND2BX1TS U92 ( .AN(n188), .B(n187), .Y(n189) );
  CLKAND2X2TS U93 ( .A(n467), .B(n466), .Y(n473) );
  NAND4XLTS U94 ( .A(n493), .B(n508), .C(n388), .D(n484), .Y(n1601) );
  INVX2TS U95 ( .A(n1593), .Y(n1592) );
  NAND4XLTS U96 ( .A(n482), .B(n1909), .C(n508), .D(n484), .Y(n1590) );
  NOR3XLTS U97 ( .A(n14), .B(n77), .C(n269), .Y(n1570) );
  NAND4XLTS U98 ( .A(n485), .B(n1914), .C(n513), .D(n388), .Y(n1559) );
  NOR3XLTS U99 ( .A(n15), .B(n180), .C(n269), .Y(n1558) );
  INVX2TS U100 ( .A(n1555), .Y(n1553) );
  NAND4XLTS U101 ( .A(n497), .B(n510), .C(n388), .D(n313), .Y(n1582) );
  INVX2TS U102 ( .A(n1577), .Y(n1575) );
  INVX2TS U103 ( .A(n1541), .Y(n1542) );
  CLKAND2X2TS U104 ( .A(n522), .B(n520), .Y(n549) );
  INVX2TS U105 ( .A(n1420), .Y(n1450) );
  INVX2TS U106 ( .A(selectBit_NORTH), .Y(n503) );
  NOR2XLTS U107 ( .A(n1629), .B(n1625), .Y(n393) );
  NOR3BXLTS U108 ( .AN(n513), .B(n450), .C(n512), .Y(n536) );
  NAND3XLTS U109 ( .A(n504), .B(n506), .C(n503), .Y(n516) );
  NAND3XLTS U110 ( .A(selectBit_NORTH), .B(n506), .C(n505), .Y(n518) );
  NOR2XLTS U111 ( .A(n1614), .B(n1610), .Y(n319) );
  NOR2XLTS U112 ( .A(n1570), .B(n1567), .Y(n226) );
  NOR2XLTS U113 ( .A(n1558), .B(n1555), .Y(n86) );
  NOR2XLTS U114 ( .A(n1600), .B(n1597), .Y(n187) );
  NAND2BXLTS U115 ( .AN(n394), .B(n393), .Y(n395) );
  XOR2XLTS U116 ( .A(n443), .B(n445), .Y(n462) );
  OAI21XLTS U117 ( .A0(n446), .A1(n1910), .B0(n445), .Y(n447) );
  NAND2BXLTS U118 ( .AN(n123), .B(selectBit_EAST), .Y(n381) );
  NAND3XLTS U119 ( .A(n19), .B(n442), .C(n387), .Y(n224) );
  XOR2X1TS U120 ( .A(n497), .B(n17), .Y(n122) );
  NOR2XLTS U121 ( .A(n131), .B(reset), .Y(n496) );
  NAND4XLTS U122 ( .A(n491), .B(n508), .C(n441), .D(n387), .Y(n1615) );
  INVX2TS U123 ( .A(n1607), .Y(n1604) );
  NOR3XLTS U124 ( .A(n312), .B(n311), .C(n381), .Y(n1610) );
  NAND4XLTS U125 ( .A(readReady), .B(n388), .C(n387), .D(n481), .Y(n1630) );
  INVX2TS U126 ( .A(n1621), .Y(n1618) );
  NOR3BXLTS U127 ( .AN(n382), .B(n381), .C(n380), .Y(n1625) );
  NOR3X1TS U128 ( .A(n180), .B(n77), .C(n379), .Y(n1589) );
  INVX2TS U129 ( .A(n1586), .Y(n1584) );
  NAND4XLTS U130 ( .A(n491), .B(n497), .C(n513), .D(n313), .Y(n1571) );
  NOR3XLTS U131 ( .A(n312), .B(n311), .C(n270), .Y(n1567) );
  INVX2TS U132 ( .A(n1552), .Y(n1551) );
  INVX2TS U133 ( .A(n1574), .Y(n1573) );
  NAND4XLTS U134 ( .A(n78), .B(n121), .C(n122), .D(selectBit_WEST), .Y(n1546)
         );
  NAND4XLTS U135 ( .A(n1909), .B(n485), .C(n469), .D(readReady), .Y(n1549) );
  INVX2TS U136 ( .A(n1420), .Y(n264) );
  INVX2TS U137 ( .A(destinationAddressIn_SOUTH[11]), .Y(n168) );
  INVX2TS U138 ( .A(destinationAddressIn_SOUTH[10]), .Y(n174) );
  INVX2TS U139 ( .A(destinationAddressIn_SOUTH[9]), .Y(n160) );
  INVX2TS U140 ( .A(destinationAddressIn_SOUTH[8]), .Y(n164) );
  CLKAND2X2TS U141 ( .A(n467), .B(n465), .Y(n472) );
  NOR2XLTS U142 ( .A(reset), .B(n438), .Y(n495) );
  AO22XLTS U143 ( .A0(n497), .A1(n496), .B0(n495), .B1(n494), .Y(n1333) );
  AO22XLTS U144 ( .A0(n491), .A1(n496), .B0(n495), .B1(n490), .Y(n1335) );
  AO22XLTS U145 ( .A0(n493), .A1(n496), .B0(n495), .B1(n492), .Y(n1334) );
  OAI21XLTS U146 ( .A0(n131), .A1(n488), .B0(n489), .Y(n1332) );
  NAND4XLTS U147 ( .A(n864), .B(n863), .C(n862), .D(n861), .Y(n1306) );
  NAND4XLTS U148 ( .A(n842), .B(n841), .C(n840), .D(n861), .Y(n1307) );
  NAND4XLTS U149 ( .A(n831), .B(n830), .C(n829), .D(n861), .Y(n1308) );
  NAND4XLTS U150 ( .A(n821), .B(n820), .C(n819), .D(n861), .Y(n1309) );
  NAND4XLTS U151 ( .A(n802), .B(n801), .C(n800), .D(n799), .Y(n1310) );
  NAND4XLTS U152 ( .A(n782), .B(n781), .C(n780), .D(n799), .Y(n1311) );
  NAND4XLTS U153 ( .A(n653), .B(n652), .C(n651), .D(n650), .Y(n1320) );
  NAND4XLTS U154 ( .A(n642), .B(n641), .C(n640), .D(n639), .Y(n1321) );
  NAND4XLTS U155 ( .A(n624), .B(n623), .C(n622), .D(n621), .Y(n1322) );
  NAND4XLTS U156 ( .A(n609), .B(n608), .C(n607), .D(n606), .Y(n1323) );
  NAND4XLTS U157 ( .A(n597), .B(n596), .C(n595), .D(n650), .Y(n1324) );
  NAND4XLTS U158 ( .A(n586), .B(n585), .C(n584), .D(n639), .Y(n1325) );
  NAND4XLTS U159 ( .A(n577), .B(n576), .C(n575), .D(n621), .Y(n1326) );
  NAND4XLTS U160 ( .A(n560), .B(n559), .C(n558), .D(n606), .Y(n1327) );
  NAND4XLTS U161 ( .A(n540), .B(n539), .C(n538), .D(n799), .Y(n1329) );
  NAND3XLTS U162 ( .A(n772), .B(n771), .C(n770), .Y(n1312) );
  NAND3XLTS U163 ( .A(n758), .B(n757), .C(n756), .Y(n1313) );
  NAND3XLTS U164 ( .A(n742), .B(n741), .C(n740), .Y(n1314) );
  NAND3XLTS U165 ( .A(n724), .B(n723), .C(n722), .Y(n1315) );
  NAND3XLTS U166 ( .A(n710), .B(n709), .C(n708), .Y(n1316) );
  NAND3XLTS U167 ( .A(n699), .B(n698), .C(n697), .Y(n1317) );
  NAND3XLTS U168 ( .A(n685), .B(n684), .C(n683), .Y(n1318) );
  NAND3XLTS U169 ( .A(n664), .B(n663), .C(n662), .Y(n1319) );
  NAND3XLTS U170 ( .A(n552), .B(n551), .C(n550), .Y(n1328) );
  NAND3XLTS U171 ( .A(n1780), .B(n1779), .C(n1778), .Y(n1158) );
  NAND3XLTS U172 ( .A(n1771), .B(n1770), .C(n1769), .Y(n1159) );
  NAND3XLTS U173 ( .A(n1765), .B(n1764), .C(n1763), .Y(n1160) );
  NAND3XLTS U174 ( .A(n1759), .B(n1758), .C(n1757), .Y(n1161) );
  NAND3XLTS U175 ( .A(n968), .B(n967), .C(n966), .Y(n1286) );
  NAND3XLTS U176 ( .A(n962), .B(n961), .C(n960), .Y(n1287) );
  NAND3XLTS U177 ( .A(n955), .B(n954), .C(n953), .Y(n1288) );
  NAND3XLTS U178 ( .A(n949), .B(n948), .C(n947), .Y(n1289) );
  NAND3XLTS U179 ( .A(n1689), .B(n1688), .C(n1687), .Y(n1194) );
  NAND3XLTS U180 ( .A(n1681), .B(n1680), .C(n1679), .Y(n1195) );
  NAND3XLTS U181 ( .A(n1673), .B(n1672), .C(n1671), .Y(n1196) );
  NAND3XLTS U182 ( .A(n1667), .B(n1666), .C(n1665), .Y(n1197) );
  NAND3XLTS U183 ( .A(n900), .B(n899), .C(n898), .Y(n1298) );
  NAND3XLTS U184 ( .A(n892), .B(n891), .C(n890), .Y(n1299) );
  NAND3XLTS U185 ( .A(n888), .B(n887), .C(n886), .Y(n1300) );
  NAND3XLTS U186 ( .A(n884), .B(n883), .C(n882), .Y(n1301) );
  NAND3XLTS U187 ( .A(n1660), .B(n1659), .C(n1658), .Y(n1206) );
  NAND3XLTS U188 ( .A(n1651), .B(n1650), .C(n1649), .Y(n1207) );
  NAND3XLTS U189 ( .A(n1642), .B(n1641), .C(n1640), .Y(n1208) );
  NAND3XLTS U190 ( .A(n1635), .B(n1634), .C(n1633), .Y(n1209) );
  NAND3XLTS U191 ( .A(n881), .B(n880), .C(n879), .Y(n1302) );
  NAND3XLTS U192 ( .A(n876), .B(n875), .C(n874), .Y(n1303) );
  NAND3XLTS U193 ( .A(n871), .B(n870), .C(n869), .Y(n1304) );
  NAND3XLTS U194 ( .A(n867), .B(n866), .C(n865), .Y(n1305) );
  NAND3XLTS U195 ( .A(n1102), .B(n1101), .C(n1100), .Y(n1262) );
  NAND3XLTS U196 ( .A(n1098), .B(n1097), .C(n1096), .Y(n1263) );
  NAND3XLTS U197 ( .A(n1091), .B(n1090), .C(n1089), .Y(n1264) );
  NAND3XLTS U198 ( .A(n1087), .B(n1086), .C(n1085), .Y(n1265) );
  NAND3XLTS U199 ( .A(n1082), .B(n1081), .C(n1080), .Y(n1266) );
  NAND3XLTS U200 ( .A(n1077), .B(n1076), .C(n1075), .Y(n1267) );
  NAND3XLTS U201 ( .A(n1419), .B(n1418), .C(n1417), .Y(n1244) );
  NAND3XLTS U202 ( .A(n1415), .B(n1414), .C(n1413), .Y(n1245) );
  NAND3XLTS U203 ( .A(n1409), .B(n1408), .C(n1407), .Y(n1246) );
  NAND3XLTS U204 ( .A(n1405), .B(n1404), .C(n1403), .Y(n1247) );
  NAND3XLTS U205 ( .A(n1401), .B(n1400), .C(n1399), .Y(n1248) );
  NAND3XLTS U206 ( .A(n1398), .B(n1397), .C(n1396), .Y(n1249) );
  NAND3XLTS U207 ( .A(n1454), .B(n1453), .C(n1452), .Y(n1238) );
  NAND3XLTS U208 ( .A(n1449), .B(n1448), .C(n1447), .Y(n1239) );
  NAND3XLTS U209 ( .A(n1442), .B(n1441), .C(n1440), .Y(n1240) );
  NAND3XLTS U210 ( .A(n1437), .B(n1436), .C(n1435), .Y(n1241) );
  NAND3XLTS U211 ( .A(n1431), .B(n1430), .C(n1429), .Y(n1242) );
  NAND3XLTS U212 ( .A(n1427), .B(n1426), .C(n1425), .Y(n1243) );
  NAND3XLTS U213 ( .A(n1888), .B(n1887), .C(n1886), .Y(n1122) );
  NAND3XLTS U214 ( .A(n1876), .B(n1875), .C(n1874), .Y(n1123) );
  NAND3XLTS U215 ( .A(n1865), .B(n1864), .C(n1863), .Y(n1124) );
  NAND3XLTS U216 ( .A(n1856), .B(n1855), .C(n1854), .Y(n1125) );
  NAND3XLTS U217 ( .A(n1046), .B(n1045), .C(n1044), .Y(n1274) );
  NAND3XLTS U218 ( .A(n1036), .B(n1035), .C(n1034), .Y(n1275) );
  NAND3XLTS U219 ( .A(n1030), .B(n1029), .C(n1028), .Y(n1276) );
  NAND3XLTS U220 ( .A(n1023), .B(n1022), .C(n1021), .Y(n1277) );
  NAND3XLTS U221 ( .A(n1845), .B(n1844), .C(n1843), .Y(n1134) );
  NAND3XLTS U222 ( .A(n1834), .B(n1833), .C(n1832), .Y(n1135) );
  NAND3XLTS U223 ( .A(n1824), .B(n1823), .C(n1822), .Y(n1136) );
  NAND3XLTS U224 ( .A(n1815), .B(n1814), .C(n1813), .Y(n1137) );
  NAND3XLTS U225 ( .A(n1016), .B(n1015), .C(n1014), .Y(n1278) );
  NAND3XLTS U226 ( .A(n1007), .B(n1006), .C(n1005), .Y(n1279) );
  NAND3XLTS U227 ( .A(n1001), .B(n1000), .C(n999), .Y(n1280) );
  NAND3XLTS U228 ( .A(n994), .B(n993), .C(n992), .Y(n1281) );
  NAND3XLTS U229 ( .A(n1752), .B(n1751), .C(n1750), .Y(n1170) );
  NAND3XLTS U230 ( .A(n1742), .B(n1741), .C(n1740), .Y(n1171) );
  NAND3XLTS U231 ( .A(n1734), .B(n1733), .C(n1732), .Y(n1172) );
  NAND3XLTS U232 ( .A(n1727), .B(n1726), .C(n1725), .Y(n1173) );
  NAND3XLTS U233 ( .A(n943), .B(n942), .C(n941), .Y(n1290) );
  NAND3XLTS U234 ( .A(n933), .B(n932), .C(n931), .Y(n1291) );
  NAND3XLTS U235 ( .A(n928), .B(n927), .C(n926), .Y(n1292) );
  NAND3XLTS U236 ( .A(n923), .B(n922), .C(n921), .Y(n1293) );
  NAND3XLTS U237 ( .A(n1719), .B(n1718), .C(n1717), .Y(n1182) );
  NAND3XLTS U238 ( .A(n1711), .B(n1710), .C(n1709), .Y(n1183) );
  NAND3XLTS U239 ( .A(n1704), .B(n1703), .C(n1702), .Y(n1184) );
  NAND3XLTS U240 ( .A(n1697), .B(n1696), .C(n1695), .Y(n1185) );
  NAND3XLTS U241 ( .A(n917), .B(n916), .C(n915), .Y(n1294) );
  NAND3XLTS U242 ( .A(n911), .B(n910), .C(n909), .Y(n1295) );
  NAND3XLTS U243 ( .A(n907), .B(n906), .C(n905), .Y(n1296) );
  NAND3XLTS U244 ( .A(n904), .B(n903), .C(n902), .Y(n1297) );
  NAND3XLTS U245 ( .A(n1360), .B(n1359), .C(n1358), .Y(n1256) );
  NAND3XLTS U246 ( .A(n1354), .B(n1353), .C(n1352), .Y(n1257) );
  NAND3XLTS U247 ( .A(n1349), .B(n1348), .C(n1347), .Y(n1258) );
  NAND3XLTS U248 ( .A(n1343), .B(n1342), .C(n1341), .Y(n1259) );
  NAND3XLTS U249 ( .A(n1338), .B(n1337), .C(n1112), .Y(n1260) );
  NAND3XLTS U250 ( .A(n1109), .B(n1108), .C(n1107), .Y(n1261) );
  NAND3XLTS U251 ( .A(n1392), .B(n1391), .C(n1390), .Y(n1250) );
  NAND3XLTS U252 ( .A(n1386), .B(n1385), .C(n1384), .Y(n1251) );
  NAND3XLTS U253 ( .A(n1380), .B(n1379), .C(n1378), .Y(n1252) );
  NAND3XLTS U254 ( .A(n1375), .B(n1374), .C(n1373), .Y(n1253) );
  NAND3XLTS U255 ( .A(n1370), .B(n1369), .C(n1368), .Y(n1254) );
  NAND3XLTS U256 ( .A(n1366), .B(n1365), .C(n1364), .Y(n1255) );
  NAND3XLTS U257 ( .A(n1493), .B(n1492), .C(n1491), .Y(n1232) );
  NAND3XLTS U258 ( .A(n1487), .B(n1486), .C(n1485), .Y(n1233) );
  NAND3XLTS U259 ( .A(n1480), .B(n1479), .C(n1478), .Y(n1234) );
  NAND3XLTS U260 ( .A(n1474), .B(n1473), .C(n1472), .Y(n1235) );
  NAND3XLTS U261 ( .A(n1468), .B(n1467), .C(n1466), .Y(n1236) );
  NAND3XLTS U262 ( .A(n1463), .B(n1462), .C(n1461), .Y(n1237) );
  NAND3XLTS U263 ( .A(n1539), .B(n1538), .C(n1537), .Y(n1226) );
  NAND3XLTS U264 ( .A(n1531), .B(n1530), .C(n1529), .Y(n1227) );
  NAND3XLTS U265 ( .A(n1524), .B(n1523), .C(n1522), .Y(n1228) );
  NAND3XLTS U266 ( .A(n1516), .B(n1515), .C(n1514), .Y(n1229) );
  NAND3XLTS U267 ( .A(n1508), .B(n1507), .C(n1506), .Y(n1230) );
  NAND3XLTS U268 ( .A(n1500), .B(n1499), .C(n1498), .Y(n1231) );
  NAND3XLTS U269 ( .A(n1805), .B(n1804), .C(n1803), .Y(n1146) );
  NAND3XLTS U270 ( .A(n1798), .B(n1797), .C(n1796), .Y(n1147) );
  NAND3XLTS U271 ( .A(n1792), .B(n1791), .C(n1790), .Y(n1148) );
  NAND3XLTS U272 ( .A(n1786), .B(n1785), .C(n1784), .Y(n1149) );
  NAND3XLTS U273 ( .A(n986), .B(n985), .C(n984), .Y(n1282) );
  NAND3XLTS U274 ( .A(n980), .B(n979), .C(n978), .Y(n1283) );
  NAND3XLTS U275 ( .A(n976), .B(n975), .C(n974), .Y(n1284) );
  NAND3XLTS U276 ( .A(n972), .B(n971), .C(n970), .Y(n1285) );
  NAND3XLTS U277 ( .A(n1072), .B(n1071), .C(n1070), .Y(n1268) );
  NAND3XLTS U278 ( .A(n1068), .B(n1067), .C(n1066), .Y(n1269) );
  NAND3XLTS U279 ( .A(n1062), .B(n1061), .C(n1060), .Y(n1270) );
  NAND3XLTS U280 ( .A(n1058), .B(n1057), .C(n1056), .Y(n1271) );
  NAND3XLTS U281 ( .A(n1054), .B(n1053), .C(n1052), .Y(n1272) );
  NAND3XLTS U282 ( .A(n1051), .B(n1050), .C(n1049), .Y(n1273) );
  OAI2BB2XLTS U283 ( .B0(n1918), .B1(n502), .A0N(n495), .A1N(n479), .Y(N2624)
         );
  AOI211XLTS U284 ( .A0(n478), .A1(n524), .B0(n477), .C0(n476), .Y(n479) );
  XOR2XLTS U285 ( .A(n523), .B(n490), .Y(n477) );
  OAI21XLTS U286 ( .A0(n478), .A1(n524), .B0(n475), .Y(n476) );
  OR2X1TS U287 ( .A(n85), .B(n1661), .Y(n1455) );
  OR2X1TS U288 ( .A(n391), .B(n1846), .Y(n1024) );
  OR2X1TS U289 ( .A(n185), .B(n1781), .Y(n973) );
  OR2X1TS U290 ( .A(n133), .B(n1753), .Y(n1361) );
  OR2X1TS U291 ( .A(n276), .B(n1720), .Y(n1393) );
  OR2X1TS U292 ( .A(n31), .B(n1654), .Y(n1494) );
  OR2X1TS U293 ( .A(n1573), .B(n279), .Y(n3) );
  OR2X1TS U294 ( .A(n1618), .B(n395), .Y(n4) );
  OR2X1TS U295 ( .A(n1574), .B(n279), .Y(n5) );
  OR2X1TS U296 ( .A(n1621), .B(n395), .Y(n6) );
  OR2X1TS U297 ( .A(n1552), .B(n89), .Y(n7) );
  OA21XLTS U298 ( .A0(n19), .A1(n446), .B0(n22), .Y(n8) );
  CLKBUFX2TS U299 ( .A(n321), .Y(n322) );
  OR2X1TS U300 ( .A(n438), .B(n1571), .Y(n10) );
  NOR3XLTS U301 ( .A(n1558), .B(n1553), .C(n87), .Y(n83) );
  NOR3XLTS U302 ( .A(n1581), .B(n1575), .C(n278), .Y(n274) );
  OR2X1TS U303 ( .A(n390), .B(n1630), .Y(n11) );
  NOR2XLTS U304 ( .A(n27), .B(n1582), .Y(n275) );
  AND3X1TS U305 ( .A(n537), .B(n1906), .C(n536), .Y(n12) );
  INVX2TS U306 ( .A(destinationAddressIn_EAST[5]), .Y(n66) );
  INVX2TS U307 ( .A(destinationAddressIn_EAST[4]), .Y(n61) );
  INVX2TS U308 ( .A(destinationAddressIn_EAST[6]), .Y(n58) );
  INVX2TS U309 ( .A(destinationAddressIn_EAST[7]), .Y(n72) );
  INVX2TS U310 ( .A(destinationAddressIn_EAST[10]), .Y(n39) );
  INVX2TS U311 ( .A(destinationAddressIn_EAST[8]), .Y(n44) );
  INVX2TS U312 ( .A(destinationAddressIn_EAST[9]), .Y(n48) );
  INVX2TS U313 ( .A(destinationAddressIn_EAST[11]), .Y(n30) );
  INVX2TS U314 ( .A(writeIn_EAST), .Y(n53) );
  CLKBUFX2TS U315 ( .A(n1910), .Y(n13) );
  INVX2TS U331 ( .A(n1916), .Y(n482) );
  INVX2TS U332 ( .A(n1913), .Y(n440) );
  ADDFX1TS U333 ( .A(selectBit_SOUTH), .B(selectBit_NORTH), .CI(selectBit_EAST), .CO(n453), .S(n449) );
  INVX2TS U334 ( .A(n15), .Y(n77) );
  INVX2TS U335 ( .A(n77), .Y(n121) );
  INVX2TS U336 ( .A(selectBit_WEST), .Y(n444) );
  INVX2TS U337 ( .A(n1546), .Y(n1548) );
  INVX2TS U338 ( .A(n1909), .Y(n448) );
  INVX2TS U339 ( .A(selectBit_SOUTH), .Y(n505) );
  INVX2TS U340 ( .A(n9), .Y(n223) );
  INVX2TS U341 ( .A(n1916), .Y(n446) );
  NAND2X1TS U342 ( .A(n18), .B(n446), .Y(n22) );
  NAND2X1TS U343 ( .A(selectBit_SOUTH), .B(n21), .Y(n20) );
  NAND2X1TS U344 ( .A(n311), .B(n380), .Y(n124) );
  INVX2TS U345 ( .A(selectBit_EAST), .Y(n509) );
  INVX2TS U346 ( .A(n509), .Y(n512) );
  INVX2TS U347 ( .A(n1915), .Y(n469) );
  INVX2TS U348 ( .A(n1914), .Y(n441) );
  AOI22X1TS U349 ( .A0(n469), .A1(n22), .B0(n125), .B1(n441), .Y(n79) );
  INVX2TS U350 ( .A(n23), .Y(n24) );
  OAI21XLTS U351 ( .A0(n25), .A1(n79), .B0(n24), .Y(n123) );
  NAND2X1TS U352 ( .A(n512), .B(n123), .Y(n270) );
  NAND2X1TS U353 ( .A(n442), .B(n125), .Y(n28) );
  INVX2TS U354 ( .A(n1916), .Y(n493) );
  INVX2TS U355 ( .A(n272), .Y(n384) );
  INVX2TS U356 ( .A(n505), .Y(n504) );
  INVX2TS U357 ( .A(n444), .Y(n511) );
  INVX2TS U358 ( .A(readReady), .Y(n128) );
  INVX2TS U359 ( .A(n128), .Y(n510) );
  NOR3XLTS U360 ( .A(n511), .B(selectBit_EAST), .C(n510), .Y(n506) );
  NAND2X1TS U361 ( .A(n537), .B(n506), .Y(n522) );
  NAND2X1TS U362 ( .A(n522), .B(n1918), .Y(n27) );
  INVX2TS U363 ( .A(n27), .Y(n126) );
  INVX2TS U364 ( .A(n27), .Y(n131) );
  INVX2TS U365 ( .A(n131), .Y(n81) );
  INVX2TS U366 ( .A(n1916), .Y(n485) );
  NAND2X1TS U367 ( .A(n31), .B(n1549), .Y(n34) );
  INVX2TS U368 ( .A(n29), .Y(n1509) );
  INVX2TS U369 ( .A(n1509), .Y(n872) );
  CLKBUFX2TS U370 ( .A(n872), .Y(n43) );
  INVX2TS U371 ( .A(n43), .Y(n65) );
  INVX2TS U372 ( .A(destinationAddressIn_EAST[11]), .Y(n245) );
  INVX2TS U373 ( .A(n126), .Y(n438) );
  OR2X1TS U374 ( .A(n1549), .B(n438), .Y(n1501) );
  INVX2TS U375 ( .A(n1501), .Y(n1654) );
  INVX2TS U376 ( .A(n1494), .Y(n49) );
  OR2X1TS U377 ( .A(n1546), .B(n34), .Y(n54) );
  INVX2TS U378 ( .A(n54), .Y(n1646) );
  INVX2TS U379 ( .A(n1646), .Y(n1502) );
  INVX2TS U380 ( .A(n1502), .Y(n32) );
  CLKBUFX2TS U381 ( .A(destinationAddressIn_WEST[11]), .Y(n412) );
  CLKBUFX2TS U382 ( .A(n412), .Y(n759) );
  AOI22X1TS U383 ( .A0(n49), .A1(\destinationAddressbuffer[7][11] ), .B0(n32), 
        .B1(n759), .Y(n38) );
  NAND2BX1TS U384 ( .AN(n34), .B(n33), .Y(n36) );
  OR2X1TS U385 ( .A(n1541), .B(n36), .Y(n55) );
  INVX2TS U386 ( .A(n55), .Y(n35) );
  INVX2TS U387 ( .A(n35), .Y(n873) );
  INVX2TS U388 ( .A(n873), .Y(n69) );
  INVX2TS U389 ( .A(n168), .Y(n762) );
  CLKBUFX2TS U390 ( .A(destinationAddressIn_NORTH[11]), .Y(n763) );
  CLKBUFX2TS U391 ( .A(n763), .Y(n332) );
  AOI22X1TS U392 ( .A0(n69), .A1(n762), .B0(n50), .B1(n332), .Y(n37) );
  OAI211XLTS U393 ( .A0(n65), .A1(n245), .B0(n38), .C0(n37), .Y(n1198) );
  INVX2TS U394 ( .A(destinationAddressIn_EAST[10]), .Y(n240) );
  INVX2TS U395 ( .A(n54), .Y(n1519) );
  CLKBUFX2TS U396 ( .A(destinationAddressIn_WEST[10]), .Y(n392) );
  CLKBUFX2TS U397 ( .A(n392), .Y(n743) );
  AOI22X1TS U398 ( .A0(n49), .A1(\destinationAddressbuffer[7][10] ), .B0(n1519), .B1(n743), .Y(n42) );
  INVX2TS U399 ( .A(n55), .Y(n868) );
  INVX2TS U400 ( .A(n174), .Y(n746) );
  INVX2TS U401 ( .A(n40), .Y(n62) );
  INVX2TS U402 ( .A(n62), .Y(n1647) );
  CLKBUFX2TS U403 ( .A(destinationAddressIn_NORTH[10]), .Y(n747) );
  CLKBUFX2TS U404 ( .A(n747), .Y(n346) );
  AOI22X1TS U405 ( .A0(n868), .A1(n746), .B0(n1647), .B1(n346), .Y(n41) );
  OAI211XLTS U406 ( .A0(n65), .A1(n240), .B0(n42), .C0(n41), .Y(n1199) );
  INVX2TS U407 ( .A(n43), .Y(n76) );
  INVX2TS U408 ( .A(destinationAddressIn_EAST[8]), .Y(n233) );
  INVX2TS U409 ( .A(n54), .Y(n45) );
  CLKBUFX2TS U410 ( .A(destinationAddressIn_WEST[8]), .Y(n400) );
  CLKBUFX2TS U411 ( .A(n400), .Y(n711) );
  AOI22X1TS U412 ( .A0(n49), .A1(\destinationAddressbuffer[7][8] ), .B0(n45), 
        .B1(n711), .Y(n47) );
  INVX2TS U413 ( .A(n164), .Y(n712) );
  CLKBUFX2TS U414 ( .A(destinationAddressIn_NORTH[8]), .Y(n713) );
  CLKBUFX2TS U415 ( .A(n713), .Y(n326) );
  AOI22X1TS U416 ( .A0(n69), .A1(n712), .B0(n50), .B1(n326), .Y(n46) );
  OAI211XLTS U417 ( .A0(n76), .A1(n233), .B0(n47), .C0(n46), .Y(n1201) );
  INVX2TS U418 ( .A(destinationAddressIn_EAST[9]), .Y(n236) );
  INVX2TS U419 ( .A(n1502), .Y(n67) );
  CLKBUFX2TS U420 ( .A(destinationAddressIn_WEST[9]), .Y(n406) );
  CLKBUFX2TS U421 ( .A(n406), .Y(n726) );
  AOI22X1TS U422 ( .A0(n49), .A1(\destinationAddressbuffer[7][9] ), .B0(n67), 
        .B1(n726), .Y(n52) );
  INVX2TS U423 ( .A(n873), .Y(n1639) );
  INVX2TS U424 ( .A(n160), .Y(n727) );
  INVX2TS U425 ( .A(n62), .Y(n50) );
  INVX2TS U426 ( .A(n50), .Y(n878) );
  INVX2TS U427 ( .A(n878), .Y(n68) );
  CLKBUFX2TS U428 ( .A(destinationAddressIn_NORTH[9]), .Y(n729) );
  CLKBUFX2TS U429 ( .A(n729), .Y(n338) );
  AOI22X1TS U430 ( .A0(n1639), .A1(n727), .B0(n68), .B1(n338), .Y(n51) );
  OAI211XLTS U431 ( .A0(n65), .A1(n236), .B0(n52), .C0(n51), .Y(n1200) );
  CLKBUFX2TS U432 ( .A(n1494), .Y(n877) );
  INVX2TS U433 ( .A(n877), .Y(n1652) );
  INVX2TS U434 ( .A(n54), .Y(n1656) );
  AOI22X1TS U435 ( .A0(n1652), .A1(writeOutbuffer[7]), .B0(n1656), .B1(
        writeIn_WEST), .Y(n57) );
  INVX2TS U436 ( .A(writeIn_SOUTH), .Y(n178) );
  INVX2TS U437 ( .A(n178), .Y(n543) );
  INVX2TS U438 ( .A(n62), .Y(n1657) );
  AOI22X1TS U439 ( .A0(n35), .A1(n543), .B0(n1657), .B1(writeIn_NORTH), .Y(n56) );
  OAI211XLTS U440 ( .A0(n76), .A1(n295), .B0(n57), .C0(n56), .Y(n1225) );
  INVX2TS U441 ( .A(destinationAddressIn_EAST[6]), .Y(n253) );
  INVX2TS U442 ( .A(n877), .Y(n73) );
  AOI22X1TS U443 ( .A0(n73), .A1(\destinationAddressbuffer[7][6] ), .B0(n1656), 
        .B1(destinationAddressIn_WEST[6]), .Y(n60) );
  INVX2TS U444 ( .A(destinationAddressIn_SOUTH[6]), .Y(n140) );
  INVX2TS U445 ( .A(n140), .Y(n688) );
  AOI22X1TS U446 ( .A0(n1639), .A1(n688), .B0(n1647), .B1(
        destinationAddressIn_NORTH[6]), .Y(n59) );
  OAI211XLTS U447 ( .A0(n76), .A1(n253), .B0(n60), .C0(n59), .Y(n1203) );
  INVX2TS U448 ( .A(destinationAddressIn_EAST[4]), .Y(n267) );
  AOI22X1TS U449 ( .A0(n73), .A1(\destinationAddressbuffer[7][4] ), .B0(n1519), 
        .B1(destinationAddressIn_WEST[4]), .Y(n64) );
  INVX2TS U450 ( .A(destinationAddressIn_SOUTH[4]), .Y(n156) );
  INVX2TS U451 ( .A(n156), .Y(n656) );
  INVX2TS U452 ( .A(n62), .Y(n1535) );
  AOI22X1TS U453 ( .A0(n868), .A1(n656), .B0(n1535), .B1(
        destinationAddressIn_NORTH[4]), .Y(n63) );
  OAI211XLTS U454 ( .A0(n65), .A1(n267), .B0(n64), .C0(n63), .Y(n1205) );
  INVX2TS U455 ( .A(destinationAddressIn_EAST[5]), .Y(n263) );
  AOI22X1TS U456 ( .A0(n73), .A1(\destinationAddressbuffer[7][5] ), .B0(n67), 
        .B1(destinationAddressIn_WEST[5]), .Y(n71) );
  INVX2TS U457 ( .A(destinationAddressIn_SOUTH[5]), .Y(n150) );
  INVX2TS U458 ( .A(n150), .Y(n668) );
  AOI22X1TS U459 ( .A0(n69), .A1(n668), .B0(n68), .B1(
        destinationAddressIn_NORTH[5]), .Y(n70) );
  OAI211XLTS U460 ( .A0(n1509), .A1(n263), .B0(n71), .C0(n70), .Y(n1204) );
  INVX2TS U461 ( .A(destinationAddressIn_EAST[7]), .Y(n257) );
  AOI22X1TS U462 ( .A0(n73), .A1(\destinationAddressbuffer[7][7] ), .B0(n45), 
        .B1(destinationAddressIn_WEST[7]), .Y(n75) );
  INVX2TS U463 ( .A(destinationAddressIn_SOUTH[7]), .Y(n145) );
  INVX2TS U464 ( .A(n145), .Y(n701) );
  AOI22X1TS U465 ( .A0(n35), .A1(n701), .B0(n1657), .B1(
        destinationAddressIn_NORTH[7]), .Y(n74) );
  OAI211XLTS U466 ( .A0(n76), .A1(n257), .B0(n75), .C0(n74), .Y(n1202) );
  INVX2TS U467 ( .A(n78), .Y(n180) );
  NAND2X1TS U468 ( .A(n122), .B(n450), .Y(n269) );
  AOI21X1TS U469 ( .A0(n223), .A1(n222), .B0(n311), .Y(n382) );
  INVX2TS U470 ( .A(n380), .Y(n312) );
  INVX2TS U471 ( .A(n312), .Y(n181) );
  NOR2XLTS U472 ( .A(n440), .B(n503), .Y(n385) );
  CLKBUFX2TS U473 ( .A(n79), .Y(n272) );
  AOI31XLTS U474 ( .A0(n469), .A1(n482), .A2(n385), .B0(n1552), .Y(n82) );
  AOI21X1TS U475 ( .A0(n86), .A1(n82), .B0(n81), .Y(n85) );
  INVX2TS U476 ( .A(n128), .Y(n513) );
  INVX2TS U477 ( .A(n1909), .Y(n388) );
  NAND2X1TS U478 ( .A(n85), .B(n1559), .Y(n87) );
  INVX2TS U479 ( .A(n83), .Y(n1469) );
  INVX2TS U480 ( .A(n1469), .Y(n896) );
  CLKBUFX2TS U481 ( .A(n896), .Y(n95) );
  INVX2TS U482 ( .A(n95), .Y(n113) );
  INVX2TS U483 ( .A(n84), .Y(n893) );
  INVX2TS U484 ( .A(n893), .Y(n1661) );
  CLKBUFX2TS U485 ( .A(n1455), .Y(n894) );
  INVX2TS U486 ( .A(n894), .Y(n101) );
  OR2X1TS U487 ( .A(n1556), .B(n87), .Y(n99) );
  INVX2TS U488 ( .A(n99), .Y(n1662) );
  AOI22X1TS U489 ( .A0(n101), .A1(\destinationAddressbuffer[6][10] ), .B0(
        n1662), .B1(n743), .Y(n92) );
  INVX2TS U490 ( .A(n7), .Y(n88) );
  INVX2TS U491 ( .A(n88), .Y(n885) );
  INVX2TS U492 ( .A(n885), .Y(n103) );
  CLKBUFX2TS U493 ( .A(n747), .Y(n397) );
  INVX2TS U494 ( .A(n90), .Y(n102) );
  INVX2TS U495 ( .A(n174), .Y(n345) );
  AOI22X1TS U496 ( .A0(n103), .A1(n397), .B0(n117), .B1(n345), .Y(n91) );
  OAI211XLTS U497 ( .A0(n113), .A1(n240), .B0(n92), .C0(n91), .Y(n1187) );
  INVX2TS U498 ( .A(n99), .Y(n1457) );
  AOI22X1TS U499 ( .A0(n101), .A1(\destinationAddressbuffer[6][8] ), .B0(n1457), .B1(n711), .Y(n94) );
  INVX2TS U500 ( .A(n7), .Y(n1686) );
  CLKBUFX2TS U501 ( .A(n713), .Y(n402) );
  INVX2TS U502 ( .A(n90), .Y(n897) );
  INVX2TS U503 ( .A(n897), .Y(n117) );
  INVX2TS U504 ( .A(n164), .Y(n325) );
  AOI22X1TS U505 ( .A0(n1686), .A1(n402), .B0(n117), .B1(n325), .Y(n93) );
  OAI211XLTS U506 ( .A0(n113), .A1(n233), .B0(n94), .C0(n93), .Y(n1189) );
  INVX2TS U507 ( .A(n95), .Y(n120) );
  INVX2TS U508 ( .A(n99), .Y(n1683) );
  AOI22X1TS U509 ( .A0(n101), .A1(\destinationAddressbuffer[6][9] ), .B0(n100), 
        .B1(n726), .Y(n98) );
  INVX2TS U510 ( .A(n885), .Y(n889) );
  CLKBUFX2TS U511 ( .A(n729), .Y(n407) );
  INVX2TS U512 ( .A(n102), .Y(n1459) );
  INVX2TS U513 ( .A(n102), .Y(n96) );
  INVX2TS U514 ( .A(n160), .Y(n337) );
  AOI22X1TS U515 ( .A0(n889), .A1(n407), .B0(n96), .B1(n337), .Y(n97) );
  OAI211XLTS U516 ( .A0(n120), .A1(n236), .B0(n98), .C0(n97), .Y(n1188) );
  INVX2TS U517 ( .A(n99), .Y(n100) );
  INVX2TS U518 ( .A(n100), .Y(n895) );
  INVX2TS U519 ( .A(n895), .Y(n110) );
  AOI22X1TS U520 ( .A0(n101), .A1(\destinationAddressbuffer[6][11] ), .B0(n110), .B1(n759), .Y(n105) );
  CLKBUFX2TS U521 ( .A(n763), .Y(n414) );
  INVX2TS U522 ( .A(n168), .Y(n330) );
  AOI22X1TS U523 ( .A0(n103), .A1(n414), .B0(n90), .B1(n330), .Y(n104) );
  OAI211XLTS U524 ( .A0(n113), .A1(n245), .B0(n105), .C0(n104), .Y(n1186) );
  INVX2TS U525 ( .A(n894), .Y(n1682) );
  AOI22X1TS U526 ( .A0(n1682), .A1(writeOutbuffer[6]), .B0(n1662), .B1(
        writeIn_WEST), .Y(n107) );
  INVX2TS U527 ( .A(n7), .Y(n1664) );
  CLKBUFX2TS U528 ( .A(writeIn_NORTH), .Y(n352) );
  CLKBUFX2TS U529 ( .A(n352), .Y(n418) );
  INVX2TS U530 ( .A(n178), .Y(n351) );
  AOI22X1TS U531 ( .A0(n1664), .A1(n418), .B0(n1678), .B1(n351), .Y(n106) );
  OAI211XLTS U532 ( .A0(n120), .A1(n295), .B0(n107), .C0(n106), .Y(n1224) );
  INVX2TS U533 ( .A(n1455), .Y(n116) );
  CLKBUFX2TS U534 ( .A(destinationAddressIn_WEST[4]), .Y(n654) );
  AOI22X1TS U535 ( .A0(n116), .A1(\destinationAddressbuffer[6][4] ), .B0(n110), 
        .B1(n654), .Y(n109) );
  CLKBUFX2TS U536 ( .A(destinationAddressIn_NORTH[4]), .Y(n375) );
  CLKBUFX2TS U537 ( .A(n375), .Y(n425) );
  INVX2TS U538 ( .A(n156), .Y(n374) );
  AOI22X1TS U539 ( .A0(n1686), .A1(n425), .B0(n90), .B1(n374), .Y(n108) );
  OAI211XLTS U540 ( .A0(n120), .A1(n267), .B0(n109), .C0(n108), .Y(n1193) );
  CLKBUFX2TS U541 ( .A(destinationAddressIn_WEST[5]), .Y(n666) );
  AOI22X1TS U542 ( .A0(n116), .A1(\destinationAddressbuffer[6][5] ), .B0(n110), 
        .B1(n666), .Y(n112) );
  INVX2TS U543 ( .A(n7), .Y(n1460) );
  CLKBUFX2TS U544 ( .A(destinationAddressIn_NORTH[5]), .Y(n368) );
  CLKBUFX2TS U545 ( .A(n368), .Y(n421) );
  INVX2TS U546 ( .A(n897), .Y(n1685) );
  INVX2TS U547 ( .A(n150), .Y(n367) );
  AOI22X1TS U548 ( .A0(n1460), .A1(n421), .B0(n1685), .B1(n367), .Y(n111) );
  OAI211XLTS U549 ( .A0(n113), .A1(n263), .B0(n112), .C0(n111), .Y(n1192) );
  CLKBUFX2TS U550 ( .A(destinationAddressIn_WEST[7]), .Y(n700) );
  AOI22X1TS U551 ( .A0(n116), .A1(\destinationAddressbuffer[6][7] ), .B0(n1457), .B1(n700), .Y(n115) );
  CLKBUFX2TS U552 ( .A(destinationAddressIn_NORTH[7]), .Y(n357) );
  CLKBUFX2TS U553 ( .A(n357), .Y(n434) );
  INVX2TS U554 ( .A(n145), .Y(n356) );
  AOI22X1TS U555 ( .A0(n1460), .A1(n434), .B0(n1459), .B1(n356), .Y(n114) );
  OAI211XLTS U556 ( .A0(n1469), .A1(n257), .B0(n115), .C0(n114), .Y(n1190) );
  CLKBUFX2TS U557 ( .A(destinationAddressIn_WEST[6]), .Y(n686) );
  AOI22X1TS U558 ( .A0(n116), .A1(\destinationAddressbuffer[6][6] ), .B0(n1683), .B1(n686), .Y(n119) );
  CLKBUFX2TS U559 ( .A(destinationAddressIn_NORTH[6]), .Y(n362) );
  CLKBUFX2TS U560 ( .A(n362), .Y(n429) );
  INVX2TS U561 ( .A(n140), .Y(n361) );
  AOI22X1TS U562 ( .A0(n889), .A1(n429), .B0(n117), .B1(n361), .Y(n118) );
  OAI211XLTS U563 ( .A0(n120), .A1(n253), .B0(n119), .C0(n118), .Y(n1191) );
  INVX2TS U564 ( .A(n1914), .Y(n481) );
  NAND2X1TS U565 ( .A(n125), .B(n481), .Y(n127) );
  INVX2TS U566 ( .A(n126), .Y(n390) );
  INVX2TS U567 ( .A(n128), .Y(n508) );
  INVX2TS U568 ( .A(n1914), .Y(n484) );
  INVX2TS U569 ( .A(n130), .Y(n958) );
  INVX2TS U570 ( .A(n958), .Y(n1762) );
  CLKBUFX2TS U571 ( .A(n1762), .Y(n146) );
  INVX2TS U572 ( .A(n146), .Y(n169) );
  INVX2TS U573 ( .A(n131), .Y(n480) );
  INVX2TS U574 ( .A(n132), .Y(n964) );
  INVX2TS U575 ( .A(n964), .Y(n1753) );
  CLKBUFX2TS U576 ( .A(n1361), .Y(n175) );
  INVX2TS U577 ( .A(n175), .Y(n152) );
  NOR3XLTS U578 ( .A(n1589), .B(n1584), .C(n136), .Y(n141) );
  INVX2TS U579 ( .A(n951), .Y(n157) );
  AOI22X1TS U580 ( .A0(n152), .A1(\destinationAddressbuffer[3][6] ), .B0(n157), 
        .B1(destinationAddressIn_EAST[6]), .Y(n139) );
  OR2X1TS U581 ( .A(n23), .B(n134), .Y(n171) );
  INVX2TS U582 ( .A(n171), .Y(n135) );
  INVX2TS U583 ( .A(n135), .Y(n142) );
  INVX2TS U584 ( .A(n137), .Y(n153) );
  INVX2TS U585 ( .A(n153), .Y(n1755) );
  CLKBUFX2TS U586 ( .A(n686), .Y(n360) );
  AOI22X1TS U587 ( .A0(n135), .A1(n362), .B0(n1755), .B1(n360), .Y(n138) );
  OAI211XLTS U588 ( .A0(n169), .A1(n140), .B0(n139), .C0(n138), .Y(n1155) );
  INVX2TS U589 ( .A(n141), .Y(n161) );
  INVX2TS U590 ( .A(n161), .Y(n1774) );
  AOI22X1TS U591 ( .A0(n152), .A1(\destinationAddressbuffer[3][7] ), .B0(n1774), .B1(destinationAddressIn_EAST[7]), .Y(n144) );
  INVX2TS U592 ( .A(n142), .Y(n1383) );
  INVX2TS U593 ( .A(n153), .Y(n1775) );
  CLKBUFX2TS U594 ( .A(n700), .Y(n355) );
  AOI22X1TS U595 ( .A0(n1383), .A1(n357), .B0(n1775), .B1(n355), .Y(n143) );
  OAI211XLTS U596 ( .A0(n169), .A1(n145), .B0(n144), .C0(n143), .Y(n1154) );
  INVX2TS U597 ( .A(n146), .Y(n179) );
  INVX2TS U598 ( .A(n161), .Y(n1767) );
  AOI22X1TS U599 ( .A0(n152), .A1(\destinationAddressbuffer[3][5] ), .B0(n1767), .B1(destinationAddressIn_EAST[5]), .Y(n149) );
  INVX2TS U600 ( .A(n171), .Y(n1777) );
  INVX2TS U601 ( .A(n142), .Y(n959) );
  INVX2TS U602 ( .A(n153), .Y(n147) );
  INVX2TS U603 ( .A(n147), .Y(n945) );
  INVX2TS U604 ( .A(n945), .Y(n165) );
  CLKBUFX2TS U605 ( .A(n666), .Y(n366) );
  AOI22X1TS U606 ( .A0(n959), .A1(n368), .B0(n165), .B1(n366), .Y(n148) );
  OAI211XLTS U607 ( .A0(n179), .A1(n150), .B0(n149), .C0(n148), .Y(n1156) );
  INVX2TS U608 ( .A(n161), .Y(n151) );
  AOI22X1TS U609 ( .A0(n152), .A1(\destinationAddressbuffer[3][4] ), .B0(n157), 
        .B1(destinationAddressIn_EAST[4]), .Y(n155) );
  INVX2TS U610 ( .A(n153), .Y(n1389) );
  CLKBUFX2TS U611 ( .A(n654), .Y(n371) );
  AOI22X1TS U612 ( .A0(n1777), .A1(n375), .B0(n1389), .B1(n371), .Y(n154) );
  OAI211XLTS U613 ( .A0(n169), .A1(n156), .B0(n155), .C0(n154), .Y(n1157) );
  INVX2TS U614 ( .A(n175), .Y(n170) );
  AOI22X1TS U615 ( .A0(n170), .A1(\destinationAddressbuffer[3][9] ), .B0(n157), 
        .B1(destinationAddressIn_EAST[9]), .Y(n159) );
  CLKBUFX2TS U616 ( .A(n406), .Y(n336) );
  AOI22X1TS U617 ( .A0(n959), .A1(n338), .B0(n137), .B1(n336), .Y(n158) );
  OAI211XLTS U618 ( .A0(n179), .A1(n160), .B0(n159), .C0(n158), .Y(n1152) );
  INVX2TS U619 ( .A(n161), .Y(n1381) );
  AOI22X1TS U620 ( .A0(n170), .A1(\destinationAddressbuffer[3][8] ), .B0(n1381), .B1(destinationAddressIn_EAST[8]), .Y(n163) );
  INVX2TS U621 ( .A(n171), .Y(n1756) );
  CLKBUFX2TS U622 ( .A(n400), .Y(n318) );
  AOI22X1TS U623 ( .A0(n1756), .A1(n326), .B0(n1755), .B1(n318), .Y(n162) );
  OAI211XLTS U624 ( .A0(n179), .A1(n164), .B0(n163), .C0(n162), .Y(n1153) );
  AOI22X1TS U625 ( .A0(n170), .A1(\destinationAddressbuffer[3][11] ), .B0(
        n1767), .B1(destinationAddressIn_EAST[11]), .Y(n167) );
  CLKBUFX2TS U626 ( .A(n412), .Y(n329) );
  AOI22X1TS U627 ( .A0(n1777), .A1(n332), .B0(n165), .B1(n329), .Y(n166) );
  OAI211XLTS U628 ( .A0(n169), .A1(n168), .B0(n167), .C0(n166), .Y(n1150) );
  AOI22X1TS U629 ( .A0(n170), .A1(\destinationAddressbuffer[3][10] ), .B0(
        n1381), .B1(destinationAddressIn_EAST[10]), .Y(n173) );
  INVX2TS U630 ( .A(n171), .Y(n1363) );
  CLKBUFX2TS U631 ( .A(n392), .Y(n342) );
  AOI22X1TS U632 ( .A0(n1363), .A1(n346), .B0(n1389), .B1(n342), .Y(n172) );
  OAI211XLTS U633 ( .A0(n958), .A1(n174), .B0(n173), .C0(n172), .Y(n1151) );
  INVX2TS U634 ( .A(n175), .Y(n1772) );
  AOI22X1TS U635 ( .A0(n1772), .A1(writeOutbuffer[3]), .B0(n1774), .B1(
        writeIn_EAST), .Y(n177) );
  CLKBUFX2TS U636 ( .A(writeIn_WEST), .Y(n541) );
  CLKBUFX2TS U637 ( .A(n541), .Y(n349) );
  AOI22X1TS U638 ( .A0(n1363), .A1(n352), .B0(n1775), .B1(n349), .Y(n176) );
  OAI211XLTS U639 ( .A0(n179), .A1(n178), .B0(n177), .C0(n176), .Y(n1221) );
  NOR3XLTS U640 ( .A(n382), .B(n181), .C(n381), .Y(n1597) );
  AOI31XLTS U641 ( .A0(n493), .A1(n385), .A2(n484), .B0(n1593), .Y(n182) );
  AOI21X1TS U642 ( .A0(n187), .A1(n182), .B0(n390), .Y(n185) );
  NAND2X1TS U643 ( .A(n185), .B(n1601), .Y(n188) );
  INVX2TS U644 ( .A(n183), .Y(n1339) );
  INVX2TS U645 ( .A(n1339), .Y(n983) );
  CLKBUFX2TS U646 ( .A(n983), .Y(n197) );
  INVX2TS U647 ( .A(n197), .Y(n213) );
  INVX2TS U648 ( .A(n184), .Y(n981) );
  INVX2TS U649 ( .A(n981), .Y(n1781) );
  INVX2TS U650 ( .A(n973), .Y(n202) );
  OR2X1TS U651 ( .A(n1598), .B(n188), .Y(n201) );
  INVX2TS U652 ( .A(n201), .Y(n186) );
  INVX2TS U653 ( .A(n186), .Y(n982) );
  INVX2TS U654 ( .A(n982), .Y(n214) );
  AOI22X1TS U655 ( .A0(n202), .A1(\destinationAddressbuffer[2][8] ), .B0(n214), 
        .B1(n318), .Y(n193) );
  INVX2TS U656 ( .A(n198), .Y(n208) );
  INVX2TS U657 ( .A(n208), .Y(n1802) );
  INVX2TS U658 ( .A(n190), .Y(n203) );
  INVX2TS U659 ( .A(n203), .Y(n191) );
  INVX2TS U660 ( .A(n191), .Y(n969) );
  INVX2TS U661 ( .A(n969), .Y(n218) );
  AOI22X1TS U662 ( .A0(n1802), .A1(n326), .B0(n218), .B1(n325), .Y(n192) );
  OAI211XLTS U663 ( .A0(n213), .A1(n233), .B0(n193), .C0(n192), .Y(n1141) );
  INVX2TS U664 ( .A(n201), .Y(n1782) );
  AOI22X1TS U665 ( .A0(n202), .A1(\destinationAddressbuffer[2][11] ), .B0(
        n1782), .B1(n329), .Y(n196) );
  INVX2TS U666 ( .A(n208), .Y(n194) );
  INVX2TS U667 ( .A(n203), .Y(n1357) );
  AOI22X1TS U668 ( .A0(n194), .A1(n332), .B0(n1357), .B1(n330), .Y(n195) );
  OAI211XLTS U669 ( .A0(n213), .A1(n245), .B0(n196), .C0(n195), .Y(n1138) );
  INVX2TS U670 ( .A(n197), .Y(n221) );
  INVX2TS U671 ( .A(n201), .Y(n1801) );
  AOI22X1TS U672 ( .A0(n202), .A1(\destinationAddressbuffer[2][9] ), .B0(n1801), .B1(n336), .Y(n200) );
  INVX2TS U673 ( .A(n198), .Y(n1111) );
  INVX2TS U674 ( .A(n1111), .Y(n977) );
  INVX2TS U675 ( .A(n203), .Y(n1105) );
  AOI22X1TS U676 ( .A0(n977), .A1(n338), .B0(n218), .B1(n337), .Y(n199) );
  INVX2TS U677 ( .A(n201), .Y(n1104) );
  AOI22X1TS U678 ( .A0(n202), .A1(\destinationAddressbuffer[2][10] ), .B0(
        n1104), .B1(n342), .Y(n205) );
  INVX2TS U679 ( .A(n203), .Y(n1346) );
  AOI22X1TS U680 ( .A0(n194), .A1(n346), .B0(n1346), .B1(n345), .Y(n204) );
  OAI211XLTS U681 ( .A0(n213), .A1(n240), .B0(n205), .C0(n204), .Y(n1139) );
  CLKBUFX2TS U682 ( .A(n973), .Y(n1602) );
  INVX2TS U683 ( .A(n1602), .Y(n1799) );
  AOI22X1TS U684 ( .A0(n1799), .A1(writeOutbuffer[2]), .B0(n214), .B1(n349), 
        .Y(n207) );
  INVX2TS U685 ( .A(n208), .Y(n1783) );
  AOI22X1TS U686 ( .A0(n1783), .A1(writeIn_NORTH), .B0(n1346), .B1(n351), .Y(
        n206) );
  OAI211XLTS U687 ( .A0(n221), .A1(n295), .B0(n207), .C0(n206), .Y(n1220) );
  INVX2TS U688 ( .A(n973), .Y(n217) );
  AOI22X1TS U689 ( .A0(n217), .A1(\destinationAddressbuffer[2][7] ), .B0(n1782), .B1(n355), .Y(n210) );
  INVX2TS U690 ( .A(n208), .Y(n1106) );
  AOI22X1TS U691 ( .A0(n1106), .A1(destinationAddressIn_NORTH[7]), .B0(n1105), 
        .B1(n356), .Y(n209) );
  OAI211XLTS U692 ( .A0(n221), .A1(n257), .B0(n210), .C0(n209), .Y(n1142) );
  AOI22X1TS U693 ( .A0(n217), .A1(\destinationAddressbuffer[2][5] ), .B0(n1104), .B1(n366), .Y(n212) );
  AOI22X1TS U694 ( .A0(n1106), .A1(destinationAddressIn_NORTH[5]), .B0(n1105), 
        .B1(n367), .Y(n211) );
  OAI211XLTS U695 ( .A0(n213), .A1(n263), .B0(n212), .C0(n211), .Y(n1144) );
  AOI22X1TS U696 ( .A0(n217), .A1(\destinationAddressbuffer[2][4] ), .B0(n214), 
        .B1(n371), .Y(n216) );
  AOI22X1TS U697 ( .A0(n1802), .A1(destinationAddressIn_NORTH[4]), .B0(n1357), 
        .B1(n374), .Y(n215) );
  OAI211XLTS U698 ( .A0(n1339), .A1(n267), .B0(n216), .C0(n215), .Y(n1145) );
  AOI22X1TS U699 ( .A0(n217), .A1(\destinationAddressbuffer[2][6] ), .B0(n186), 
        .B1(n360), .Y(n220) );
  AOI22X1TS U700 ( .A0(n977), .A1(destinationAddressIn_NORTH[6]), .B0(n218), 
        .B1(n361), .Y(n219) );
  OAI211XLTS U701 ( .A0(n221), .A1(n253), .B0(n220), .C0(n219), .Y(n1143) );
  INVX2TS U702 ( .A(n1912), .Y(n387) );
  INVX2TS U703 ( .A(n1913), .Y(n491) );
  INVX2TS U704 ( .A(n1912), .Y(n313) );
  NAND2X1TS U705 ( .A(n225), .B(n1571), .Y(n227) );
  INVX2TS U706 ( .A(n1), .Y(n1432) );
  INVX2TS U707 ( .A(n1432), .Y(n914) );
  CLKBUFX2TS U708 ( .A(n914), .Y(n237) );
  INVX2TS U709 ( .A(n237), .Y(n258) );
  INVX2TS U710 ( .A(n10), .Y(n1690) );
  OR2X1TS U711 ( .A(n225), .B(n1690), .Y(n1420) );
  CLKBUFX2TS U712 ( .A(n1420), .Y(n912) );
  INVX2TS U713 ( .A(n912), .Y(n241) );
  OR2X1TS U714 ( .A(n1568), .B(n227), .Y(n246) );
  INVX2TS U715 ( .A(n246), .Y(n1421) );
  AOI22X1TS U716 ( .A0(n241), .A1(\destinationAddressbuffer[5][8] ), .B0(n1421), .B1(n711), .Y(n232) );
  INVX2TS U717 ( .A(n1561), .Y(n1564) );
  NAND2BX1TS U718 ( .AN(n227), .B(n226), .Y(n229) );
  INVX2TS U719 ( .A(n254), .Y(n1424) );
  OR2X1TS U720 ( .A(n1561), .B(n229), .Y(n248) );
  INVX2TS U721 ( .A(n248), .Y(n230) );
  INVX2TS U722 ( .A(n230), .Y(n901) );
  INVX2TS U723 ( .A(n901), .Y(n242) );
  AOI22X1TS U724 ( .A0(n1434), .A1(n402), .B0(n242), .B1(n325), .Y(n231) );
  OAI211XLTS U725 ( .A0(n258), .A1(n233), .B0(n232), .C0(n231), .Y(n1177) );
  INVX2TS U726 ( .A(n246), .Y(n1715) );
  AOI22X1TS U727 ( .A0(n241), .A1(\destinationAddressbuffer[5][9] ), .B0(n247), 
        .B1(n726), .Y(n235) );
  INVX2TS U728 ( .A(n248), .Y(n1693) );
  AOI22X1TS U729 ( .A0(n1424), .A1(n407), .B0(n1693), .B1(n337), .Y(n234) );
  OAI211XLTS U730 ( .A0(n258), .A1(n236), .B0(n235), .C0(n234), .Y(n1176) );
  INVX2TS U731 ( .A(n237), .Y(n268) );
  INVX2TS U732 ( .A(n246), .Y(n1692) );
  AOI22X1TS U733 ( .A0(n241), .A1(\destinationAddressbuffer[5][10] ), .B0(
        n1692), .B1(n743), .Y(n239) );
  INVX2TS U734 ( .A(n254), .Y(n1694) );
  INVX2TS U735 ( .A(n1694), .Y(n260) );
  INVX2TS U736 ( .A(n260), .Y(n908) );
  INVX2TS U737 ( .A(n248), .Y(n1444) );
  AOI22X1TS U738 ( .A0(n908), .A1(n397), .B0(n1444), .B1(n345), .Y(n238) );
  OAI211XLTS U739 ( .A0(n268), .A1(n240), .B0(n239), .C0(n238), .Y(n1175) );
  AOI22X1TS U740 ( .A0(n241), .A1(\destinationAddressbuffer[5][11] ), .B0(n259), .B1(n759), .Y(n244) );
  INVX2TS U741 ( .A(n254), .Y(n1446) );
  AOI22X1TS U742 ( .A0(n1446), .A1(n414), .B0(n242), .B1(n330), .Y(n243) );
  OAI211XLTS U743 ( .A0(n258), .A1(n245), .B0(n244), .C0(n243), .Y(n1174) );
  INVX2TS U744 ( .A(n912), .Y(n1712) );
  INVX2TS U745 ( .A(n246), .Y(n247) );
  INVX2TS U746 ( .A(n247), .Y(n913) );
  INVX2TS U747 ( .A(n913), .Y(n259) );
  AOI22X1TS U748 ( .A0(n1712), .A1(writeOutbuffer[5]), .B0(n259), .B1(n541), 
        .Y(n250) );
  INVX2TS U749 ( .A(n248), .Y(n1422) );
  AOI22X1TS U750 ( .A0(n1424), .A1(n418), .B0(n1422), .B1(n351), .Y(n249) );
  OAI211XLTS U751 ( .A0(n268), .A1(n295), .B0(n250), .C0(n249), .Y(n1223) );
  AOI22X1TS U752 ( .A0(n264), .A1(\destinationAddressbuffer[5][6] ), .B0(n1715), .B1(n686), .Y(n252) );
  AOI22X1TS U753 ( .A0(n1694), .A1(n429), .B0(n230), .B1(n361), .Y(n251) );
  OAI211XLTS U754 ( .A0(n268), .A1(n253), .B0(n252), .C0(n251), .Y(n1179) );
  AOI22X1TS U755 ( .A0(n264), .A1(\destinationAddressbuffer[5][7] ), .B0(n1421), .B1(n700), .Y(n256) );
  INVX2TS U756 ( .A(n254), .Y(n1434) );
  AOI22X1TS U757 ( .A0(n1434), .A1(n434), .B0(n1422), .B1(n356), .Y(n255) );
  OAI211XLTS U758 ( .A0(n258), .A1(n257), .B0(n256), .C0(n255), .Y(n1178) );
  AOI22X1TS U759 ( .A0(n264), .A1(\destinationAddressbuffer[5][5] ), .B0(n259), 
        .B1(n666), .Y(n262) );
  INVX2TS U760 ( .A(n260), .Y(n1701) );
  AOI22X1TS U761 ( .A0(n1701), .A1(n421), .B0(n1444), .B1(n367), .Y(n261) );
  OAI211XLTS U762 ( .A0(n1432), .A1(n263), .B0(n262), .C0(n261), .Y(n1180) );
  AOI22X1TS U763 ( .A0(n264), .A1(\destinationAddressbuffer[5][4] ), .B0(n1692), .B1(n654), .Y(n266) );
  AOI22X1TS U764 ( .A0(n1446), .A1(n425), .B0(n242), .B1(n374), .Y(n265) );
  OAI211XLTS U765 ( .A0(n268), .A1(n267), .B0(n266), .C0(n265), .Y(n1181) );
  AOI31XLTS U766 ( .A0(n442), .A1(n385), .A2(n313), .B0(n1574), .Y(n273) );
  AOI21X1TS U767 ( .A0(n277), .A1(n273), .B0(n27), .Y(n276) );
  NAND2X1TS U768 ( .A(n276), .B(n1582), .Y(n278) );
  INVX2TS U769 ( .A(n274), .Y(n1402) );
  INVX2TS U770 ( .A(n1402), .Y(n937) );
  CLKBUFX2TS U771 ( .A(n937), .Y(n287) );
  INVX2TS U772 ( .A(n287), .Y(n304) );
  INVX2TS U773 ( .A(n275), .Y(n934) );
  INVX2TS U774 ( .A(n934), .Y(n1720) );
  CLKBUFX2TS U775 ( .A(n1393), .Y(n935) );
  INVX2TS U776 ( .A(n935), .Y(n292) );
  OR2X1TS U777 ( .A(n1578), .B(n278), .Y(n291) );
  INVX2TS U778 ( .A(n291), .Y(n1394) );
  AOI22X1TS U779 ( .A0(n292), .A1(\destinationAddressbuffer[4][10] ), .B0(
        n1394), .B1(n342), .Y(n282) );
  INVX2TS U780 ( .A(n5), .Y(n280) );
  INVX2TS U781 ( .A(n280), .Y(n919) );
  INVX2TS U782 ( .A(n919), .Y(n288) );
  AOI22X1TS U783 ( .A0(n284), .A1(n746), .B0(n288), .B1(n397), .Y(n281) );
  OAI211XLTS U784 ( .A0(n304), .A1(n39), .B0(n282), .C0(n281), .Y(n1163) );
  INVX2TS U785 ( .A(n287), .Y(n307) );
  INVX2TS U786 ( .A(n291), .Y(n283) );
  INVX2TS U787 ( .A(n283), .Y(n936) );
  INVX2TS U788 ( .A(n936), .Y(n298) );
  AOI22X1TS U789 ( .A0(n292), .A1(\destinationAddressbuffer[4][8] ), .B0(n298), 
        .B1(n318), .Y(n286) );
  INVX2TS U790 ( .A(n3), .Y(n284) );
  INVX2TS U791 ( .A(n284), .Y(n939) );
  INVX2TS U792 ( .A(n939), .Y(n301) );
  INVX2TS U793 ( .A(n5), .Y(n1723) );
  AOI22X1TS U794 ( .A0(n301), .A1(n712), .B0(n1723), .B1(n402), .Y(n285) );
  OAI211XLTS U795 ( .A0(n307), .A1(n44), .B0(n286), .C0(n285), .Y(n1165) );
  INVX2TS U796 ( .A(n291), .Y(n1722) );
  AOI22X1TS U797 ( .A0(n292), .A1(\destinationAddressbuffer[4][11] ), .B0(
        n1722), .B1(n329), .Y(n290) );
  INVX2TS U798 ( .A(n3), .Y(n1739) );
  AOI22X1TS U799 ( .A0(n1739), .A1(n762), .B0(n288), .B1(n414), .Y(n289) );
  OAI211XLTS U800 ( .A0(n304), .A1(n30), .B0(n290), .C0(n289), .Y(n1162) );
  INVX2TS U801 ( .A(n291), .Y(n1747) );
  AOI22X1TS U802 ( .A0(n292), .A1(\destinationAddressbuffer[4][9] ), .B0(n1747), .B1(n336), .Y(n294) );
  INVX2TS U803 ( .A(n3), .Y(n1749) );
  INVX2TS U804 ( .A(n5), .Y(n1748) );
  AOI22X1TS U805 ( .A0(n1749), .A1(n727), .B0(n280), .B1(n407), .Y(n293) );
  OAI211XLTS U806 ( .A0(n304), .A1(n48), .B0(n294), .C0(n293), .Y(n1164) );
  INVX2TS U807 ( .A(n935), .Y(n1743) );
  AOI22X1TS U808 ( .A0(n1743), .A1(writeOutbuffer[4]), .B0(n298), .B1(n349), 
        .Y(n297) );
  INVX2TS U809 ( .A(n3), .Y(n1412) );
  INVX2TS U810 ( .A(n5), .Y(n1395) );
  AOI22X1TS U811 ( .A0(n1412), .A1(n543), .B0(n1395), .B1(n418), .Y(n296) );
  OAI211XLTS U812 ( .A0(n307), .A1(n53), .B0(n297), .C0(n296), .Y(n1222) );
  INVX2TS U813 ( .A(n1393), .Y(n308) );
  AOI22X1TS U814 ( .A0(n308), .A1(\destinationAddressbuffer[4][4] ), .B0(n298), 
        .B1(n371), .Y(n300) );
  AOI22X1TS U815 ( .A0(n284), .A1(n656), .B0(n1723), .B1(n425), .Y(n299) );
  OAI211XLTS U816 ( .A0(n307), .A1(n61), .B0(n300), .C0(n299), .Y(n1169) );
  AOI22X1TS U817 ( .A0(n308), .A1(\destinationAddressbuffer[4][6] ), .B0(n283), 
        .B1(n360), .Y(n303) );
  AOI22X1TS U818 ( .A0(n301), .A1(n688), .B0(n280), .B1(n429), .Y(n302) );
  OAI211XLTS U819 ( .A0(n304), .A1(n58), .B0(n303), .C0(n302), .Y(n1167) );
  AOI22X1TS U820 ( .A0(n308), .A1(\destinationAddressbuffer[4][7] ), .B0(n1722), .B1(n355), .Y(n306) );
  AOI22X1TS U821 ( .A0(n284), .A1(n701), .B0(n1395), .B1(n434), .Y(n305) );
  OAI211XLTS U822 ( .A0(n307), .A1(n72), .B0(n306), .C0(n305), .Y(n1166) );
  AOI22X1TS U823 ( .A0(n308), .A1(\destinationAddressbuffer[4][5] ), .B0(n1394), .B1(n366), .Y(n310) );
  AOI22X1TS U824 ( .A0(n1412), .A1(n668), .B0(n288), .B1(n421), .Y(n309) );
  OAI211XLTS U825 ( .A0(n1402), .A1(n66), .B0(n310), .C0(n309), .Y(n1168) );
  AOI31XLTS U826 ( .A0(n19), .A1(n313), .A2(n441), .B0(n1607), .Y(n314) );
  AOI21X1TS U827 ( .A0(n319), .A1(n314), .B0(n438), .Y(n316) );
  NAND2X1TS U828 ( .A(n316), .B(n1615), .Y(n320) );
  INVX2TS U829 ( .A(n315), .Y(n1083) );
  INVX2TS U830 ( .A(n1083), .Y(n1009) );
  CLKBUFX2TS U831 ( .A(n1009), .Y(n335) );
  INVX2TS U832 ( .A(n335), .Y(n365) );
  OR2X1TS U833 ( .A(n480), .B(n1615), .Y(n1078) );
  INVX2TS U834 ( .A(n1078), .Y(n1836) );
  OR2X1TS U835 ( .A(n316), .B(n1836), .Y(n995) );
  INVX2TS U836 ( .A(n995), .Y(n343) );
  OR2X1TS U837 ( .A(n1611), .B(n320), .Y(n341) );
  INVX2TS U838 ( .A(n341), .Y(n317) );
  INVX2TS U839 ( .A(n317), .Y(n1008) );
  INVX2TS U840 ( .A(n1008), .Y(n372) );
  AOI22X1TS U841 ( .A0(n343), .A1(\destinationAddressbuffer[1][8] ), .B0(n372), 
        .B1(n318), .Y(n328) );
  INVX2TS U842 ( .A(n344), .Y(n1095) );
  OR2X1TS U843 ( .A(n1604), .B(n323), .Y(n350) );
  INVX2TS U844 ( .A(n350), .Y(n324) );
  INVX2TS U845 ( .A(n324), .Y(n989) );
  INVX2TS U846 ( .A(n989), .Y(n331) );
  AOI22X1TS U847 ( .A0(n1095), .A1(n326), .B0(n331), .B1(n325), .Y(n327) );
  OAI211XLTS U848 ( .A0(n365), .A1(n44), .B0(n328), .C0(n327), .Y(n1129) );
  INVX2TS U849 ( .A(n341), .Y(n1808) );
  AOI22X1TS U850 ( .A0(n343), .A1(\destinationAddressbuffer[1][11] ), .B0(
        n1808), .B1(n329), .Y(n334) );
  INVX2TS U851 ( .A(n344), .Y(n1812) );
  AOI22X1TS U852 ( .A0(n1812), .A1(n332), .B0(n331), .B1(n330), .Y(n333) );
  OAI211XLTS U853 ( .A0(n365), .A1(n30), .B0(n334), .C0(n333), .Y(n1126) );
  INVX2TS U854 ( .A(n335), .Y(n378) );
  INVX2TS U855 ( .A(n341), .Y(n1839) );
  AOI22X1TS U856 ( .A0(n343), .A1(\destinationAddressbuffer[1][9] ), .B0(n1839), .B1(n336), .Y(n340) );
  INVX2TS U857 ( .A(n344), .Y(n1011) );
  INVX2TS U858 ( .A(n350), .Y(n1810) );
  AOI22X1TS U859 ( .A0(n1011), .A1(n338), .B0(n1810), .B1(n337), .Y(n339) );
  OAI211XLTS U860 ( .A0(n378), .A1(n48), .B0(n340), .C0(n339), .Y(n1128) );
  INVX2TS U861 ( .A(n341), .Y(n1073) );
  AOI22X1TS U862 ( .A0(n343), .A1(\destinationAddressbuffer[1][10] ), .B0(
        n1073), .B1(n342), .Y(n348) );
  INVX2TS U863 ( .A(n344), .Y(n1084) );
  INVX2TS U864 ( .A(n350), .Y(n1094) );
  AOI22X1TS U865 ( .A0(n322), .A1(n346), .B0(n1094), .B1(n345), .Y(n347) );
  OAI211XLTS U866 ( .A0(n365), .A1(n39), .B0(n348), .C0(n347), .Y(n1127) );
  CLKBUFX2TS U867 ( .A(n995), .Y(n1616) );
  INVX2TS U868 ( .A(n1616), .Y(n1835) );
  AOI22X1TS U869 ( .A0(n1835), .A1(writeOutbuffer[1]), .B0(n372), .B1(n349), 
        .Y(n354) );
  INVX2TS U870 ( .A(n350), .Y(n1074) );
  AOI22X1TS U871 ( .A0(n1095), .A1(n352), .B0(n1074), .B1(n351), .Y(n353) );
  OAI211XLTS U872 ( .A0(n378), .A1(n53), .B0(n354), .C0(n353), .Y(n1219) );
  INVX2TS U873 ( .A(n995), .Y(n373) );
  AOI22X1TS U874 ( .A0(n373), .A1(\destinationAddressbuffer[1][7] ), .B0(n1808), .B1(n355), .Y(n359) );
  AOI22X1TS U875 ( .A0(n1011), .A1(n357), .B0(n1074), .B1(n356), .Y(n358) );
  OAI211XLTS U876 ( .A0(n378), .A1(n72), .B0(n359), .C0(n358), .Y(n1130) );
  AOI22X1TS U877 ( .A0(n373), .A1(\destinationAddressbuffer[1][6] ), .B0(n317), 
        .B1(n360), .Y(n364) );
  AOI22X1TS U878 ( .A0(n1084), .A1(n362), .B0(n324), .B1(n361), .Y(n363) );
  OAI211XLTS U879 ( .A0(n365), .A1(n58), .B0(n364), .C0(n363), .Y(n1131) );
  AOI22X1TS U880 ( .A0(n373), .A1(\destinationAddressbuffer[1][5] ), .B0(n1073), .B1(n366), .Y(n370) );
  AOI22X1TS U881 ( .A0(n321), .A1(n368), .B0(n1094), .B1(n367), .Y(n369) );
  OAI211XLTS U882 ( .A0(n1083), .A1(n66), .B0(n370), .C0(n369), .Y(n1132) );
  AOI22X1TS U883 ( .A0(n373), .A1(\destinationAddressbuffer[1][4] ), .B0(n372), 
        .B1(n371), .Y(n377) );
  AOI22X1TS U884 ( .A0(n1095), .A1(n375), .B0(n331), .B1(n374), .Y(n376) );
  OAI211XLTS U885 ( .A0(n378), .A1(n61), .B0(n377), .C0(n376), .Y(n1133) );
  AOI31XLTS U886 ( .A0(n385), .A1(n387), .A2(n481), .B0(n1621), .Y(n386) );
  AOI21X1TS U887 ( .A0(n393), .A1(n386), .B0(n480), .Y(n391) );
  NAND2X1TS U888 ( .A(n391), .B(n1630), .Y(n394) );
  INVX2TS U889 ( .A(n389), .Y(n1055) );
  INVX2TS U890 ( .A(n1055), .Y(n1039) );
  CLKBUFX2TS U891 ( .A(n1039), .Y(n405) );
  INVX2TS U892 ( .A(n405), .Y(n428) );
  INVX2TS U893 ( .A(n11), .Y(n1846) );
  CLKBUFX2TS U894 ( .A(n1024), .Y(n1037) );
  INVX2TS U895 ( .A(n1037), .Y(n413) );
  OR2X1TS U896 ( .A(n1626), .B(n394), .Y(n410) );
  INVX2TS U897 ( .A(n410), .Y(n1849) );
  AOI22X1TS U898 ( .A0(n413), .A1(\destinationAddressbuffer[0][10] ), .B0(
        n1849), .B1(n392), .Y(n399) );
  INVX2TS U899 ( .A(n6), .Y(n396) );
  INVX2TS U900 ( .A(n396), .Y(n1018) );
  INVX2TS U901 ( .A(n1018), .Y(n415) );
  AOI22X1TS U902 ( .A0(n401), .A1(n746), .B0(n415), .B1(n397), .Y(n398) );
  OAI211XLTS U903 ( .A0(n428), .A1(n39), .B0(n399), .C0(n398), .Y(n1115) );
  INVX2TS U904 ( .A(n410), .Y(n1047) );
  AOI22X1TS U905 ( .A0(n413), .A1(\destinationAddressbuffer[0][8] ), .B0(n1047), .B1(n400), .Y(n404) );
  INVX2TS U906 ( .A(n4), .Y(n401) );
  INVX2TS U907 ( .A(n401), .Y(n1041) );
  INVX2TS U908 ( .A(n1041), .Y(n430) );
  INVX2TS U909 ( .A(n6), .Y(n1851) );
  AOI22X1TS U910 ( .A0(n430), .A1(n712), .B0(n1851), .B1(n402), .Y(n403) );
  OAI211XLTS U911 ( .A0(n428), .A1(n44), .B0(n404), .C0(n403), .Y(n1117) );
  INVX2TS U912 ( .A(n405), .Y(n437) );
  INVX2TS U913 ( .A(n410), .Y(n1881) );
  AOI22X1TS U914 ( .A0(n413), .A1(\destinationAddressbuffer[0][9] ), .B0(n411), 
        .B1(n406), .Y(n409) );
  INVX2TS U915 ( .A(n4), .Y(n1885) );
  INVX2TS U916 ( .A(n6), .Y(n1883) );
  AOI22X1TS U917 ( .A0(n1885), .A1(n727), .B0(n1883), .B1(n407), .Y(n408) );
  OAI211XLTS U918 ( .A0(n437), .A1(n48), .B0(n409), .C0(n408), .Y(n1116) );
  INVX2TS U919 ( .A(n410), .Y(n411) );
  INVX2TS U920 ( .A(n411), .Y(n1038) );
  INVX2TS U921 ( .A(n1038), .Y(n424) );
  AOI22X1TS U922 ( .A0(n413), .A1(\destinationAddressbuffer[0][11] ), .B0(n424), .B1(n412), .Y(n417) );
  INVX2TS U923 ( .A(n4), .Y(n1873) );
  AOI22X1TS U924 ( .A0(n1873), .A1(n762), .B0(n415), .B1(n414), .Y(n416) );
  OAI211XLTS U925 ( .A0(n428), .A1(n30), .B0(n417), .C0(n416), .Y(n1114) );
  INVX2TS U926 ( .A(n1024), .Y(n1877) );
  AOI22X1TS U927 ( .A0(n1877), .A1(writeOutbuffer[0]), .B0(n1849), .B1(
        writeIn_WEST), .Y(n420) );
  INVX2TS U928 ( .A(n4), .Y(n1065) );
  INVX2TS U929 ( .A(n6), .Y(n1048) );
  AOI22X1TS U930 ( .A0(n1065), .A1(n543), .B0(n1048), .B1(n418), .Y(n419) );
  OAI211XLTS U931 ( .A0(n437), .A1(n53), .B0(n420), .C0(n419), .Y(n1218) );
  INVX2TS U932 ( .A(n1024), .Y(n433) );
  AOI22X1TS U933 ( .A0(n433), .A1(\destinationAddressbuffer[0][5] ), .B0(n1881), .B1(destinationAddressIn_WEST[5]), .Y(n423) );
  AOI22X1TS U934 ( .A0(n1065), .A1(n668), .B0(n415), .B1(n421), .Y(n422) );
  OAI211XLTS U935 ( .A0(n437), .A1(n66), .B0(n423), .C0(n422), .Y(n1120) );
  AOI22X1TS U936 ( .A0(n433), .A1(\destinationAddressbuffer[0][4] ), .B0(n424), 
        .B1(destinationAddressIn_WEST[4]), .Y(n427) );
  AOI22X1TS U937 ( .A0(n401), .A1(n656), .B0(n1851), .B1(n425), .Y(n426) );
  OAI211XLTS U938 ( .A0(n428), .A1(n61), .B0(n427), .C0(n426), .Y(n1121) );
  AOI22X1TS U939 ( .A0(n433), .A1(\destinationAddressbuffer[0][6] ), .B0(n1047), .B1(destinationAddressIn_WEST[6]), .Y(n432) );
  AOI22X1TS U940 ( .A0(n430), .A1(n688), .B0(n396), .B1(n429), .Y(n431) );
  OAI211XLTS U941 ( .A0(n1055), .A1(n58), .B0(n432), .C0(n431), .Y(n1119) );
  AOI22X1TS U942 ( .A0(n433), .A1(\destinationAddressbuffer[0][7] ), .B0(n424), 
        .B1(destinationAddressIn_WEST[7]), .Y(n436) );
  AOI22X1TS U943 ( .A0(n401), .A1(n701), .B0(n1048), .B1(n434), .Y(n435) );
  OAI211XLTS U944 ( .A0(n437), .A1(n72), .B0(n436), .C0(n435), .Y(n1118) );
  INVX2TS U945 ( .A(reset), .Y(n489) );
  NAND2X1TS U946 ( .A(n489), .B(n1906), .Y(n502) );
  INVX2TS U947 ( .A(n1910), .Y(n529) );
  INVX2TS U948 ( .A(n1912), .Y(n451) );
  INVX2TS U949 ( .A(n1904), .Y(n439) );
  NAND2X1TS U950 ( .A(n440), .B(n439), .Y(n454) );
  INVX2TS U951 ( .A(n1915), .Y(n442) );
  INVX2TS U952 ( .A(n1907), .Y(n525) );
  INVX2TS U953 ( .A(n1908), .Y(n528) );
  AOI22X1TS U954 ( .A0(n442), .A1(n525), .B0(n528), .B1(n441), .Y(n445) );
  INVX2TS U955 ( .A(n444), .Y(n450) );
  INVX2TS U956 ( .A(n1917), .Y(n526) );
  AOI21X1TS U957 ( .A0(n526), .A1(n448), .B0(n447), .Y(n460) );
  ADDFX2TS U958 ( .A(n450), .B(n510), .CI(n449), .CO(n452), .S(n465) );
  ADDHX1TS U959 ( .A(n453), .B(n452), .CO(n464), .S(n466) );
  INVX2TS U960 ( .A(n466), .Y(n455) );
  OAI21XLTS U961 ( .A0(n491), .A1(n1917), .B0(n454), .Y(n486) );
  AOI21X1TS U962 ( .A0(n456), .A1(n455), .B0(n486), .Y(n458) );
  OAI22X1TS U963 ( .A0(n456), .A1(n455), .B0(n462), .B1(n461), .Y(n457) );
  AOI21X1TS U964 ( .A0(n465), .A1(n458), .B0(n457), .Y(n459) );
  AOI211X1TS U965 ( .A0(n462), .A1(n461), .B0(n460), .C0(n459), .Y(n463) );
  INVX2TS U966 ( .A(n463), .Y(n467) );
  NAND2X1TS U967 ( .A(n467), .B(n464), .Y(n471) );
  XNOR2X1TS U968 ( .A(n469), .B(n468), .Y(n470) );
  INVX2TS U969 ( .A(n494), .Y(n478) );
  INVX2TS U970 ( .A(n1908), .Y(n524) );
  INVX2TS U971 ( .A(n1917), .Y(n523) );
  ADDHXLTS U972 ( .A(n440), .B(n472), .CO(n474), .S(n490) );
  XNOR2X1TS U973 ( .A(n1911), .B(n492), .Y(n475) );
  NAND2X1TS U974 ( .A(n523), .B(n529), .Y(n527) );
  OAI21XLTS U975 ( .A0(n526), .A1(n1911), .B0(n527), .Y(n501) );
  INVX2TS U976 ( .A(n1907), .Y(n530) );
  NOR2XLTS U977 ( .A(n527), .B(n525), .Y(n832) );
  CLKBUFX2TS U978 ( .A(n832), .Y(n792) );
  CLKBUFX2TS U979 ( .A(n792), .Y(n812) );
  AOI21X1TS U980 ( .A0(n527), .A1(n530), .B0(n812), .Y(n498) );
  OAI22X1TS U981 ( .A0(n482), .A1(n501), .B0(n481), .B1(n498), .Y(n483) );
  AOI221XLTS U982 ( .A0(n501), .A1(n485), .B0(n484), .B1(n498), .C0(n483), .Y(
        n487) );
  AOI21X1TS U983 ( .A0(n487), .A1(n486), .B0(n1906), .Y(n488) );
  CLKBUFX2TS U984 ( .A(n1905), .Y(n638) );
  CLKBUFX2TS U985 ( .A(n638), .Y(n605) );
  NAND2X1TS U986 ( .A(n489), .B(n605), .Y(n500) );
  AOI22X1TS U987 ( .A0(n1904), .A1(n502), .B0(n500), .B1(n439), .Y(n1336) );
  INVX2TS U988 ( .A(n498), .Y(n499) );
  OAI22X1TS U989 ( .A0(n530), .A1(n502), .B0(n499), .B1(n500), .Y(n1331) );
  OAI22X1TS U990 ( .A0(n13), .A1(n502), .B0(n501), .B1(n500), .Y(n1330) );
  CLKBUFX2TS U991 ( .A(readIn_SOUTH), .Y(n1620) );
  CLKBUFX2TS U992 ( .A(n1620), .Y(n1563) );
  CLKBUFX2TS U993 ( .A(n1905), .Y(n838) );
  CLKBUFX2TS U994 ( .A(n542), .Y(n844) );
  CLKBUFX2TS U995 ( .A(readIn_WEST), .Y(n1628) );
  CLKBUFX2TS U996 ( .A(n1628), .Y(n1613) );
  INVX2TS U997 ( .A(n1905), .Y(n519) );
  NOR4XLTS U998 ( .A(n513), .B(n512), .C(n444), .D(n507), .Y(n611) );
  CLKBUFX2TS U999 ( .A(n611), .Y(n625) );
  CLKBUFX2TS U1000 ( .A(n625), .Y(n805) );
  CLKBUFX2TS U1001 ( .A(n805), .Y(n562) );
  AOI22X1TS U1002 ( .A0(n1563), .A1(n844), .B0(n1613), .B1(n562), .Y(n540) );
  CLKBUFX2TS U1003 ( .A(readIn_NORTH), .Y(n1619) );
  CLKBUFX2TS U1004 ( .A(n1619), .Y(n1562) );
  CLKBUFX2TS U1005 ( .A(n687), .Y(n561) );
  NOR4XLTS U1006 ( .A(n511), .B(n508), .C(n509), .D(n507), .Y(n587) );
  CLKBUFX2TS U1007 ( .A(n587), .Y(n598) );
  CLKBUFX2TS U1008 ( .A(n598), .Y(n773) );
  CLKBUFX2TS U1009 ( .A(n773), .Y(n822) );
  AOI22X1TS U1010 ( .A0(n1562), .A1(n561), .B0(readIn_EAST), .B1(n822), .Y(
        n539) );
  NOR3XLTS U1011 ( .A(n512), .B(readReady), .C(n444), .Y(n515) );
  NOR3XLTS U1012 ( .A(n511), .B(n510), .C(n509), .Y(n514) );
  NAND4XLTS U1013 ( .A(n519), .B(n518), .C(n517), .D(n516), .Y(n730) );
  INVX2TS U1014 ( .A(n730), .Y(n520) );
  INVX2TS U1015 ( .A(n520), .Y(n578) );
  INVX2TS U1016 ( .A(n578), .Y(n521) );
  NOR3XLTS U1017 ( .A(n523), .B(n524), .C(n1910), .Y(n714) );
  CLKBUFX2TS U1018 ( .A(n714), .Y(n626) );
  CLKBUFX2TS U1019 ( .A(n626), .Y(n564) );
  NOR3XLTS U1020 ( .A(n526), .B(n1911), .C(n524), .Y(n689) );
  CLKBUFX2TS U1021 ( .A(n689), .Y(n627) );
  CLKBUFX2TS U1022 ( .A(n627), .Y(n563) );
  AOI22X1TS U1023 ( .A0(readOutbuffer[2]), .A1(n564), .B0(readOutbuffer[0]), 
        .B1(n563), .Y(n534) );
  NOR3XLTS U1024 ( .A(n523), .B(n13), .C(n525), .Y(n715) );
  CLKBUFX2TS U1025 ( .A(n715), .Y(n628) );
  CLKBUFX2TS U1026 ( .A(n628), .Y(n566) );
  NOR3XLTS U1027 ( .A(n526), .B(n529), .C(n530), .Y(n690) );
  CLKBUFX2TS U1028 ( .A(n690), .Y(n629) );
  CLKBUFX2TS U1029 ( .A(n629), .Y(n565) );
  AOI22X1TS U1030 ( .A0(readOutbuffer[6]), .A1(n566), .B0(readOutbuffer[4]), 
        .B1(n565), .Y(n533) );
  NOR2XLTS U1031 ( .A(n528), .B(n527), .Y(n716) );
  CLKBUFX2TS U1032 ( .A(n716), .Y(n630) );
  CLKBUFX2TS U1033 ( .A(n630), .Y(n568) );
  NOR3XLTS U1034 ( .A(n529), .B(n528), .C(n1917), .Y(n691) );
  CLKBUFX2TS U1035 ( .A(n691), .Y(n631) );
  CLKBUFX2TS U1036 ( .A(n631), .Y(n567) );
  AOI22X1TS U1037 ( .A0(readOutbuffer[3]), .A1(n568), .B0(readOutbuffer[1]), 
        .B1(n567), .Y(n532) );
  CLKBUFX2TS U1038 ( .A(n832), .Y(n853) );
  NOR3XLTS U1039 ( .A(n1911), .B(n439), .C(n530), .Y(n854) );
  CLKBUFX2TS U1040 ( .A(n854), .Y(n632) );
  CLKBUFX2TS U1041 ( .A(n632), .Y(n569) );
  AOI22X1TS U1042 ( .A0(readOutbuffer[7]), .A1(n853), .B0(readOutbuffer[5]), 
        .B1(n569), .Y(n531) );
  NAND4XLTS U1043 ( .A(n534), .B(n533), .C(n532), .D(n531), .Y(n535) );
  AOI22X1TS U1044 ( .A0(readOut), .A1(n549), .B0(n605), .B1(n535), .Y(n538) );
  INVX2TS U1045 ( .A(n12), .Y(n799) );
  CLKBUFX2TS U1046 ( .A(n773), .Y(n744) );
  AOI22X1TS U1047 ( .A0(writeIn_EAST), .A1(n744), .B0(n541), .B1(n562), .Y(
        n552) );
  CLKBUFX2TS U1048 ( .A(n542), .Y(n667) );
  CLKBUFX2TS U1049 ( .A(n667), .Y(n761) );
  AOI22X1TS U1050 ( .A0(writeIn_NORTH), .A1(n561), .B0(n543), .B1(n761), .Y(
        n551) );
  AOI22X1TS U1051 ( .A0(writeOutbuffer[2]), .A1(n564), .B0(writeOutbuffer[0]), 
        .B1(n563), .Y(n547) );
  AOI22X1TS U1052 ( .A0(writeOutbuffer[6]), .A1(n566), .B0(writeOutbuffer[4]), 
        .B1(n565), .Y(n546) );
  AOI22X1TS U1053 ( .A0(writeOutbuffer[3]), .A1(n568), .B0(writeOutbuffer[1]), 
        .B1(n567), .Y(n545) );
  AOI22X1TS U1054 ( .A0(writeOutbuffer[7]), .A1(n853), .B0(writeOutbuffer[5]), 
        .B1(n569), .Y(n544) );
  NAND4XLTS U1055 ( .A(n547), .B(n546), .C(n545), .D(n544), .Y(n548) );
  AOI22X1TS U1056 ( .A0(writeOut), .A1(n549), .B0(n605), .B1(n548), .Y(n550)
         );
  CLKBUFX2TS U1057 ( .A(requesterAddressIn_NORTH[0]), .Y(n1019) );
  CLKBUFX2TS U1058 ( .A(n1019), .Y(n990) );
  CLKBUFX2TS U1059 ( .A(requesterAddressIn_EAST[0]), .Y(n1017) );
  CLKBUFX2TS U1060 ( .A(n1017), .Y(n988) );
  AOI22X1TS U1061 ( .A0(n990), .A1(n561), .B0(n988), .B1(n598), .Y(n560) );
  CLKBUFX2TS U1062 ( .A(requesterAddressIn_SOUTH[0]), .Y(n1020) );
  CLKBUFX2TS U1063 ( .A(n1020), .Y(n991) );
  CLKBUFX2TS U1064 ( .A(n667), .Y(n655) );
  CLKBUFX2TS U1065 ( .A(requesterAddressIn_WEST[0]), .Y(n918) );
  CLKBUFX2TS U1066 ( .A(n918), .Y(n946) );
  AOI22X1TS U1067 ( .A0(n991), .A1(n655), .B0(n946), .B1(n562), .Y(n559) );
  INVX2TS U1068 ( .A(n730), .Y(n682) );
  CLKBUFX2TS U1069 ( .A(n638), .Y(n593) );
  AOI22X1TS U1070 ( .A0(\requesterAddressbuffer[2][0] ), .A1(n564), .B0(
        \requesterAddressbuffer[0][0] ), .B1(n563), .Y(n556) );
  AOI22X1TS U1071 ( .A0(\requesterAddressbuffer[6][0] ), .A1(n566), .B0(
        \requesterAddressbuffer[4][0] ), .B1(n565), .Y(n555) );
  AOI22X1TS U1072 ( .A0(\requesterAddressbuffer[3][0] ), .A1(n568), .B0(
        \requesterAddressbuffer[1][0] ), .B1(n567), .Y(n554) );
  CLKBUFX2TS U1073 ( .A(n792), .Y(n748) );
  CLKBUFX2TS U1074 ( .A(n748), .Y(n599) );
  AOI22X1TS U1075 ( .A0(\requesterAddressbuffer[7][0] ), .A1(n599), .B0(
        \requesterAddressbuffer[5][0] ), .B1(n569), .Y(n553) );
  NAND4XLTS U1076 ( .A(n556), .B(n555), .C(n554), .D(n553), .Y(n557) );
  AOI22X1TS U1077 ( .A0(requesterAddressOut[0]), .A1(n682), .B0(n593), .B1(
        n557), .Y(n558) );
  INVX2TS U1078 ( .A(readRequesterAddress[0]), .Y(n944) );
  INVX2TS U1079 ( .A(n944), .Y(n987) );
  INVX2TS U1080 ( .A(n799), .Y(n594) );
  NAND2X1TS U1081 ( .A(n987), .B(n594), .Y(n606) );
  CLKBUFX2TS U1082 ( .A(requesterAddressIn_NORTH[1]), .Y(n1026) );
  CLKBUFX2TS U1083 ( .A(n1026), .Y(n997) );
  CLKBUFX2TS U1084 ( .A(requesterAddressIn_EAST[1]), .Y(n1025) );
  CLKBUFX2TS U1085 ( .A(n1025), .Y(n996) );
  AOI22X1TS U1086 ( .A0(n997), .A1(n561), .B0(n996), .B1(n587), .Y(n577) );
  CLKBUFX2TS U1087 ( .A(requesterAddressIn_SOUTH[1]), .Y(n1027) );
  CLKBUFX2TS U1088 ( .A(n1027), .Y(n998) );
  CLKBUFX2TS U1089 ( .A(n542), .Y(n803) );
  CLKBUFX2TS U1090 ( .A(requesterAddressIn_WEST[1]), .Y(n924) );
  CLKBUFX2TS U1091 ( .A(n924), .Y(n952) );
  AOI22X1TS U1092 ( .A0(n998), .A1(n803), .B0(n952), .B1(n562), .Y(n576) );
  INVX2TS U1093 ( .A(n730), .Y(n779) );
  AOI22X1TS U1094 ( .A0(\requesterAddressbuffer[2][1] ), .A1(n564), .B0(
        \requesterAddressbuffer[0][1] ), .B1(n563), .Y(n573) );
  AOI22X1TS U1095 ( .A0(\requesterAddressbuffer[6][1] ), .A1(n566), .B0(
        \requesterAddressbuffer[4][1] ), .B1(n565), .Y(n572) );
  AOI22X1TS U1096 ( .A0(\requesterAddressbuffer[3][1] ), .A1(n568), .B0(
        \requesterAddressbuffer[1][1] ), .B1(n567), .Y(n571) );
  AOI22X1TS U1097 ( .A0(\requesterAddressbuffer[7][1] ), .A1(n599), .B0(
        \requesterAddressbuffer[5][1] ), .B1(n569), .Y(n570) );
  NAND4XLTS U1098 ( .A(n573), .B(n572), .C(n571), .D(n570), .Y(n574) );
  AOI22X1TS U1099 ( .A0(requesterAddressOut[1]), .A1(n779), .B0(n593), .B1(
        n574), .Y(n575) );
  INVX2TS U1100 ( .A(readRequesterAddress[1]), .Y(n950) );
  INVX2TS U1101 ( .A(n950), .Y(n1636) );
  NAND2X1TS U1102 ( .A(n1636), .B(n594), .Y(n621) );
  CLKBUFX2TS U1103 ( .A(requesterAddressIn_NORTH[2]), .Y(n1032) );
  CLKBUFX2TS U1104 ( .A(n1032), .Y(n1003) );
  CLKBUFX2TS U1105 ( .A(n687), .Y(n610) );
  CLKBUFX2TS U1106 ( .A(requesterAddressIn_EAST[2]), .Y(n1031) );
  CLKBUFX2TS U1107 ( .A(n1031), .Y(n1002) );
  AOI22X1TS U1108 ( .A0(n1003), .A1(n610), .B0(n1002), .B1(n587), .Y(n586) );
  CLKBUFX2TS U1109 ( .A(requesterAddressIn_SOUTH[2]), .Y(n1033) );
  CLKBUFX2TS U1110 ( .A(n1033), .Y(n1004) );
  CLKBUFX2TS U1111 ( .A(requesterAddressIn_WEST[2]), .Y(n929) );
  CLKBUFX2TS U1112 ( .A(n929), .Y(n957) );
  AOI22X1TS U1113 ( .A0(n1004), .A1(n655), .B0(n957), .B1(n625), .Y(n585) );
  INVX2TS U1114 ( .A(n578), .Y(n755) );
  CLKBUFX2TS U1115 ( .A(n626), .Y(n612) );
  AOI22X1TS U1116 ( .A0(\requesterAddressbuffer[2][2] ), .A1(n612), .B0(
        \requesterAddressbuffer[0][2] ), .B1(n689), .Y(n582) );
  CLKBUFX2TS U1117 ( .A(n628), .Y(n613) );
  AOI22X1TS U1118 ( .A0(\requesterAddressbuffer[6][2] ), .A1(n613), .B0(
        \requesterAddressbuffer[4][2] ), .B1(n690), .Y(n581) );
  CLKBUFX2TS U1119 ( .A(n630), .Y(n614) );
  AOI22X1TS U1120 ( .A0(\requesterAddressbuffer[3][2] ), .A1(n614), .B0(
        \requesterAddressbuffer[1][2] ), .B1(n691), .Y(n580) );
  CLKBUFX2TS U1121 ( .A(n632), .Y(n615) );
  AOI22X1TS U1122 ( .A0(\requesterAddressbuffer[7][2] ), .A1(n599), .B0(
        \requesterAddressbuffer[5][2] ), .B1(n615), .Y(n579) );
  NAND4XLTS U1123 ( .A(n582), .B(n581), .C(n580), .D(n579), .Y(n583) );
  AOI22X1TS U1124 ( .A0(requesterAddressOut[2]), .A1(n755), .B0(n593), .B1(
        n583), .Y(n584) );
  INVX2TS U1125 ( .A(readRequesterAddress[2]), .Y(n956) );
  INVX2TS U1126 ( .A(n956), .Y(n1644) );
  NAND2X1TS U1127 ( .A(n1644), .B(n594), .Y(n639) );
  CLKBUFX2TS U1128 ( .A(requesterAddressIn_NORTH[3]), .Y(n1042) );
  CLKBUFX2TS U1129 ( .A(n1042), .Y(n1012) );
  CLKBUFX2TS U1130 ( .A(requesterAddressIn_EAST[3]), .Y(n1040) );
  CLKBUFX2TS U1131 ( .A(n1040), .Y(n1010) );
  AOI22X1TS U1132 ( .A0(n1012), .A1(n610), .B0(n1010), .B1(n587), .Y(n597) );
  CLKBUFX2TS U1133 ( .A(requesterAddressIn_SOUTH[3]), .Y(n1043) );
  CLKBUFX2TS U1134 ( .A(n1043), .Y(n1013) );
  CLKBUFX2TS U1135 ( .A(requesterAddressIn_WEST[3]), .Y(n938) );
  CLKBUFX2TS U1136 ( .A(n938), .Y(n965) );
  AOI22X1TS U1137 ( .A0(n1013), .A1(n803), .B0(n965), .B1(n611), .Y(n596) );
  AOI22X1TS U1138 ( .A0(\requesterAddressbuffer[2][3] ), .A1(n612), .B0(
        \requesterAddressbuffer[0][3] ), .B1(n689), .Y(n591) );
  AOI22X1TS U1139 ( .A0(\requesterAddressbuffer[6][3] ), .A1(n613), .B0(
        \requesterAddressbuffer[4][3] ), .B1(n690), .Y(n590) );
  AOI22X1TS U1140 ( .A0(\requesterAddressbuffer[3][3] ), .A1(n614), .B0(
        \requesterAddressbuffer[1][3] ), .B1(n691), .Y(n589) );
  CLKBUFX2TS U1141 ( .A(n748), .Y(n644) );
  AOI22X1TS U1142 ( .A0(\requesterAddressbuffer[7][3] ), .A1(n644), .B0(
        \requesterAddressbuffer[5][3] ), .B1(n615), .Y(n588) );
  NAND4XLTS U1143 ( .A(n591), .B(n590), .C(n589), .D(n588), .Y(n592) );
  AOI22X1TS U1144 ( .A0(requesterAddressOut[3]), .A1(n521), .B0(n593), .B1(
        n592), .Y(n595) );
  INVX2TS U1145 ( .A(readRequesterAddress[3]), .Y(n963) );
  INVX2TS U1146 ( .A(n963), .Y(n1653) );
  NAND2X1TS U1147 ( .A(n1653), .B(n594), .Y(n650) );
  CLKBUFX2TS U1148 ( .A(destinationAddressIn_NORTH[0]), .Y(n1663) );
  CLKBUFX2TS U1149 ( .A(destinationAddressIn_EAST[0]), .Y(n1807) );
  CLKBUFX2TS U1150 ( .A(n1807), .Y(n1691) );
  CLKBUFX2TS U1151 ( .A(n598), .Y(n643) );
  AOI22X1TS U1152 ( .A0(n1663), .A1(n610), .B0(n1691), .B1(n643), .Y(n609) );
  CLKBUFX2TS U1153 ( .A(destinationAddressIn_WEST[0]), .Y(n1848) );
  AOI22X1TS U1154 ( .A0(destinationAddressIn_SOUTH[0]), .A1(n655), .B0(n1848), 
        .B1(n611), .Y(n608) );
  AOI22X1TS U1155 ( .A0(\destinationAddressbuffer[2][0] ), .A1(n612), .B0(
        \destinationAddressbuffer[0][0] ), .B1(n627), .Y(n603) );
  AOI22X1TS U1156 ( .A0(\destinationAddressbuffer[6][0] ), .A1(n613), .B0(
        \destinationAddressbuffer[4][0] ), .B1(n629), .Y(n602) );
  AOI22X1TS U1157 ( .A0(\destinationAddressbuffer[3][0] ), .A1(n614), .B0(
        \destinationAddressbuffer[1][0] ), .B1(n631), .Y(n601) );
  AOI22X1TS U1158 ( .A0(\destinationAddressbuffer[7][0] ), .A1(n599), .B0(
        \destinationAddressbuffer[5][0] ), .B1(n615), .Y(n600) );
  NAND4XLTS U1159 ( .A(n603), .B(n602), .C(n601), .D(n600), .Y(n604) );
  AOI22X1TS U1160 ( .A0(destinationAddressOut[0]), .A1(n682), .B0(n605), .B1(
        n604), .Y(n607) );
  CLKBUFX2TS U1161 ( .A(destinationAddressIn_NORTH[1]), .Y(n1670) );
  CLKBUFX2TS U1162 ( .A(destinationAddressIn_EAST[1]), .Y(n1818) );
  CLKBUFX2TS U1163 ( .A(n1818), .Y(n1699) );
  AOI22X1TS U1164 ( .A0(n1670), .A1(n610), .B0(n1699), .B1(n643), .Y(n624) );
  CLKBUFX2TS U1165 ( .A(destinationAddressIn_WEST[1]), .Y(n1860) );
  AOI22X1TS U1166 ( .A0(destinationAddressIn_SOUTH[1]), .A1(n803), .B0(n1860), 
        .B1(n611), .Y(n623) );
  AOI22X1TS U1167 ( .A0(\destinationAddressbuffer[2][1] ), .A1(n612), .B0(
        \destinationAddressbuffer[0][1] ), .B1(n627), .Y(n619) );
  AOI22X1TS U1168 ( .A0(\destinationAddressbuffer[6][1] ), .A1(n613), .B0(
        \destinationAddressbuffer[4][1] ), .B1(n629), .Y(n618) );
  AOI22X1TS U1169 ( .A0(\destinationAddressbuffer[3][1] ), .A1(n614), .B0(
        \destinationAddressbuffer[1][1] ), .B1(n631), .Y(n617) );
  AOI22X1TS U1170 ( .A0(\destinationAddressbuffer[7][1] ), .A1(n644), .B0(
        \destinationAddressbuffer[5][1] ), .B1(n615), .Y(n616) );
  NAND4XLTS U1171 ( .A(n619), .B(n618), .C(n617), .D(n616), .Y(n620) );
  AOI22X1TS U1172 ( .A0(destinationAddressOut[1]), .A1(n682), .B0(n638), .B1(
        n620), .Y(n622) );
  CLKBUFX2TS U1173 ( .A(destinationAddressIn_NORTH[2]), .Y(n1677) );
  CLKBUFX2TS U1174 ( .A(n687), .Y(n669) );
  CLKBUFX2TS U1175 ( .A(destinationAddressIn_EAST[2]), .Y(n1828) );
  CLKBUFX2TS U1176 ( .A(n1828), .Y(n1707) );
  AOI22X1TS U1177 ( .A0(n1677), .A1(n669), .B0(n1707), .B1(n643), .Y(n642) );
  CLKBUFX2TS U1178 ( .A(n542), .Y(n783) );
  CLKBUFX2TS U1179 ( .A(destinationAddressIn_WEST[2]), .Y(n1870) );
  CLKBUFX2TS U1180 ( .A(n625), .Y(n665) );
  AOI22X1TS U1181 ( .A0(destinationAddressIn_SOUTH[2]), .A1(n783), .B0(n1870), 
        .B1(n665), .Y(n641) );
  CLKBUFX2TS U1182 ( .A(n626), .Y(n671) );
  CLKBUFX2TS U1183 ( .A(n627), .Y(n670) );
  AOI22X1TS U1184 ( .A0(\destinationAddressbuffer[2][2] ), .A1(n671), .B0(
        \destinationAddressbuffer[0][2] ), .B1(n670), .Y(n636) );
  CLKBUFX2TS U1185 ( .A(n628), .Y(n673) );
  CLKBUFX2TS U1186 ( .A(n629), .Y(n672) );
  AOI22X1TS U1187 ( .A0(\destinationAddressbuffer[6][2] ), .A1(n673), .B0(
        \destinationAddressbuffer[4][2] ), .B1(n672), .Y(n635) );
  CLKBUFX2TS U1188 ( .A(n630), .Y(n675) );
  CLKBUFX2TS U1189 ( .A(n631), .Y(n674) );
  AOI22X1TS U1190 ( .A0(\destinationAddressbuffer[3][2] ), .A1(n675), .B0(
        \destinationAddressbuffer[1][2] ), .B1(n674), .Y(n634) );
  CLKBUFX2TS U1191 ( .A(n632), .Y(n676) );
  AOI22X1TS U1192 ( .A0(\destinationAddressbuffer[7][2] ), .A1(n644), .B0(
        \destinationAddressbuffer[5][2] ), .B1(n676), .Y(n633) );
  NAND4XLTS U1193 ( .A(n636), .B(n635), .C(n634), .D(n633), .Y(n637) );
  AOI22X1TS U1194 ( .A0(destinationAddressOut[2]), .A1(n521), .B0(n638), .B1(
        n637), .Y(n640) );
  CLKBUFX2TS U1195 ( .A(destinationAddressIn_NORTH[3]), .Y(n1684) );
  CLKBUFX2TS U1196 ( .A(destinationAddressIn_EAST[3]), .Y(n1838) );
  CLKBUFX2TS U1197 ( .A(n1838), .Y(n1714) );
  AOI22X1TS U1198 ( .A0(n1684), .A1(n669), .B0(n1714), .B1(n643), .Y(n653) );
  CLKBUFX2TS U1199 ( .A(destinationAddressIn_WEST[3]), .Y(n1880) );
  AOI22X1TS U1200 ( .A0(destinationAddressIn_SOUTH[3]), .A1(n783), .B0(n1880), 
        .B1(n665), .Y(n652) );
  AOI22X1TS U1201 ( .A0(\destinationAddressbuffer[2][3] ), .A1(n671), .B0(
        \destinationAddressbuffer[0][3] ), .B1(n670), .Y(n648) );
  AOI22X1TS U1202 ( .A0(\destinationAddressbuffer[6][3] ), .A1(n673), .B0(
        \destinationAddressbuffer[4][3] ), .B1(n672), .Y(n647) );
  AOI22X1TS U1203 ( .A0(\destinationAddressbuffer[3][3] ), .A1(n675), .B0(
        \destinationAddressbuffer[1][3] ), .B1(n674), .Y(n646) );
  AOI22X1TS U1204 ( .A0(\destinationAddressbuffer[7][3] ), .A1(n644), .B0(
        \destinationAddressbuffer[5][3] ), .B1(n676), .Y(n645) );
  NAND4XLTS U1205 ( .A(n648), .B(n647), .C(n646), .D(n645), .Y(n649) );
  AOI22X1TS U1206 ( .A0(destinationAddressOut[3]), .A1(n755), .B0(n1905), .B1(
        n649), .Y(n651) );
  AOI22X1TS U1207 ( .A0(destinationAddressIn_EAST[4]), .A1(n744), .B0(n654), 
        .B1(n665), .Y(n664) );
  AOI22X1TS U1208 ( .A0(destinationAddressIn_NORTH[4]), .A1(n669), .B0(n656), 
        .B1(n655), .Y(n663) );
  INVX2TS U1209 ( .A(n1906), .Y(n764) );
  CLKBUFX2TS U1210 ( .A(n764), .Y(n860) );
  AOI22X1TS U1211 ( .A0(\destinationAddressbuffer[2][4] ), .A1(n671), .B0(
        \destinationAddressbuffer[0][4] ), .B1(n670), .Y(n660) );
  AOI22X1TS U1212 ( .A0(\destinationAddressbuffer[6][4] ), .A1(n673), .B0(
        \destinationAddressbuffer[4][4] ), .B1(n672), .Y(n659) );
  AOI22X1TS U1213 ( .A0(\destinationAddressbuffer[3][4] ), .A1(n675), .B0(
        \destinationAddressbuffer[1][4] ), .B1(n674), .Y(n658) );
  CLKBUFX2TS U1214 ( .A(n748), .Y(n702) );
  AOI22X1TS U1215 ( .A0(\destinationAddressbuffer[7][4] ), .A1(n702), .B0(
        \destinationAddressbuffer[5][4] ), .B1(n676), .Y(n657) );
  NAND4XLTS U1216 ( .A(n660), .B(n659), .C(n658), .D(n657), .Y(n661) );
  AOI22X1TS U1217 ( .A0(destinationAddressOut[4]), .A1(n779), .B0(n860), .B1(
        n661), .Y(n662) );
  CLKBUFX2TS U1218 ( .A(n773), .Y(n760) );
  AOI22X1TS U1219 ( .A0(destinationAddressIn_EAST[5]), .A1(n760), .B0(n666), 
        .B1(n665), .Y(n685) );
  CLKBUFX2TS U1220 ( .A(n667), .Y(n745) );
  AOI22X1TS U1221 ( .A0(destinationAddressIn_NORTH[5]), .A1(n669), .B0(n668), 
        .B1(n745), .Y(n684) );
  AOI22X1TS U1222 ( .A0(\destinationAddressbuffer[2][5] ), .A1(n671), .B0(
        \destinationAddressbuffer[0][5] ), .B1(n670), .Y(n680) );
  AOI22X1TS U1223 ( .A0(\destinationAddressbuffer[6][5] ), .A1(n673), .B0(
        \destinationAddressbuffer[4][5] ), .B1(n672), .Y(n679) );
  AOI22X1TS U1224 ( .A0(\destinationAddressbuffer[3][5] ), .A1(n675), .B0(
        \destinationAddressbuffer[1][5] ), .B1(n674), .Y(n678) );
  AOI22X1TS U1225 ( .A0(\destinationAddressbuffer[7][5] ), .A1(n702), .B0(
        \destinationAddressbuffer[5][5] ), .B1(n676), .Y(n677) );
  NAND4XLTS U1226 ( .A(n680), .B(n679), .C(n678), .D(n677), .Y(n681) );
  AOI22X1TS U1227 ( .A0(destinationAddressOut[5]), .A1(n682), .B0(n860), .B1(
        n681), .Y(n683) );
  CLKBUFX2TS U1228 ( .A(n805), .Y(n725) );
  AOI22X1TS U1229 ( .A0(destinationAddressIn_EAST[6]), .A1(n760), .B0(n686), 
        .B1(n725), .Y(n699) );
  CLKBUFX2TS U1230 ( .A(n687), .Y(n804) );
  CLKBUFX2TS U1231 ( .A(n804), .Y(n728) );
  AOI22X1TS U1232 ( .A0(destinationAddressIn_NORTH[6]), .A1(n728), .B0(n688), 
        .B1(n745), .Y(n698) );
  CLKBUFX2TS U1233 ( .A(n689), .Y(n806) );
  CLKBUFX2TS U1234 ( .A(n806), .Y(n731) );
  AOI22X1TS U1235 ( .A0(\destinationAddressbuffer[2][6] ), .A1(n714), .B0(
        \destinationAddressbuffer[0][6] ), .B1(n731), .Y(n695) );
  CLKBUFX2TS U1236 ( .A(n690), .Y(n808) );
  CLKBUFX2TS U1237 ( .A(n808), .Y(n732) );
  AOI22X1TS U1238 ( .A0(\destinationAddressbuffer[6][6] ), .A1(n715), .B0(
        \destinationAddressbuffer[4][6] ), .B1(n732), .Y(n694) );
  CLKBUFX2TS U1239 ( .A(n691), .Y(n810) );
  CLKBUFX2TS U1240 ( .A(n810), .Y(n733) );
  AOI22X1TS U1241 ( .A0(\destinationAddressbuffer[3][6] ), .A1(n716), .B0(
        \destinationAddressbuffer[1][6] ), .B1(n733), .Y(n693) );
  CLKBUFX2TS U1242 ( .A(n854), .Y(n823) );
  CLKBUFX2TS U1243 ( .A(n823), .Y(n734) );
  AOI22X1TS U1244 ( .A0(\destinationAddressbuffer[7][6] ), .A1(n702), .B0(
        \destinationAddressbuffer[5][6] ), .B1(n734), .Y(n692) );
  NAND4XLTS U1245 ( .A(n695), .B(n694), .C(n693), .D(n692), .Y(n696) );
  AOI22X1TS U1246 ( .A0(destinationAddressOut[6]), .A1(n779), .B0(n860), .B1(
        n696), .Y(n697) );
  AOI22X1TS U1247 ( .A0(destinationAddressIn_EAST[7]), .A1(n822), .B0(n700), 
        .B1(n725), .Y(n710) );
  AOI22X1TS U1248 ( .A0(destinationAddressIn_NORTH[7]), .A1(n728), .B0(n701), 
        .B1(n761), .Y(n709) );
  CLKBUFX2TS U1249 ( .A(n764), .Y(n754) );
  AOI22X1TS U1250 ( .A0(\destinationAddressbuffer[2][7] ), .A1(n714), .B0(
        \destinationAddressbuffer[0][7] ), .B1(n731), .Y(n706) );
  AOI22X1TS U1251 ( .A0(\destinationAddressbuffer[6][7] ), .A1(n715), .B0(
        \destinationAddressbuffer[4][7] ), .B1(n732), .Y(n705) );
  AOI22X1TS U1252 ( .A0(\destinationAddressbuffer[3][7] ), .A1(n716), .B0(
        \destinationAddressbuffer[1][7] ), .B1(n733), .Y(n704) );
  AOI22X1TS U1253 ( .A0(\destinationAddressbuffer[7][7] ), .A1(n702), .B0(
        \destinationAddressbuffer[5][7] ), .B1(n734), .Y(n703) );
  NAND4XLTS U1254 ( .A(n706), .B(n705), .C(n704), .D(n703), .Y(n707) );
  AOI22X1TS U1255 ( .A0(destinationAddressOut[7]), .A1(n520), .B0(n754), .B1(
        n707), .Y(n708) );
  AOI22X1TS U1256 ( .A0(destinationAddressIn_EAST[8]), .A1(n744), .B0(n711), 
        .B1(n725), .Y(n724) );
  AOI22X1TS U1257 ( .A0(n713), .A1(n728), .B0(n712), .B1(n745), .Y(n723) );
  CLKBUFX2TS U1258 ( .A(n714), .Y(n807) );
  AOI22X1TS U1259 ( .A0(\destinationAddressbuffer[2][8] ), .A1(n807), .B0(
        \destinationAddressbuffer[0][8] ), .B1(n731), .Y(n720) );
  CLKBUFX2TS U1260 ( .A(n715), .Y(n809) );
  AOI22X1TS U1261 ( .A0(\destinationAddressbuffer[6][8] ), .A1(n809), .B0(
        \destinationAddressbuffer[4][8] ), .B1(n732), .Y(n719) );
  CLKBUFX2TS U1262 ( .A(n716), .Y(n811) );
  AOI22X1TS U1263 ( .A0(\destinationAddressbuffer[3][8] ), .A1(n811), .B0(
        \destinationAddressbuffer[1][8] ), .B1(n733), .Y(n718) );
  AOI22X1TS U1264 ( .A0(\destinationAddressbuffer[7][8] ), .A1(n812), .B0(
        \destinationAddressbuffer[5][8] ), .B1(n734), .Y(n717) );
  NAND4XLTS U1265 ( .A(n720), .B(n719), .C(n718), .D(n717), .Y(n721) );
  AOI22X1TS U1266 ( .A0(destinationAddressOut[8]), .A1(n755), .B0(n754), .B1(
        n721), .Y(n722) );
  AOI22X1TS U1267 ( .A0(destinationAddressIn_EAST[9]), .A1(n760), .B0(n726), 
        .B1(n725), .Y(n742) );
  AOI22X1TS U1268 ( .A0(n729), .A1(n728), .B0(n727), .B1(n761), .Y(n741) );
  INVX2TS U1269 ( .A(n730), .Y(n839) );
  AOI22X1TS U1270 ( .A0(\destinationAddressbuffer[2][9] ), .A1(n807), .B0(
        \destinationAddressbuffer[0][9] ), .B1(n731), .Y(n738) );
  AOI22X1TS U1271 ( .A0(\destinationAddressbuffer[6][9] ), .A1(n809), .B0(
        \destinationAddressbuffer[4][9] ), .B1(n732), .Y(n737) );
  AOI22X1TS U1272 ( .A0(\destinationAddressbuffer[3][9] ), .A1(n811), .B0(
        \destinationAddressbuffer[1][9] ), .B1(n733), .Y(n736) );
  AOI22X1TS U1273 ( .A0(\destinationAddressbuffer[7][9] ), .A1(n812), .B0(
        \destinationAddressbuffer[5][9] ), .B1(n734), .Y(n735) );
  NAND4XLTS U1274 ( .A(n738), .B(n737), .C(n736), .D(n735), .Y(n739) );
  AOI22X1TS U1275 ( .A0(destinationAddressOut[9]), .A1(n839), .B0(n754), .B1(
        n739), .Y(n740) );
  CLKBUFX2TS U1276 ( .A(n805), .Y(n784) );
  AOI22X1TS U1277 ( .A0(destinationAddressIn_EAST[10]), .A1(n744), .B0(n743), 
        .B1(n784), .Y(n758) );
  CLKBUFX2TS U1278 ( .A(n804), .Y(n785) );
  AOI22X1TS U1279 ( .A0(n747), .A1(n785), .B0(n746), .B1(n745), .Y(n757) );
  CLKBUFX2TS U1280 ( .A(n807), .Y(n786) );
  CLKBUFX2TS U1281 ( .A(n806), .Y(n787) );
  AOI22X1TS U1282 ( .A0(\destinationAddressbuffer[2][10] ), .A1(n786), .B0(
        \destinationAddressbuffer[0][10] ), .B1(n787), .Y(n752) );
  CLKBUFX2TS U1283 ( .A(n809), .Y(n788) );
  CLKBUFX2TS U1284 ( .A(n808), .Y(n789) );
  AOI22X1TS U1285 ( .A0(\destinationAddressbuffer[6][10] ), .A1(n788), .B0(
        \destinationAddressbuffer[4][10] ), .B1(n789), .Y(n751) );
  CLKBUFX2TS U1286 ( .A(n811), .Y(n790) );
  CLKBUFX2TS U1287 ( .A(n810), .Y(n791) );
  AOI22X1TS U1288 ( .A0(\destinationAddressbuffer[3][10] ), .A1(n790), .B0(
        \destinationAddressbuffer[1][10] ), .B1(n791), .Y(n750) );
  CLKBUFX2TS U1289 ( .A(n823), .Y(n793) );
  AOI22X1TS U1290 ( .A0(\destinationAddressbuffer[7][10] ), .A1(n748), .B0(
        \destinationAddressbuffer[5][10] ), .B1(n793), .Y(n749) );
  NAND4XLTS U1291 ( .A(n752), .B(n751), .C(n750), .D(n749), .Y(n753) );
  AOI22X1TS U1292 ( .A0(destinationAddressOut[10]), .A1(n755), .B0(n754), .B1(
        n753), .Y(n756) );
  AOI22X1TS U1293 ( .A0(destinationAddressIn_EAST[11]), .A1(n760), .B0(n759), 
        .B1(n784), .Y(n772) );
  AOI22X1TS U1294 ( .A0(n763), .A1(n785), .B0(n762), .B1(n761), .Y(n771) );
  CLKBUFX2TS U1295 ( .A(n764), .Y(n818) );
  AOI22X1TS U1296 ( .A0(\destinationAddressbuffer[2][11] ), .A1(n786), .B0(
        \destinationAddressbuffer[0][11] ), .B1(n787), .Y(n768) );
  AOI22X1TS U1297 ( .A0(\destinationAddressbuffer[6][11] ), .A1(n788), .B0(
        \destinationAddressbuffer[4][11] ), .B1(n789), .Y(n767) );
  AOI22X1TS U1298 ( .A0(\destinationAddressbuffer[3][11] ), .A1(n790), .B0(
        \destinationAddressbuffer[1][11] ), .B1(n791), .Y(n766) );
  AOI22X1TS U1299 ( .A0(\destinationAddressbuffer[7][11] ), .A1(n792), .B0(
        \destinationAddressbuffer[5][11] ), .B1(n793), .Y(n765) );
  NAND4XLTS U1300 ( .A(n768), .B(n767), .C(n766), .D(n765), .Y(n769) );
  AOI22X1TS U1301 ( .A0(destinationAddressOut[11]), .A1(n520), .B0(n818), .B1(
        n769), .Y(n770) );
  CLKBUFX2TS U1302 ( .A(dataIn_SOUTH[0]), .Y(n1497) );
  CLKBUFX2TS U1303 ( .A(dataIn_EAST[0]), .Y(n1456) );
  CLKBUFX2TS U1304 ( .A(n1456), .Y(n1103) );
  CLKBUFX2TS U1305 ( .A(n773), .Y(n843) );
  AOI22X1TS U1306 ( .A0(n1497), .A1(n783), .B0(n1103), .B1(n843), .Y(n782) );
  CLKBUFX2TS U1307 ( .A(dataIn_WEST[0]), .Y(n1362) );
  AOI22X1TS U1308 ( .A0(dataIn_NORTH[0]), .A1(n785), .B0(n1362), .B1(n784), 
        .Y(n781) );
  AOI22X1TS U1309 ( .A0(\dataoutbuffer[0][0] ), .A1(n787), .B0(
        \dataoutbuffer[2][0] ), .B1(n786), .Y(n777) );
  AOI22X1TS U1310 ( .A0(\dataoutbuffer[4][0] ), .A1(n789), .B0(
        \dataoutbuffer[6][0] ), .B1(n788), .Y(n776) );
  AOI22X1TS U1311 ( .A0(\dataoutbuffer[1][0] ), .A1(n791), .B0(
        \dataoutbuffer[3][0] ), .B1(n790), .Y(n775) );
  AOI22X1TS U1312 ( .A0(\dataoutbuffer[5][0] ), .A1(n793), .B0(
        \dataoutbuffer[7][0] ), .B1(n853), .Y(n774) );
  NAND4XLTS U1313 ( .A(n777), .B(n776), .C(n775), .D(n774), .Y(n778) );
  AOI22X1TS U1314 ( .A0(dataOut[0]), .A1(n779), .B0(n818), .B1(n778), .Y(n780)
         );
  CLKBUFX2TS U1315 ( .A(dataIn_SOUTH[1]), .Y(n1505) );
  CLKBUFX2TS U1316 ( .A(dataIn_EAST[1]), .Y(n1464) );
  CLKBUFX2TS U1317 ( .A(n1464), .Y(n1110) );
  AOI22X1TS U1318 ( .A0(n1505), .A1(n783), .B0(n1110), .B1(n822), .Y(n802) );
  CLKBUFX2TS U1319 ( .A(dataIn_WEST[1]), .Y(n1367) );
  AOI22X1TS U1320 ( .A0(dataIn_NORTH[1]), .A1(n785), .B0(n1367), .B1(n784), 
        .Y(n801) );
  AOI22X1TS U1321 ( .A0(\dataoutbuffer[0][1] ), .A1(n787), .B0(
        \dataoutbuffer[2][1] ), .B1(n786), .Y(n797) );
  AOI22X1TS U1322 ( .A0(\dataoutbuffer[4][1] ), .A1(n789), .B0(
        \dataoutbuffer[6][1] ), .B1(n788), .Y(n796) );
  AOI22X1TS U1323 ( .A0(\dataoutbuffer[1][1] ), .A1(n791), .B0(
        \dataoutbuffer[3][1] ), .B1(n790), .Y(n795) );
  AOI22X1TS U1324 ( .A0(\dataoutbuffer[5][1] ), .A1(n793), .B0(
        \dataoutbuffer[7][1] ), .B1(n792), .Y(n794) );
  NAND4XLTS U1325 ( .A(n797), .B(n796), .C(n795), .D(n794), .Y(n798) );
  AOI22X1TS U1326 ( .A0(dataOut[1]), .A1(n521), .B0(n818), .B1(n798), .Y(n800)
         );
  CLKBUFX2TS U1327 ( .A(dataIn_SOUTH[2]), .Y(n1512) );
  CLKBUFX2TS U1328 ( .A(dataIn_EAST[2]), .Y(n1470) );
  CLKBUFX2TS U1329 ( .A(n1470), .Y(n1340) );
  AOI22X1TS U1330 ( .A0(n1512), .A1(n803), .B0(n1340), .B1(n843), .Y(n821) );
  CLKBUFX2TS U1331 ( .A(n804), .Y(n846) );
  CLKBUFX2TS U1332 ( .A(dataIn_WEST[2]), .Y(n1371) );
  CLKBUFX2TS U1333 ( .A(n805), .Y(n845) );
  AOI22X1TS U1334 ( .A0(dataIn_NORTH[2]), .A1(n846), .B0(n1371), .B1(n845), 
        .Y(n820) );
  CLKBUFX2TS U1335 ( .A(n806), .Y(n848) );
  CLKBUFX2TS U1336 ( .A(n807), .Y(n847) );
  AOI22X1TS U1337 ( .A0(\dataoutbuffer[0][2] ), .A1(n848), .B0(
        \dataoutbuffer[2][2] ), .B1(n847), .Y(n816) );
  CLKBUFX2TS U1338 ( .A(n808), .Y(n850) );
  CLKBUFX2TS U1339 ( .A(n809), .Y(n849) );
  AOI22X1TS U1340 ( .A0(\dataoutbuffer[4][2] ), .A1(n850), .B0(
        \dataoutbuffer[6][2] ), .B1(n849), .Y(n815) );
  CLKBUFX2TS U1341 ( .A(n810), .Y(n852) );
  CLKBUFX2TS U1342 ( .A(n811), .Y(n851) );
  AOI22X1TS U1343 ( .A0(\dataoutbuffer[1][2] ), .A1(n852), .B0(
        \dataoutbuffer[3][2] ), .B1(n851), .Y(n814) );
  AOI22X1TS U1344 ( .A0(\dataoutbuffer[5][2] ), .A1(n823), .B0(
        \dataoutbuffer[7][2] ), .B1(n812), .Y(n813) );
  NAND4XLTS U1345 ( .A(n816), .B(n815), .C(n814), .D(n813), .Y(n817) );
  AOI22X1TS U1346 ( .A0(dataOut[2]), .A1(n839), .B0(n818), .B1(n817), .Y(n819)
         );
  INVX2TS U1347 ( .A(n12), .Y(n861) );
  CLKBUFX2TS U1348 ( .A(dataIn_SOUTH[3]), .Y(n1521) );
  CLKBUFX2TS U1349 ( .A(dataIn_EAST[3]), .Y(n1476) );
  CLKBUFX2TS U1350 ( .A(n1476), .Y(n1345) );
  AOI22X1TS U1351 ( .A0(n1521), .A1(n844), .B0(n1345), .B1(n822), .Y(n831) );
  CLKBUFX2TS U1352 ( .A(dataIn_WEST[3]), .Y(n1377) );
  AOI22X1TS U1353 ( .A0(dataIn_NORTH[3]), .A1(n846), .B0(n1377), .B1(n845), 
        .Y(n830) );
  AOI22X1TS U1354 ( .A0(\dataoutbuffer[0][3] ), .A1(n848), .B0(
        \dataoutbuffer[2][3] ), .B1(n847), .Y(n827) );
  AOI22X1TS U1355 ( .A0(\dataoutbuffer[4][3] ), .A1(n850), .B0(
        \dataoutbuffer[6][3] ), .B1(n849), .Y(n826) );
  AOI22X1TS U1356 ( .A0(\dataoutbuffer[1][3] ), .A1(n852), .B0(
        \dataoutbuffer[3][3] ), .B1(n851), .Y(n825) );
  AOI22X1TS U1357 ( .A0(\dataoutbuffer[5][3] ), .A1(n823), .B0(
        \dataoutbuffer[7][3] ), .B1(n832), .Y(n824) );
  NAND4XLTS U1358 ( .A(n827), .B(n826), .C(n825), .D(n824), .Y(n828) );
  AOI22X1TS U1359 ( .A0(dataOut[3]), .A1(n839), .B0(n838), .B1(n828), .Y(n829)
         );
  CLKBUFX2TS U1360 ( .A(dataIn_SOUTH[4]), .Y(n1528) );
  CLKBUFX2TS U1361 ( .A(dataIn_EAST[4]), .Y(n1481) );
  CLKBUFX2TS U1362 ( .A(n1481), .Y(n1350) );
  AOI22X1TS U1363 ( .A0(n1528), .A1(n844), .B0(n1350), .B1(n843), .Y(n842) );
  CLKBUFX2TS U1364 ( .A(dataIn_WEST[4]), .Y(n1382) );
  AOI22X1TS U1365 ( .A0(dataIn_NORTH[4]), .A1(n846), .B0(n1382), .B1(n845), 
        .Y(n841) );
  AOI22X1TS U1366 ( .A0(\dataoutbuffer[0][4] ), .A1(n848), .B0(
        \dataoutbuffer[2][4] ), .B1(n847), .Y(n836) );
  AOI22X1TS U1367 ( .A0(\dataoutbuffer[4][4] ), .A1(n850), .B0(
        \dataoutbuffer[6][4] ), .B1(n849), .Y(n835) );
  AOI22X1TS U1368 ( .A0(\dataoutbuffer[1][4] ), .A1(n852), .B0(
        \dataoutbuffer[3][4] ), .B1(n851), .Y(n834) );
  AOI22X1TS U1369 ( .A0(\dataoutbuffer[5][4] ), .A1(n854), .B0(
        \dataoutbuffer[7][4] ), .B1(n832), .Y(n833) );
  NAND4XLTS U1370 ( .A(n836), .B(n835), .C(n834), .D(n833), .Y(n837) );
  AOI22X1TS U1371 ( .A0(dataOut[4]), .A1(n839), .B0(n838), .B1(n837), .Y(n840)
         );
  CLKBUFX2TS U1372 ( .A(dataIn_SOUTH[5]), .Y(n1536) );
  CLKBUFX2TS U1373 ( .A(dataIn_EAST[5]), .Y(n1489) );
  CLKBUFX2TS U1374 ( .A(n1489), .Y(n1356) );
  AOI22X1TS U1375 ( .A0(n1536), .A1(n844), .B0(n1356), .B1(n843), .Y(n864) );
  CLKBUFX2TS U1376 ( .A(dataIn_WEST[5]), .Y(n1388) );
  AOI22X1TS U1377 ( .A0(dataIn_NORTH[5]), .A1(n846), .B0(n1388), .B1(n845), 
        .Y(n863) );
  AOI22X1TS U1378 ( .A0(\dataoutbuffer[0][5] ), .A1(n848), .B0(
        \dataoutbuffer[2][5] ), .B1(n847), .Y(n858) );
  AOI22X1TS U1379 ( .A0(\dataoutbuffer[4][5] ), .A1(n850), .B0(
        \dataoutbuffer[6][5] ), .B1(n849), .Y(n857) );
  AOI22X1TS U1380 ( .A0(\dataoutbuffer[1][5] ), .A1(n852), .B0(
        \dataoutbuffer[3][5] ), .B1(n851), .Y(n856) );
  AOI22X1TS U1381 ( .A0(\dataoutbuffer[5][5] ), .A1(n854), .B0(
        \dataoutbuffer[7][5] ), .B1(n853), .Y(n855) );
  NAND4XLTS U1382 ( .A(n858), .B(n857), .C(n856), .D(n855), .Y(n859) );
  AOI22X1TS U1383 ( .A0(dataOut[5]), .A1(n521), .B0(n860), .B1(n859), .Y(n862)
         );
  INVX2TS U1384 ( .A(n944), .Y(n1754) );
  INVX2TS U1385 ( .A(n1501), .Y(n1525) );
  AOI22X1TS U1386 ( .A0(n1754), .A1(n1525), .B0(n1652), .B1(
        \requesterAddressbuffer[7][0] ), .Y(n867) );
  INVX2TS U1387 ( .A(n1509), .Y(n1638) );
  AOI22X1TS U1388 ( .A0(n32), .A1(n946), .B0(n1638), .B1(
        requesterAddressIn_EAST[0]), .Y(n866) );
  CLKBUFX2TS U1389 ( .A(n1020), .Y(n920) );
  AOI22X1TS U1390 ( .A0(n868), .A1(n920), .B0(n1535), .B1(n990), .Y(n865) );
  INVX2TS U1391 ( .A(n1501), .Y(n1645) );
  INVX2TS U1392 ( .A(n1494), .Y(n1532) );
  AOI22X1TS U1393 ( .A0(n1645), .A1(n1636), .B0(n1532), .B1(
        \requesterAddressbuffer[7][1] ), .Y(n871) );
  AOI22X1TS U1394 ( .A0(n1656), .A1(n952), .B0(n872), .B1(
        requesterAddressIn_EAST[1]), .Y(n870) );
  CLKBUFX2TS U1395 ( .A(n1027), .Y(n925) );
  AOI22X1TS U1396 ( .A0(n868), .A1(n925), .B0(n50), .B1(n997), .Y(n869) );
  AOI22X1TS U1397 ( .A0(n1654), .A1(n1644), .B0(n1532), .B1(
        \requesterAddressbuffer[7][2] ), .Y(n876) );
  AOI22X1TS U1398 ( .A0(n1519), .A1(n957), .B0(n872), .B1(
        requesterAddressIn_EAST[2]), .Y(n875) );
  INVX2TS U1399 ( .A(n873), .Y(n1513) );
  CLKBUFX2TS U1400 ( .A(n1033), .Y(n930) );
  AOI22X1TS U1401 ( .A0(n1513), .A1(n930), .B0(n1535), .B1(n1003), .Y(n874) );
  INVX2TS U1402 ( .A(n877), .Y(n1643) );
  AOI22X1TS U1403 ( .A0(n1525), .A1(n1653), .B0(n1643), .B1(
        \requesterAddressbuffer[7][3] ), .Y(n881) );
  INVX2TS U1404 ( .A(n1509), .Y(n1655) );
  AOI22X1TS U1405 ( .A0(n1646), .A1(n965), .B0(n1655), .B1(
        requesterAddressIn_EAST[3]), .Y(n880) );
  CLKBUFX2TS U1406 ( .A(n1043), .Y(n940) );
  INVX2TS U1407 ( .A(n878), .Y(n1632) );
  AOI22X1TS U1408 ( .A0(n1513), .A1(n940), .B0(n1632), .B1(n1012), .Y(n879) );
  INVX2TS U1409 ( .A(n944), .Y(n1806) );
  AOI22X1TS U1410 ( .A0(n1806), .A1(n1661), .B0(n1682), .B1(
        \requesterAddressbuffer[6][0] ), .Y(n884) );
  INVX2TS U1411 ( .A(n1469), .Y(n1669) );
  AOI22X1TS U1412 ( .A0(n918), .A1(n1683), .B0(n1017), .B1(n1669), .Y(n883) );
  AOI22X1TS U1413 ( .A0(n920), .A1(n1459), .B0(n990), .B1(n1460), .Y(n882) );
  INVX2TS U1414 ( .A(n950), .Y(n1729) );
  INVX2TS U1415 ( .A(n893), .Y(n1668) );
  INVX2TS U1416 ( .A(n1455), .Y(n1488) );
  AOI22X1TS U1417 ( .A0(n1729), .A1(n1668), .B0(n1488), .B1(
        \requesterAddressbuffer[6][1] ), .Y(n888) );
  INVX2TS U1418 ( .A(n1469), .Y(n1676) );
  AOI22X1TS U1419 ( .A0(n924), .A1(n1482), .B0(n1025), .B1(n1676), .Y(n887) );
  INVX2TS U1420 ( .A(n102), .Y(n1484) );
  AOI22X1TS U1421 ( .A0(n925), .A1(n1484), .B0(n997), .B1(n103), .Y(n886) );
  INVX2TS U1422 ( .A(n956), .Y(n1736) );
  INVX2TS U1423 ( .A(n893), .Y(n1675) );
  AOI22X1TS U1424 ( .A0(n1736), .A1(n1675), .B0(n1488), .B1(
        \requesterAddressbuffer[6][2] ), .Y(n892) );
  AOI22X1TS U1425 ( .A0(n929), .A1(n1457), .B0(n1031), .B1(n896), .Y(n891) );
  AOI22X1TS U1426 ( .A0(n930), .A1(n96), .B0(n1003), .B1(n889), .Y(n890) );
  INVX2TS U1427 ( .A(n963), .Y(n1745) );
  INVX2TS U1428 ( .A(n894), .Y(n1674) );
  AOI22X1TS U1429 ( .A0(n1745), .A1(n1661), .B0(n1674), .B1(
        \requesterAddressbuffer[6][3] ), .Y(n900) );
  INVX2TS U1430 ( .A(n895), .Y(n1482) );
  AOI22X1TS U1431 ( .A0(n938), .A1(n1482), .B0(n1040), .B1(n896), .Y(n899) );
  INVX2TS U1432 ( .A(n897), .Y(n1678) );
  AOI22X1TS U1433 ( .A0(n940), .A1(n1678), .B0(n1012), .B1(n1664), .Y(n898) );
  AOI22X1TS U1434 ( .A0(n987), .A1(n1690), .B0(n1712), .B1(
        \requesterAddressbuffer[5][0] ), .Y(n904) );
  INVX2TS U1435 ( .A(n1432), .Y(n1700) );
  AOI22X1TS U1436 ( .A0(n918), .A1(n1715), .B0(n1017), .B1(n1700), .Y(n903) );
  INVX2TS U1437 ( .A(n901), .Y(n1716) );
  AOI22X1TS U1438 ( .A0(n920), .A1(n1716), .B0(requesterAddressIn_NORTH[0]), 
        .B1(n1434), .Y(n902) );
  INVX2TS U1439 ( .A(n10), .Y(n1698) );
  AOI22X1TS U1440 ( .A0(n1636), .A1(n1698), .B0(n1450), .B1(
        \requesterAddressbuffer[5][1] ), .Y(n907) );
  INVX2TS U1441 ( .A(n1432), .Y(n1708) );
  AOI22X1TS U1442 ( .A0(n924), .A1(n1443), .B0(n1025), .B1(n1708), .Y(n906) );
  AOI22X1TS U1443 ( .A0(n925), .A1(n1693), .B0(requesterAddressIn_NORTH[1]), 
        .B1(n1694), .Y(n905) );
  INVX2TS U1444 ( .A(n10), .Y(n1706) );
  AOI22X1TS U1445 ( .A0(n1644), .A1(n1706), .B0(n1450), .B1(
        \requesterAddressbuffer[5][2] ), .Y(n911) );
  AOI22X1TS U1446 ( .A0(n929), .A1(n1421), .B0(n1031), .B1(n914), .Y(n910) );
  AOI22X1TS U1447 ( .A0(n930), .A1(n1422), .B0(requesterAddressIn_NORTH[2]), 
        .B1(n908), .Y(n909) );
  INVX2TS U1448 ( .A(n10), .Y(n1713) );
  INVX2TS U1449 ( .A(n912), .Y(n1705) );
  AOI22X1TS U1450 ( .A0(n1653), .A1(n1713), .B0(n1705), .B1(
        \requesterAddressbuffer[5][3] ), .Y(n917) );
  INVX2TS U1451 ( .A(n913), .Y(n1443) );
  AOI22X1TS U1452 ( .A0(n938), .A1(n1443), .B0(n1040), .B1(n914), .Y(n916) );
  AOI22X1TS U1453 ( .A0(n940), .A1(n230), .B0(requesterAddressIn_NORTH[3]), 
        .B1(n1446), .Y(n915) );
  AOI22X1TS U1454 ( .A0(n987), .A1(n1720), .B0(n1743), .B1(
        \requesterAddressbuffer[4][0] ), .Y(n923) );
  INVX2TS U1455 ( .A(n1402), .Y(n1730) );
  AOI22X1TS U1456 ( .A0(n918), .A1(n1747), .B0(requesterAddressIn_EAST[0]), 
        .B1(n1730), .Y(n922) );
  INVX2TS U1457 ( .A(n919), .Y(n1411) );
  AOI22X1TS U1458 ( .A0(n920), .A1(n1739), .B0(requesterAddressIn_NORTH[0]), 
        .B1(n1411), .Y(n921) );
  INVX2TS U1459 ( .A(n950), .Y(n1858) );
  INVX2TS U1460 ( .A(n934), .Y(n1728) );
  INVX2TS U1461 ( .A(n1393), .Y(n1416) );
  AOI22X1TS U1462 ( .A0(n1858), .A1(n1728), .B0(n1416), .B1(
        \requesterAddressbuffer[4][1] ), .Y(n928) );
  INVX2TS U1463 ( .A(n1402), .Y(n1737) );
  AOI22X1TS U1464 ( .A0(n924), .A1(n1410), .B0(requesterAddressIn_EAST[1]), 
        .B1(n1737), .Y(n927) );
  AOI22X1TS U1465 ( .A0(n925), .A1(n1412), .B0(requesterAddressIn_NORTH[1]), 
        .B1(n1748), .Y(n926) );
  INVX2TS U1466 ( .A(n956), .Y(n1868) );
  AOI22X1TS U1467 ( .A0(n1868), .A1(n1720), .B0(n1416), .B1(
        \requesterAddressbuffer[4][2] ), .Y(n933) );
  AOI22X1TS U1468 ( .A0(n929), .A1(n1394), .B0(requesterAddressIn_EAST[2]), 
        .B1(n937), .Y(n932) );
  AOI22X1TS U1469 ( .A0(n930), .A1(n1749), .B0(requesterAddressIn_NORTH[2]), 
        .B1(n1748), .Y(n931) );
  INVX2TS U1470 ( .A(n963), .Y(n1879) );
  INVX2TS U1471 ( .A(n934), .Y(n1744) );
  INVX2TS U1472 ( .A(n935), .Y(n1735) );
  AOI22X1TS U1473 ( .A0(n1879), .A1(n1744), .B0(n1735), .B1(
        \requesterAddressbuffer[4][3] ), .Y(n943) );
  INVX2TS U1474 ( .A(n936), .Y(n1410) );
  AOI22X1TS U1475 ( .A0(n938), .A1(n1410), .B0(requesterAddressIn_EAST[3]), 
        .B1(n937), .Y(n942) );
  INVX2TS U1476 ( .A(n939), .Y(n1724) );
  AOI22X1TS U1477 ( .A0(n940), .A1(n1724), .B0(requesterAddressIn_NORTH[3]), 
        .B1(n1395), .Y(n941) );
  INVX2TS U1478 ( .A(n944), .Y(n1847) );
  AOI22X1TS U1479 ( .A0(n1847), .A1(n1753), .B0(n1772), .B1(
        \requesterAddressbuffer[3][0] ), .Y(n949) );
  INVX2TS U1480 ( .A(n945), .Y(n1372) );
  AOI22X1TS U1481 ( .A0(n946), .A1(n1372), .B0(n988), .B1(n151), .Y(n948) );
  INVX2TS U1482 ( .A(n958), .Y(n1768) );
  AOI22X1TS U1483 ( .A0(n991), .A1(n1768), .B0(n1019), .B1(n1363), .Y(n947) );
  INVX2TS U1484 ( .A(n950), .Y(n1817) );
  INVX2TS U1485 ( .A(n964), .Y(n1760) );
  INVX2TS U1486 ( .A(n1361), .Y(n1387) );
  AOI22X1TS U1487 ( .A0(n1817), .A1(n1760), .B0(n1387), .B1(
        \requesterAddressbuffer[3][1] ), .Y(n955) );
  INVX2TS U1488 ( .A(n951), .Y(n1761) );
  AOI22X1TS U1489 ( .A0(n952), .A1(n137), .B0(n996), .B1(n1761), .Y(n954) );
  INVX2TS U1490 ( .A(n958), .Y(n1776) );
  AOI22X1TS U1491 ( .A0(n998), .A1(n1776), .B0(n1026), .B1(n959), .Y(n953) );
  INVX2TS U1492 ( .A(n956), .Y(n1827) );
  AOI22X1TS U1493 ( .A0(n1827), .A1(n1753), .B0(n1387), .B1(
        \requesterAddressbuffer[3][2] ), .Y(n962) );
  AOI22X1TS U1494 ( .A0(n957), .A1(n1389), .B0(n1002), .B1(n1381), .Y(n961) );
  AOI22X1TS U1495 ( .A0(n1004), .A1(n130), .B0(n1032), .B1(n959), .Y(n960) );
  INVX2TS U1496 ( .A(n963), .Y(n1837) );
  INVX2TS U1497 ( .A(n964), .Y(n1773) );
  INVX2TS U1498 ( .A(n1361), .Y(n1766) );
  AOI22X1TS U1499 ( .A0(n1837), .A1(n1773), .B0(n1766), .B1(
        \requesterAddressbuffer[3][3] ), .Y(n968) );
  AOI22X1TS U1500 ( .A0(n965), .A1(n1372), .B0(n1010), .B1(n1774), .Y(n967) );
  AOI22X1TS U1501 ( .A0(n1013), .A1(n1768), .B0(n1042), .B1(n1756), .Y(n966)
         );
  AOI22X1TS U1502 ( .A0(n1754), .A1(n1781), .B0(n1799), .B1(
        \requesterAddressbuffer[2][0] ), .Y(n972) );
  INVX2TS U1503 ( .A(n1339), .Y(n1788) );
  AOI22X1TS U1504 ( .A0(requesterAddressIn_WEST[0]), .A1(n1801), .B0(n988), 
        .B1(n1788), .Y(n971) );
  INVX2TS U1505 ( .A(n969), .Y(n1795) );
  AOI22X1TS U1506 ( .A0(n991), .A1(n1795), .B0(n1019), .B1(n1106), .Y(n970) );
  INVX2TS U1507 ( .A(n981), .Y(n1787) );
  INVX2TS U1508 ( .A(n973), .Y(n1355) );
  AOI22X1TS U1509 ( .A0(n1858), .A1(n1787), .B0(n1355), .B1(
        \requesterAddressbuffer[2][1] ), .Y(n976) );
  INVX2TS U1510 ( .A(n1339), .Y(n1794) );
  AOI22X1TS U1511 ( .A0(requesterAddressIn_WEST[1]), .A1(n1351), .B0(n996), 
        .B1(n1794), .Y(n975) );
  AOI22X1TS U1512 ( .A0(n998), .A1(n191), .B0(n1026), .B1(n1789), .Y(n974) );
  AOI22X1TS U1513 ( .A0(n1868), .A1(n1781), .B0(n1355), .B1(
        \requesterAddressbuffer[2][2] ), .Y(n980) );
  AOI22X1TS U1514 ( .A0(requesterAddressIn_WEST[2]), .A1(n1104), .B0(n1002), 
        .B1(n983), .Y(n979) );
  AOI22X1TS U1515 ( .A0(n1004), .A1(n1105), .B0(n1032), .B1(n977), .Y(n978) );
  INVX2TS U1516 ( .A(n981), .Y(n1800) );
  INVX2TS U1517 ( .A(n1602), .Y(n1793) );
  AOI22X1TS U1518 ( .A0(n1879), .A1(n1800), .B0(n1793), .B1(
        \requesterAddressbuffer[2][3] ), .Y(n986) );
  INVX2TS U1519 ( .A(n982), .Y(n1351) );
  AOI22X1TS U1520 ( .A0(requesterAddressIn_WEST[3]), .A1(n1351), .B0(n1010), 
        .B1(n983), .Y(n985) );
  AOI22X1TS U1521 ( .A0(n1013), .A1(n1346), .B0(n1042), .B1(n1783), .Y(n984)
         );
  INVX2TS U1522 ( .A(n1078), .Y(n1092) );
  AOI22X1TS U1523 ( .A0(n987), .A1(n1092), .B0(n1835), .B1(
        \requesterAddressbuffer[1][0] ), .Y(n994) );
  INVX2TS U1524 ( .A(n1083), .Y(n1819) );
  AOI22X1TS U1525 ( .A0(requesterAddressIn_WEST[0]), .A1(n1839), .B0(n988), 
        .B1(n1819), .Y(n993) );
  INVX2TS U1526 ( .A(n989), .Y(n1841) );
  AOI22X1TS U1527 ( .A0(n991), .A1(n1841), .B0(n990), .B1(n1812), .Y(n992) );
  INVX2TS U1528 ( .A(n1078), .Y(n1826) );
  INVX2TS U1529 ( .A(n995), .Y(n1099) );
  AOI22X1TS U1530 ( .A0(n1729), .A1(n1826), .B0(n1099), .B1(
        \requesterAddressbuffer[1][1] ), .Y(n1001) );
  INVX2TS U1531 ( .A(n1083), .Y(n1829) );
  AOI22X1TS U1532 ( .A0(requesterAddressIn_WEST[1]), .A1(n1093), .B0(n996), 
        .B1(n1829), .Y(n1000) );
  AOI22X1TS U1533 ( .A0(n998), .A1(n1810), .B0(n997), .B1(n1084), .Y(n999) );
  AOI22X1TS U1534 ( .A0(n1736), .A1(n1836), .B0(n1099), .B1(
        \requesterAddressbuffer[1][2] ), .Y(n1007) );
  AOI22X1TS U1535 ( .A0(requesterAddressIn_WEST[2]), .A1(n1073), .B0(n1002), 
        .B1(n1009), .Y(n1006) );
  AOI22X1TS U1536 ( .A0(n1004), .A1(n1074), .B0(n1003), .B1(n322), .Y(n1005)
         );
  INVX2TS U1537 ( .A(n1616), .Y(n1825) );
  AOI22X1TS U1538 ( .A0(n1745), .A1(n1092), .B0(n1825), .B1(
        \requesterAddressbuffer[1][3] ), .Y(n1016) );
  INVX2TS U1539 ( .A(n1008), .Y(n1093) );
  AOI22X1TS U1540 ( .A0(requesterAddressIn_WEST[3]), .A1(n1093), .B0(n1010), 
        .B1(n1009), .Y(n1015) );
  AOI22X1TS U1541 ( .A0(n1013), .A1(n324), .B0(n1012), .B1(n1011), .Y(n1014)
         );
  AOI22X1TS U1542 ( .A0(readRequesterAddress[0]), .A1(n1846), .B0(n1877), .B1(
        \requesterAddressbuffer[0][0] ), .Y(n1023) );
  INVX2TS U1543 ( .A(n1055), .Y(n1859) );
  AOI22X1TS U1544 ( .A0(requesterAddressIn_WEST[0]), .A1(n1881), .B0(n1017), 
        .B1(n1859), .Y(n1022) );
  INVX2TS U1545 ( .A(n1018), .Y(n1064) );
  AOI22X1TS U1546 ( .A0(n1020), .A1(n1873), .B0(n1019), .B1(n1064), .Y(n1021)
         );
  INVX2TS U1547 ( .A(n11), .Y(n1857) );
  INVX2TS U1548 ( .A(n1024), .Y(n1069) );
  AOI22X1TS U1549 ( .A0(n1817), .A1(n1857), .B0(n1069), .B1(
        \requesterAddressbuffer[0][1] ), .Y(n1030) );
  INVX2TS U1550 ( .A(n1055), .Y(n1869) );
  AOI22X1TS U1551 ( .A0(requesterAddressIn_WEST[1]), .A1(n1063), .B0(n1025), 
        .B1(n1869), .Y(n1029) );
  AOI22X1TS U1552 ( .A0(n1027), .A1(n1065), .B0(n1026), .B1(n1064), .Y(n1028)
         );
  INVX2TS U1553 ( .A(n11), .Y(n1867) );
  AOI22X1TS U1554 ( .A0(n1827), .A1(n1867), .B0(n1069), .B1(
        \requesterAddressbuffer[0][2] ), .Y(n1036) );
  AOI22X1TS U1555 ( .A0(requesterAddressIn_WEST[2]), .A1(n1047), .B0(n1031), 
        .B1(n1039), .Y(n1035) );
  AOI22X1TS U1556 ( .A0(n1033), .A1(n1885), .B0(n1032), .B1(n1883), .Y(n1034)
         );
  INVX2TS U1557 ( .A(n11), .Y(n1878) );
  INVX2TS U1558 ( .A(n1037), .Y(n1866) );
  AOI22X1TS U1559 ( .A0(n1837), .A1(n1878), .B0(n1866), .B1(
        \requesterAddressbuffer[0][3] ), .Y(n1046) );
  INVX2TS U1560 ( .A(n1038), .Y(n1063) );
  AOI22X1TS U1561 ( .A0(requesterAddressIn_WEST[3]), .A1(n1063), .B0(n1040), 
        .B1(n1039), .Y(n1045) );
  INVX2TS U1562 ( .A(n1041), .Y(n1853) );
  AOI22X1TS U1563 ( .A0(n1043), .A1(n1853), .B0(n1042), .B1(n1048), .Y(n1044)
         );
  INVX2TS U1564 ( .A(n1037), .Y(n1059) );
  AOI21X1TS U1565 ( .A0(n1059), .A1(\dataoutbuffer[0][0] ), .B0(n1857), .Y(
        n1051) );
  AOI22X1TS U1566 ( .A0(n1047), .A1(dataIn_WEST[0]), .B0(n1859), .B1(n1103), 
        .Y(n1050) );
  AOI22X1TS U1567 ( .A0(n1853), .A1(n1497), .B0(n1048), .B1(dataIn_NORTH[0]), 
        .Y(n1049) );
  AOI21X1TS U1568 ( .A0(n1059), .A1(\dataoutbuffer[0][1] ), .B0(n1867), .Y(
        n1054) );
  AOI22X1TS U1569 ( .A0(n411), .A1(dataIn_WEST[1]), .B0(n1869), .B1(n1110), 
        .Y(n1053) );
  AOI22X1TS U1570 ( .A0(n1873), .A1(n1505), .B0(n396), .B1(dataIn_NORTH[1]), 
        .Y(n1052) );
  AOI21X1TS U1571 ( .A0(n1059), .A1(\dataoutbuffer[0][2] ), .B0(n1878), .Y(
        n1058) );
  AOI22X1TS U1572 ( .A0(n1063), .A1(dataIn_WEST[2]), .B0(n389), .B1(n1340), 
        .Y(n1057) );
  AOI22X1TS U1573 ( .A0(n1885), .A1(n1512), .B0(n1064), .B1(dataIn_NORTH[2]), 
        .Y(n1056) );
  AOI21X1TS U1574 ( .A0(n1059), .A1(\dataoutbuffer[0][3] ), .B0(n1857), .Y(
        n1062) );
  AOI22X1TS U1575 ( .A0(n1849), .A1(dataIn_WEST[3]), .B0(n1859), .B1(n1345), 
        .Y(n1061) );
  AOI22X1TS U1576 ( .A0(n430), .A1(n1521), .B0(n1851), .B1(dataIn_NORTH[3]), 
        .Y(n1060) );
  AOI21X1TS U1577 ( .A0(n1069), .A1(\dataoutbuffer[0][4] ), .B0(n1867), .Y(
        n1068) );
  AOI22X1TS U1578 ( .A0(n1063), .A1(dataIn_WEST[4]), .B0(n1869), .B1(n1350), 
        .Y(n1067) );
  AOI22X1TS U1579 ( .A0(n1065), .A1(n1528), .B0(n1064), .B1(dataIn_NORTH[4]), 
        .Y(n1066) );
  AOI21X1TS U1580 ( .A0(n1069), .A1(\dataoutbuffer[0][5] ), .B0(n1878), .Y(
        n1072) );
  AOI22X1TS U1581 ( .A0(n411), .A1(dataIn_WEST[5]), .B0(n389), .B1(n1356), .Y(
        n1071) );
  AOI22X1TS U1582 ( .A0(n1853), .A1(n1536), .B0(n396), .B1(dataIn_NORTH[5]), 
        .Y(n1070) );
  INVX2TS U1583 ( .A(n1616), .Y(n1088) );
  AOI21X1TS U1584 ( .A0(n1088), .A1(\dataoutbuffer[1][0] ), .B0(n1092), .Y(
        n1077) );
  AOI22X1TS U1585 ( .A0(n1073), .A1(n1362), .B0(n1819), .B1(n1103), .Y(n1076)
         );
  CLKBUFX2TS U1586 ( .A(dataIn_NORTH[0]), .Y(n1423) );
  CLKBUFX2TS U1587 ( .A(n1423), .Y(n1496) );
  CLKBUFX2TS U1588 ( .A(n1497), .Y(n1458) );
  AOI22X1TS U1589 ( .A0(n1079), .A1(n1496), .B0(n1074), .B1(n1458), .Y(n1075)
         );
  INVX2TS U1590 ( .A(n1078), .Y(n1816) );
  AOI21X1TS U1591 ( .A0(n1088), .A1(\dataoutbuffer[1][1] ), .B0(n1816), .Y(
        n1082) );
  AOI22X1TS U1592 ( .A0(n317), .A1(n1367), .B0(n1829), .B1(n1110), .Y(n1081)
         );
  CLKBUFX2TS U1593 ( .A(dataIn_NORTH[1]), .Y(n1428) );
  CLKBUFX2TS U1594 ( .A(n1428), .Y(n1504) );
  CLKBUFX2TS U1595 ( .A(n1505), .Y(n1465) );
  AOI22X1TS U1596 ( .A0(n1079), .A1(n1504), .B0(n331), .B1(n1465), .Y(n1080)
         );
  AOI21X1TS U1597 ( .A0(n1088), .A1(\dataoutbuffer[1][2] ), .B0(n1826), .Y(
        n1087) );
  AOI22X1TS U1598 ( .A0(n1093), .A1(n1371), .B0(n315), .B1(n1340), .Y(n1086)
         );
  CLKBUFX2TS U1599 ( .A(dataIn_NORTH[2]), .Y(n1433) );
  CLKBUFX2TS U1600 ( .A(n1433), .Y(n1511) );
  CLKBUFX2TS U1601 ( .A(n1512), .Y(n1471) );
  AOI22X1TS U1602 ( .A0(n1084), .A1(n1511), .B0(n1094), .B1(n1471), .Y(n1085)
         );
  AOI21X1TS U1603 ( .A0(n1088), .A1(\dataoutbuffer[1][3] ), .B0(n1836), .Y(
        n1091) );
  AOI22X1TS U1604 ( .A0(n1808), .A1(n1377), .B0(n1819), .B1(n1345), .Y(n1090)
         );
  CLKBUFX2TS U1605 ( .A(dataIn_NORTH[3]), .Y(n1439) );
  CLKBUFX2TS U1606 ( .A(n1439), .Y(n1520) );
  CLKBUFX2TS U1607 ( .A(n1521), .Y(n1477) );
  AOI22X1TS U1608 ( .A0(n322), .A1(n1520), .B0(n1810), .B1(n1477), .Y(n1089)
         );
  AOI21X1TS U1609 ( .A0(n1099), .A1(\dataoutbuffer[1][4] ), .B0(n1092), .Y(
        n1098) );
  AOI22X1TS U1610 ( .A0(n1093), .A1(n1382), .B0(n1829), .B1(n1350), .Y(n1097)
         );
  CLKBUFX2TS U1611 ( .A(dataIn_NORTH[4]), .Y(n1445) );
  CLKBUFX2TS U1612 ( .A(n1445), .Y(n1527) );
  CLKBUFX2TS U1613 ( .A(n1528), .Y(n1483) );
  AOI22X1TS U1614 ( .A0(n1095), .A1(n1527), .B0(n1094), .B1(n1483), .Y(n1096)
         );
  AOI21X1TS U1615 ( .A0(n1099), .A1(\dataoutbuffer[1][5] ), .B0(n1816), .Y(
        n1102) );
  AOI22X1TS U1616 ( .A0(n317), .A1(n1388), .B0(n315), .B1(n1356), .Y(n1101) );
  CLKBUFX2TS U1617 ( .A(dataIn_NORTH[5]), .Y(n1451) );
  CLKBUFX2TS U1618 ( .A(n1451), .Y(n1534) );
  CLKBUFX2TS U1619 ( .A(n1536), .Y(n1490) );
  AOI22X1TS U1620 ( .A0(n1079), .A1(n1534), .B0(n324), .B1(n1490), .Y(n1100)
         );
  INVX2TS U1621 ( .A(n1602), .Y(n1344) );
  AOI21X1TS U1622 ( .A0(n1344), .A1(\dataoutbuffer[2][0] ), .B0(n1787), .Y(
        n1109) );
  AOI22X1TS U1623 ( .A0(n1104), .A1(n1362), .B0(n1788), .B1(n1103), .Y(n1108)
         );
  AOI22X1TS U1624 ( .A0(n1106), .A1(n1496), .B0(n1105), .B1(dataIn_SOUTH[0]), 
        .Y(n1107) );
  AOI21X1TS U1625 ( .A0(n1344), .A1(\dataoutbuffer[2][1] ), .B0(n184), .Y(
        n1338) );
  AOI22X1TS U1626 ( .A0(n186), .A1(n1367), .B0(n1794), .B1(n1110), .Y(n1337)
         );
  INVX2TS U1627 ( .A(n1111), .Y(n1789) );
  AOI22X1TS U1628 ( .A0(n1789), .A1(n1504), .B0(n1357), .B1(dataIn_SOUTH[1]), 
        .Y(n1112) );
  AOI21X1TS U1629 ( .A0(n1344), .A1(\dataoutbuffer[2][2] ), .B0(n1800), .Y(
        n1343) );
  AOI22X1TS U1630 ( .A0(n1351), .A1(n1371), .B0(n183), .B1(n1340), .Y(n1342)
         );
  AOI22X1TS U1631 ( .A0(n977), .A1(n1511), .B0(n1795), .B1(dataIn_SOUTH[2]), 
        .Y(n1341) );
  AOI21X1TS U1632 ( .A0(n1344), .A1(\dataoutbuffer[2][3] ), .B0(n1787), .Y(
        n1349) );
  AOI22X1TS U1633 ( .A0(n1782), .A1(n1377), .B0(n1788), .B1(n1345), .Y(n1348)
         );
  AOI22X1TS U1634 ( .A0(n1783), .A1(n1520), .B0(n1346), .B1(dataIn_SOUTH[3]), 
        .Y(n1347) );
  AOI21X1TS U1635 ( .A0(n1355), .A1(\dataoutbuffer[2][4] ), .B0(n184), .Y(
        n1354) );
  AOI22X1TS U1636 ( .A0(n1351), .A1(n1382), .B0(n1794), .B1(n1350), .Y(n1353)
         );
  AOI22X1TS U1637 ( .A0(n194), .A1(n1527), .B0(n218), .B1(dataIn_SOUTH[4]), 
        .Y(n1352) );
  AOI21X1TS U1638 ( .A0(n1355), .A1(\dataoutbuffer[2][5] ), .B0(n1800), .Y(
        n1360) );
  AOI22X1TS U1639 ( .A0(n186), .A1(n1388), .B0(n183), .B1(n1356), .Y(n1359) );
  AOI22X1TS U1640 ( .A0(n1789), .A1(n1534), .B0(n1357), .B1(dataIn_SOUTH[5]), 
        .Y(n1358) );
  INVX2TS U1641 ( .A(n175), .Y(n1376) );
  AOI21X1TS U1642 ( .A0(n1376), .A1(\dataoutbuffer[3][0] ), .B0(n1760), .Y(
        n1366) );
  AOI22X1TS U1643 ( .A0(n1372), .A1(n1362), .B0(n1767), .B1(dataIn_EAST[0]), 
        .Y(n1365) );
  AOI22X1TS U1644 ( .A0(n1363), .A1(n1423), .B0(n146), .B1(n1458), .Y(n1364)
         );
  AOI21X1TS U1645 ( .A0(n1376), .A1(\dataoutbuffer[3][1] ), .B0(n132), .Y(
        n1370) );
  AOI22X1TS U1646 ( .A0(n147), .A1(n1367), .B0(n1761), .B1(dataIn_EAST[1]), 
        .Y(n1369) );
  AOI22X1TS U1647 ( .A0(n135), .A1(n1428), .B0(n1768), .B1(n1465), .Y(n1368)
         );
  AOI21X1TS U1648 ( .A0(n1376), .A1(\dataoutbuffer[3][2] ), .B0(n1773), .Y(
        n1375) );
  AOI22X1TS U1649 ( .A0(n1372), .A1(n1371), .B0(n157), .B1(dataIn_EAST[2]), 
        .Y(n1374) );
  AOI22X1TS U1650 ( .A0(n1383), .A1(n1433), .B0(n1776), .B1(n1471), .Y(n1373)
         );
  AOI21X1TS U1651 ( .A0(n1376), .A1(\dataoutbuffer[3][3] ), .B0(n1760), .Y(
        n1380) );
  AOI22X1TS U1652 ( .A0(n1755), .A1(n1377), .B0(n151), .B1(dataIn_EAST[3]), 
        .Y(n1379) );
  AOI22X1TS U1653 ( .A0(n1756), .A1(n1439), .B0(n1762), .B1(n1477), .Y(n1378)
         );
  AOI21X1TS U1654 ( .A0(n1387), .A1(\dataoutbuffer[3][4] ), .B0(n132), .Y(
        n1386) );
  AOI22X1TS U1655 ( .A0(n147), .A1(n1382), .B0(n1381), .B1(dataIn_EAST[4]), 
        .Y(n1385) );
  AOI22X1TS U1656 ( .A0(n1383), .A1(n1445), .B0(n1776), .B1(n1483), .Y(n1384)
         );
  AOI21X1TS U1657 ( .A0(n1387), .A1(\dataoutbuffer[3][5] ), .B0(n1773), .Y(
        n1392) );
  AOI22X1TS U1658 ( .A0(n1389), .A1(n1388), .B0(n1761), .B1(dataIn_EAST[5]), 
        .Y(n1391) );
  AOI22X1TS U1659 ( .A0(n1383), .A1(n1451), .B0(n130), .B1(n1490), .Y(n1390)
         );
  INVX2TS U1660 ( .A(n935), .Y(n1406) );
  AOI21X1TS U1661 ( .A0(n1406), .A1(\dataoutbuffer[4][0] ), .B0(n1728), .Y(
        n1398) );
  CLKBUFX2TS U1662 ( .A(dataIn_WEST[0]), .Y(n1495) );
  AOI22X1TS U1663 ( .A0(n1394), .A1(n1495), .B0(n1730), .B1(dataIn_EAST[0]), 
        .Y(n1397) );
  AOI22X1TS U1664 ( .A0(n1724), .A1(dataIn_SOUTH[0]), .B0(n1395), .B1(n1496), 
        .Y(n1396) );
  AOI21X1TS U1665 ( .A0(n1406), .A1(\dataoutbuffer[4][1] ), .B0(n275), .Y(
        n1401) );
  CLKBUFX2TS U1666 ( .A(dataIn_WEST[1]), .Y(n1503) );
  AOI22X1TS U1667 ( .A0(n283), .A1(n1503), .B0(n1737), .B1(dataIn_EAST[1]), 
        .Y(n1400) );
  AOI22X1TS U1668 ( .A0(n1739), .A1(dataIn_SOUTH[1]), .B0(n288), .B1(n1504), 
        .Y(n1399) );
  AOI21X1TS U1669 ( .A0(n1406), .A1(\dataoutbuffer[4][2] ), .B0(n1744), .Y(
        n1405) );
  CLKBUFX2TS U1670 ( .A(dataIn_WEST[2]), .Y(n1510) );
  AOI22X1TS U1671 ( .A0(n1410), .A1(n1510), .B0(n274), .B1(dataIn_EAST[2]), 
        .Y(n1404) );
  AOI22X1TS U1672 ( .A0(n1749), .A1(dataIn_SOUTH[2]), .B0(n1411), .B1(n1511), 
        .Y(n1403) );
  AOI21X1TS U1673 ( .A0(n1406), .A1(\dataoutbuffer[4][3] ), .B0(n1728), .Y(
        n1409) );
  CLKBUFX2TS U1674 ( .A(dataIn_WEST[3]), .Y(n1518) );
  AOI22X1TS U1675 ( .A0(n1722), .A1(n1518), .B0(n1730), .B1(dataIn_EAST[3]), 
        .Y(n1408) );
  AOI22X1TS U1676 ( .A0(n301), .A1(dataIn_SOUTH[3]), .B0(n1723), .B1(n1520), 
        .Y(n1407) );
  AOI21X1TS U1677 ( .A0(n1416), .A1(\dataoutbuffer[4][4] ), .B0(n275), .Y(
        n1415) );
  CLKBUFX2TS U1678 ( .A(dataIn_WEST[4]), .Y(n1526) );
  AOI22X1TS U1679 ( .A0(n1410), .A1(n1526), .B0(n1737), .B1(dataIn_EAST[4]), 
        .Y(n1414) );
  AOI22X1TS U1680 ( .A0(n1412), .A1(dataIn_SOUTH[4]), .B0(n1411), .B1(n1527), 
        .Y(n1413) );
  AOI21X1TS U1681 ( .A0(n1416), .A1(\dataoutbuffer[4][5] ), .B0(n1744), .Y(
        n1419) );
  CLKBUFX2TS U1682 ( .A(dataIn_WEST[5]), .Y(n1533) );
  AOI22X1TS U1683 ( .A0(n283), .A1(n1533), .B0(n274), .B1(dataIn_EAST[5]), .Y(
        n1418) );
  AOI22X1TS U1684 ( .A0(n1724), .A1(dataIn_SOUTH[5]), .B0(n280), .B1(n1534), 
        .Y(n1417) );
  INVX2TS U1685 ( .A(n912), .Y(n1438) );
  AOI21X1TS U1686 ( .A0(n1438), .A1(\dataoutbuffer[5][0] ), .B0(n1698), .Y(
        n1427) );
  AOI22X1TS U1687 ( .A0(n1421), .A1(n1495), .B0(n1700), .B1(n1456), .Y(n1426)
         );
  AOI22X1TS U1688 ( .A0(n1424), .A1(n1423), .B0(n1422), .B1(n1458), .Y(n1425)
         );
  AOI21X1TS U1689 ( .A0(n1438), .A1(\dataoutbuffer[5][1] ), .B0(n1706), .Y(
        n1431) );
  AOI22X1TS U1690 ( .A0(n247), .A1(n1503), .B0(n1708), .B1(n1464), .Y(n1430)
         );
  AOI22X1TS U1691 ( .A0(n1701), .A1(n1428), .B0(n1716), .B1(n1465), .Y(n1429)
         );
  AOI21X1TS U1692 ( .A0(n1438), .A1(\dataoutbuffer[5][2] ), .B0(n1713), .Y(
        n1437) );
  AOI22X1TS U1693 ( .A0(n1443), .A1(n1510), .B0(n1), .B1(n1470), .Y(n1436) );
  AOI22X1TS U1694 ( .A0(n1434), .A1(n1433), .B0(n1444), .B1(n1471), .Y(n1435)
         );
  AOI21X1TS U1695 ( .A0(n1438), .A1(\dataoutbuffer[5][3] ), .B0(n1698), .Y(
        n1442) );
  AOI22X1TS U1696 ( .A0(n1692), .A1(n1518), .B0(n1700), .B1(n1476), .Y(n1441)
         );
  AOI22X1TS U1697 ( .A0(n228), .A1(n1439), .B0(n1693), .B1(n1477), .Y(n1440)
         );
  AOI21X1TS U1698 ( .A0(n1450), .A1(\dataoutbuffer[5][4] ), .B0(n1706), .Y(
        n1449) );
  AOI22X1TS U1699 ( .A0(n1443), .A1(n1526), .B0(n1708), .B1(n1481), .Y(n1448)
         );
  AOI22X1TS U1700 ( .A0(n1446), .A1(n1445), .B0(n1444), .B1(n1483), .Y(n1447)
         );
  AOI21X1TS U1701 ( .A0(n1450), .A1(\dataoutbuffer[5][5] ), .B0(n1713), .Y(
        n1454) );
  AOI22X1TS U1702 ( .A0(n247), .A1(n1533), .B0(n1), .B1(n1489), .Y(n1453) );
  AOI22X1TS U1703 ( .A0(n1701), .A1(n1451), .B0(n242), .B1(n1490), .Y(n1452)
         );
  INVX2TS U1704 ( .A(n894), .Y(n1475) );
  AOI21X1TS U1705 ( .A0(n1475), .A1(\dataoutbuffer[6][0] ), .B0(n1668), .Y(
        n1463) );
  AOI22X1TS U1706 ( .A0(n1457), .A1(n1495), .B0(n1669), .B1(n1456), .Y(n1462)
         );
  AOI22X1TS U1707 ( .A0(n1460), .A1(dataIn_NORTH[0]), .B0(n1459), .B1(n1458), 
        .Y(n1461) );
  AOI21X1TS U1708 ( .A0(n1475), .A1(\dataoutbuffer[6][1] ), .B0(n1675), .Y(
        n1468) );
  AOI22X1TS U1709 ( .A0(n100), .A1(n1503), .B0(n1676), .B1(n1464), .Y(n1467)
         );
  AOI22X1TS U1710 ( .A0(n889), .A1(dataIn_NORTH[1]), .B0(n1484), .B1(n1465), 
        .Y(n1466) );
  AOI21X1TS U1711 ( .A0(n1475), .A1(\dataoutbuffer[6][2] ), .B0(n84), .Y(n1474) );
  AOI22X1TS U1712 ( .A0(n1482), .A1(n1510), .B0(n83), .B1(n1470), .Y(n1473) );
  AOI22X1TS U1713 ( .A0(n88), .A1(dataIn_NORTH[2]), .B0(n1484), .B1(n1471), 
        .Y(n1472) );
  AOI21X1TS U1714 ( .A0(n1475), .A1(\dataoutbuffer[6][3] ), .B0(n1668), .Y(
        n1480) );
  AOI22X1TS U1715 ( .A0(n1662), .A1(n1518), .B0(n1669), .B1(n1476), .Y(n1479)
         );
  AOI22X1TS U1716 ( .A0(n1664), .A1(dataIn_NORTH[3]), .B0(n96), .B1(n1477), 
        .Y(n1478) );
  AOI21X1TS U1717 ( .A0(n1488), .A1(\dataoutbuffer[6][4] ), .B0(n1675), .Y(
        n1487) );
  AOI22X1TS U1718 ( .A0(n1482), .A1(n1526), .B0(n1676), .B1(n1481), .Y(n1486)
         );
  AOI22X1TS U1719 ( .A0(n88), .A1(dataIn_NORTH[4]), .B0(n1484), .B1(n1483), 
        .Y(n1485) );
  AOI21X1TS U1720 ( .A0(n1488), .A1(\dataoutbuffer[6][5] ), .B0(n84), .Y(n1493) );
  AOI22X1TS U1721 ( .A0(n100), .A1(n1533), .B0(n83), .B1(n1489), .Y(n1492) );
  AOI22X1TS U1722 ( .A0(n103), .A1(dataIn_NORTH[5]), .B0(n117), .B1(n1490), 
        .Y(n1491) );
  INVX2TS U1723 ( .A(n877), .Y(n1517) );
  AOI21X1TS U1724 ( .A0(n1517), .A1(\dataoutbuffer[7][0] ), .B0(n1525), .Y(
        n1500) );
  AOI22X1TS U1725 ( .A0(n45), .A1(n1495), .B0(n1655), .B1(dataIn_EAST[0]), .Y(
        n1499) );
  AOI22X1TS U1726 ( .A0(n1513), .A1(n1497), .B0(n68), .B1(n1496), .Y(n1498) );
  INVX2TS U1727 ( .A(n1501), .Y(n1637) );
  AOI21X1TS U1728 ( .A0(n1517), .A1(\dataoutbuffer[7][1] ), .B0(n1637), .Y(
        n1508) );
  AOI22X1TS U1729 ( .A0(n67), .A1(n1503), .B0(n1638), .B1(dataIn_EAST[1]), .Y(
        n1507) );
  INVX2TS U1730 ( .A(n873), .Y(n1648) );
  AOI22X1TS U1731 ( .A0(n1648), .A1(n1505), .B0(n1647), .B1(n1504), .Y(n1506)
         );
  AOI21X1TS U1732 ( .A0(n1517), .A1(\dataoutbuffer[7][2] ), .B0(n1645), .Y(
        n1516) );
  AOI22X1TS U1733 ( .A0(n45), .A1(n1510), .B0(n29), .B1(dataIn_EAST[2]), .Y(
        n1515) );
  AOI22X1TS U1734 ( .A0(n1513), .A1(n1512), .B0(n1632), .B1(n1511), .Y(n1514)
         );
  AOI21X1TS U1735 ( .A0(n1517), .A1(\dataoutbuffer[7][3] ), .B0(n1654), .Y(
        n1524) );
  AOI22X1TS U1736 ( .A0(n1519), .A1(n1518), .B0(n1655), .B1(dataIn_EAST[3]), 
        .Y(n1523) );
  AOI22X1TS U1737 ( .A0(n69), .A1(n1521), .B0(n1632), .B1(n1520), .Y(n1522) );
  AOI21X1TS U1738 ( .A0(n1532), .A1(\dataoutbuffer[7][4] ), .B0(n1525), .Y(
        n1531) );
  AOI22X1TS U1739 ( .A0(n1646), .A1(n1526), .B0(n1638), .B1(dataIn_EAST[4]), 
        .Y(n1530) );
  AOI22X1TS U1740 ( .A0(n1639), .A1(n1528), .B0(n1657), .B1(n1527), .Y(n1529)
         );
  AOI21X1TS U1741 ( .A0(n1532), .A1(\dataoutbuffer[7][5] ), .B0(n1637), .Y(
        n1539) );
  AOI22X1TS U1742 ( .A0(n32), .A1(n1533), .B0(n29), .B1(dataIn_EAST[5]), .Y(
        n1538) );
  AOI22X1TS U1743 ( .A0(n1648), .A1(n1536), .B0(n1535), .B1(n1534), .Y(n1537)
         );
  CLKBUFX2TS U1744 ( .A(n1628), .Y(n1580) );
  INVX2TS U1745 ( .A(n1540), .Y(n1624) );
  AOI22X1TS U1746 ( .A0(n1542), .A1(n1563), .B0(n1562), .B1(n1541), .Y(n1544)
         );
  AOI22X1TS U1747 ( .A0(n1545), .A1(n1624), .B0(n1544), .B1(n1543), .Y(n1547)
         );
  AOI22X1TS U1748 ( .A0(n1548), .A1(n1580), .B0(n1547), .B1(n1546), .Y(n1550)
         );
  AOI32X1TS U1749 ( .A0(n1550), .A1(n1494), .A2(n1549), .B0(n1652), .B1(n1919), 
        .Y(n1217) );
  INVX2TS U1750 ( .A(n1540), .Y(n1596) );
  AOI22X1TS U1751 ( .A0(n1552), .A1(n1563), .B0(n1562), .B1(n1551), .Y(n1554)
         );
  AOI22X1TS U1752 ( .A0(n1555), .A1(n1596), .B0(n1554), .B1(n1553), .Y(n1557)
         );
  AOI22X1TS U1753 ( .A0(n1558), .A1(n1580), .B0(n1557), .B1(n1556), .Y(n1560)
         );
  AOI32X1TS U1754 ( .A0(n1560), .A1(n1455), .A2(n1559), .B0(n1682), .B1(n1920), 
        .Y(n1216) );
  AOI22X1TS U1755 ( .A0(n1564), .A1(n1563), .B0(n1562), .B1(n1561), .Y(n1566)
         );
  AOI22X1TS U1756 ( .A0(n1567), .A1(n1596), .B0(n1566), .B1(n1565), .Y(n1569)
         );
  AOI22X1TS U1757 ( .A0(n1570), .A1(n1580), .B0(n1569), .B1(n1568), .Y(n1572)
         );
  AOI32X1TS U1758 ( .A0(n1572), .A1(n1420), .A2(n1571), .B0(n1712), .B1(n1921), 
        .Y(n1215) );
  CLKBUFX2TS U1759 ( .A(n1620), .Y(n1606) );
  CLKBUFX2TS U1760 ( .A(n1619), .Y(n1605) );
  AOI22X1TS U1761 ( .A0(n1574), .A1(n1606), .B0(n1605), .B1(n1573), .Y(n1576)
         );
  AOI22X1TS U1762 ( .A0(n1577), .A1(n1624), .B0(n1576), .B1(n1575), .Y(n1579)
         );
  AOI22X1TS U1763 ( .A0(n1581), .A1(n1580), .B0(n1579), .B1(n1578), .Y(n1583)
         );
  AOI32X1TS U1764 ( .A0(n1583), .A1(n1393), .A2(n1582), .B0(n1743), .B1(n1922), 
        .Y(n1214) );
  AOI22X1TS U1765 ( .A0(n23), .A1(n1606), .B0(n1605), .B1(n24), .Y(n1585) );
  AOI22X1TS U1766 ( .A0(n1586), .A1(n1596), .B0(n1585), .B1(n1584), .Y(n1588)
         );
  AOI22X1TS U1767 ( .A0(n1589), .A1(n1628), .B0(n1588), .B1(n1587), .Y(n1591)
         );
  AOI32X1TS U1768 ( .A0(n1591), .A1(n1361), .A2(n1590), .B0(n1772), .B1(n1923), 
        .Y(n1213) );
  AOI22X1TS U1769 ( .A0(n1593), .A1(n1606), .B0(n1605), .B1(n1592), .Y(n1595)
         );
  AOI22X1TS U1770 ( .A0(n1597), .A1(n1596), .B0(n1595), .B1(n1594), .Y(n1599)
         );
  AOI22X1TS U1771 ( .A0(n1600), .A1(n1613), .B0(n1599), .B1(n1598), .Y(n1603)
         );
  AOI32X1TS U1772 ( .A0(n1603), .A1(n1602), .A2(n1601), .B0(n1799), .B1(n1924), 
        .Y(n1212) );
  AOI22X1TS U1773 ( .A0(n1607), .A1(n1606), .B0(n1605), .B1(n1604), .Y(n1609)
         );
  AOI22X1TS U1774 ( .A0(n1610), .A1(n1624), .B0(n1609), .B1(n1608), .Y(n1612)
         );
  AOI22X1TS U1775 ( .A0(n1614), .A1(n1613), .B0(n1612), .B1(n1611), .Y(n1617)
         );
  AOI32X1TS U1776 ( .A0(n1617), .A1(n1616), .A2(n1615), .B0(n1835), .B1(n1925), 
        .Y(n1211) );
  AOI22X1TS U1777 ( .A0(n1621), .A1(n1620), .B0(n1619), .B1(n1618), .Y(n1623)
         );
  AOI22X1TS U1778 ( .A0(n1625), .A1(n1624), .B0(n1623), .B1(n1622), .Y(n1627)
         );
  AOI22X1TS U1779 ( .A0(n1629), .A1(n1628), .B0(n1627), .B1(n1626), .Y(n1631)
         );
  AOI32X1TS U1780 ( .A0(n1631), .A1(n1037), .A2(n1630), .B0(n1877), .B1(n1926), 
        .Y(n1210) );
  AOI22X1TS U1781 ( .A0(n1806), .A1(n1637), .B0(n1643), .B1(
        \destinationAddressbuffer[7][0] ), .Y(n1635) );
  CLKBUFX2TS U1782 ( .A(destinationAddressIn_WEST[0]), .Y(n1721) );
  AOI22X1TS U1783 ( .A0(n67), .A1(n1721), .B0(n872), .B1(n1691), .Y(n1634) );
  CLKBUFX2TS U1784 ( .A(n1663), .Y(n1811) );
  AOI22X1TS U1785 ( .A0(n1648), .A1(destinationAddressIn_SOUTH[0]), .B0(n1632), 
        .B1(n1811), .Y(n1633) );
  AOI22X1TS U1786 ( .A0(n1637), .A1(n1636), .B0(n1643), .B1(
        \destinationAddressbuffer[7][1] ), .Y(n1642) );
  CLKBUFX2TS U1787 ( .A(destinationAddressIn_WEST[1]), .Y(n1731) );
  AOI22X1TS U1788 ( .A0(n32), .A1(n1731), .B0(n1638), .B1(n1699), .Y(n1641) );
  CLKBUFX2TS U1789 ( .A(n1670), .Y(n1821) );
  AOI22X1TS U1790 ( .A0(n1639), .A1(destinationAddressIn_SOUTH[1]), .B0(n40), 
        .B1(n1821), .Y(n1640) );
  AOI22X1TS U1791 ( .A0(n1645), .A1(n1644), .B0(n1643), .B1(
        \destinationAddressbuffer[7][2] ), .Y(n1651) );
  CLKBUFX2TS U1792 ( .A(destinationAddressIn_WEST[2]), .Y(n1738) );
  AOI22X1TS U1793 ( .A0(n1646), .A1(n1738), .B0(n29), .B1(n1707), .Y(n1650) );
  CLKBUFX2TS U1794 ( .A(n1677), .Y(n1831) );
  AOI22X1TS U1795 ( .A0(n1648), .A1(destinationAddressIn_SOUTH[2]), .B0(n1647), 
        .B1(n1831), .Y(n1649) );
  AOI22X1TS U1796 ( .A0(n1654), .A1(n1653), .B0(n1652), .B1(
        \destinationAddressbuffer[7][3] ), .Y(n1660) );
  CLKBUFX2TS U1797 ( .A(destinationAddressIn_WEST[3]), .Y(n1746) );
  AOI22X1TS U1798 ( .A0(n1656), .A1(n1746), .B0(n1655), .B1(n1714), .Y(n1659)
         );
  CLKBUFX2TS U1799 ( .A(n1684), .Y(n1842) );
  AOI22X1TS U1800 ( .A0(n35), .A1(destinationAddressIn_SOUTH[3]), .B0(n1657), 
        .B1(n1842), .Y(n1658) );
  AOI22X1TS U1801 ( .A0(n1847), .A1(n1661), .B0(n1674), .B1(
        \destinationAddressbuffer[6][0] ), .Y(n1667) );
  AOI22X1TS U1802 ( .A0(n1662), .A1(n1721), .B0(n95), .B1(n1691), .Y(n1666) );
  CLKBUFX2TS U1803 ( .A(n1663), .Y(n1850) );
  CLKBUFX2TS U1804 ( .A(destinationAddressIn_SOUTH[0]), .Y(n1852) );
  CLKBUFX2TS U1805 ( .A(n1852), .Y(n1809) );
  AOI22X1TS U1806 ( .A0(n1664), .A1(n1850), .B0(n1685), .B1(n1809), .Y(n1665)
         );
  AOI22X1TS U1807 ( .A0(n1729), .A1(n1668), .B0(n1674), .B1(
        \destinationAddressbuffer[6][1] ), .Y(n1673) );
  AOI22X1TS U1808 ( .A0(n110), .A1(n1731), .B0(n1669), .B1(n1699), .Y(n1672)
         );
  CLKBUFX2TS U1809 ( .A(n1670), .Y(n1861) );
  CLKBUFX2TS U1810 ( .A(destinationAddressIn_SOUTH[1]), .Y(n1862) );
  CLKBUFX2TS U1811 ( .A(n1862), .Y(n1820) );
  AOI22X1TS U1812 ( .A0(n88), .A1(n1861), .B0(n1678), .B1(n1820), .Y(n1671) );
  AOI22X1TS U1813 ( .A0(n1736), .A1(n1675), .B0(n1674), .B1(
        \destinationAddressbuffer[6][2] ), .Y(n1681) );
  AOI22X1TS U1814 ( .A0(n1683), .A1(n1738), .B0(n1676), .B1(n1707), .Y(n1680)
         );
  CLKBUFX2TS U1815 ( .A(n1677), .Y(n1871) );
  CLKBUFX2TS U1816 ( .A(destinationAddressIn_SOUTH[2]), .Y(n1872) );
  CLKBUFX2TS U1817 ( .A(n1872), .Y(n1830) );
  AOI22X1TS U1818 ( .A0(n1686), .A1(n1871), .B0(n1678), .B1(n1830), .Y(n1679)
         );
  AOI22X1TS U1819 ( .A0(n1745), .A1(n84), .B0(n1682), .B1(
        \destinationAddressbuffer[6][3] ), .Y(n1689) );
  AOI22X1TS U1820 ( .A0(n1683), .A1(n1746), .B0(n896), .B1(n1714), .Y(n1688)
         );
  CLKBUFX2TS U1821 ( .A(n1684), .Y(n1882) );
  CLKBUFX2TS U1822 ( .A(destinationAddressIn_SOUTH[3]), .Y(n1884) );
  CLKBUFX2TS U1823 ( .A(n1884), .Y(n1840) );
  AOI22X1TS U1824 ( .A0(n1686), .A1(n1882), .B0(n1685), .B1(n1840), .Y(n1687)
         );
  AOI22X1TS U1825 ( .A0(n1847), .A1(n1690), .B0(n1705), .B1(
        \destinationAddressbuffer[5][0] ), .Y(n1697) );
  AOI22X1TS U1826 ( .A0(n1692), .A1(n1721), .B0(n914), .B1(n1691), .Y(n1696)
         );
  AOI22X1TS U1827 ( .A0(n1694), .A1(n1850), .B0(n1693), .B1(
        destinationAddressIn_SOUTH[0]), .Y(n1695) );
  AOI22X1TS U1828 ( .A0(readRequesterAddress[1]), .A1(n1698), .B0(n1705), .B1(
        \destinationAddressbuffer[5][1] ), .Y(n1704) );
  AOI22X1TS U1829 ( .A0(n259), .A1(n1731), .B0(n1700), .B1(n1699), .Y(n1703)
         );
  AOI22X1TS U1830 ( .A0(n1701), .A1(n1861), .B0(n230), .B1(
        destinationAddressIn_SOUTH[1]), .Y(n1702) );
  AOI22X1TS U1831 ( .A0(readRequesterAddress[2]), .A1(n1706), .B0(n1705), .B1(
        \destinationAddressbuffer[5][2] ), .Y(n1711) );
  AOI22X1TS U1832 ( .A0(n1715), .A1(n1738), .B0(n1708), .B1(n1707), .Y(n1710)
         );
  AOI22X1TS U1833 ( .A0(n1424), .A1(n1871), .B0(n1716), .B1(
        destinationAddressIn_SOUTH[2]), .Y(n1709) );
  AOI22X1TS U1834 ( .A0(readRequesterAddress[3]), .A1(n1713), .B0(n1712), .B1(
        \destinationAddressbuffer[5][3] ), .Y(n1719) );
  AOI22X1TS U1835 ( .A0(n1715), .A1(n1746), .B0(n1), .B1(n1714), .Y(n1718) );
  AOI22X1TS U1836 ( .A0(n228), .A1(n1882), .B0(n1716), .B1(
        destinationAddressIn_SOUTH[3]), .Y(n1717) );
  AOI22X1TS U1837 ( .A0(n1754), .A1(n1720), .B0(n1735), .B1(
        \destinationAddressbuffer[4][0] ), .Y(n1727) );
  AOI22X1TS U1838 ( .A0(n1722), .A1(n1721), .B0(n937), .B1(
        destinationAddressIn_EAST[0]), .Y(n1726) );
  AOI22X1TS U1839 ( .A0(n1724), .A1(n1852), .B0(n1723), .B1(n1850), .Y(n1725)
         );
  AOI22X1TS U1840 ( .A0(n1729), .A1(n1728), .B0(n1735), .B1(
        \destinationAddressbuffer[4][1] ), .Y(n1734) );
  AOI22X1TS U1841 ( .A0(n298), .A1(n1731), .B0(n1730), .B1(
        destinationAddressIn_EAST[1]), .Y(n1733) );
  AOI22X1TS U1842 ( .A0(n301), .A1(n1862), .B0(n1411), .B1(n1861), .Y(n1732)
         );
  AOI22X1TS U1843 ( .A0(n1736), .A1(n275), .B0(n1735), .B1(
        \destinationAddressbuffer[4][2] ), .Y(n1742) );
  AOI22X1TS U1844 ( .A0(n1747), .A1(n1738), .B0(n1737), .B1(
        destinationAddressIn_EAST[2]), .Y(n1741) );
  AOI22X1TS U1845 ( .A0(n1739), .A1(n1872), .B0(n1748), .B1(n1871), .Y(n1740)
         );
  AOI22X1TS U1846 ( .A0(n1745), .A1(n1744), .B0(n1743), .B1(
        \destinationAddressbuffer[4][3] ), .Y(n1752) );
  AOI22X1TS U1847 ( .A0(n1747), .A1(n1746), .B0(n274), .B1(
        destinationAddressIn_EAST[3]), .Y(n1751) );
  AOI22X1TS U1848 ( .A0(n1749), .A1(n1884), .B0(n1748), .B1(n1882), .Y(n1750)
         );
  AOI22X1TS U1849 ( .A0(n1754), .A1(n1753), .B0(n1766), .B1(
        \destinationAddressbuffer[3][0] ), .Y(n1759) );
  AOI22X1TS U1850 ( .A0(n1755), .A1(destinationAddressIn_WEST[0]), .B0(n151), 
        .B1(destinationAddressIn_EAST[0]), .Y(n1758) );
  AOI22X1TS U1851 ( .A0(n1756), .A1(n1811), .B0(n1762), .B1(n1809), .Y(n1757)
         );
  AOI22X1TS U1852 ( .A0(n1817), .A1(n1760), .B0(n1766), .B1(
        \destinationAddressbuffer[3][1] ), .Y(n1765) );
  AOI22X1TS U1853 ( .A0(n1775), .A1(destinationAddressIn_WEST[1]), .B0(n1761), 
        .B1(destinationAddressIn_EAST[1]), .Y(n1764) );
  AOI22X1TS U1854 ( .A0(n1777), .A1(n1821), .B0(n1762), .B1(n1820), .Y(n1763)
         );
  AOI22X1TS U1855 ( .A0(n1827), .A1(n132), .B0(n1766), .B1(
        \destinationAddressbuffer[3][2] ), .Y(n1771) );
  AOI22X1TS U1856 ( .A0(n165), .A1(destinationAddressIn_WEST[2]), .B0(n1767), 
        .B1(destinationAddressIn_EAST[2]), .Y(n1770) );
  AOI22X1TS U1857 ( .A0(n135), .A1(n1831), .B0(n1768), .B1(n1830), .Y(n1769)
         );
  AOI22X1TS U1858 ( .A0(n1837), .A1(n1773), .B0(n1772), .B1(
        \destinationAddressbuffer[3][3] ), .Y(n1780) );
  AOI22X1TS U1859 ( .A0(n1775), .A1(destinationAddressIn_WEST[3]), .B0(n1774), 
        .B1(destinationAddressIn_EAST[3]), .Y(n1779) );
  AOI22X1TS U1860 ( .A0(n1777), .A1(n1842), .B0(n1776), .B1(n1840), .Y(n1778)
         );
  AOI22X1TS U1861 ( .A0(n1806), .A1(n1781), .B0(n1793), .B1(
        \destinationAddressbuffer[2][0] ), .Y(n1786) );
  AOI22X1TS U1862 ( .A0(n1782), .A1(n1848), .B0(n197), .B1(n1807), .Y(n1785)
         );
  AOI22X1TS U1863 ( .A0(n1783), .A1(n1811), .B0(n190), .B1(n1809), .Y(n1784)
         );
  AOI22X1TS U1864 ( .A0(n1858), .A1(n1787), .B0(n1793), .B1(
        \destinationAddressbuffer[2][1] ), .Y(n1792) );
  AOI22X1TS U1865 ( .A0(n214), .A1(n1860), .B0(n1788), .B1(n1818), .Y(n1791)
         );
  AOI22X1TS U1866 ( .A0(n1789), .A1(n1821), .B0(n1795), .B1(n1820), .Y(n1790)
         );
  AOI22X1TS U1867 ( .A0(n1868), .A1(n184), .B0(n1793), .B1(
        \destinationAddressbuffer[2][2] ), .Y(n1798) );
  AOI22X1TS U1868 ( .A0(n1801), .A1(n1870), .B0(n1794), .B1(n1828), .Y(n1797)
         );
  AOI22X1TS U1869 ( .A0(n1802), .A1(n1831), .B0(n1795), .B1(n1830), .Y(n1796)
         );
  AOI22X1TS U1870 ( .A0(n1879), .A1(n1800), .B0(n1799), .B1(
        \destinationAddressbuffer[2][3] ), .Y(n1805) );
  AOI22X1TS U1871 ( .A0(n1801), .A1(n1880), .B0(n983), .B1(n1838), .Y(n1804)
         );
  AOI22X1TS U1872 ( .A0(n1802), .A1(n1842), .B0(n190), .B1(n1840), .Y(n1803)
         );
  AOI22X1TS U1873 ( .A0(n1806), .A1(n1816), .B0(n1825), .B1(
        \destinationAddressbuffer[1][0] ), .Y(n1815) );
  AOI22X1TS U1874 ( .A0(n1808), .A1(n1848), .B0(n335), .B1(n1807), .Y(n1814)
         );
  AOI22X1TS U1875 ( .A0(n1812), .A1(n1811), .B0(n1810), .B1(n1809), .Y(n1813)
         );
  AOI22X1TS U1876 ( .A0(n1817), .A1(n1816), .B0(n1825), .B1(
        \destinationAddressbuffer[1][1] ), .Y(n1824) );
  AOI22X1TS U1877 ( .A0(n372), .A1(n1860), .B0(n1819), .B1(n1818), .Y(n1823)
         );
  AOI22X1TS U1878 ( .A0(n1079), .A1(n1821), .B0(n1841), .B1(n1820), .Y(n1822)
         );
  AOI22X1TS U1879 ( .A0(n1827), .A1(n1826), .B0(n1825), .B1(
        \destinationAddressbuffer[1][2] ), .Y(n1834) );
  AOI22X1TS U1880 ( .A0(n1839), .A1(n1870), .B0(n1829), .B1(n1828), .Y(n1833)
         );
  AOI22X1TS U1881 ( .A0(n1011), .A1(n1831), .B0(n1841), .B1(n1830), .Y(n1832)
         );
  AOI22X1TS U1882 ( .A0(n1837), .A1(n1836), .B0(n1835), .B1(
        \destinationAddressbuffer[1][3] ), .Y(n1845) );
  AOI22X1TS U1883 ( .A0(n1839), .A1(n1880), .B0(n1009), .B1(n1838), .Y(n1844)
         );
  AOI22X1TS U1884 ( .A0(n1812), .A1(n1842), .B0(n1841), .B1(n1840), .Y(n1843)
         );
  AOI22X1TS U1885 ( .A0(n1847), .A1(n1846), .B0(n1866), .B1(
        \destinationAddressbuffer[0][0] ), .Y(n1856) );
  AOI22X1TS U1886 ( .A0(n1849), .A1(n1848), .B0(n405), .B1(
        destinationAddressIn_EAST[0]), .Y(n1855) );
  AOI22X1TS U1887 ( .A0(n1853), .A1(n1852), .B0(n1851), .B1(n1850), .Y(n1854)
         );
  AOI22X1TS U1888 ( .A0(n1858), .A1(n1857), .B0(n1866), .B1(
        \destinationAddressbuffer[0][1] ), .Y(n1865) );
  AOI22X1TS U1889 ( .A0(n424), .A1(n1860), .B0(n1859), .B1(
        destinationAddressIn_EAST[1]), .Y(n1864) );
  AOI22X1TS U1890 ( .A0(n430), .A1(n1862), .B0(n415), .B1(n1861), .Y(n1863) );
  AOI22X1TS U1891 ( .A0(n1868), .A1(n1867), .B0(n1866), .B1(
        \destinationAddressbuffer[0][2] ), .Y(n1876) );
  AOI22X1TS U1892 ( .A0(n1881), .A1(n1870), .B0(n1869), .B1(
        destinationAddressIn_EAST[2]), .Y(n1875) );
  AOI22X1TS U1893 ( .A0(n1873), .A1(n1872), .B0(n1883), .B1(n1871), .Y(n1874)
         );
  AOI22X1TS U1894 ( .A0(n1879), .A1(n1878), .B0(n1877), .B1(
        \destinationAddressbuffer[0][3] ), .Y(n1888) );
  AOI22X1TS U1895 ( .A0(n1881), .A1(n1880), .B0(n1039), .B1(
        destinationAddressIn_EAST[3]), .Y(n1887) );
  AOI22X1TS U1896 ( .A0(n1885), .A1(n1884), .B0(n1883), .B1(n1882), .Y(n1886)
         );
endmodule


module outputPortArbiter_1 ( clk, reset, selectBit_NORTH, 
        destinationAddressIn_NORTH, requesterAddressIn_NORTH, readIn_NORTH, 
        writeIn_NORTH, dataIn_NORTH, selectBit_SOUTH, 
        destinationAddressIn_SOUTH, requesterAddressIn_SOUTH, readIn_SOUTH, 
        writeIn_SOUTH, dataIn_SOUTH, selectBit_EAST, destinationAddressIn_EAST, 
        requesterAddressIn_EAST, readIn_EAST, writeIn_EAST, dataIn_EAST, 
        selectBit_WEST, destinationAddressIn_WEST, requesterAddressIn_WEST, 
        readIn_WEST, writeIn_WEST, dataIn_WEST, readReady, 
        readRequesterAddress, cacheDataOut, destinationAddressOut, 
        requesterAddressOut, readOut, writeOut, dataOut );
  input [11:0] destinationAddressIn_NORTH;
  input [3:0] requesterAddressIn_NORTH;
  input [5:0] dataIn_NORTH;
  input [11:0] destinationAddressIn_SOUTH;
  input [3:0] requesterAddressIn_SOUTH;
  input [5:0] dataIn_SOUTH;
  input [11:0] destinationAddressIn_EAST;
  input [3:0] requesterAddressIn_EAST;
  input [5:0] dataIn_EAST;
  input [11:0] destinationAddressIn_WEST;
  input [3:0] requesterAddressIn_WEST;
  input [5:0] dataIn_WEST;
  input [3:0] readRequesterAddress;
  input [5:0] cacheDataOut;
  output [11:0] destinationAddressOut;
  output [3:0] requesterAddressOut;
  output [5:0] dataOut;
  input clk, reset, selectBit_NORTH, readIn_NORTH, writeIn_NORTH,
         selectBit_SOUTH, readIn_SOUTH, writeIn_SOUTH, selectBit_EAST,
         readIn_EAST, writeIn_EAST, selectBit_WEST, readIn_WEST, writeIn_WEST,
         readReady;
  output readOut, writeOut;
  wire   \requesterAddressbuffer[0][3] , \requesterAddressbuffer[0][2] ,
         \requesterAddressbuffer[0][1] , \requesterAddressbuffer[0][0] ,
         \requesterAddressbuffer[1][3] , \requesterAddressbuffer[1][2] ,
         \requesterAddressbuffer[1][1] , \requesterAddressbuffer[1][0] ,
         \requesterAddressbuffer[2][3] , \requesterAddressbuffer[2][2] ,
         \requesterAddressbuffer[2][1] , \requesterAddressbuffer[2][0] ,
         \requesterAddressbuffer[3][3] , \requesterAddressbuffer[3][2] ,
         \requesterAddressbuffer[3][1] , \requesterAddressbuffer[3][0] ,
         \requesterAddressbuffer[4][3] , \requesterAddressbuffer[4][2] ,
         \requesterAddressbuffer[4][1] , \requesterAddressbuffer[4][0] ,
         \requesterAddressbuffer[5][3] , \requesterAddressbuffer[5][2] ,
         \requesterAddressbuffer[5][1] , \requesterAddressbuffer[5][0] ,
         \requesterAddressbuffer[6][3] , \requesterAddressbuffer[6][2] ,
         \requesterAddressbuffer[6][1] , \requesterAddressbuffer[6][0] ,
         \requesterAddressbuffer[7][3] , \requesterAddressbuffer[7][2] ,
         \requesterAddressbuffer[7][1] , \requesterAddressbuffer[7][0] ,
         \destinationAddressbuffer[0][11] , \destinationAddressbuffer[0][10] ,
         \destinationAddressbuffer[0][9] , \destinationAddressbuffer[0][8] ,
         \destinationAddressbuffer[0][7] , \destinationAddressbuffer[0][6] ,
         \destinationAddressbuffer[0][5] , \destinationAddressbuffer[0][4] ,
         \destinationAddressbuffer[0][3] , \destinationAddressbuffer[0][2] ,
         \destinationAddressbuffer[0][1] , \destinationAddressbuffer[0][0] ,
         \destinationAddressbuffer[1][11] , \destinationAddressbuffer[1][10] ,
         \destinationAddressbuffer[1][9] , \destinationAddressbuffer[1][8] ,
         \destinationAddressbuffer[1][7] , \destinationAddressbuffer[1][6] ,
         \destinationAddressbuffer[1][5] , \destinationAddressbuffer[1][4] ,
         \destinationAddressbuffer[1][3] , \destinationAddressbuffer[1][2] ,
         \destinationAddressbuffer[1][1] , \destinationAddressbuffer[1][0] ,
         \destinationAddressbuffer[2][11] , \destinationAddressbuffer[2][10] ,
         \destinationAddressbuffer[2][9] , \destinationAddressbuffer[2][8] ,
         \destinationAddressbuffer[2][7] , \destinationAddressbuffer[2][6] ,
         \destinationAddressbuffer[2][5] , \destinationAddressbuffer[2][4] ,
         \destinationAddressbuffer[2][3] , \destinationAddressbuffer[2][2] ,
         \destinationAddressbuffer[2][1] , \destinationAddressbuffer[2][0] ,
         \destinationAddressbuffer[3][11] , \destinationAddressbuffer[3][10] ,
         \destinationAddressbuffer[3][9] , \destinationAddressbuffer[3][8] ,
         \destinationAddressbuffer[3][7] , \destinationAddressbuffer[3][6] ,
         \destinationAddressbuffer[3][5] , \destinationAddressbuffer[3][4] ,
         \destinationAddressbuffer[3][3] , \destinationAddressbuffer[3][2] ,
         \destinationAddressbuffer[3][1] , \destinationAddressbuffer[3][0] ,
         \destinationAddressbuffer[4][11] , \destinationAddressbuffer[4][10] ,
         \destinationAddressbuffer[4][9] , \destinationAddressbuffer[4][8] ,
         \destinationAddressbuffer[4][7] , \destinationAddressbuffer[4][6] ,
         \destinationAddressbuffer[4][5] , \destinationAddressbuffer[4][4] ,
         \destinationAddressbuffer[4][3] , \destinationAddressbuffer[4][2] ,
         \destinationAddressbuffer[4][1] , \destinationAddressbuffer[4][0] ,
         \destinationAddressbuffer[5][11] , \destinationAddressbuffer[5][10] ,
         \destinationAddressbuffer[5][9] , \destinationAddressbuffer[5][8] ,
         \destinationAddressbuffer[5][7] , \destinationAddressbuffer[5][6] ,
         \destinationAddressbuffer[5][5] , \destinationAddressbuffer[5][4] ,
         \destinationAddressbuffer[5][3] , \destinationAddressbuffer[5][2] ,
         \destinationAddressbuffer[5][1] , \destinationAddressbuffer[5][0] ,
         \destinationAddressbuffer[6][11] , \destinationAddressbuffer[6][10] ,
         \destinationAddressbuffer[6][9] , \destinationAddressbuffer[6][8] ,
         \destinationAddressbuffer[6][7] , \destinationAddressbuffer[6][6] ,
         \destinationAddressbuffer[6][5] , \destinationAddressbuffer[6][4] ,
         \destinationAddressbuffer[6][3] , \destinationAddressbuffer[6][2] ,
         \destinationAddressbuffer[6][1] , \destinationAddressbuffer[6][0] ,
         \destinationAddressbuffer[7][11] , \destinationAddressbuffer[7][10] ,
         \destinationAddressbuffer[7][9] , \destinationAddressbuffer[7][8] ,
         \destinationAddressbuffer[7][7] , \destinationAddressbuffer[7][6] ,
         \destinationAddressbuffer[7][5] , \destinationAddressbuffer[7][4] ,
         \destinationAddressbuffer[7][3] , \destinationAddressbuffer[7][2] ,
         \destinationAddressbuffer[7][1] , \destinationAddressbuffer[7][0] ,
         \dataoutbuffer[7][5] , \dataoutbuffer[7][4] , \dataoutbuffer[7][3] ,
         \dataoutbuffer[7][2] , \dataoutbuffer[7][1] , \dataoutbuffer[7][0] ,
         \dataoutbuffer[6][5] , \dataoutbuffer[6][4] , \dataoutbuffer[6][3] ,
         \dataoutbuffer[6][2] , \dataoutbuffer[6][1] , \dataoutbuffer[6][0] ,
         \dataoutbuffer[5][5] , \dataoutbuffer[5][4] , \dataoutbuffer[5][3] ,
         \dataoutbuffer[5][2] , \dataoutbuffer[5][1] , \dataoutbuffer[5][0] ,
         \dataoutbuffer[4][5] , \dataoutbuffer[4][4] , \dataoutbuffer[4][3] ,
         \dataoutbuffer[4][2] , \dataoutbuffer[4][1] , \dataoutbuffer[4][0] ,
         \dataoutbuffer[3][5] , \dataoutbuffer[3][4] , \dataoutbuffer[3][3] ,
         \dataoutbuffer[3][2] , \dataoutbuffer[3][1] , \dataoutbuffer[3][0] ,
         \dataoutbuffer[2][5] , \dataoutbuffer[2][4] , \dataoutbuffer[2][3] ,
         \dataoutbuffer[2][2] , \dataoutbuffer[2][1] , \dataoutbuffer[2][0] ,
         \dataoutbuffer[1][5] , \dataoutbuffer[1][4] , \dataoutbuffer[1][3] ,
         \dataoutbuffer[1][2] , \dataoutbuffer[1][1] , \dataoutbuffer[1][0] ,
         \dataoutbuffer[0][5] , \dataoutbuffer[0][4] , \dataoutbuffer[0][3] ,
         \dataoutbuffer[0][2] , \dataoutbuffer[0][1] , \dataoutbuffer[0][0] ,
         N2624, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155;
  wire   [0:7] writeOutbuffer;
  wire   [0:7] readOutbuffer;

  DFFNSRX1TS full_reg_reg ( .D(N2624), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(
        n1924) );
  DFFNSRX1TS \dataoutbuffer_reg[0][0]  ( .D(n1996), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][1]  ( .D(n1997), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][2]  ( .D(n1998), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][3]  ( .D(n1999), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][4]  ( .D(n2000), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][5]  ( .D(n2001), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][5] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[2][0]  ( .D(n1984), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[2][1]  ( .D(n1985), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[2][2]  ( .D(n1986), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[2][3]  ( .D(n1987), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][0]  ( .D(n2120), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][1]  ( .D(n2121), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][2]  ( .D(n2122), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][3]  ( .D(n2123), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][3] ) );
  DFFNSRX1TS \writeOutbuffer_reg[7]  ( .D(n2044), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[7]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][4]  ( .D(n2064), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][5]  ( .D(n2065), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][6]  ( .D(n2066), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][7]  ( .D(n2067), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][8]  ( .D(n2068), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][9]  ( .D(n2069), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][11]  ( .D(n2071), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[6]  ( .D(n2045), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[6]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][4]  ( .D(n2076), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][5]  ( .D(n2077), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][6]  ( .D(n2078), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][7]  ( .D(n2079), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][8]  ( .D(n2080), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][9]  ( .D(n2081), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][10]  ( .D(n2082), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][11]  ( .D(n2083), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[3]  ( .D(n2048), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[3]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][4]  ( .D(n2112), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][5]  ( .D(n2113), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][6]  ( .D(n2114), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][7]  ( .D(n2115), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][8]  ( .D(n2116), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][9]  ( .D(n2117), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][10]  ( .D(n2118), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][11]  ( .D(n2119), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[2]  ( .D(n2049), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[2]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][4]  ( .D(n2124), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][5]  ( .D(n2125), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][6]  ( .D(n2126), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][7]  ( .D(n2127), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][8]  ( .D(n2128), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][9]  ( .D(n2129), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][10]  ( .D(n2130), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][11]  ( .D(n2131), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][11] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][0]  ( .D(n2038), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][1]  ( .D(n2039), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][2]  ( .D(n2040), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][3]  ( .D(n2041), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][4]  ( .D(n2042), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][5]  ( .D(n2043), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][0]  ( .D(n2032), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][1]  ( .D(n2033), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][2]  ( .D(n2034), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][3]  ( .D(n2035), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][4]  ( .D(n2036), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][5]  ( .D(n2037), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][0]  ( .D(n2014), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][1]  ( .D(n2015), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][2]  ( .D(n2016), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][3]  ( .D(n2017), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][4]  ( .D(n2018), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][5]  ( .D(n2019), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][0]  ( .D(n2008), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][1]  ( .D(n2009), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][2]  ( .D(n2010), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][3]  ( .D(n2011), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][4]  ( .D(n2012), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][5]  ( .D(n2013), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][5] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[5][0]  ( .D(n1972), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[5][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[5][1]  ( .D(n1973), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[5][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[5][2]  ( .D(n1974), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[5][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[5][3]  ( .D(n1975), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[5][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][0]  ( .D(n2084), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][1]  ( .D(n2085), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][2]  ( .D(n2086), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][3]  ( .D(n2087), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[4][0]  ( .D(n1976), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[4][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[4][1]  ( .D(n1977), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[4][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[4][2]  ( .D(n1978), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[4][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[4][3]  ( .D(n1979), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[4][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][0]  ( .D(n2096), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][1]  ( .D(n2097), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][2]  ( .D(n2098), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][3]  ( .D(n2099), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[1][0]  ( .D(n1988), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[1][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[1][1]  ( .D(n1989), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[1][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[1][2]  ( .D(n1990), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[1][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[1][3]  ( .D(n1991), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[1][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][0]  ( .D(n2132), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][1]  ( .D(n2133), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][2]  ( .D(n2134), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][3]  ( .D(n2135), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[0][0]  ( .D(n1992), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[0][1]  ( .D(n1993), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[0][2]  ( .D(n1994), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[0][3]  ( .D(n1995), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][0]  ( .D(n2144), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][1]  ( .D(n2145), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][2]  ( .D(n2146), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][3]  ( .D(n2147), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][0]  ( .D(n2026), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][1]  ( .D(n2027), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][2]  ( .D(n2028), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][3]  ( .D(n2029), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][4]  ( .D(n2030), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][5]  ( .D(n2031), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][0]  ( .D(n2020), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][1]  ( .D(n2021), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][2]  ( .D(n2022), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][3]  ( .D(n2023), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][4]  ( .D(n2024), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][5]  ( .D(n2025), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][0]  ( .D(n2002), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][1]  ( .D(n2003), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][2]  ( .D(n2004), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][3]  ( .D(n2005), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][4]  ( .D(n2006), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][5]  ( .D(n2007), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][5] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[7][0]  ( .D(n1964), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[7][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[7][1]  ( .D(n1965), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[7][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[7][2]  ( .D(n1966), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[7][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[7][3]  ( .D(n1967), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[7][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][0]  ( .D(n2060), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][1]  ( .D(n2061), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][2]  ( .D(n2062), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][3]  ( .D(n2063), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[6][0]  ( .D(n1968), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[6][1]  ( .D(n1969), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[6][2]  ( .D(n1970), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[6][3]  ( .D(n1971), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][0]  ( .D(n2072), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][1]  ( .D(n2073), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][2]  ( .D(n2074), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][3]  ( .D(n2075), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[3][0]  ( .D(n1980), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[3][1]  ( .D(n1981), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[3][2]  ( .D(n1982), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[3][3]  ( .D(n1983), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][0]  ( .D(n2108), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][1]  ( .D(n2109), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][2]  ( .D(n2110), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][3]  ( .D(n2111), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][3] ) );
  DFFNSRX1TS \writeOutbuffer_reg[5]  ( .D(n2046), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[5]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][4]  ( .D(n2088), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][5]  ( .D(n2089), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][6]  ( .D(n2090), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][7]  ( .D(n2091), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][8]  ( .D(n2092), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][9]  ( .D(n2093), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][10]  ( .D(n2094), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][11]  ( .D(n2095), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[4]  ( .D(n2047), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[4]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][4]  ( .D(n2100), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][5]  ( .D(n2101), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][6]  ( .D(n2102), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][7]  ( .D(n2103), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][8]  ( .D(n2104), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][9]  ( .D(n2105), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][10]  ( .D(n2106), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][11]  ( .D(n2107), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[1]  ( .D(n2050), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[1]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][4]  ( .D(n2136), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][5]  ( .D(n2137), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][6]  ( .D(n2138), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][7]  ( .D(n2139), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][8]  ( .D(n2140), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][9]  ( .D(n2141), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][10]  ( .D(n2142), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][11]  ( .D(n2143), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[0]  ( .D(n2051), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[0]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][4]  ( .D(n2148), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][5]  ( .D(n2149), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][6]  ( .D(n2150), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][7]  ( .D(n2151), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][8]  ( .D(n2152), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][9]  ( .D(n2153), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][10]  ( .D(n2154), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][11]  ( .D(n2155), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][11] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][10]  ( .D(n2070), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][10] ) );
  DFFNSRX1TS writeOut_reg ( .D(n1941), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        writeOut) );
  DFFNSRX1TS \destinationAddressOut_reg[4]  ( .D(n1950), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[4]) );
  DFFNSRX1TS \destinationAddressOut_reg[5]  ( .D(n1951), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[5]) );
  DFFNSRX1TS \destinationAddressOut_reg[6]  ( .D(n1952), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[6]) );
  DFFNSRX1TS \destinationAddressOut_reg[7]  ( .D(n1953), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[7]) );
  DFFNSRX1TS \destinationAddressOut_reg[8]  ( .D(n1954), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[8]) );
  DFFNSRX1TS \destinationAddressOut_reg[9]  ( .D(n1955), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[9]) );
  DFFNSRX1TS \destinationAddressOut_reg[10]  ( .D(n1956), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[10]) );
  DFFNSRX1TS \destinationAddressOut_reg[11]  ( .D(n1957), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[11]) );
  DFFNSRX1TS readOut_reg ( .D(n1940), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        readOut) );
  DFFNSRX1TS \requesterAddressOut_reg[0]  ( .D(n1942), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[0]) );
  DFFNSRX1TS \requesterAddressOut_reg[1]  ( .D(n1943), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[1]) );
  DFFNSRX1TS \requesterAddressOut_reg[2]  ( .D(n1944), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[2]) );
  DFFNSRX1TS \requesterAddressOut_reg[3]  ( .D(n1945), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[3]) );
  DFFNSRX1TS \destinationAddressOut_reg[0]  ( .D(n1946), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[0]) );
  DFFNSRX1TS \destinationAddressOut_reg[1]  ( .D(n1947), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[1]) );
  DFFNSRX1TS \destinationAddressOut_reg[2]  ( .D(n1948), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[2]) );
  DFFNSRX1TS \destinationAddressOut_reg[3]  ( .D(n1949), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[3]) );
  DFFNSRX1TS \dataOut_reg[0]  ( .D(n1958), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[0]) );
  DFFNSRX1TS \dataOut_reg[1]  ( .D(n1959), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[1]) );
  DFFNSRX1TS \dataOut_reg[2]  ( .D(n1960), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[2]) );
  DFFNSRX1TS \dataOut_reg[3]  ( .D(n1961), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[3]) );
  DFFNSRX1TS \dataOut_reg[4]  ( .D(n1962), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[4]) );
  DFFNSRX1TS \dataOut_reg[5]  ( .D(n1963), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[5]) );
  DFFNSRX1TS \read_reg_reg[1]  ( .D(n1939), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1917), .QN(n1916) );
  DFFNSRX1TS \write_reg_reg[0]  ( .D(n1934), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1915), .QN(n1919) );
  DFFNSRX1TS \write_reg_reg[2]  ( .D(n1936), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1920), .QN(n1921) );
  DFFNSRX1TS \read_reg_reg[0]  ( .D(n1933), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1910), .QN(n1922) );
  DFFNSRX1TS \read_reg_reg[2]  ( .D(n1938), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1913), .QN(n1914) );
  DFFNSRX1TS empty_reg_reg ( .D(n1937), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        n1912), .QN(n1911) );
  DFFNSRX1TS \readOutbuffer_reg[0]  ( .D(n2059), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[0]), .QN(n1932) );
  DFFNSRX1TS \readOutbuffer_reg[3]  ( .D(n2056), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[3]), .QN(n1929) );
  DFFNSRX1TS \readOutbuffer_reg[7]  ( .D(n2052), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[7]), .QN(n1925) );
  DFFNSRX1TS \readOutbuffer_reg[1]  ( .D(n2058), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[1]), .QN(n1931) );
  DFFNSRX1TS \readOutbuffer_reg[2]  ( .D(n2057), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[2]), .QN(n1930) );
  DFFNSRX1TS \readOutbuffer_reg[4]  ( .D(n2055), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[4]), .QN(n1928) );
  DFFNSRX1TS \readOutbuffer_reg[6]  ( .D(n2053), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[6]), .QN(n1926) );
  DFFNSRX1TS \readOutbuffer_reg[5]  ( .D(n2054), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[5]), .QN(n1927) );
  DFFNSRX1TS \write_reg_reg[1]  ( .D(n1935), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1918), .QN(n1923) );
  XNOR2X2TS U3 ( .A(n479), .B(n478), .Y(n480) );
  CLKBUFX2TS U4 ( .A(n14), .Y(n82) );
  CMPR32X2TS U5 ( .A(n530), .B(n461), .C(n460), .CO(n452), .S(n466) );
  CLKBUFX2TS U6 ( .A(n20), .Y(n84) );
  CMPR32X2TS U7 ( .A(selectBit_SOUTH), .B(selectBit_NORTH), .C(selectBit_EAST), 
        .CO(n463), .S(n458) );
  OR2X1TS U8 ( .A(n21), .B(n507), .Y(n8) );
  INVX2TS U9 ( .A(n22), .Y(n130) );
  OAI31X1TS U10 ( .A0(n516), .A1(n515), .A2(n537), .B0(n538), .Y(n518) );
  NOR3XLTS U11 ( .A(n29), .B(n85), .C(n8), .Y(n1609) );
  NOR3XLTS U12 ( .A(n29), .B(n84), .C(n19), .Y(n1596) );
  NOR2XLTS U13 ( .A(n1551), .B(n1548), .Y(n36) );
  NOR2XLTS U14 ( .A(n129), .B(n385), .Y(n1589) );
  NAND2X1TS U15 ( .A(n538), .B(n520), .Y(n509) );
  NOR2XLTS U16 ( .A(n839), .B(n517), .Y(n543) );
  NOR2XLTS U17 ( .A(n839), .B(n519), .Y(n688) );
  INVX2TS U18 ( .A(n1580), .Y(n1578) );
  INVX2TS U19 ( .A(n1599), .Y(n1597) );
  INVX2TS U20 ( .A(n1555), .Y(n1554) );
  INVX2TS U21 ( .A(n1548), .Y(n1546) );
  INVX2TS U22 ( .A(n1628), .Y(n1625) );
  NOR3XLTS U23 ( .A(n14), .B(n81), .C(n271), .Y(n1573) );
  INVX2TS U24 ( .A(n1602), .Y(n1600) );
  AOI31XLTS U25 ( .A0(n134), .A1(n27), .A2(n132), .B0(n316), .Y(n137) );
  INVX2TS U26 ( .A(n1632), .Y(n1629) );
  NOR2XLTS U27 ( .A(n1544), .B(n38), .Y(n46) );
  NOR2XLTS U28 ( .A(n1606), .B(n324), .Y(n325) );
  NOR2XLTS U29 ( .A(n449), .B(n1585), .Y(n277) );
  NOR2XLTS U30 ( .A(n1567), .B(n231), .Y(n230) );
  NOR2XLTS U31 ( .A(n440), .B(n1593), .Y(n136) );
  NOR2XLTS U32 ( .A(n226), .B(n1562), .Y(n88) );
  NOR2XLTS U33 ( .A(n1552), .B(n316), .Y(n34) );
  NOR2XLTS U34 ( .A(n1590), .B(n140), .Y(n141) );
  NOR2XLTS U35 ( .A(n1554), .B(n94), .Y(n95) );
  NOR3XLTS U36 ( .A(n1551), .B(n1546), .C(n37), .Y(n32) );
  NOR2XLTS U37 ( .A(n316), .B(n1603), .Y(n185) );
  NOR2XLTS U38 ( .A(n1595), .B(n189), .Y(n190) );
  INVX2TS U39 ( .A(n440), .Y(n389) );
  INVX2TS U40 ( .A(n276), .Y(n1402) );
  NOR2X1TS U41 ( .A(n1596), .B(n189), .Y(n193) );
  NOR2X1TS U42 ( .A(n1609), .B(n324), .Y(n346) );
  NAND2BX1TS U43 ( .AN(n140), .B(n134), .Y(n138) );
  NAND2BXLTS U44 ( .AN(n281), .B(n280), .Y(n283) );
  NAND2BXLTS U45 ( .AN(n397), .B(n396), .Y(n398) );
  NAND2BXLTS U46 ( .AN(n92), .B(n91), .Y(n94) );
  NOR3X1TS U47 ( .A(n1561), .B(n1556), .C(n92), .Y(n87) );
  NAND2BX1TS U48 ( .AN(n37), .B(n36), .Y(n38) );
  AOI31X1TS U49 ( .A0(n228), .A1(n1564), .A2(n224), .B0(n440), .Y(n227) );
  AOI31X1TS U50 ( .A0(n36), .A1(n31), .A2(n1544), .B0(n226), .Y(n35) );
  NOR2X1TS U51 ( .A(n1592), .B(n1589), .Y(n134) );
  INVX1TS U52 ( .A(n1570), .Y(n1568) );
  INVX1TS U53 ( .A(n1558), .Y(n1556) );
  INVX1TS U54 ( .A(n1613), .Y(n1610) );
  NOR2X1TS U55 ( .A(n129), .B(n273), .Y(n1548) );
  ADDFX1TS U56 ( .A(n485), .B(n484), .CI(n483), .CO(n478), .S(n494) );
  NAND3X1TS U57 ( .A(n29), .B(n223), .C(n19), .Y(n1564) );
  NAND3X1TS U58 ( .A(n484), .B(n29), .C(n223), .Y(n1544) );
  INVX1TS U59 ( .A(n1577), .Y(n1576) );
  INVX1TS U60 ( .A(n1561), .Y(n1559) );
  INVX1TS U61 ( .A(n1592), .Y(n1590) );
  NOR2X1TS U62 ( .A(n223), .B(n83), .Y(n313) );
  OAI21X1TS U63 ( .A0(selectBit_SOUTH), .A1(n21), .B0(n84), .Y(n272) );
  NOR3X1TS U64 ( .A(n24), .B(n85), .C(n20), .Y(n1624) );
  NOR3X1TS U65 ( .A(n126), .B(n182), .C(n271), .Y(n1561) );
  INVX1TS U66 ( .A(n1617), .Y(n1614) );
  NOR2X1TS U67 ( .A(selectBit_NORTH), .B(n505), .Y(n538) );
  ADDFX1TS U68 ( .A(n463), .B(n484), .CI(n16), .CO(n17), .S(n14) );
  CLKBUFX2TS U69 ( .A(n56), .Y(n297) );
  OR2X2TS U70 ( .A(n457), .B(n504), .Y(n2) );
  CLKBUFX2TS U71 ( .A(readIn_EAST), .Y(n1543) );
  INVX1TS U72 ( .A(n1921), .Y(n275) );
  CLKINVX1TS U73 ( .A(n1584), .Y(n1581) );
  NAND2X2TS U74 ( .A(n127), .B(n506), .Y(n271) );
  CMPR22X2TS U75 ( .A(n446), .B(n458), .CO(n16), .S(n15) );
  OAI21X1TS U76 ( .A0(n315), .A1(n495), .B0(n22), .Y(n19) );
  NOR2X1TS U77 ( .A(n26), .B(n138), .Y(n135) );
  INVX2TS U78 ( .A(selectBit_NORTH), .Y(n504) );
  NOR2XLTS U79 ( .A(n1632), .B(n1628), .Y(n396) );
  NOR2XLTS U80 ( .A(n1617), .B(n1613), .Y(n321) );
  NOR2XLTS U81 ( .A(n1602), .B(n1599), .Y(n187) );
  NAND2BX1TS U82 ( .AN(n322), .B(n321), .Y(n324) );
  INVX2TS U83 ( .A(n230), .Y(n256) );
  NAND2X1TS U84 ( .A(n137), .B(n1593), .Y(n140) );
  NAND2BX1TS U85 ( .AN(n188), .B(n187), .Y(n189) );
  NAND4XLTS U86 ( .A(n444), .B(n451), .C(n513), .D(n392), .Y(n1562) );
  NAND4XLTS U87 ( .A(n275), .B(n511), .C(n392), .D(n387), .Y(n1585) );
  NOR3XLTS U88 ( .A(n82), .B(n15), .C(n271), .Y(n1584) );
  NAND4XLTS U89 ( .A(n495), .B(n510), .C(n392), .D(n441), .Y(n1603) );
  NOR3X1TS U90 ( .A(n15), .B(n182), .C(n383), .Y(n1602) );
  INVX2TS U91 ( .A(n1596), .Y(n1595) );
  NOR3X1TS U92 ( .A(n82), .B(n81), .C(n383), .Y(n1617) );
  INVX2TS U93 ( .A(n1609), .Y(n1606) );
  NAND4XLTS U94 ( .A(n1915), .B(n455), .C(n451), .D(n511), .Y(n1552) );
  NAND4XLTS U95 ( .A(n455), .B(n1915), .C(n510), .D(n443), .Y(n1593) );
  NOR3X1TS U96 ( .A(n82), .B(n15), .C(n383), .Y(n1632) );
  CLKAND2X2TS U97 ( .A(n523), .B(n521), .Y(n550) );
  CLKAND2X2TS U98 ( .A(n477), .B(n475), .Y(n482) );
  NOR2XLTS U99 ( .A(reset), .B(n449), .Y(n497) );
  NOR2XLTS U100 ( .A(n1584), .B(n1580), .Y(n280) );
  AO21X2TS U101 ( .A0(n457), .A1(n504), .B0(n315), .Y(n21) );
  OAI21XLTS U102 ( .A0(n28), .A1(n25), .B0(n27), .Y(n128) );
  NOR3BXLTS U103 ( .AN(readReady), .B(selectBit_WEST), .C(n514), .Y(n537) );
  NAND3XLTS U104 ( .A(n505), .B(n508), .C(n504), .Y(n517) );
  NAND3XLTS U105 ( .A(selectBit_NORTH), .B(n508), .C(n507), .Y(n519) );
  AOI21X1TS U106 ( .A0(n321), .A1(n317), .B0(n316), .Y(n319) );
  NOR2XLTS U107 ( .A(n1573), .B(n1570), .Y(n228) );
  NOR2XLTS U108 ( .A(n1561), .B(n1558), .Y(n91) );
  AOI21X1TS U109 ( .A0(n187), .A1(n183), .B0(n226), .Y(n186) );
  AOI21X1TS U110 ( .A0(n396), .A1(n390), .B0(n30), .Y(n394) );
  XOR2XLTS U111 ( .A(n452), .B(n454), .Y(n472) );
  OAI21XLTS U112 ( .A0(n455), .A1(n1916), .B0(n454), .Y(n456) );
  NAND3XLTS U113 ( .A(n315), .B(n479), .C(n387), .Y(n224) );
  XOR2X1TS U114 ( .A(n275), .B(n17), .Y(n127) );
  NOR2X1TS U115 ( .A(n8), .B(n83), .Y(n28) );
  NAND2BX1TS U116 ( .AN(n127), .B(n506), .Y(n383) );
  NAND2BX1TS U117 ( .AN(n128), .B(n514), .Y(n385) );
  CLKAND2X2TS U118 ( .A(n477), .B(n476), .Y(n483) );
  NOR2XLTS U119 ( .A(n389), .B(reset), .Y(n498) );
  NAND4XLTS U120 ( .A(n493), .B(n275), .C(readReady), .D(n391), .Y(n1574) );
  INVX2TS U121 ( .A(n1573), .Y(n1571) );
  NOR3XLTS U122 ( .A(n314), .B(n313), .C(n273), .Y(n1570) );
  NOR3XLTS U123 ( .A(n85), .B(n84), .C(n23), .Y(n1577) );
  NOR3BXLTS U124 ( .AN(n386), .B(n273), .C(n272), .Y(n1580) );
  NAND4XLTS U125 ( .A(n493), .B(n510), .C(n450), .D(n391), .Y(n1618) );
  NOR3XLTS U126 ( .A(n314), .B(n313), .C(n385), .Y(n1613) );
  NAND4XLTS U127 ( .A(n14), .B(n126), .C(n127), .D(n459), .Y(n1549) );
  INVX2TS U128 ( .A(n1544), .Y(n1545) );
  NOR3X1TS U129 ( .A(n182), .B(n81), .C(n383), .Y(n1592) );
  INVX2TS U130 ( .A(n1589), .Y(n1587) );
  NAND4XLTS U131 ( .A(n511), .B(n392), .C(n391), .D(n443), .Y(n1633) );
  INVX2TS U132 ( .A(n1624), .Y(n1621) );
  NOR3BXLTS U133 ( .AN(n386), .B(n385), .C(n384), .Y(n1628) );
  INVX2TS U134 ( .A(destinationAddressIn_SOUTH[11]), .Y(n164) );
  INVX2TS U135 ( .A(destinationAddressIn_SOUTH[10]), .Y(n171) );
  INVX2TS U136 ( .A(destinationAddressIn_SOUTH[9]), .Y(n176) );
  INVX2TS U137 ( .A(destinationAddressIn_SOUTH[8]), .Y(n167) );
  AO22XLTS U138 ( .A0(n1920), .A1(n498), .B0(n497), .B1(n496), .Y(n1936) );
  AO22XLTS U139 ( .A0(n493), .A1(n498), .B0(n497), .B1(n492), .Y(n1934) );
  AO22XLTS U140 ( .A0(n495), .A1(n498), .B0(n497), .B1(n494), .Y(n1935) );
  OAI21XLTS U141 ( .A0(n389), .A1(n448), .B0(n491), .Y(n1937) );
  NAND4XLTS U142 ( .A(n865), .B(n864), .C(n863), .D(n862), .Y(n1963) );
  NAND4XLTS U143 ( .A(n843), .B(n842), .C(n841), .D(n862), .Y(n1962) );
  NAND4XLTS U144 ( .A(n832), .B(n831), .C(n830), .D(n862), .Y(n1961) );
  NAND4XLTS U145 ( .A(n822), .B(n821), .C(n820), .D(n862), .Y(n1960) );
  NAND4XLTS U146 ( .A(n803), .B(n802), .C(n801), .D(n800), .Y(n1959) );
  NAND4XLTS U147 ( .A(n783), .B(n782), .C(n781), .D(n800), .Y(n1958) );
  NAND4XLTS U148 ( .A(n654), .B(n653), .C(n652), .D(n651), .Y(n1949) );
  NAND4XLTS U149 ( .A(n643), .B(n642), .C(n641), .D(n640), .Y(n1948) );
  NAND4XLTS U150 ( .A(n625), .B(n624), .C(n623), .D(n622), .Y(n1947) );
  NAND4XLTS U151 ( .A(n610), .B(n609), .C(n608), .D(n607), .Y(n1946) );
  NAND4XLTS U152 ( .A(n598), .B(n597), .C(n596), .D(n651), .Y(n1945) );
  NAND4XLTS U153 ( .A(n587), .B(n586), .C(n585), .D(n640), .Y(n1944) );
  NAND4XLTS U154 ( .A(n578), .B(n577), .C(n576), .D(n622), .Y(n1943) );
  NAND4XLTS U155 ( .A(n561), .B(n560), .C(n559), .D(n607), .Y(n1942) );
  NAND4XLTS U156 ( .A(n541), .B(n540), .C(n539), .D(n800), .Y(n1940) );
  NAND3XLTS U157 ( .A(n773), .B(n772), .C(n771), .Y(n1957) );
  NAND3XLTS U158 ( .A(n759), .B(n758), .C(n757), .Y(n1956) );
  NAND3XLTS U159 ( .A(n743), .B(n742), .C(n741), .Y(n1955) );
  NAND3XLTS U160 ( .A(n725), .B(n724), .C(n723), .Y(n1954) );
  NAND3XLTS U161 ( .A(n711), .B(n710), .C(n709), .Y(n1953) );
  NAND3XLTS U162 ( .A(n700), .B(n699), .C(n698), .Y(n1952) );
  NAND3XLTS U163 ( .A(n686), .B(n685), .C(n684), .Y(n1951) );
  NAND3XLTS U164 ( .A(n665), .B(n664), .C(n663), .Y(n1950) );
  NAND3XLTS U165 ( .A(n553), .B(n552), .C(n551), .Y(n1941) );
  NAND3XLTS U166 ( .A(n1788), .B(n1787), .C(n1786), .Y(n2111) );
  NAND3XLTS U167 ( .A(n1779), .B(n1778), .C(n1777), .Y(n2110) );
  NAND3XLTS U168 ( .A(n1771), .B(n1770), .C(n1769), .Y(n2109) );
  NAND3XLTS U169 ( .A(n1765), .B(n1764), .C(n1763), .Y(n2108) );
  NAND3XLTS U170 ( .A(n977), .B(n976), .C(n975), .Y(n1983) );
  NAND3XLTS U171 ( .A(n970), .B(n969), .C(n968), .Y(n1982) );
  NAND3XLTS U172 ( .A(n962), .B(n961), .C(n960), .Y(n1981) );
  NAND3XLTS U173 ( .A(n955), .B(n954), .C(n953), .Y(n1980) );
  NAND3XLTS U174 ( .A(n1693), .B(n1692), .C(n1691), .Y(n2075) );
  NAND3XLTS U175 ( .A(n1684), .B(n1683), .C(n1682), .Y(n2074) );
  NAND3XLTS U176 ( .A(n1677), .B(n1676), .C(n1675), .Y(n2073) );
  NAND3XLTS U177 ( .A(n1670), .B(n1669), .C(n1668), .Y(n2072) );
  NAND3XLTS U178 ( .A(n900), .B(n899), .C(n898), .Y(n1971) );
  NAND3XLTS U179 ( .A(n892), .B(n891), .C(n890), .Y(n1970) );
  NAND3XLTS U180 ( .A(n889), .B(n888), .C(n887), .Y(n1969) );
  NAND3XLTS U181 ( .A(n885), .B(n884), .C(n883), .Y(n1968) );
  NAND3XLTS U182 ( .A(n1663), .B(n1662), .C(n1661), .Y(n2063) );
  NAND3XLTS U183 ( .A(n1654), .B(n1653), .C(n1652), .Y(n2062) );
  NAND3XLTS U184 ( .A(n1646), .B(n1645), .C(n1644), .Y(n2061) );
  NAND3XLTS U185 ( .A(n1639), .B(n1638), .C(n1637), .Y(n2060) );
  NAND3XLTS U186 ( .A(n882), .B(n881), .C(n880), .Y(n1967) );
  NAND3XLTS U187 ( .A(n875), .B(n874), .C(n873), .Y(n1966) );
  NAND3XLTS U188 ( .A(n872), .B(n871), .C(n870), .Y(n1965) );
  NAND3XLTS U189 ( .A(n868), .B(n867), .C(n866), .Y(n1964) );
  NAND3XLTS U190 ( .A(n1107), .B(n1106), .C(n1105), .Y(n2007) );
  NAND3XLTS U191 ( .A(n1102), .B(n1101), .C(n1100), .Y(n2006) );
  NAND3XLTS U192 ( .A(n1097), .B(n1096), .C(n1095), .Y(n2005) );
  NAND3XLTS U193 ( .A(n1092), .B(n1091), .C(n1090), .Y(n2004) );
  NAND3XLTS U194 ( .A(n1088), .B(n1087), .C(n1086), .Y(n2003) );
  NAND3XLTS U195 ( .A(n1083), .B(n1082), .C(n1081), .Y(n2002) );
  NAND3XLTS U196 ( .A(n1423), .B(n1422), .C(n1421), .Y(n2025) );
  NAND3XLTS U197 ( .A(n1418), .B(n1417), .C(n1416), .Y(n2024) );
  NAND3XLTS U198 ( .A(n1411), .B(n1410), .C(n1409), .Y(n2023) );
  NAND3XLTS U199 ( .A(n1406), .B(n1405), .C(n1404), .Y(n2022) );
  NAND3XLTS U200 ( .A(n1401), .B(n1400), .C(n1399), .Y(n2021) );
  NAND3XLTS U201 ( .A(n1397), .B(n1396), .C(n1395), .Y(n2020) );
  NAND3XLTS U202 ( .A(n1458), .B(n1457), .C(n1456), .Y(n2031) );
  NAND3XLTS U203 ( .A(n1453), .B(n1452), .C(n1451), .Y(n2030) );
  NAND3XLTS U204 ( .A(n1446), .B(n1445), .C(n1444), .Y(n2029) );
  NAND3XLTS U205 ( .A(n1441), .B(n1440), .C(n1439), .Y(n2028) );
  NAND3XLTS U206 ( .A(n1435), .B(n1434), .C(n1433), .Y(n2027) );
  NAND3XLTS U207 ( .A(n1431), .B(n1430), .C(n1429), .Y(n2026) );
  NAND3XLTS U208 ( .A(n1894), .B(n1893), .C(n1892), .Y(n2147) );
  NAND3XLTS U209 ( .A(n1883), .B(n1882), .C(n1881), .Y(n2146) );
  NAND3XLTS U210 ( .A(n1873), .B(n1872), .C(n1871), .Y(n2145) );
  NAND3XLTS U211 ( .A(n1864), .B(n1863), .C(n1862), .Y(n2144) );
  NAND3XLTS U212 ( .A(n1051), .B(n1050), .C(n1049), .Y(n1995) );
  NAND3XLTS U213 ( .A(n1042), .B(n1041), .C(n1040), .Y(n1994) );
  NAND3XLTS U214 ( .A(n1037), .B(n1036), .C(n1035), .Y(n1993) );
  NAND3XLTS U215 ( .A(n1030), .B(n1029), .C(n1028), .Y(n1992) );
  NAND3XLTS U216 ( .A(n1854), .B(n1853), .C(n1852), .Y(n2135) );
  NAND3XLTS U217 ( .A(n1843), .B(n1842), .C(n1841), .Y(n2134) );
  NAND3XLTS U218 ( .A(n1832), .B(n1831), .C(n1830), .Y(n2133) );
  NAND3XLTS U219 ( .A(n1822), .B(n1821), .C(n1820), .Y(n2132) );
  NAND3XLTS U220 ( .A(n1025), .B(n1024), .C(n1023), .Y(n1991) );
  NAND3XLTS U221 ( .A(n1016), .B(n1015), .C(n1014), .Y(n1990) );
  NAND3XLTS U222 ( .A(n1009), .B(n1008), .C(n1007), .Y(n1989) );
  NAND3XLTS U223 ( .A(n1002), .B(n1001), .C(n1000), .Y(n1988) );
  NAND3XLTS U224 ( .A(n1756), .B(n1755), .C(n1754), .Y(n2099) );
  NAND3XLTS U225 ( .A(n1747), .B(n1746), .C(n1745), .Y(n2098) );
  NAND3XLTS U226 ( .A(n1740), .B(n1739), .C(n1738), .Y(n2097) );
  NAND3XLTS U227 ( .A(n1734), .B(n1733), .C(n1732), .Y(n2096) );
  NAND3XLTS U228 ( .A(n947), .B(n946), .C(n945), .Y(n1979) );
  NAND3XLTS U229 ( .A(n936), .B(n935), .C(n934), .Y(n1978) );
  NAND3XLTS U230 ( .A(n930), .B(n929), .C(n928), .Y(n1977) );
  NAND3XLTS U231 ( .A(n924), .B(n923), .C(n922), .Y(n1976) );
  NAND3XLTS U232 ( .A(n1727), .B(n1726), .C(n1725), .Y(n2087) );
  NAND3XLTS U233 ( .A(n1718), .B(n1717), .C(n1716), .Y(n2086) );
  NAND3XLTS U234 ( .A(n1710), .B(n1709), .C(n1708), .Y(n2085) );
  NAND3XLTS U235 ( .A(n1702), .B(n1701), .C(n1700), .Y(n2084) );
  NAND3XLTS U236 ( .A(n917), .B(n916), .C(n915), .Y(n1975) );
  NAND3XLTS U237 ( .A(n911), .B(n910), .C(n909), .Y(n1974) );
  NAND3XLTS U238 ( .A(n907), .B(n906), .C(n905), .Y(n1973) );
  NAND3XLTS U239 ( .A(n904), .B(n903), .C(n902), .Y(n1972) );
  NAND3XLTS U240 ( .A(n1365), .B(n1364), .C(n1363), .Y(n2013) );
  NAND3XLTS U241 ( .A(n1359), .B(n1358), .C(n1357), .Y(n2012) );
  NAND3XLTS U242 ( .A(n1354), .B(n1353), .C(n1352), .Y(n2011) );
  NAND3XLTS U243 ( .A(n1348), .B(n1347), .C(n1346), .Y(n2010) );
  NAND3XLTS U244 ( .A(n1343), .B(n1342), .C(n1341), .Y(n2009) );
  NAND3XLTS U245 ( .A(n1338), .B(n1337), .C(n1112), .Y(n2008) );
  NAND3XLTS U246 ( .A(n1390), .B(n1389), .C(n1388), .Y(n2019) );
  NAND3XLTS U247 ( .A(n1385), .B(n1384), .C(n1383), .Y(n2018) );
  NAND3XLTS U248 ( .A(n1380), .B(n1379), .C(n1378), .Y(n2017) );
  NAND3XLTS U249 ( .A(n1376), .B(n1375), .C(n1374), .Y(n2016) );
  NAND3XLTS U250 ( .A(n1372), .B(n1371), .C(n1370), .Y(n2015) );
  NAND3XLTS U251 ( .A(n1369), .B(n1368), .C(n1367), .Y(n2014) );
  NAND3XLTS U252 ( .A(n1497), .B(n1496), .C(n1495), .Y(n2037) );
  NAND3XLTS U253 ( .A(n1491), .B(n1490), .C(n1489), .Y(n2036) );
  NAND3XLTS U254 ( .A(n1484), .B(n1483), .C(n1482), .Y(n2035) );
  NAND3XLTS U255 ( .A(n1478), .B(n1477), .C(n1476), .Y(n2034) );
  NAND3XLTS U256 ( .A(n1472), .B(n1471), .C(n1470), .Y(n2033) );
  NAND3XLTS U257 ( .A(n1467), .B(n1466), .C(n1465), .Y(n2032) );
  NAND3XLTS U258 ( .A(n1542), .B(n1541), .C(n1540), .Y(n2043) );
  NAND3XLTS U259 ( .A(n1534), .B(n1533), .C(n1532), .Y(n2042) );
  NAND3XLTS U260 ( .A(n1526), .B(n1525), .C(n1524), .Y(n2041) );
  NAND3XLTS U261 ( .A(n1518), .B(n1517), .C(n1516), .Y(n2040) );
  NAND3XLTS U262 ( .A(n1512), .B(n1511), .C(n1510), .Y(n2039) );
  NAND3XLTS U263 ( .A(n1504), .B(n1503), .C(n1502), .Y(n2038) );
  NAND3XLTS U264 ( .A(n1813), .B(n1812), .C(n1811), .Y(n2123) );
  NAND3XLTS U265 ( .A(n1807), .B(n1806), .C(n1805), .Y(n2122) );
  NAND3XLTS U266 ( .A(n1800), .B(n1799), .C(n1798), .Y(n2121) );
  NAND3XLTS U267 ( .A(n1794), .B(n1793), .C(n1792), .Y(n2120) );
  NAND3XLTS U268 ( .A(n995), .B(n994), .C(n993), .Y(n1987) );
  NAND3XLTS U269 ( .A(n988), .B(n987), .C(n986), .Y(n1986) );
  NAND3XLTS U270 ( .A(n984), .B(n983), .C(n982), .Y(n1985) );
  NAND3XLTS U271 ( .A(n980), .B(n979), .C(n978), .Y(n1984) );
  NAND3XLTS U272 ( .A(n1077), .B(n1076), .C(n1075), .Y(n2001) );
  NAND3XLTS U273 ( .A(n1073), .B(n1072), .C(n1071), .Y(n2000) );
  NAND3XLTS U274 ( .A(n1068), .B(n1067), .C(n1066), .Y(n1999) );
  NAND3XLTS U275 ( .A(n1064), .B(n1063), .C(n1062), .Y(n1998) );
  NAND3XLTS U276 ( .A(n1060), .B(n1059), .C(n1058), .Y(n1997) );
  NAND3XLTS U277 ( .A(n1056), .B(n1055), .C(n1054), .Y(n1996) );
  AOI211XLTS U278 ( .A0(n489), .A1(n525), .B0(n488), .C0(n487), .Y(n490) );
  XOR2XLTS U279 ( .A(n524), .B(n492), .Y(n488) );
  OR2X1TS U280 ( .A(n35), .B(n1635), .Y(n1498) );
  OR2X1TS U281 ( .A(n186), .B(n1789), .Y(n981) );
  OR2X1TS U282 ( .A(n394), .B(n1855), .Y(n1031) );
  OR2X1TS U283 ( .A(n137), .B(n1757), .Y(n1366) );
  OR2X1TS U284 ( .A(n278), .B(n1728), .Y(n1391) );
  OR2X1TS U285 ( .A(n89), .B(n1664), .Y(n1459) );
  NAND2X1TS U286 ( .A(n28), .B(n25), .Y(n26) );
  NAND2X1TS U287 ( .A(n523), .B(n1924), .Y(n30) );
  OR3X1TS U288 ( .A(n1592), .B(n1587), .C(n140), .Y(n3) );
  OR2X1TS U289 ( .A(n1576), .B(n283), .Y(n4) );
  OR2X1TS U290 ( .A(n1577), .B(n283), .Y(n5) );
  OR2X1TS U291 ( .A(n1624), .B(n398), .Y(n6) );
  OR2X1TS U292 ( .A(n1555), .B(n94), .Y(n7) );
  OR2X1TS U293 ( .A(n226), .B(n1574), .Y(n9) );
  OR2X1TS U294 ( .A(n1621), .B(n398), .Y(n10) );
  OR2X1TS U295 ( .A(n227), .B(n1694), .Y(n1424) );
  NOR3XLTS U296 ( .A(n1573), .B(n1568), .C(n229), .Y(n225) );
  NOR3XLTS U297 ( .A(n1584), .B(n1578), .C(n281), .Y(n276) );
  NOR3XLTS U298 ( .A(n1602), .B(n1597), .C(n188), .Y(n184) );
  NOR3XLTS U299 ( .A(n1617), .B(n1610), .C(n322), .Y(n318) );
  NOR3XLTS U300 ( .A(n1632), .B(n1625), .C(n397), .Y(n393) );
  INVX2TS U301 ( .A(n25), .Y(n29) );
  OR2X1TS U302 ( .A(n30), .B(n1633), .Y(n11) );
  AND3X1TS U303 ( .A(n538), .B(n1912), .C(n537), .Y(n12) );
  INVX2TS U304 ( .A(destinationAddressIn_EAST[9]), .Y(n45) );
  INVX2TS U305 ( .A(destinationAddressIn_EAST[11]), .Y(n49) );
  INVX2TS U306 ( .A(destinationAddressIn_EAST[10]), .Y(n41) );
  INVX2TS U307 ( .A(destinationAddressIn_EAST[8]), .Y(n33) );
  INVX2TS U308 ( .A(writeIn_EAST), .Y(n56) );
  INVX2TS U309 ( .A(destinationAddressIn_EAST[5]), .Y(n71) );
  INVX2TS U310 ( .A(destinationAddressIn_EAST[6]), .Y(n66) );
  INVX2TS U311 ( .A(destinationAddressIn_EAST[4]), .Y(n75) );
  INVX2TS U312 ( .A(destinationAddressIn_EAST[7]), .Y(n62) );
  CLKBUFX2TS U313 ( .A(n1916), .Y(n13) );
  INVX2TS U329 ( .A(n1923), .Y(n484) );
  INVX2TS U330 ( .A(n1919), .Y(n446) );
  INVX2TS U331 ( .A(n15), .Y(n81) );
  INVX2TS U332 ( .A(n81), .Y(n126) );
  INVX2TS U333 ( .A(selectBit_WEST), .Y(n453) );
  INVX2TS U334 ( .A(n1549), .Y(n1551) );
  INVX2TS U335 ( .A(n1915), .Y(n457) );
  INVX2TS U336 ( .A(n2), .Y(n315) );
  INVX2TS U337 ( .A(selectBit_SOUTH), .Y(n507) );
  INVX2TS U338 ( .A(n8), .Y(n223) );
  INVX2TS U339 ( .A(n1923), .Y(n495) );
  INVX2TS U340 ( .A(n2), .Y(n18) );
  INVX2TS U341 ( .A(n1923), .Y(n444) );
  NAND2X1TS U342 ( .A(n18), .B(n444), .Y(n22) );
  INVX2TS U343 ( .A(n19), .Y(n85) );
  INVX2TS U344 ( .A(n85), .Y(n83) );
  NAND2X1TS U345 ( .A(selectBit_SOUTH), .B(n21), .Y(n20) );
  NAND2X1TS U346 ( .A(n313), .B(n272), .Y(n129) );
  INVX2TS U347 ( .A(n1921), .Y(n479) );
  INVX2TS U348 ( .A(n1920), .Y(n450) );
  AOI22X1TS U349 ( .A0(n479), .A1(n22), .B0(n130), .B1(n450), .Y(n23) );
  INVX2TS U350 ( .A(n23), .Y(n24) );
  INVX2TS U351 ( .A(n24), .Y(n25) );
  INVX2TS U352 ( .A(n26), .Y(n125) );
  INVX2TS U353 ( .A(n125), .Y(n27) );
  NAND2X1TS U354 ( .A(selectBit_EAST), .B(n128), .Y(n273) );
  NAND2X1TS U355 ( .A(n479), .B(n130), .Y(n31) );
  INVX2TS U356 ( .A(n507), .Y(n505) );
  INVX2TS U357 ( .A(n453), .Y(n506) );
  INVX2TS U358 ( .A(readReady), .Y(n133) );
  INVX2TS U359 ( .A(n133), .Y(n513) );
  NOR3XLTS U360 ( .A(n506), .B(selectBit_EAST), .C(n513), .Y(n508) );
  NAND2X1TS U361 ( .A(n538), .B(n508), .Y(n523) );
  INVX2TS U362 ( .A(n30), .Y(n131) );
  INVX2TS U363 ( .A(n131), .Y(n226) );
  INVX2TS U364 ( .A(n1923), .Y(n455) );
  INVX2TS U365 ( .A(n133), .Y(n511) );
  NAND2X1TS U366 ( .A(n35), .B(n1552), .Y(n37) );
  INVX2TS U367 ( .A(n32), .Y(n878) );
  INVX2TS U368 ( .A(n878), .Y(n1649) );
  CLKBUFX2TS U369 ( .A(n1649), .Y(n44) );
  INVX2TS U370 ( .A(n44), .Y(n70) );
  INVX2TS U371 ( .A(destinationAddressIn_EAST[8]), .Y(n240) );
  INVX2TS U372 ( .A(n131), .Y(n440) );
  INVX2TS U373 ( .A(n34), .Y(n876) );
  INVX2TS U374 ( .A(n876), .Y(n1635) );
  INVX2TS U375 ( .A(n1498), .Y(n52) );
  OR2X1TS U376 ( .A(n1549), .B(n37), .Y(n50) );
  INVX2TS U377 ( .A(n50), .Y(n1659) );
  CLKBUFX2TS U378 ( .A(destinationAddressIn_WEST[8]), .Y(n413) );
  CLKBUFX2TS U379 ( .A(n413), .Y(n712) );
  AOI22X1TS U380 ( .A0(n52), .A1(\destinationAddressbuffer[7][8] ), .B0(n1659), 
        .B1(n712), .Y(n40) );
  INVX2TS U381 ( .A(n46), .Y(n57) );
  INVX2TS U382 ( .A(n57), .Y(n1643) );
  INVX2TS U383 ( .A(n167), .Y(n713) );
  OR2X1TS U384 ( .A(n1545), .B(n38), .Y(n59) );
  INVX2TS U385 ( .A(n59), .Y(n1530) );
  CLKBUFX2TS U386 ( .A(destinationAddressIn_NORTH[8]), .Y(n714) );
  CLKBUFX2TS U387 ( .A(n714), .Y(n334) );
  AOI22X1TS U388 ( .A0(n1643), .A1(n713), .B0(n1530), .B1(n334), .Y(n39) );
  OAI211XLTS U389 ( .A0(n70), .A1(n240), .B0(n40), .C0(n39), .Y(n2068) );
  INVX2TS U390 ( .A(destinationAddressIn_EAST[10]), .Y(n249) );
  INVX2TS U391 ( .A(n50), .Y(n1650) );
  CLKBUFX2TS U392 ( .A(destinationAddressIn_WEST[10]), .Y(n408) );
  CLKBUFX2TS U393 ( .A(n408), .Y(n744) );
  AOI22X1TS U394 ( .A0(n52), .A1(\destinationAddressbuffer[7][10] ), .B0(n1650), .B1(n744), .Y(n43) );
  INVX2TS U395 ( .A(n57), .Y(n1660) );
  INVX2TS U396 ( .A(n171), .Y(n747) );
  INVX2TS U397 ( .A(n59), .Y(n869) );
  CLKBUFX2TS U398 ( .A(destinationAddressIn_NORTH[10]), .Y(n748) );
  CLKBUFX2TS U399 ( .A(n748), .Y(n327) );
  AOI22X1TS U400 ( .A0(n1660), .A1(n747), .B0(n869), .B1(n327), .Y(n42) );
  OAI211XLTS U401 ( .A0(n70), .A1(n249), .B0(n43), .C0(n42), .Y(n2070) );
  INVX2TS U402 ( .A(n44), .Y(n80) );
  INVX2TS U403 ( .A(destinationAddressIn_EAST[9]), .Y(n244) );
  INVX2TS U404 ( .A(n50), .Y(n1528) );
  INVX2TS U405 ( .A(n1528), .Y(n1505) );
  INVX2TS U406 ( .A(n1505), .Y(n67) );
  CLKBUFX2TS U407 ( .A(destinationAddressIn_WEST[9]), .Y(n395) );
  CLKBUFX2TS U408 ( .A(n395), .Y(n727) );
  AOI22X1TS U409 ( .A0(n52), .A1(\destinationAddressbuffer[7][9] ), .B0(n67), 
        .B1(n727), .Y(n48) );
  INVX2TS U410 ( .A(n176), .Y(n728) );
  INVX2TS U411 ( .A(n1530), .Y(n1507) );
  INVX2TS U412 ( .A(n1507), .Y(n1642) );
  CLKBUFX2TS U413 ( .A(destinationAddressIn_NORTH[9]), .Y(n730) );
  CLKBUFX2TS U414 ( .A(n730), .Y(n349) );
  AOI22X1TS U415 ( .A0(n58), .A1(n728), .B0(n1642), .B1(n349), .Y(n47) );
  OAI211XLTS U416 ( .A0(n80), .A1(n244), .B0(n48), .C0(n47), .Y(n2069) );
  INVX2TS U417 ( .A(destinationAddressIn_EAST[11]), .Y(n235) );
  INVX2TS U418 ( .A(n50), .Y(n51) );
  CLKBUFX2TS U419 ( .A(destinationAddressIn_WEST[11]), .Y(n403) );
  CLKBUFX2TS U420 ( .A(n403), .Y(n760) );
  AOI22X1TS U421 ( .A0(n52), .A1(\destinationAddressbuffer[7][11] ), .B0(n51), 
        .B1(n760), .Y(n55) );
  INVX2TS U422 ( .A(n57), .Y(n1523) );
  INVX2TS U423 ( .A(n164), .Y(n763) );
  INVX2TS U424 ( .A(n59), .Y(n53) );
  INVX2TS U425 ( .A(n1507), .Y(n72) );
  CLKBUFX2TS U426 ( .A(destinationAddressIn_NORTH[11]), .Y(n764) );
  CLKBUFX2TS U427 ( .A(n764), .Y(n340) );
  AOI22X1TS U428 ( .A0(n1523), .A1(n763), .B0(n72), .B1(n340), .Y(n54) );
  OAI211XLTS U429 ( .A0(n70), .A1(n235), .B0(n55), .C0(n54), .Y(n2071) );
  CLKBUFX2TS U430 ( .A(n1498), .Y(n877) );
  INVX2TS U431 ( .A(n877), .Y(n1655) );
  AOI22X1TS U432 ( .A0(n1655), .A1(writeOutbuffer[7]), .B0(n1650), .B1(
        writeIn_WEST), .Y(n61) );
  INVX2TS U433 ( .A(n57), .Y(n58) );
  INVX2TS U434 ( .A(n58), .Y(n879) );
  INVX2TS U435 ( .A(n879), .Y(n63) );
  INVX2TS U436 ( .A(writeIn_SOUTH), .Y(n181) );
  INVX2TS U437 ( .A(n181), .Y(n544) );
  AOI22X1TS U438 ( .A0(n63), .A1(n544), .B0(n53), .B1(writeIn_NORTH), .Y(n60)
         );
  OAI211XLTS U439 ( .A0(n80), .A1(n297), .B0(n61), .C0(n60), .Y(n2044) );
  INVX2TS U440 ( .A(destinationAddressIn_EAST[7]), .Y(n259) );
  INVX2TS U441 ( .A(n877), .Y(n77) );
  AOI22X1TS U442 ( .A0(n77), .A1(\destinationAddressbuffer[7][7] ), .B0(n1659), 
        .B1(destinationAddressIn_WEST[7]), .Y(n65) );
  INVX2TS U443 ( .A(destinationAddressIn_SOUTH[7]), .Y(n154) );
  INVX2TS U444 ( .A(n154), .Y(n702) );
  AOI22X1TS U445 ( .A0(n63), .A1(n702), .B0(n53), .B1(
        destinationAddressIn_NORTH[7]), .Y(n64) );
  OAI211XLTS U446 ( .A0(n80), .A1(n259), .B0(n65), .C0(n64), .Y(n2067) );
  INVX2TS U447 ( .A(destinationAddressIn_EAST[6]), .Y(n255) );
  AOI22X1TS U448 ( .A0(n77), .A1(\destinationAddressbuffer[7][6] ), .B0(n67), 
        .B1(destinationAddressIn_WEST[6]), .Y(n69) );
  INVX2TS U449 ( .A(destinationAddressIn_SOUTH[6]), .Y(n144) );
  INVX2TS U450 ( .A(n144), .Y(n689) );
  AOI22X1TS U451 ( .A0(n1660), .A1(n689), .B0(n1642), .B1(
        destinationAddressIn_NORTH[6]), .Y(n68) );
  OAI211XLTS U452 ( .A0(n70), .A1(n255), .B0(n69), .C0(n68), .Y(n2066) );
  INVX2TS U453 ( .A(destinationAddressIn_EAST[5]), .Y(n269) );
  AOI22X1TS U454 ( .A0(n77), .A1(\destinationAddressbuffer[7][5] ), .B0(n51), 
        .B1(destinationAddressIn_WEST[5]), .Y(n74) );
  INVX2TS U455 ( .A(destinationAddressIn_SOUTH[5]), .Y(n160) );
  INVX2TS U456 ( .A(n160), .Y(n669) );
  AOI22X1TS U457 ( .A0(n1643), .A1(n669), .B0(n72), .B1(
        destinationAddressIn_NORTH[5]), .Y(n73) );
  OAI211XLTS U458 ( .A0(n878), .A1(n269), .B0(n74), .C0(n73), .Y(n2065) );
  INVX2TS U459 ( .A(destinationAddressIn_EAST[4]), .Y(n264) );
  INVX2TS U460 ( .A(n1505), .Y(n76) );
  AOI22X1TS U461 ( .A0(n77), .A1(\destinationAddressbuffer[7][4] ), .B0(n76), 
        .B1(destinationAddressIn_WEST[4]), .Y(n79) );
  INVX2TS U462 ( .A(destinationAddressIn_SOUTH[4]), .Y(n149) );
  INVX2TS U463 ( .A(n149), .Y(n657) );
  AOI22X1TS U464 ( .A0(n1523), .A1(n657), .B0(n869), .B1(
        destinationAddressIn_NORTH[4]), .Y(n78) );
  OAI211XLTS U465 ( .A0(n80), .A1(n264), .B0(n79), .C0(n78), .Y(n2064) );
  INVX2TS U466 ( .A(n82), .Y(n182) );
  AOI21X1TS U467 ( .A0(n223), .A1(n83), .B0(n313), .Y(n386) );
  NOR3XLTS U468 ( .A(n386), .B(n273), .C(n272), .Y(n1558) );
  NOR2XLTS U469 ( .A(n446), .B(n504), .Y(n388) );
  NOR3XLTS U470 ( .A(n23), .B(n84), .C(n83), .Y(n1555) );
  AOI31XLTS U471 ( .A0(n451), .A1(n444), .A2(n388), .B0(n1555), .Y(n86) );
  INVX2TS U472 ( .A(n131), .Y(n449) );
  AOI21X1TS U473 ( .A0(n91), .A1(n86), .B0(n449), .Y(n89) );
  INVX2TS U474 ( .A(n1915), .Y(n392) );
  NAND2X1TS U475 ( .A(n89), .B(n1562), .Y(n92) );
  INVX2TS U476 ( .A(n87), .Y(n1473) );
  INVX2TS U477 ( .A(n1473), .Y(n896) );
  CLKBUFX2TS U478 ( .A(n896), .Y(n101) );
  INVX2TS U479 ( .A(n101), .Y(n118) );
  INVX2TS U480 ( .A(n88), .Y(n893) );
  INVX2TS U481 ( .A(n893), .Y(n1664) );
  CLKBUFX2TS U482 ( .A(n1459), .Y(n894) );
  INVX2TS U483 ( .A(n894), .Y(n106) );
  OR2X1TS U484 ( .A(n1559), .B(n92), .Y(n105) );
  INVX2TS U485 ( .A(n105), .Y(n90) );
  INVX2TS U486 ( .A(n90), .Y(n895) );
  INVX2TS U487 ( .A(n895), .Y(n115) );
  AOI22X1TS U488 ( .A0(n106), .A1(\destinationAddressbuffer[6][11] ), .B0(n115), .B1(n760), .Y(n97) );
  INVX2TS U489 ( .A(n7), .Y(n93) );
  INVX2TS U490 ( .A(n93), .Y(n886) );
  INVX2TS U491 ( .A(n886), .Y(n102) );
  CLKBUFX2TS U492 ( .A(n764), .Y(n404) );
  INVX2TS U493 ( .A(n95), .Y(n107) );
  INVX2TS U494 ( .A(n164), .Y(n339) );
  AOI22X1TS U495 ( .A0(n102), .A1(n404), .B0(n95), .B1(n339), .Y(n96) );
  OAI211XLTS U496 ( .A0(n118), .A1(n235), .B0(n97), .C0(n96), .Y(n2083) );
  INVX2TS U497 ( .A(n105), .Y(n1687) );
  AOI22X1TS U498 ( .A0(n106), .A1(\destinationAddressbuffer[6][9] ), .B0(n90), 
        .B1(n727), .Y(n100) );
  CLKBUFX2TS U499 ( .A(n730), .Y(n399) );
  INVX2TS U500 ( .A(n107), .Y(n1463) );
  INVX2TS U501 ( .A(n107), .Y(n98) );
  INVX2TS U502 ( .A(n176), .Y(n348) );
  AOI22X1TS U503 ( .A0(n93), .A1(n399), .B0(n98), .B1(n348), .Y(n99) );
  OAI211XLTS U504 ( .A0(n118), .A1(n244), .B0(n100), .C0(n99), .Y(n2081) );
  INVX2TS U505 ( .A(n101), .Y(n124) );
  INVX2TS U506 ( .A(n105), .Y(n1665) );
  AOI22X1TS U507 ( .A0(n106), .A1(\destinationAddressbuffer[6][10] ), .B0(
        n1665), .B1(n744), .Y(n104) );
  CLKBUFX2TS U508 ( .A(n748), .Y(n409) );
  INVX2TS U509 ( .A(n171), .Y(n326) );
  AOI22X1TS U510 ( .A0(n102), .A1(n409), .B0(n112), .B1(n326), .Y(n103) );
  OAI211XLTS U511 ( .A0(n124), .A1(n249), .B0(n104), .C0(n103), .Y(n2082) );
  INVX2TS U512 ( .A(n105), .Y(n1461) );
  AOI22X1TS U513 ( .A0(n106), .A1(\destinationAddressbuffer[6][8] ), .B0(n1461), .B1(n712), .Y(n109) );
  INVX2TS U514 ( .A(n7), .Y(n1690) );
  CLKBUFX2TS U515 ( .A(n714), .Y(n416) );
  INVX2TS U516 ( .A(n95), .Y(n897) );
  INVX2TS U517 ( .A(n897), .Y(n112) );
  INVX2TS U518 ( .A(n167), .Y(n333) );
  AOI22X1TS U519 ( .A0(n1690), .A1(n416), .B0(n112), .B1(n333), .Y(n108) );
  OAI211XLTS U520 ( .A0(n118), .A1(n240), .B0(n109), .C0(n108), .Y(n2080) );
  INVX2TS U521 ( .A(n894), .Y(n1685) );
  AOI22X1TS U522 ( .A0(n1685), .A1(writeOutbuffer[6]), .B0(n1665), .B1(
        writeIn_WEST), .Y(n111) );
  INVX2TS U523 ( .A(n7), .Y(n1667) );
  CLKBUFX2TS U524 ( .A(writeIn_NORTH), .Y(n354) );
  CLKBUFX2TS U525 ( .A(n354), .Y(n419) );
  INVX2TS U526 ( .A(n181), .Y(n353) );
  AOI22X1TS U527 ( .A0(n1667), .A1(n419), .B0(n1681), .B1(n353), .Y(n110) );
  OAI211XLTS U528 ( .A0(n124), .A1(n297), .B0(n111), .C0(n110), .Y(n2045) );
  INVX2TS U529 ( .A(n1459), .Y(n121) );
  AOI22X1TS U530 ( .A0(n121), .A1(\destinationAddressbuffer[6][6] ), .B0(n1687), .B1(destinationAddressIn_WEST[6]), .Y(n114) );
  INVX2TS U531 ( .A(n886), .Y(n1674) );
  CLKBUFX2TS U532 ( .A(destinationAddressIn_NORTH[6]), .Y(n366) );
  CLKBUFX2TS U533 ( .A(n366), .Y(n427) );
  INVX2TS U534 ( .A(n144), .Y(n364) );
  AOI22X1TS U535 ( .A0(n1674), .A1(n427), .B0(n112), .B1(n364), .Y(n113) );
  OAI211XLTS U536 ( .A0(n124), .A1(n255), .B0(n114), .C0(n113), .Y(n2078) );
  AOI22X1TS U537 ( .A0(n121), .A1(\destinationAddressbuffer[6][5] ), .B0(n115), 
        .B1(destinationAddressIn_WEST[5]), .Y(n117) );
  INVX2TS U538 ( .A(n7), .Y(n1464) );
  CLKBUFX2TS U539 ( .A(destinationAddressIn_NORTH[5]), .Y(n373) );
  CLKBUFX2TS U540 ( .A(n373), .Y(n423) );
  INVX2TS U541 ( .A(n107), .Y(n1689) );
  INVX2TS U542 ( .A(n160), .Y(n372) );
  AOI22X1TS U543 ( .A0(n1464), .A1(n423), .B0(n1689), .B1(n372), .Y(n116) );
  OAI211XLTS U544 ( .A0(n118), .A1(n269), .B0(n117), .C0(n116), .Y(n2077) );
  AOI22X1TS U545 ( .A0(n121), .A1(\destinationAddressbuffer[6][4] ), .B0(n115), 
        .B1(destinationAddressIn_WEST[4]), .Y(n120) );
  CLKBUFX2TS U546 ( .A(destinationAddressIn_NORTH[4]), .Y(n360) );
  CLKBUFX2TS U547 ( .A(n360), .Y(n431) );
  INVX2TS U548 ( .A(n149), .Y(n359) );
  AOI22X1TS U549 ( .A0(n1690), .A1(n431), .B0(n95), .B1(n359), .Y(n119) );
  OAI211XLTS U550 ( .A0(n1473), .A1(n264), .B0(n120), .C0(n119), .Y(n2076) );
  AOI22X1TS U551 ( .A0(n121), .A1(\destinationAddressbuffer[6][7] ), .B0(n1461), .B1(destinationAddressIn_WEST[7]), .Y(n123) );
  CLKBUFX2TS U552 ( .A(destinationAddressIn_NORTH[7]), .Y(n379) );
  CLKBUFX2TS U553 ( .A(n379), .Y(n436) );
  INVX2TS U554 ( .A(n154), .Y(n378) );
  AOI22X1TS U555 ( .A0(n1464), .A1(n436), .B0(n1463), .B1(n378), .Y(n122) );
  OAI211XLTS U556 ( .A0(n124), .A1(n259), .B0(n123), .C0(n122), .Y(n2079) );
  INVX2TS U557 ( .A(selectBit_EAST), .Y(n512) );
  INVX2TS U558 ( .A(n512), .Y(n514) );
  INVX2TS U559 ( .A(n1920), .Y(n441) );
  NAND2X1TS U560 ( .A(n130), .B(n441), .Y(n132) );
  INVX2TS U561 ( .A(n131), .Y(n316) );
  INVX2TS U562 ( .A(n133), .Y(n510) );
  INVX2TS U563 ( .A(n1920), .Y(n443) );
  INVX2TS U564 ( .A(n135), .Y(n965) );
  INVX2TS U565 ( .A(n965), .Y(n1768) );
  CLKBUFX2TS U566 ( .A(n1768), .Y(n150) );
  INVX2TS U567 ( .A(n150), .Y(n172) );
  INVX2TS U568 ( .A(n136), .Y(n972) );
  INVX2TS U569 ( .A(n972), .Y(n1757) );
  CLKBUFX2TS U570 ( .A(n1366), .Y(n178) );
  INVX2TS U571 ( .A(n178), .Y(n155) );
  AOI22X1TS U572 ( .A0(n155), .A1(\destinationAddressbuffer[3][6] ), .B0(n145), 
        .B1(destinationAddressIn_EAST[6]), .Y(n143) );
  OR2X1TS U573 ( .A(n125), .B(n138), .Y(n168) );
  INVX2TS U574 ( .A(n168), .Y(n139) );
  INVX2TS U575 ( .A(n139), .Y(n151) );
  INVX2TS U576 ( .A(n151), .Y(n958) );
  INVX2TS U577 ( .A(n141), .Y(n156) );
  INVX2TS U578 ( .A(n156), .Y(n1761) );
  CLKBUFX2TS U579 ( .A(destinationAddressIn_WEST[6]), .Y(n687) );
  CLKBUFX2TS U580 ( .A(n687), .Y(n363) );
  AOI22X1TS U581 ( .A0(n958), .A1(n366), .B0(n1761), .B1(n363), .Y(n142) );
  OAI211XLTS U582 ( .A0(n172), .A1(n144), .B0(n143), .C0(n142), .Y(n2114) );
  INVX2TS U583 ( .A(n150), .Y(n177) );
  INVX2TS U584 ( .A(n3), .Y(n145) );
  INVX2TS U585 ( .A(n145), .Y(n950) );
  INVX2TS U586 ( .A(n950), .Y(n146) );
  AOI22X1TS U587 ( .A0(n155), .A1(\destinationAddressbuffer[3][4] ), .B0(n146), 
        .B1(destinationAddressIn_EAST[4]), .Y(n148) );
  INVX2TS U588 ( .A(n156), .Y(n1387) );
  CLKBUFX2TS U589 ( .A(destinationAddressIn_WEST[4]), .Y(n655) );
  CLKBUFX2TS U590 ( .A(n655), .Y(n357) );
  AOI22X1TS U591 ( .A0(n1382), .A1(n360), .B0(n1387), .B1(n357), .Y(n147) );
  OAI211XLTS U592 ( .A0(n177), .A1(n149), .B0(n148), .C0(n147), .Y(n2112) );
  INVX2TS U593 ( .A(n3), .Y(n1782) );
  AOI22X1TS U594 ( .A0(n155), .A1(\destinationAddressbuffer[3][7] ), .B0(n1782), .B1(destinationAddressIn_EAST[7]), .Y(n153) );
  INVX2TS U595 ( .A(n151), .Y(n1382) );
  INVX2TS U596 ( .A(n156), .Y(n1784) );
  CLKBUFX2TS U597 ( .A(destinationAddressIn_WEST[7]), .Y(n701) );
  CLKBUFX2TS U598 ( .A(n701), .Y(n376) );
  AOI22X1TS U599 ( .A0(n1382), .A1(n379), .B0(n1784), .B1(n376), .Y(n152) );
  OAI211XLTS U600 ( .A0(n172), .A1(n154), .B0(n153), .C0(n152), .Y(n2115) );
  INVX2TS U601 ( .A(n3), .Y(n1773) );
  AOI22X1TS U602 ( .A0(n155), .A1(\destinationAddressbuffer[3][5] ), .B0(n1773), .B1(destinationAddressIn_EAST[5]), .Y(n159) );
  INVX2TS U603 ( .A(n151), .Y(n966) );
  INVX2TS U604 ( .A(n156), .Y(n157) );
  INVX2TS U605 ( .A(n157), .Y(n949) );
  INVX2TS U606 ( .A(n949), .Y(n161) );
  CLKBUFX2TS U607 ( .A(destinationAddressIn_WEST[5]), .Y(n667) );
  CLKBUFX2TS U608 ( .A(n667), .Y(n370) );
  AOI22X1TS U609 ( .A0(n966), .A1(n373), .B0(n161), .B1(n370), .Y(n158) );
  OAI211XLTS U610 ( .A0(n172), .A1(n160), .B0(n159), .C0(n158), .Y(n2113) );
  INVX2TS U611 ( .A(n178), .Y(n173) );
  AOI22X1TS U612 ( .A0(n173), .A1(\destinationAddressbuffer[3][11] ), .B0(
        n1773), .B1(destinationAddressIn_EAST[11]), .Y(n163) );
  CLKBUFX2TS U613 ( .A(n403), .Y(n338) );
  AOI22X1TS U614 ( .A0(n958), .A1(n340), .B0(n161), .B1(n338), .Y(n162) );
  OAI211XLTS U615 ( .A0(n177), .A1(n164), .B0(n163), .C0(n162), .Y(n2119) );
  INVX2TS U616 ( .A(n3), .Y(n1381) );
  AOI22X1TS U617 ( .A0(n173), .A1(\destinationAddressbuffer[3][8] ), .B0(n1381), .B1(destinationAddressIn_EAST[8]), .Y(n166) );
  INVX2TS U618 ( .A(n168), .Y(n1762) );
  CLKBUFX2TS U619 ( .A(n413), .Y(n331) );
  AOI22X1TS U620 ( .A0(n1762), .A1(n334), .B0(n1761), .B1(n331), .Y(n165) );
  OAI211XLTS U621 ( .A0(n965), .A1(n167), .B0(n166), .C0(n165), .Y(n2116) );
  AOI22X1TS U622 ( .A0(n173), .A1(\destinationAddressbuffer[3][10] ), .B0(
        n1381), .B1(destinationAddressIn_EAST[10]), .Y(n170) );
  CLKBUFX2TS U623 ( .A(n408), .Y(n320) );
  AOI22X1TS U624 ( .A0(n139), .A1(n327), .B0(n1387), .B1(n320), .Y(n169) );
  OAI211XLTS U625 ( .A0(n172), .A1(n171), .B0(n170), .C0(n169), .Y(n2118) );
  AOI22X1TS U626 ( .A0(n173), .A1(\destinationAddressbuffer[3][9] ), .B0(n145), 
        .B1(destinationAddressIn_EAST[9]), .Y(n175) );
  CLKBUFX2TS U627 ( .A(n395), .Y(n344) );
  AOI22X1TS U628 ( .A0(n966), .A1(n349), .B0(n141), .B1(n344), .Y(n174) );
  OAI211XLTS U629 ( .A0(n177), .A1(n176), .B0(n175), .C0(n174), .Y(n2117) );
  INVX2TS U630 ( .A(n178), .Y(n1780) );
  AOI22X1TS U631 ( .A0(n1780), .A1(writeOutbuffer[3]), .B0(n1782), .B1(
        writeIn_EAST), .Y(n180) );
  CLKBUFX2TS U632 ( .A(writeIn_WEST), .Y(n542) );
  CLKBUFX2TS U633 ( .A(n542), .Y(n352) );
  AOI22X1TS U634 ( .A0(n139), .A1(n354), .B0(n1784), .B1(n352), .Y(n179) );
  OAI211XLTS U635 ( .A0(n177), .A1(n181), .B0(n180), .C0(n179), .Y(n2048) );
  INVX2TS U636 ( .A(n272), .Y(n314) );
  INVX2TS U637 ( .A(n314), .Y(n384) );
  NOR3XLTS U638 ( .A(n386), .B(n384), .C(n385), .Y(n1599) );
  AOI31XLTS U639 ( .A0(n495), .A1(n388), .A2(n450), .B0(n1596), .Y(n183) );
  NAND2X1TS U640 ( .A(n186), .B(n1603), .Y(n188) );
  INVX2TS U641 ( .A(n184), .Y(n1344) );
  INVX2TS U642 ( .A(n1344), .Y(n991) );
  CLKBUFX2TS U643 ( .A(n991), .Y(n197) );
  INVX2TS U644 ( .A(n197), .Y(n215) );
  INVX2TS U645 ( .A(n185), .Y(n989) );
  INVX2TS U646 ( .A(n989), .Y(n1789) );
  INVX2TS U647 ( .A(n981), .Y(n203) );
  OR2X1TS U648 ( .A(n1600), .B(n188), .Y(n202) );
  INVX2TS U649 ( .A(n202), .Y(n1809) );
  AOI22X1TS U650 ( .A0(n203), .A1(\destinationAddressbuffer[2][9] ), .B0(n1809), .B1(n344), .Y(n192) );
  INVX2TS U651 ( .A(n193), .Y(n1340) );
  INVX2TS U652 ( .A(n1340), .Y(n985) );
  INVX2TS U653 ( .A(n190), .Y(n204) );
  INVX2TS U654 ( .A(n204), .Y(n1110) );
  AOI22X1TS U655 ( .A0(n985), .A1(n349), .B0(n212), .B1(n348), .Y(n191) );
  OAI211XLTS U656 ( .A0(n215), .A1(n244), .B0(n192), .C0(n191), .Y(n2129) );
  INVX2TS U657 ( .A(n202), .Y(n1109) );
  AOI22X1TS U658 ( .A0(n203), .A1(\destinationAddressbuffer[2][10] ), .B0(
        n1109), .B1(n320), .Y(n196) );
  INVX2TS U659 ( .A(n193), .Y(n216) );
  INVX2TS U660 ( .A(n216), .Y(n194) );
  INVX2TS U661 ( .A(n204), .Y(n1351) );
  AOI22X1TS U662 ( .A0(n194), .A1(n327), .B0(n1351), .B1(n326), .Y(n195) );
  OAI211XLTS U663 ( .A0(n215), .A1(n249), .B0(n196), .C0(n195), .Y(n2130) );
  INVX2TS U664 ( .A(n197), .Y(n222) );
  INVX2TS U665 ( .A(n202), .Y(n198) );
  INVX2TS U666 ( .A(n198), .Y(n990) );
  INVX2TS U667 ( .A(n990), .Y(n209) );
  AOI22X1TS U668 ( .A0(n203), .A1(\destinationAddressbuffer[2][8] ), .B0(n209), 
        .B1(n331), .Y(n201) );
  INVX2TS U669 ( .A(n216), .Y(n1810) );
  INVX2TS U670 ( .A(n204), .Y(n199) );
  INVX2TS U671 ( .A(n199), .Y(n992) );
  INVX2TS U672 ( .A(n992), .Y(n212) );
  AOI22X1TS U673 ( .A0(n1810), .A1(n334), .B0(n212), .B1(n333), .Y(n200) );
  OAI211XLTS U674 ( .A0(n222), .A1(n240), .B0(n201), .C0(n200), .Y(n2128) );
  INVX2TS U675 ( .A(n202), .Y(n1790) );
  AOI22X1TS U676 ( .A0(n203), .A1(\destinationAddressbuffer[2][11] ), .B0(
        n1790), .B1(n338), .Y(n206) );
  INVX2TS U677 ( .A(n204), .Y(n1362) );
  AOI22X1TS U678 ( .A0(n194), .A1(n340), .B0(n1362), .B1(n339), .Y(n205) );
  OAI211XLTS U679 ( .A0(n215), .A1(n235), .B0(n206), .C0(n205), .Y(n2131) );
  CLKBUFX2TS U680 ( .A(n981), .Y(n1604) );
  INVX2TS U681 ( .A(n1604), .Y(n1808) );
  AOI22X1TS U682 ( .A0(n1808), .A1(writeOutbuffer[2]), .B0(n209), .B1(n352), 
        .Y(n208) );
  INVX2TS U683 ( .A(n216), .Y(n1791) );
  AOI22X1TS U684 ( .A0(n1791), .A1(writeIn_NORTH), .B0(n1351), .B1(n353), .Y(
        n207) );
  OAI211XLTS U685 ( .A0(n222), .A1(n297), .B0(n208), .C0(n207), .Y(n2049) );
  INVX2TS U686 ( .A(n981), .Y(n219) );
  AOI22X1TS U687 ( .A0(n219), .A1(\destinationAddressbuffer[2][4] ), .B0(n209), 
        .B1(n357), .Y(n211) );
  AOI22X1TS U688 ( .A0(n1810), .A1(destinationAddressIn_NORTH[4]), .B0(n1362), 
        .B1(n359), .Y(n210) );
  OAI211XLTS U689 ( .A0(n222), .A1(n264), .B0(n211), .C0(n210), .Y(n2124) );
  AOI22X1TS U690 ( .A0(n219), .A1(\destinationAddressbuffer[2][6] ), .B0(n198), 
        .B1(n363), .Y(n214) );
  AOI22X1TS U691 ( .A0(n985), .A1(destinationAddressIn_NORTH[6]), .B0(n212), 
        .B1(n364), .Y(n213) );
  OAI211XLTS U692 ( .A0(n215), .A1(n255), .B0(n214), .C0(n213), .Y(n2126) );
  AOI22X1TS U693 ( .A0(n219), .A1(\destinationAddressbuffer[2][5] ), .B0(n1109), .B1(n370), .Y(n218) );
  INVX2TS U694 ( .A(n216), .Y(n1111) );
  AOI22X1TS U695 ( .A0(n1111), .A1(destinationAddressIn_NORTH[5]), .B0(n1110), 
        .B1(n372), .Y(n217) );
  OAI211XLTS U696 ( .A0(n1344), .A1(n269), .B0(n218), .C0(n217), .Y(n2125) );
  AOI22X1TS U697 ( .A0(n219), .A1(\destinationAddressbuffer[2][7] ), .B0(n1790), .B1(n376), .Y(n221) );
  AOI22X1TS U698 ( .A0(n1111), .A1(destinationAddressIn_NORTH[7]), .B0(n1110), 
        .B1(n378), .Y(n220) );
  OAI211XLTS U699 ( .A0(n222), .A1(n259), .B0(n221), .C0(n220), .Y(n2127) );
  INVX2TS U700 ( .A(n1918), .Y(n387) );
  INVX2TS U701 ( .A(n1919), .Y(n493) );
  INVX2TS U702 ( .A(n1918), .Y(n391) );
  NAND2X1TS U703 ( .A(n227), .B(n1574), .Y(n229) );
  INVX2TS U704 ( .A(n225), .Y(n1436) );
  INVX2TS U705 ( .A(n1436), .Y(n914) );
  CLKBUFX2TS U706 ( .A(n914), .Y(n241) );
  INVX2TS U707 ( .A(n241), .Y(n260) );
  INVX2TS U708 ( .A(n9), .Y(n1694) );
  CLKBUFX2TS U709 ( .A(n1424), .Y(n912) );
  INVX2TS U710 ( .A(n912), .Y(n246) );
  OR2X1TS U711 ( .A(n1571), .B(n229), .Y(n245) );
  INVX2TS U712 ( .A(n245), .Y(n1697) );
  AOI22X1TS U713 ( .A0(n246), .A1(\destinationAddressbuffer[5][11] ), .B0(
        n1697), .B1(n760), .Y(n234) );
  INVX2TS U714 ( .A(n1564), .Y(n1567) );
  NAND2BX1TS U715 ( .AN(n229), .B(n228), .Y(n231) );
  INVX2TS U716 ( .A(n256), .Y(n1450) );
  OR2X1TS U717 ( .A(n1564), .B(n231), .Y(n250) );
  INVX2TS U718 ( .A(n250), .Y(n232) );
  INVX2TS U719 ( .A(n232), .Y(n901) );
  INVX2TS U720 ( .A(n901), .Y(n237) );
  AOI22X1TS U721 ( .A0(n1450), .A1(n404), .B0(n237), .B1(n339), .Y(n233) );
  OAI211XLTS U722 ( .A0(n260), .A1(n235), .B0(n234), .C0(n233), .Y(n2095) );
  INVX2TS U723 ( .A(n245), .Y(n236) );
  INVX2TS U724 ( .A(n236), .Y(n913) );
  INVX2TS U725 ( .A(n913), .Y(n261) );
  AOI22X1TS U726 ( .A0(n246), .A1(\destinationAddressbuffer[5][8] ), .B0(n261), 
        .B1(n712), .Y(n239) );
  INVX2TS U727 ( .A(n256), .Y(n1428) );
  AOI22X1TS U728 ( .A0(n1450), .A1(n416), .B0(n237), .B1(n333), .Y(n238) );
  OAI211XLTS U729 ( .A0(n260), .A1(n240), .B0(n239), .C0(n238), .Y(n2092) );
  INVX2TS U730 ( .A(n241), .Y(n270) );
  INVX2TS U731 ( .A(n245), .Y(n1723) );
  AOI22X1TS U732 ( .A0(n246), .A1(\destinationAddressbuffer[5][9] ), .B0(n1723), .B1(n727), .Y(n243) );
  INVX2TS U733 ( .A(n250), .Y(n1698) );
  AOI22X1TS U734 ( .A0(n1428), .A1(n399), .B0(n1698), .B1(n348), .Y(n242) );
  OAI211XLTS U735 ( .A0(n270), .A1(n244), .B0(n243), .C0(n242), .Y(n2093) );
  INVX2TS U736 ( .A(n245), .Y(n1425) );
  AOI22X1TS U737 ( .A0(n246), .A1(\destinationAddressbuffer[5][10] ), .B0(
        n1425), .B1(n744), .Y(n248) );
  INVX2TS U738 ( .A(n256), .Y(n1699) );
  INVX2TS U739 ( .A(n1699), .Y(n266) );
  INVX2TS U740 ( .A(n266), .Y(n908) );
  INVX2TS U741 ( .A(n250), .Y(n1448) );
  AOI22X1TS U742 ( .A0(n908), .A1(n409), .B0(n1448), .B1(n326), .Y(n247) );
  OAI211XLTS U743 ( .A0(n260), .A1(n249), .B0(n248), .C0(n247), .Y(n2094) );
  INVX2TS U744 ( .A(n912), .Y(n1719) );
  AOI22X1TS U745 ( .A0(n1719), .A1(writeOutbuffer[5]), .B0(n261), .B1(n542), 
        .Y(n252) );
  INVX2TS U746 ( .A(n250), .Y(n1426) );
  AOI22X1TS U747 ( .A0(n1428), .A1(n419), .B0(n1426), .B1(n353), .Y(n251) );
  OAI211XLTS U748 ( .A0(n270), .A1(n297), .B0(n252), .C0(n251), .Y(n2046) );
  INVX2TS U749 ( .A(n1424), .Y(n265) );
  AOI22X1TS U750 ( .A0(n265), .A1(\destinationAddressbuffer[5][6] ), .B0(n236), 
        .B1(n687), .Y(n254) );
  AOI22X1TS U751 ( .A0(n1699), .A1(n427), .B0(n232), .B1(n364), .Y(n253) );
  OAI211XLTS U752 ( .A0(n270), .A1(n255), .B0(n254), .C0(n253), .Y(n2090) );
  AOI22X1TS U753 ( .A0(n265), .A1(\destinationAddressbuffer[5][7] ), .B0(n1697), .B1(n701), .Y(n258) );
  INVX2TS U754 ( .A(n256), .Y(n1438) );
  AOI22X1TS U755 ( .A0(n1438), .A1(n436), .B0(n1426), .B1(n378), .Y(n257) );
  OAI211XLTS U756 ( .A0(n260), .A1(n259), .B0(n258), .C0(n257), .Y(n2091) );
  AOI22X1TS U757 ( .A0(n265), .A1(\destinationAddressbuffer[5][4] ), .B0(n261), 
        .B1(n655), .Y(n263) );
  AOI22X1TS U758 ( .A0(n1438), .A1(n431), .B0(n237), .B1(n359), .Y(n262) );
  OAI211XLTS U759 ( .A0(n1436), .A1(n264), .B0(n263), .C0(n262), .Y(n2088) );
  AOI22X1TS U760 ( .A0(n265), .A1(\destinationAddressbuffer[5][5] ), .B0(n1425), .B1(n667), .Y(n268) );
  INVX2TS U761 ( .A(n266), .Y(n1707) );
  AOI22X1TS U762 ( .A0(n1707), .A1(n423), .B0(n1448), .B1(n372), .Y(n267) );
  OAI211XLTS U763 ( .A0(n270), .A1(n269), .B0(n268), .C0(n267), .Y(n2089) );
  AOI31XLTS U764 ( .A0(n275), .A1(n388), .A2(n387), .B0(n1577), .Y(n274) );
  AOI21X1TS U765 ( .A0(n280), .A1(n274), .B0(n440), .Y(n278) );
  NAND2X1TS U766 ( .A(n278), .B(n1585), .Y(n281) );
  INVX2TS U767 ( .A(n1402), .Y(n940) );
  CLKBUFX2TS U768 ( .A(n940), .Y(n289) );
  INVX2TS U769 ( .A(n289), .Y(n305) );
  INVX2TS U770 ( .A(n277), .Y(n937) );
  INVX2TS U771 ( .A(n937), .Y(n1728) );
  CLKBUFX2TS U772 ( .A(n1391), .Y(n938) );
  INVX2TS U773 ( .A(n938), .Y(n293) );
  OR2X1TS U774 ( .A(n1581), .B(n281), .Y(n292) );
  INVX2TS U775 ( .A(n292), .Y(n279) );
  INVX2TS U776 ( .A(n279), .Y(n939) );
  INVX2TS U777 ( .A(n939), .Y(n309) );
  AOI22X1TS U778 ( .A0(n293), .A1(\destinationAddressbuffer[4][8] ), .B0(n309), 
        .B1(n331), .Y(n285) );
  INVX2TS U779 ( .A(n4), .Y(n282) );
  INVX2TS U780 ( .A(n282), .Y(n943) );
  INVX2TS U781 ( .A(n943), .Y(n302) );
  INVX2TS U782 ( .A(n5), .Y(n1730) );
  AOI22X1TS U783 ( .A0(n302), .A1(n713), .B0(n1730), .B1(n416), .Y(n284) );
  OAI211XLTS U784 ( .A0(n305), .A1(n33), .B0(n285), .C0(n284), .Y(n2104) );
  INVX2TS U785 ( .A(n289), .Y(n308) );
  INVX2TS U786 ( .A(n292), .Y(n1729) );
  AOI22X1TS U787 ( .A0(n293), .A1(\destinationAddressbuffer[4][11] ), .B0(
        n1729), .B1(n338), .Y(n288) );
  INVX2TS U788 ( .A(n4), .Y(n1744) );
  INVX2TS U789 ( .A(n5), .Y(n286) );
  INVX2TS U790 ( .A(n286), .Y(n294) );
  INVX2TS U791 ( .A(n294), .Y(n1414) );
  AOI22X1TS U792 ( .A0(n1744), .A1(n763), .B0(n1414), .B1(n404), .Y(n287) );
  OAI211XLTS U793 ( .A0(n308), .A1(n49), .B0(n288), .C0(n287), .Y(n2107) );
  INVX2TS U794 ( .A(n292), .Y(n1751) );
  AOI22X1TS U795 ( .A0(n293), .A1(\destinationAddressbuffer[4][9] ), .B0(n1751), .B1(n344), .Y(n291) );
  INVX2TS U796 ( .A(n4), .Y(n1753) );
  INVX2TS U797 ( .A(n5), .Y(n1752) );
  AOI22X1TS U798 ( .A0(n1753), .A1(n728), .B0(n286), .B1(n399), .Y(n290) );
  OAI211XLTS U799 ( .A0(n305), .A1(n45), .B0(n291), .C0(n290), .Y(n2105) );
  INVX2TS U800 ( .A(n292), .Y(n1393) );
  AOI22X1TS U801 ( .A0(n293), .A1(\destinationAddressbuffer[4][10] ), .B0(
        n1393), .B1(n320), .Y(n296) );
  INVX2TS U802 ( .A(n294), .Y(n920) );
  AOI22X1TS U803 ( .A0(n302), .A1(n747), .B0(n920), .B1(n409), .Y(n295) );
  OAI211XLTS U804 ( .A0(n305), .A1(n41), .B0(n296), .C0(n295), .Y(n2106) );
  INVX2TS U805 ( .A(n938), .Y(n1748) );
  AOI22X1TS U806 ( .A0(n1748), .A1(writeOutbuffer[4]), .B0(n309), .B1(n352), 
        .Y(n299) );
  INVX2TS U807 ( .A(n4), .Y(n1415) );
  INVX2TS U808 ( .A(n5), .Y(n1394) );
  AOI22X1TS U809 ( .A0(n1415), .A1(n544), .B0(n1394), .B1(n419), .Y(n298) );
  OAI211XLTS U810 ( .A0(n308), .A1(n56), .B0(n299), .C0(n298), .Y(n2047) );
  INVX2TS U811 ( .A(n1391), .Y(n310) );
  AOI22X1TS U812 ( .A0(n310), .A1(\destinationAddressbuffer[4][7] ), .B0(n1729), .B1(n376), .Y(n301) );
  AOI22X1TS U813 ( .A0(n282), .A1(n702), .B0(n1394), .B1(n436), .Y(n300) );
  OAI211XLTS U814 ( .A0(n308), .A1(n62), .B0(n301), .C0(n300), .Y(n2103) );
  AOI22X1TS U815 ( .A0(n310), .A1(\destinationAddressbuffer[4][6] ), .B0(n279), 
        .B1(n363), .Y(n304) );
  AOI22X1TS U816 ( .A0(n302), .A1(n689), .B0(n286), .B1(n427), .Y(n303) );
  OAI211XLTS U817 ( .A0(n305), .A1(n66), .B0(n304), .C0(n303), .Y(n2102) );
  AOI22X1TS U818 ( .A0(n310), .A1(\destinationAddressbuffer[4][5] ), .B0(n1393), .B1(n370), .Y(n307) );
  AOI22X1TS U819 ( .A0(n1415), .A1(n669), .B0(n920), .B1(n423), .Y(n306) );
  OAI211XLTS U820 ( .A0(n308), .A1(n71), .B0(n307), .C0(n306), .Y(n2101) );
  AOI22X1TS U821 ( .A0(n310), .A1(\destinationAddressbuffer[4][4] ), .B0(n309), 
        .B1(n357), .Y(n312) );
  AOI22X1TS U822 ( .A0(n282), .A1(n657), .B0(n1730), .B1(n431), .Y(n311) );
  OAI211XLTS U823 ( .A0(n1402), .A1(n75), .B0(n312), .C0(n311), .Y(n2100) );
  AOI31XLTS U824 ( .A0(n315), .A1(n391), .A2(n441), .B0(n1609), .Y(n317) );
  NAND2X1TS U825 ( .A(n319), .B(n1618), .Y(n322) );
  INVX2TS U826 ( .A(n318), .Y(n1089) );
  INVX2TS U827 ( .A(n1089), .Y(n1018) );
  CLKBUFX2TS U828 ( .A(n1018), .Y(n337) );
  INVX2TS U829 ( .A(n337), .Y(n369) );
  OR2X1TS U830 ( .A(n449), .B(n1618), .Y(n1084) );
  INVX2TS U831 ( .A(n1084), .Y(n1845) );
  OR2X1TS U832 ( .A(n319), .B(n1845), .Y(n1003) );
  INVX2TS U833 ( .A(n1003), .Y(n345) );
  OR2X1TS U834 ( .A(n1614), .B(n322), .Y(n343) );
  INVX2TS U835 ( .A(n343), .Y(n1078) );
  AOI22X1TS U836 ( .A0(n345), .A1(\destinationAddressbuffer[1][10] ), .B0(
        n1078), .B1(n320), .Y(n329) );
  INVX2TS U837 ( .A(n346), .Y(n371) );
  INVX2TS U838 ( .A(n371), .Y(n323) );
  INVX2TS U839 ( .A(n325), .Y(n347) );
  INVX2TS U840 ( .A(n347), .Y(n1094) );
  AOI22X1TS U841 ( .A0(n323), .A1(n327), .B0(n1094), .B1(n326), .Y(n328) );
  OAI211XLTS U842 ( .A0(n369), .A1(n41), .B0(n329), .C0(n328), .Y(n2142) );
  INVX2TS U843 ( .A(n343), .Y(n330) );
  INVX2TS U844 ( .A(n330), .Y(n1017) );
  INVX2TS U845 ( .A(n1017), .Y(n358) );
  AOI22X1TS U846 ( .A0(n345), .A1(\destinationAddressbuffer[1][8] ), .B0(n358), 
        .B1(n331), .Y(n336) );
  INVX2TS U847 ( .A(n371), .Y(n1851) );
  INVX2TS U848 ( .A(n347), .Y(n332) );
  INVX2TS U849 ( .A(n332), .Y(n1020) );
  INVX2TS U850 ( .A(n1020), .Y(n365) );
  AOI22X1TS U851 ( .A0(n1851), .A1(n334), .B0(n365), .B1(n333), .Y(n335) );
  OAI211XLTS U852 ( .A0(n369), .A1(n33), .B0(n336), .C0(n335), .Y(n2140) );
  INVX2TS U853 ( .A(n337), .Y(n382) );
  INVX2TS U854 ( .A(n343), .Y(n1816) );
  AOI22X1TS U855 ( .A0(n345), .A1(\destinationAddressbuffer[1][11] ), .B0(
        n1816), .B1(n338), .Y(n342) );
  INVX2TS U856 ( .A(n347), .Y(n1104) );
  AOI22X1TS U857 ( .A0(n323), .A1(n340), .B0(n1104), .B1(n339), .Y(n341) );
  OAI211XLTS U858 ( .A0(n382), .A1(n49), .B0(n342), .C0(n341), .Y(n2143) );
  INVX2TS U859 ( .A(n343), .Y(n1848) );
  AOI22X1TS U860 ( .A0(n345), .A1(\destinationAddressbuffer[1][9] ), .B0(n1848), .B1(n344), .Y(n351) );
  INVX2TS U861 ( .A(n346), .Y(n1085) );
  INVX2TS U862 ( .A(n1085), .Y(n1011) );
  INVX2TS U863 ( .A(n347), .Y(n1079) );
  AOI22X1TS U864 ( .A0(n1011), .A1(n349), .B0(n365), .B1(n348), .Y(n350) );
  OAI211XLTS U865 ( .A0(n369), .A1(n45), .B0(n351), .C0(n350), .Y(n2141) );
  CLKBUFX2TS U866 ( .A(n1003), .Y(n1619) );
  INVX2TS U867 ( .A(n1619), .Y(n1844) );
  AOI22X1TS U868 ( .A0(n1844), .A1(writeOutbuffer[1]), .B0(n358), .B1(n352), 
        .Y(n356) );
  INVX2TS U869 ( .A(n371), .Y(n1819) );
  AOI22X1TS U870 ( .A0(n1819), .A1(n354), .B0(n1094), .B1(n353), .Y(n355) );
  OAI211XLTS U871 ( .A0(n382), .A1(n56), .B0(n356), .C0(n355), .Y(n2050) );
  INVX2TS U872 ( .A(n1003), .Y(n377) );
  AOI22X1TS U873 ( .A0(n377), .A1(\destinationAddressbuffer[1][4] ), .B0(n358), 
        .B1(n357), .Y(n362) );
  AOI22X1TS U874 ( .A0(n1851), .A1(n360), .B0(n1104), .B1(n359), .Y(n361) );
  OAI211XLTS U875 ( .A0(n382), .A1(n75), .B0(n362), .C0(n361), .Y(n2136) );
  AOI22X1TS U876 ( .A0(n377), .A1(\destinationAddressbuffer[1][6] ), .B0(n330), 
        .B1(n363), .Y(n368) );
  AOI22X1TS U877 ( .A0(n1011), .A1(n366), .B0(n365), .B1(n364), .Y(n367) );
  OAI211XLTS U878 ( .A0(n369), .A1(n66), .B0(n368), .C0(n367), .Y(n2138) );
  AOI22X1TS U879 ( .A0(n377), .A1(\destinationAddressbuffer[1][5] ), .B0(n1078), .B1(n370), .Y(n375) );
  INVX2TS U880 ( .A(n371), .Y(n1080) );
  AOI22X1TS U881 ( .A0(n1080), .A1(n373), .B0(n1079), .B1(n372), .Y(n374) );
  OAI211XLTS U882 ( .A0(n1089), .A1(n71), .B0(n375), .C0(n374), .Y(n2137) );
  AOI22X1TS U883 ( .A0(n377), .A1(\destinationAddressbuffer[1][7] ), .B0(n1816), .B1(n376), .Y(n381) );
  AOI22X1TS U884 ( .A0(n1080), .A1(n379), .B0(n1079), .B1(n378), .Y(n380) );
  OAI211XLTS U885 ( .A0(n382), .A1(n62), .B0(n381), .C0(n380), .Y(n2139) );
  AOI31XLTS U886 ( .A0(n388), .A1(n387), .A2(n443), .B0(n1624), .Y(n390) );
  NAND2X1TS U887 ( .A(n394), .B(n1633), .Y(n397) );
  INVX2TS U888 ( .A(n393), .Y(n1061) );
  INVX2TS U889 ( .A(n1061), .Y(n1045) );
  CLKBUFX2TS U890 ( .A(n1045), .Y(n407) );
  INVX2TS U891 ( .A(n407), .Y(n430) );
  INVX2TS U892 ( .A(n11), .Y(n1855) );
  CLKBUFX2TS U893 ( .A(n1031), .Y(n1043) );
  INVX2TS U894 ( .A(n1043), .Y(n414) );
  OR2X1TS U895 ( .A(n1629), .B(n397), .Y(n412) );
  INVX2TS U896 ( .A(n412), .Y(n1887) );
  AOI22X1TS U897 ( .A0(n414), .A1(\destinationAddressbuffer[0][9] ), .B0(n402), 
        .B1(n395), .Y(n401) );
  INVX2TS U898 ( .A(n10), .Y(n1891) );
  INVX2TS U899 ( .A(n6), .Y(n1889) );
  INVX2TS U900 ( .A(n1889), .Y(n1057) );
  INVX2TS U901 ( .A(n1057), .Y(n1033) );
  AOI22X1TS U902 ( .A0(n1891), .A1(n728), .B0(n1033), .B1(n399), .Y(n400) );
  OAI211XLTS U903 ( .A0(n430), .A1(n45), .B0(n401), .C0(n400), .Y(n2153) );
  INVX2TS U904 ( .A(n407), .Y(n434) );
  INVX2TS U905 ( .A(n412), .Y(n402) );
  INVX2TS U906 ( .A(n402), .Y(n1044) );
  INVX2TS U907 ( .A(n1044), .Y(n422) );
  AOI22X1TS U908 ( .A0(n414), .A1(\destinationAddressbuffer[0][11] ), .B0(n422), .B1(n403), .Y(n406) );
  INVX2TS U909 ( .A(n10), .Y(n1880) );
  AOI22X1TS U910 ( .A0(n1880), .A1(n763), .B0(n424), .B1(n404), .Y(n405) );
  OAI211XLTS U911 ( .A0(n434), .A1(n49), .B0(n406), .C0(n405), .Y(n2155) );
  INVX2TS U912 ( .A(n412), .Y(n1857) );
  AOI22X1TS U913 ( .A0(n414), .A1(\destinationAddressbuffer[0][10] ), .B0(
        n1857), .B1(n408), .Y(n411) );
  INVX2TS U914 ( .A(n1047), .Y(n437) );
  AOI22X1TS U915 ( .A0(n437), .A1(n747), .B0(n424), .B1(n409), .Y(n410) );
  OAI211XLTS U916 ( .A0(n430), .A1(n41), .B0(n411), .C0(n410), .Y(n2154) );
  INVX2TS U917 ( .A(n412), .Y(n1052) );
  AOI22X1TS U918 ( .A0(n414), .A1(\destinationAddressbuffer[0][8] ), .B0(n1052), .B1(n413), .Y(n418) );
  INVX2TS U919 ( .A(n10), .Y(n415) );
  INVX2TS U920 ( .A(n415), .Y(n1047) );
  INVX2TS U921 ( .A(n6), .Y(n1859) );
  AOI22X1TS U922 ( .A0(n437), .A1(n713), .B0(n1859), .B1(n416), .Y(n417) );
  OAI211XLTS U923 ( .A0(n430), .A1(n33), .B0(n418), .C0(n417), .Y(n2152) );
  INVX2TS U924 ( .A(n1031), .Y(n1884) );
  AOI22X1TS U925 ( .A0(n1884), .A1(writeOutbuffer[0]), .B0(n1857), .B1(
        writeIn_WEST), .Y(n421) );
  INVX2TS U926 ( .A(n10), .Y(n1070) );
  INVX2TS U927 ( .A(n6), .Y(n1053) );
  AOI22X1TS U928 ( .A0(n1070), .A1(n544), .B0(n1053), .B1(n419), .Y(n420) );
  OAI211XLTS U929 ( .A0(n434), .A1(n56), .B0(n421), .C0(n420), .Y(n2051) );
  INVX2TS U930 ( .A(n1031), .Y(n435) );
  AOI22X1TS U931 ( .A0(n435), .A1(\destinationAddressbuffer[0][5] ), .B0(n422), 
        .B1(destinationAddressIn_WEST[5]), .Y(n426) );
  INVX2TS U932 ( .A(n1057), .Y(n424) );
  AOI22X1TS U933 ( .A0(n1070), .A1(n669), .B0(n424), .B1(n423), .Y(n425) );
  OAI211XLTS U934 ( .A0(n434), .A1(n71), .B0(n426), .C0(n425), .Y(n2149) );
  AOI22X1TS U935 ( .A0(n435), .A1(\destinationAddressbuffer[0][6] ), .B0(n1887), .B1(destinationAddressIn_WEST[6]), .Y(n429) );
  AOI22X1TS U936 ( .A0(n1861), .A1(n689), .B0(n1033), .B1(n427), .Y(n428) );
  OAI211XLTS U937 ( .A0(n430), .A1(n66), .B0(n429), .C0(n428), .Y(n2150) );
  AOI22X1TS U938 ( .A0(n435), .A1(\destinationAddressbuffer[0][4] ), .B0(n422), 
        .B1(destinationAddressIn_WEST[4]), .Y(n433) );
  AOI22X1TS U939 ( .A0(n437), .A1(n657), .B0(n1859), .B1(n431), .Y(n432) );
  OAI211XLTS U940 ( .A0(n434), .A1(n75), .B0(n433), .C0(n432), .Y(n2148) );
  AOI22X1TS U941 ( .A0(n435), .A1(\destinationAddressbuffer[0][7] ), .B0(n1052), .B1(destinationAddressIn_WEST[7]), .Y(n439) );
  AOI22X1TS U942 ( .A0(n437), .A1(n702), .B0(n1053), .B1(n436), .Y(n438) );
  OAI211XLTS U943 ( .A0(n1061), .A1(n62), .B0(n439), .C0(n438), .Y(n2151) );
  INVX2TS U944 ( .A(n1922), .Y(n527) );
  INVX2TS U945 ( .A(n1922), .Y(n524) );
  INVX2TS U946 ( .A(n1916), .Y(n530) );
  NAND2X1TS U947 ( .A(n524), .B(n530), .Y(n528) );
  OAI21XLTS U948 ( .A0(n527), .A1(n1917), .B0(n528), .Y(n502) );
  INVX2TS U949 ( .A(n1913), .Y(n531) );
  INVX2TS U950 ( .A(n1913), .Y(n526) );
  NOR2XLTS U951 ( .A(n528), .B(n526), .Y(n833) );
  CLKBUFX2TS U952 ( .A(n833), .Y(n793) );
  CLKBUFX2TS U953 ( .A(n793), .Y(n813) );
  AOI21X1TS U954 ( .A0(n528), .A1(n531), .B0(n813), .Y(n499) );
  OAI22X1TS U955 ( .A0(n455), .A1(n502), .B0(n441), .B1(n499), .Y(n442) );
  AOI221XLTS U956 ( .A0(n502), .A1(n444), .B0(n443), .B1(n499), .C0(n442), .Y(
        n447) );
  INVX2TS U957 ( .A(n1910), .Y(n445) );
  NAND2X1TS U958 ( .A(n446), .B(n445), .Y(n460) );
  OAI21XLTS U959 ( .A0(n493), .A1(n1922), .B0(n460), .Y(n464) );
  AOI21X1TS U960 ( .A0(n447), .A1(n464), .B0(n1912), .Y(n448) );
  INVX2TS U961 ( .A(reset), .Y(n491) );
  NAND2X1TS U962 ( .A(n491), .B(n1912), .Y(n503) );
  INVX2TS U963 ( .A(n1918), .Y(n461) );
  INVX2TS U964 ( .A(n1921), .Y(n451) );
  INVX2TS U965 ( .A(n1914), .Y(n529) );
  AOI22X1TS U966 ( .A0(n451), .A1(n526), .B0(n529), .B1(n450), .Y(n454) );
  INVX2TS U967 ( .A(n453), .Y(n459) );
  INVX2TS U968 ( .A(n474), .Y(n471) );
  AOI21X1TS U969 ( .A0(n527), .A1(n457), .B0(n456), .Y(n470) );
  ADDFHX1TS U970 ( .A(n459), .B(n513), .CI(n458), .CO(n462), .S(n475) );
  ADDHXLTS U971 ( .A(n463), .B(n462), .CO(n474), .S(n476) );
  INVX2TS U972 ( .A(n476), .Y(n465) );
  AOI21X1TS U973 ( .A0(n466), .A1(n465), .B0(n464), .Y(n468) );
  OAI22X1TS U974 ( .A0(n466), .A1(n465), .B0(n472), .B1(n471), .Y(n467) );
  AOI21X1TS U975 ( .A0(n475), .A1(n468), .B0(n467), .Y(n469) );
  AOI211X1TS U976 ( .A0(n472), .A1(n471), .B0(n470), .C0(n469), .Y(n473) );
  INVX2TS U977 ( .A(n473), .Y(n477) );
  NAND2X1TS U978 ( .A(n477), .B(n474), .Y(n481) );
  XOR2X2TS U979 ( .A(n481), .B(n480), .Y(n496) );
  INVX2TS U980 ( .A(n496), .Y(n489) );
  INVX2TS U981 ( .A(n1914), .Y(n525) );
  ADDHXLTS U982 ( .A(n446), .B(n482), .CO(n485), .S(n492) );
  XNOR2X1TS U983 ( .A(n1917), .B(n494), .Y(n486) );
  OAI21X1TS U984 ( .A0(n489), .A1(n525), .B0(n486), .Y(n487) );
  OAI2BB2XLTS U985 ( .B0(n1924), .B1(n503), .A0N(n497), .A1N(n490), .Y(N2624)
         );
  CLKBUFX2TS U986 ( .A(n1911), .Y(n639) );
  CLKBUFX2TS U987 ( .A(n639), .Y(n606) );
  NAND2X1TS U988 ( .A(n491), .B(n606), .Y(n501) );
  AOI22X1TS U989 ( .A0(n1910), .A1(n503), .B0(n501), .B1(n445), .Y(n1933) );
  INVX2TS U990 ( .A(n499), .Y(n500) );
  OAI22X1TS U991 ( .A0(n531), .A1(n503), .B0(n500), .B1(n501), .Y(n1938) );
  OAI22X1TS U992 ( .A0(n13), .A1(n503), .B0(n502), .B1(n501), .Y(n1939) );
  CLKBUFX2TS U993 ( .A(readIn_SOUTH), .Y(n1623) );
  CLKBUFX2TS U994 ( .A(n1623), .Y(n1566) );
  CLKBUFX2TS U995 ( .A(n1911), .Y(n839) );
  CLKBUFX2TS U996 ( .A(n543), .Y(n845) );
  CLKBUFX2TS U997 ( .A(readIn_WEST), .Y(n1631) );
  CLKBUFX2TS U998 ( .A(n1631), .Y(n1616) );
  INVX2TS U999 ( .A(n1911), .Y(n520) );
  NOR4XLTS U1000 ( .A(readReady), .B(n514), .C(n453), .D(n509), .Y(n612) );
  CLKBUFX2TS U1001 ( .A(n612), .Y(n626) );
  CLKBUFX2TS U1002 ( .A(n626), .Y(n806) );
  CLKBUFX2TS U1003 ( .A(n806), .Y(n563) );
  AOI22X1TS U1004 ( .A0(n1566), .A1(n845), .B0(n1616), .B1(n563), .Y(n541) );
  CLKBUFX2TS U1005 ( .A(readIn_NORTH), .Y(n1622) );
  CLKBUFX2TS U1006 ( .A(n1622), .Y(n1565) );
  CLKBUFX2TS U1007 ( .A(n688), .Y(n562) );
  NOR4XLTS U1008 ( .A(n459), .B(n510), .C(n512), .D(n509), .Y(n588) );
  CLKBUFX2TS U1009 ( .A(n588), .Y(n599) );
  CLKBUFX2TS U1010 ( .A(n599), .Y(n774) );
  CLKBUFX2TS U1011 ( .A(n774), .Y(n823) );
  AOI22X1TS U1012 ( .A0(n1565), .A1(n562), .B0(readIn_EAST), .B1(n823), .Y(
        n540) );
  NOR3XLTS U1013 ( .A(n514), .B(n511), .C(n453), .Y(n516) );
  NOR3XLTS U1014 ( .A(selectBit_WEST), .B(n513), .C(n512), .Y(n515) );
  NAND4XLTS U1015 ( .A(n520), .B(n519), .C(n518), .D(n517), .Y(n731) );
  INVX2TS U1016 ( .A(n731), .Y(n521) );
  INVX2TS U1017 ( .A(n521), .Y(n579) );
  INVX2TS U1018 ( .A(n579), .Y(n522) );
  NOR3XLTS U1019 ( .A(n524), .B(n525), .C(n1916), .Y(n715) );
  CLKBUFX2TS U1020 ( .A(n715), .Y(n627) );
  CLKBUFX2TS U1021 ( .A(n627), .Y(n565) );
  NOR3XLTS U1022 ( .A(n527), .B(n1917), .C(n525), .Y(n690) );
  CLKBUFX2TS U1023 ( .A(n690), .Y(n628) );
  CLKBUFX2TS U1024 ( .A(n628), .Y(n564) );
  AOI22X1TS U1025 ( .A0(readOutbuffer[2]), .A1(n565), .B0(readOutbuffer[0]), 
        .B1(n564), .Y(n535) );
  NOR3XLTS U1026 ( .A(n524), .B(n13), .C(n526), .Y(n716) );
  CLKBUFX2TS U1027 ( .A(n716), .Y(n629) );
  CLKBUFX2TS U1028 ( .A(n629), .Y(n567) );
  NOR3XLTS U1029 ( .A(n527), .B(n530), .C(n531), .Y(n691) );
  CLKBUFX2TS U1030 ( .A(n691), .Y(n630) );
  CLKBUFX2TS U1031 ( .A(n630), .Y(n566) );
  AOI22X1TS U1032 ( .A0(readOutbuffer[6]), .A1(n567), .B0(readOutbuffer[4]), 
        .B1(n566), .Y(n534) );
  NOR2XLTS U1033 ( .A(n529), .B(n528), .Y(n717) );
  CLKBUFX2TS U1034 ( .A(n717), .Y(n631) );
  CLKBUFX2TS U1035 ( .A(n631), .Y(n569) );
  NOR3XLTS U1036 ( .A(n530), .B(n529), .C(n1922), .Y(n692) );
  CLKBUFX2TS U1037 ( .A(n692), .Y(n632) );
  CLKBUFX2TS U1038 ( .A(n632), .Y(n568) );
  AOI22X1TS U1039 ( .A0(readOutbuffer[3]), .A1(n569), .B0(readOutbuffer[1]), 
        .B1(n568), .Y(n533) );
  CLKBUFX2TS U1040 ( .A(n833), .Y(n854) );
  NOR3XLTS U1041 ( .A(n1917), .B(n445), .C(n531), .Y(n855) );
  CLKBUFX2TS U1042 ( .A(n855), .Y(n633) );
  CLKBUFX2TS U1043 ( .A(n633), .Y(n570) );
  AOI22X1TS U1044 ( .A0(readOutbuffer[7]), .A1(n854), .B0(readOutbuffer[5]), 
        .B1(n570), .Y(n532) );
  NAND4XLTS U1045 ( .A(n535), .B(n534), .C(n533), .D(n532), .Y(n536) );
  AOI22X1TS U1046 ( .A0(readOut), .A1(n550), .B0(n606), .B1(n536), .Y(n539) );
  INVX2TS U1047 ( .A(n12), .Y(n800) );
  CLKBUFX2TS U1048 ( .A(n774), .Y(n745) );
  AOI22X1TS U1049 ( .A0(writeIn_EAST), .A1(n745), .B0(n542), .B1(n563), .Y(
        n553) );
  CLKBUFX2TS U1050 ( .A(n543), .Y(n668) );
  CLKBUFX2TS U1051 ( .A(n668), .Y(n762) );
  AOI22X1TS U1052 ( .A0(writeIn_NORTH), .A1(n562), .B0(n544), .B1(n762), .Y(
        n552) );
  AOI22X1TS U1053 ( .A0(writeOutbuffer[2]), .A1(n565), .B0(writeOutbuffer[0]), 
        .B1(n564), .Y(n548) );
  AOI22X1TS U1054 ( .A0(writeOutbuffer[6]), .A1(n567), .B0(writeOutbuffer[4]), 
        .B1(n566), .Y(n547) );
  AOI22X1TS U1055 ( .A0(writeOutbuffer[3]), .A1(n569), .B0(writeOutbuffer[1]), 
        .B1(n568), .Y(n546) );
  AOI22X1TS U1056 ( .A0(writeOutbuffer[7]), .A1(n854), .B0(writeOutbuffer[5]), 
        .B1(n570), .Y(n545) );
  NAND4XLTS U1057 ( .A(n548), .B(n547), .C(n546), .D(n545), .Y(n549) );
  AOI22X1TS U1058 ( .A0(writeOut), .A1(n550), .B0(n606), .B1(n549), .Y(n551)
         );
  CLKBUFX2TS U1059 ( .A(requesterAddressIn_NORTH[0]), .Y(n998) );
  CLKBUFX2TS U1060 ( .A(requesterAddressIn_EAST[0]), .Y(n1026) );
  CLKBUFX2TS U1061 ( .A(n1026), .Y(n997) );
  AOI22X1TS U1062 ( .A0(n998), .A1(n562), .B0(n997), .B1(n599), .Y(n561) );
  CLKBUFX2TS U1063 ( .A(requesterAddressIn_SOUTH[0]), .Y(n1027) );
  CLKBUFX2TS U1064 ( .A(n1027), .Y(n999) );
  CLKBUFX2TS U1065 ( .A(n668), .Y(n656) );
  CLKBUFX2TS U1066 ( .A(requesterAddressIn_WEST[0]), .Y(n919) );
  CLKBUFX2TS U1067 ( .A(n919), .Y(n951) );
  AOI22X1TS U1068 ( .A0(n999), .A1(n656), .B0(n951), .B1(n563), .Y(n560) );
  INVX2TS U1069 ( .A(n731), .Y(n683) );
  CLKBUFX2TS U1070 ( .A(n639), .Y(n594) );
  AOI22X1TS U1071 ( .A0(\requesterAddressbuffer[2][0] ), .A1(n565), .B0(
        \requesterAddressbuffer[0][0] ), .B1(n564), .Y(n557) );
  AOI22X1TS U1072 ( .A0(\requesterAddressbuffer[6][0] ), .A1(n567), .B0(
        \requesterAddressbuffer[4][0] ), .B1(n566), .Y(n556) );
  AOI22X1TS U1073 ( .A0(\requesterAddressbuffer[3][0] ), .A1(n569), .B0(
        \requesterAddressbuffer[1][0] ), .B1(n568), .Y(n555) );
  CLKBUFX2TS U1074 ( .A(n793), .Y(n749) );
  CLKBUFX2TS U1075 ( .A(n749), .Y(n600) );
  AOI22X1TS U1076 ( .A0(\requesterAddressbuffer[7][0] ), .A1(n600), .B0(
        \requesterAddressbuffer[5][0] ), .B1(n570), .Y(n554) );
  NAND4XLTS U1077 ( .A(n557), .B(n556), .C(n555), .D(n554), .Y(n558) );
  AOI22X1TS U1078 ( .A0(requesterAddressOut[0]), .A1(n683), .B0(n594), .B1(
        n558), .Y(n559) );
  INVX2TS U1079 ( .A(readRequesterAddress[0]), .Y(n948) );
  INVX2TS U1080 ( .A(n948), .Y(n996) );
  INVX2TS U1081 ( .A(n800), .Y(n595) );
  NAND2X1TS U1082 ( .A(n996), .B(n595), .Y(n607) );
  CLKBUFX2TS U1083 ( .A(requesterAddressIn_NORTH[1]), .Y(n1005) );
  CLKBUFX2TS U1084 ( .A(requesterAddressIn_EAST[1]), .Y(n1032) );
  CLKBUFX2TS U1085 ( .A(n1032), .Y(n1004) );
  AOI22X1TS U1086 ( .A0(n1005), .A1(n562), .B0(n1004), .B1(n588), .Y(n578) );
  CLKBUFX2TS U1087 ( .A(requesterAddressIn_SOUTH[1]), .Y(n1034) );
  CLKBUFX2TS U1088 ( .A(n1034), .Y(n1006) );
  CLKBUFX2TS U1089 ( .A(n543), .Y(n804) );
  CLKBUFX2TS U1090 ( .A(requesterAddressIn_WEST[1]), .Y(n926) );
  CLKBUFX2TS U1091 ( .A(n926), .Y(n957) );
  AOI22X1TS U1092 ( .A0(n1006), .A1(n804), .B0(n957), .B1(n563), .Y(n577) );
  INVX2TS U1093 ( .A(n731), .Y(n780) );
  AOI22X1TS U1094 ( .A0(\requesterAddressbuffer[2][1] ), .A1(n565), .B0(
        \requesterAddressbuffer[0][1] ), .B1(n564), .Y(n574) );
  AOI22X1TS U1095 ( .A0(\requesterAddressbuffer[6][1] ), .A1(n567), .B0(
        \requesterAddressbuffer[4][1] ), .B1(n566), .Y(n573) );
  AOI22X1TS U1096 ( .A0(\requesterAddressbuffer[3][1] ), .A1(n569), .B0(
        \requesterAddressbuffer[1][1] ), .B1(n568), .Y(n572) );
  AOI22X1TS U1097 ( .A0(\requesterAddressbuffer[7][1] ), .A1(n600), .B0(
        \requesterAddressbuffer[5][1] ), .B1(n570), .Y(n571) );
  NAND4XLTS U1098 ( .A(n574), .B(n573), .C(n572), .D(n571), .Y(n575) );
  AOI22X1TS U1099 ( .A0(requesterAddressOut[1]), .A1(n780), .B0(n594), .B1(
        n575), .Y(n576) );
  INVX2TS U1100 ( .A(readRequesterAddress[1]), .Y(n956) );
  INVX2TS U1101 ( .A(n956), .Y(n1640) );
  NAND2X1TS U1102 ( .A(n1640), .B(n595), .Y(n622) );
  CLKBUFX2TS U1103 ( .A(requesterAddressIn_NORTH[2]), .Y(n1012) );
  CLKBUFX2TS U1104 ( .A(n688), .Y(n611) );
  CLKBUFX2TS U1105 ( .A(requesterAddressIn_EAST[2]), .Y(n1038) );
  CLKBUFX2TS U1106 ( .A(n1038), .Y(n1010) );
  AOI22X1TS U1107 ( .A0(n1012), .A1(n611), .B0(n1010), .B1(n588), .Y(n587) );
  CLKBUFX2TS U1108 ( .A(requesterAddressIn_SOUTH[2]), .Y(n1039) );
  CLKBUFX2TS U1109 ( .A(n1039), .Y(n1013) );
  CLKBUFX2TS U1110 ( .A(requesterAddressIn_WEST[2]), .Y(n932) );
  CLKBUFX2TS U1111 ( .A(n932), .Y(n964) );
  AOI22X1TS U1112 ( .A0(n1013), .A1(n656), .B0(n964), .B1(n626), .Y(n586) );
  INVX2TS U1113 ( .A(n579), .Y(n756) );
  CLKBUFX2TS U1114 ( .A(n627), .Y(n613) );
  AOI22X1TS U1115 ( .A0(\requesterAddressbuffer[2][2] ), .A1(n613), .B0(
        \requesterAddressbuffer[0][2] ), .B1(n690), .Y(n583) );
  CLKBUFX2TS U1116 ( .A(n629), .Y(n614) );
  AOI22X1TS U1117 ( .A0(\requesterAddressbuffer[6][2] ), .A1(n614), .B0(
        \requesterAddressbuffer[4][2] ), .B1(n691), .Y(n582) );
  CLKBUFX2TS U1118 ( .A(n631), .Y(n615) );
  AOI22X1TS U1119 ( .A0(\requesterAddressbuffer[3][2] ), .A1(n615), .B0(
        \requesterAddressbuffer[1][2] ), .B1(n692), .Y(n581) );
  CLKBUFX2TS U1120 ( .A(n633), .Y(n616) );
  AOI22X1TS U1121 ( .A0(\requesterAddressbuffer[7][2] ), .A1(n600), .B0(
        \requesterAddressbuffer[5][2] ), .B1(n616), .Y(n580) );
  NAND4XLTS U1122 ( .A(n583), .B(n582), .C(n581), .D(n580), .Y(n584) );
  AOI22X1TS U1123 ( .A0(requesterAddressOut[2]), .A1(n756), .B0(n594), .B1(
        n584), .Y(n585) );
  INVX2TS U1124 ( .A(readRequesterAddress[2]), .Y(n963) );
  INVX2TS U1125 ( .A(n963), .Y(n1648) );
  NAND2X1TS U1126 ( .A(n1648), .B(n595), .Y(n640) );
  CLKBUFX2TS U1127 ( .A(requesterAddressIn_NORTH[3]), .Y(n1021) );
  CLKBUFX2TS U1128 ( .A(requesterAddressIn_EAST[3]), .Y(n1046) );
  CLKBUFX2TS U1129 ( .A(n1046), .Y(n1019) );
  AOI22X1TS U1130 ( .A0(n1021), .A1(n611), .B0(n1019), .B1(n588), .Y(n598) );
  CLKBUFX2TS U1131 ( .A(requesterAddressIn_SOUTH[3]), .Y(n1048) );
  CLKBUFX2TS U1132 ( .A(n1048), .Y(n1022) );
  CLKBUFX2TS U1133 ( .A(requesterAddressIn_WEST[3]), .Y(n942) );
  CLKBUFX2TS U1134 ( .A(n942), .Y(n973) );
  AOI22X1TS U1135 ( .A0(n1022), .A1(n804), .B0(n973), .B1(n612), .Y(n597) );
  AOI22X1TS U1136 ( .A0(\requesterAddressbuffer[2][3] ), .A1(n613), .B0(
        \requesterAddressbuffer[0][3] ), .B1(n690), .Y(n592) );
  AOI22X1TS U1137 ( .A0(\requesterAddressbuffer[6][3] ), .A1(n614), .B0(
        \requesterAddressbuffer[4][3] ), .B1(n691), .Y(n591) );
  AOI22X1TS U1138 ( .A0(\requesterAddressbuffer[3][3] ), .A1(n615), .B0(
        \requesterAddressbuffer[1][3] ), .B1(n692), .Y(n590) );
  CLKBUFX2TS U1139 ( .A(n749), .Y(n645) );
  AOI22X1TS U1140 ( .A0(\requesterAddressbuffer[7][3] ), .A1(n645), .B0(
        \requesterAddressbuffer[5][3] ), .B1(n616), .Y(n589) );
  NAND4XLTS U1141 ( .A(n592), .B(n591), .C(n590), .D(n589), .Y(n593) );
  AOI22X1TS U1142 ( .A0(requesterAddressOut[3]), .A1(n522), .B0(n594), .B1(
        n593), .Y(n596) );
  INVX2TS U1143 ( .A(readRequesterAddress[3]), .Y(n971) );
  INVX2TS U1144 ( .A(n971), .Y(n1656) );
  NAND2X1TS U1145 ( .A(n1656), .B(n595), .Y(n651) );
  CLKBUFX2TS U1146 ( .A(destinationAddressIn_NORTH[0]), .Y(n1666) );
  CLKBUFX2TS U1147 ( .A(destinationAddressIn_EAST[0]), .Y(n1815) );
  CLKBUFX2TS U1148 ( .A(n1815), .Y(n1695) );
  CLKBUFX2TS U1149 ( .A(n599), .Y(n644) );
  AOI22X1TS U1150 ( .A0(n1666), .A1(n611), .B0(n1695), .B1(n644), .Y(n610) );
  CLKBUFX2TS U1151 ( .A(destinationAddressIn_WEST[0]), .Y(n1696) );
  CLKBUFX2TS U1152 ( .A(n1696), .Y(n1760) );
  AOI22X1TS U1153 ( .A0(destinationAddressIn_SOUTH[0]), .A1(n656), .B0(n1760), 
        .B1(n612), .Y(n609) );
  AOI22X1TS U1154 ( .A0(\destinationAddressbuffer[2][0] ), .A1(n613), .B0(
        \destinationAddressbuffer[0][0] ), .B1(n628), .Y(n604) );
  AOI22X1TS U1155 ( .A0(\destinationAddressbuffer[6][0] ), .A1(n614), .B0(
        \destinationAddressbuffer[4][0] ), .B1(n630), .Y(n603) );
  AOI22X1TS U1156 ( .A0(\destinationAddressbuffer[3][0] ), .A1(n615), .B0(
        \destinationAddressbuffer[1][0] ), .B1(n632), .Y(n602) );
  AOI22X1TS U1157 ( .A0(\destinationAddressbuffer[7][0] ), .A1(n600), .B0(
        \destinationAddressbuffer[5][0] ), .B1(n616), .Y(n601) );
  NAND4XLTS U1158 ( .A(n604), .B(n603), .C(n602), .D(n601), .Y(n605) );
  AOI22X1TS U1159 ( .A0(destinationAddressOut[0]), .A1(n683), .B0(n606), .B1(
        n605), .Y(n608) );
  CLKBUFX2TS U1160 ( .A(destinationAddressIn_NORTH[1]), .Y(n1673) );
  CLKBUFX2TS U1161 ( .A(destinationAddressIn_EAST[1]), .Y(n1825) );
  CLKBUFX2TS U1162 ( .A(n1825), .Y(n1704) );
  AOI22X1TS U1163 ( .A0(n1673), .A1(n611), .B0(n1704), .B1(n644), .Y(n625) );
  CLKBUFX2TS U1164 ( .A(destinationAddressIn_WEST[1]), .Y(n1706) );
  CLKBUFX2TS U1165 ( .A(n1706), .Y(n1767) );
  AOI22X1TS U1166 ( .A0(destinationAddressIn_SOUTH[1]), .A1(n804), .B0(n1767), 
        .B1(n612), .Y(n624) );
  AOI22X1TS U1167 ( .A0(\destinationAddressbuffer[2][1] ), .A1(n613), .B0(
        \destinationAddressbuffer[0][1] ), .B1(n628), .Y(n620) );
  AOI22X1TS U1168 ( .A0(\destinationAddressbuffer[6][1] ), .A1(n614), .B0(
        \destinationAddressbuffer[4][1] ), .B1(n630), .Y(n619) );
  AOI22X1TS U1169 ( .A0(\destinationAddressbuffer[3][1] ), .A1(n615), .B0(
        \destinationAddressbuffer[1][1] ), .B1(n632), .Y(n618) );
  AOI22X1TS U1170 ( .A0(\destinationAddressbuffer[7][1] ), .A1(n645), .B0(
        \destinationAddressbuffer[5][1] ), .B1(n616), .Y(n617) );
  NAND4XLTS U1171 ( .A(n620), .B(n619), .C(n618), .D(n617), .Y(n621) );
  AOI22X1TS U1172 ( .A0(destinationAddressOut[1]), .A1(n683), .B0(n639), .B1(
        n621), .Y(n623) );
  CLKBUFX2TS U1173 ( .A(destinationAddressIn_NORTH[2]), .Y(n1680) );
  CLKBUFX2TS U1174 ( .A(n688), .Y(n670) );
  CLKBUFX2TS U1175 ( .A(destinationAddressIn_EAST[2]), .Y(n1836) );
  CLKBUFX2TS U1176 ( .A(n1836), .Y(n1713) );
  AOI22X1TS U1177 ( .A0(n1680), .A1(n670), .B0(n1713), .B1(n644), .Y(n643) );
  CLKBUFX2TS U1178 ( .A(n543), .Y(n784) );
  CLKBUFX2TS U1179 ( .A(destinationAddressIn_WEST[2]), .Y(n1715) );
  CLKBUFX2TS U1180 ( .A(n1715), .Y(n1774) );
  CLKBUFX2TS U1181 ( .A(n626), .Y(n666) );
  AOI22X1TS U1182 ( .A0(destinationAddressIn_SOUTH[2]), .A1(n784), .B0(n1774), 
        .B1(n666), .Y(n642) );
  CLKBUFX2TS U1183 ( .A(n627), .Y(n672) );
  CLKBUFX2TS U1184 ( .A(n628), .Y(n671) );
  AOI22X1TS U1185 ( .A0(\destinationAddressbuffer[2][2] ), .A1(n672), .B0(
        \destinationAddressbuffer[0][2] ), .B1(n671), .Y(n637) );
  CLKBUFX2TS U1186 ( .A(n629), .Y(n674) );
  CLKBUFX2TS U1187 ( .A(n630), .Y(n673) );
  AOI22X1TS U1188 ( .A0(\destinationAddressbuffer[6][2] ), .A1(n674), .B0(
        \destinationAddressbuffer[4][2] ), .B1(n673), .Y(n636) );
  CLKBUFX2TS U1189 ( .A(n631), .Y(n676) );
  CLKBUFX2TS U1190 ( .A(n632), .Y(n675) );
  AOI22X1TS U1191 ( .A0(\destinationAddressbuffer[3][2] ), .A1(n676), .B0(
        \destinationAddressbuffer[1][2] ), .B1(n675), .Y(n635) );
  CLKBUFX2TS U1192 ( .A(n633), .Y(n677) );
  AOI22X1TS U1193 ( .A0(\destinationAddressbuffer[7][2] ), .A1(n645), .B0(
        \destinationAddressbuffer[5][2] ), .B1(n677), .Y(n634) );
  NAND4XLTS U1194 ( .A(n637), .B(n636), .C(n635), .D(n634), .Y(n638) );
  AOI22X1TS U1195 ( .A0(destinationAddressOut[2]), .A1(n522), .B0(n639), .B1(
        n638), .Y(n641) );
  CLKBUFX2TS U1196 ( .A(destinationAddressIn_NORTH[3]), .Y(n1688) );
  CLKBUFX2TS U1197 ( .A(destinationAddressIn_EAST[3]), .Y(n1847) );
  CLKBUFX2TS U1198 ( .A(n1847), .Y(n1721) );
  AOI22X1TS U1199 ( .A0(n1688), .A1(n670), .B0(n1721), .B1(n644), .Y(n654) );
  CLKBUFX2TS U1200 ( .A(destinationAddressIn_WEST[3]), .Y(n1722) );
  CLKBUFX2TS U1201 ( .A(n1722), .Y(n1783) );
  AOI22X1TS U1202 ( .A0(destinationAddressIn_SOUTH[3]), .A1(n784), .B0(n1783), 
        .B1(n666), .Y(n653) );
  AOI22X1TS U1203 ( .A0(\destinationAddressbuffer[2][3] ), .A1(n672), .B0(
        \destinationAddressbuffer[0][3] ), .B1(n671), .Y(n649) );
  AOI22X1TS U1204 ( .A0(\destinationAddressbuffer[6][3] ), .A1(n674), .B0(
        \destinationAddressbuffer[4][3] ), .B1(n673), .Y(n648) );
  AOI22X1TS U1205 ( .A0(\destinationAddressbuffer[3][3] ), .A1(n676), .B0(
        \destinationAddressbuffer[1][3] ), .B1(n675), .Y(n647) );
  AOI22X1TS U1206 ( .A0(\destinationAddressbuffer[7][3] ), .A1(n645), .B0(
        \destinationAddressbuffer[5][3] ), .B1(n677), .Y(n646) );
  NAND4XLTS U1207 ( .A(n649), .B(n648), .C(n647), .D(n646), .Y(n650) );
  AOI22X1TS U1208 ( .A0(destinationAddressOut[3]), .A1(n756), .B0(n1911), .B1(
        n650), .Y(n652) );
  AOI22X1TS U1209 ( .A0(destinationAddressIn_EAST[4]), .A1(n745), .B0(n655), 
        .B1(n666), .Y(n665) );
  AOI22X1TS U1210 ( .A0(destinationAddressIn_NORTH[4]), .A1(n670), .B0(n657), 
        .B1(n656), .Y(n664) );
  INVX2TS U1211 ( .A(n1912), .Y(n765) );
  CLKBUFX2TS U1212 ( .A(n765), .Y(n861) );
  AOI22X1TS U1213 ( .A0(\destinationAddressbuffer[2][4] ), .A1(n672), .B0(
        \destinationAddressbuffer[0][4] ), .B1(n671), .Y(n661) );
  AOI22X1TS U1214 ( .A0(\destinationAddressbuffer[6][4] ), .A1(n674), .B0(
        \destinationAddressbuffer[4][4] ), .B1(n673), .Y(n660) );
  AOI22X1TS U1215 ( .A0(\destinationAddressbuffer[3][4] ), .A1(n676), .B0(
        \destinationAddressbuffer[1][4] ), .B1(n675), .Y(n659) );
  CLKBUFX2TS U1216 ( .A(n749), .Y(n703) );
  AOI22X1TS U1217 ( .A0(\destinationAddressbuffer[7][4] ), .A1(n703), .B0(
        \destinationAddressbuffer[5][4] ), .B1(n677), .Y(n658) );
  NAND4XLTS U1218 ( .A(n661), .B(n660), .C(n659), .D(n658), .Y(n662) );
  AOI22X1TS U1219 ( .A0(destinationAddressOut[4]), .A1(n780), .B0(n861), .B1(
        n662), .Y(n663) );
  CLKBUFX2TS U1220 ( .A(n774), .Y(n761) );
  AOI22X1TS U1221 ( .A0(destinationAddressIn_EAST[5]), .A1(n761), .B0(n667), 
        .B1(n666), .Y(n686) );
  CLKBUFX2TS U1222 ( .A(n668), .Y(n746) );
  AOI22X1TS U1223 ( .A0(destinationAddressIn_NORTH[5]), .A1(n670), .B0(n669), 
        .B1(n746), .Y(n685) );
  AOI22X1TS U1224 ( .A0(\destinationAddressbuffer[2][5] ), .A1(n672), .B0(
        \destinationAddressbuffer[0][5] ), .B1(n671), .Y(n681) );
  AOI22X1TS U1225 ( .A0(\destinationAddressbuffer[6][5] ), .A1(n674), .B0(
        \destinationAddressbuffer[4][5] ), .B1(n673), .Y(n680) );
  AOI22X1TS U1226 ( .A0(\destinationAddressbuffer[3][5] ), .A1(n676), .B0(
        \destinationAddressbuffer[1][5] ), .B1(n675), .Y(n679) );
  AOI22X1TS U1227 ( .A0(\destinationAddressbuffer[7][5] ), .A1(n703), .B0(
        \destinationAddressbuffer[5][5] ), .B1(n677), .Y(n678) );
  NAND4XLTS U1228 ( .A(n681), .B(n680), .C(n679), .D(n678), .Y(n682) );
  AOI22X1TS U1229 ( .A0(destinationAddressOut[5]), .A1(n683), .B0(n861), .B1(
        n682), .Y(n684) );
  CLKBUFX2TS U1230 ( .A(n806), .Y(n726) );
  AOI22X1TS U1231 ( .A0(destinationAddressIn_EAST[6]), .A1(n761), .B0(n687), 
        .B1(n726), .Y(n700) );
  CLKBUFX2TS U1232 ( .A(n688), .Y(n805) );
  CLKBUFX2TS U1233 ( .A(n805), .Y(n729) );
  AOI22X1TS U1234 ( .A0(destinationAddressIn_NORTH[6]), .A1(n729), .B0(n689), 
        .B1(n746), .Y(n699) );
  CLKBUFX2TS U1235 ( .A(n690), .Y(n807) );
  CLKBUFX2TS U1236 ( .A(n807), .Y(n732) );
  AOI22X1TS U1237 ( .A0(\destinationAddressbuffer[2][6] ), .A1(n715), .B0(
        \destinationAddressbuffer[0][6] ), .B1(n732), .Y(n696) );
  CLKBUFX2TS U1238 ( .A(n691), .Y(n809) );
  CLKBUFX2TS U1239 ( .A(n809), .Y(n733) );
  AOI22X1TS U1240 ( .A0(\destinationAddressbuffer[6][6] ), .A1(n716), .B0(
        \destinationAddressbuffer[4][6] ), .B1(n733), .Y(n695) );
  CLKBUFX2TS U1241 ( .A(n692), .Y(n811) );
  CLKBUFX2TS U1242 ( .A(n811), .Y(n734) );
  AOI22X1TS U1243 ( .A0(\destinationAddressbuffer[3][6] ), .A1(n717), .B0(
        \destinationAddressbuffer[1][6] ), .B1(n734), .Y(n694) );
  CLKBUFX2TS U1244 ( .A(n855), .Y(n824) );
  CLKBUFX2TS U1245 ( .A(n824), .Y(n735) );
  AOI22X1TS U1246 ( .A0(\destinationAddressbuffer[7][6] ), .A1(n703), .B0(
        \destinationAddressbuffer[5][6] ), .B1(n735), .Y(n693) );
  NAND4XLTS U1247 ( .A(n696), .B(n695), .C(n694), .D(n693), .Y(n697) );
  AOI22X1TS U1248 ( .A0(destinationAddressOut[6]), .A1(n780), .B0(n861), .B1(
        n697), .Y(n698) );
  AOI22X1TS U1249 ( .A0(destinationAddressIn_EAST[7]), .A1(n823), .B0(n701), 
        .B1(n726), .Y(n711) );
  AOI22X1TS U1250 ( .A0(destinationAddressIn_NORTH[7]), .A1(n729), .B0(n702), 
        .B1(n762), .Y(n710) );
  CLKBUFX2TS U1251 ( .A(n765), .Y(n755) );
  AOI22X1TS U1252 ( .A0(\destinationAddressbuffer[2][7] ), .A1(n715), .B0(
        \destinationAddressbuffer[0][7] ), .B1(n732), .Y(n707) );
  AOI22X1TS U1253 ( .A0(\destinationAddressbuffer[6][7] ), .A1(n716), .B0(
        \destinationAddressbuffer[4][7] ), .B1(n733), .Y(n706) );
  AOI22X1TS U1254 ( .A0(\destinationAddressbuffer[3][7] ), .A1(n717), .B0(
        \destinationAddressbuffer[1][7] ), .B1(n734), .Y(n705) );
  AOI22X1TS U1255 ( .A0(\destinationAddressbuffer[7][7] ), .A1(n703), .B0(
        \destinationAddressbuffer[5][7] ), .B1(n735), .Y(n704) );
  NAND4XLTS U1256 ( .A(n707), .B(n706), .C(n705), .D(n704), .Y(n708) );
  AOI22X1TS U1257 ( .A0(destinationAddressOut[7]), .A1(n521), .B0(n755), .B1(
        n708), .Y(n709) );
  AOI22X1TS U1258 ( .A0(destinationAddressIn_EAST[8]), .A1(n745), .B0(n712), 
        .B1(n726), .Y(n725) );
  AOI22X1TS U1259 ( .A0(n714), .A1(n729), .B0(n713), .B1(n746), .Y(n724) );
  CLKBUFX2TS U1260 ( .A(n715), .Y(n808) );
  AOI22X1TS U1261 ( .A0(\destinationAddressbuffer[2][8] ), .A1(n808), .B0(
        \destinationAddressbuffer[0][8] ), .B1(n732), .Y(n721) );
  CLKBUFX2TS U1262 ( .A(n716), .Y(n810) );
  AOI22X1TS U1263 ( .A0(\destinationAddressbuffer[6][8] ), .A1(n810), .B0(
        \destinationAddressbuffer[4][8] ), .B1(n733), .Y(n720) );
  CLKBUFX2TS U1264 ( .A(n717), .Y(n812) );
  AOI22X1TS U1265 ( .A0(\destinationAddressbuffer[3][8] ), .A1(n812), .B0(
        \destinationAddressbuffer[1][8] ), .B1(n734), .Y(n719) );
  AOI22X1TS U1266 ( .A0(\destinationAddressbuffer[7][8] ), .A1(n813), .B0(
        \destinationAddressbuffer[5][8] ), .B1(n735), .Y(n718) );
  NAND4XLTS U1267 ( .A(n721), .B(n720), .C(n719), .D(n718), .Y(n722) );
  AOI22X1TS U1268 ( .A0(destinationAddressOut[8]), .A1(n756), .B0(n755), .B1(
        n722), .Y(n723) );
  AOI22X1TS U1269 ( .A0(destinationAddressIn_EAST[9]), .A1(n761), .B0(n727), 
        .B1(n726), .Y(n743) );
  AOI22X1TS U1270 ( .A0(n730), .A1(n729), .B0(n728), .B1(n762), .Y(n742) );
  INVX2TS U1271 ( .A(n731), .Y(n840) );
  AOI22X1TS U1272 ( .A0(\destinationAddressbuffer[2][9] ), .A1(n808), .B0(
        \destinationAddressbuffer[0][9] ), .B1(n732), .Y(n739) );
  AOI22X1TS U1273 ( .A0(\destinationAddressbuffer[6][9] ), .A1(n810), .B0(
        \destinationAddressbuffer[4][9] ), .B1(n733), .Y(n738) );
  AOI22X1TS U1274 ( .A0(\destinationAddressbuffer[3][9] ), .A1(n812), .B0(
        \destinationAddressbuffer[1][9] ), .B1(n734), .Y(n737) );
  AOI22X1TS U1275 ( .A0(\destinationAddressbuffer[7][9] ), .A1(n813), .B0(
        \destinationAddressbuffer[5][9] ), .B1(n735), .Y(n736) );
  NAND4XLTS U1276 ( .A(n739), .B(n738), .C(n737), .D(n736), .Y(n740) );
  AOI22X1TS U1277 ( .A0(destinationAddressOut[9]), .A1(n840), .B0(n755), .B1(
        n740), .Y(n741) );
  CLKBUFX2TS U1278 ( .A(n806), .Y(n785) );
  AOI22X1TS U1279 ( .A0(destinationAddressIn_EAST[10]), .A1(n745), .B0(n744), 
        .B1(n785), .Y(n759) );
  CLKBUFX2TS U1280 ( .A(n805), .Y(n786) );
  AOI22X1TS U1281 ( .A0(n748), .A1(n786), .B0(n747), .B1(n746), .Y(n758) );
  CLKBUFX2TS U1282 ( .A(n808), .Y(n787) );
  CLKBUFX2TS U1283 ( .A(n807), .Y(n788) );
  AOI22X1TS U1284 ( .A0(\destinationAddressbuffer[2][10] ), .A1(n787), .B0(
        \destinationAddressbuffer[0][10] ), .B1(n788), .Y(n753) );
  CLKBUFX2TS U1285 ( .A(n810), .Y(n789) );
  CLKBUFX2TS U1286 ( .A(n809), .Y(n790) );
  AOI22X1TS U1287 ( .A0(\destinationAddressbuffer[6][10] ), .A1(n789), .B0(
        \destinationAddressbuffer[4][10] ), .B1(n790), .Y(n752) );
  CLKBUFX2TS U1288 ( .A(n812), .Y(n791) );
  CLKBUFX2TS U1289 ( .A(n811), .Y(n792) );
  AOI22X1TS U1290 ( .A0(\destinationAddressbuffer[3][10] ), .A1(n791), .B0(
        \destinationAddressbuffer[1][10] ), .B1(n792), .Y(n751) );
  CLKBUFX2TS U1291 ( .A(n824), .Y(n794) );
  AOI22X1TS U1292 ( .A0(\destinationAddressbuffer[7][10] ), .A1(n749), .B0(
        \destinationAddressbuffer[5][10] ), .B1(n794), .Y(n750) );
  NAND4XLTS U1293 ( .A(n753), .B(n752), .C(n751), .D(n750), .Y(n754) );
  AOI22X1TS U1294 ( .A0(destinationAddressOut[10]), .A1(n756), .B0(n755), .B1(
        n754), .Y(n757) );
  AOI22X1TS U1295 ( .A0(destinationAddressIn_EAST[11]), .A1(n761), .B0(n760), 
        .B1(n785), .Y(n773) );
  AOI22X1TS U1296 ( .A0(n764), .A1(n786), .B0(n763), .B1(n762), .Y(n772) );
  CLKBUFX2TS U1297 ( .A(n765), .Y(n819) );
  AOI22X1TS U1298 ( .A0(\destinationAddressbuffer[2][11] ), .A1(n787), .B0(
        \destinationAddressbuffer[0][11] ), .B1(n788), .Y(n769) );
  AOI22X1TS U1299 ( .A0(\destinationAddressbuffer[6][11] ), .A1(n789), .B0(
        \destinationAddressbuffer[4][11] ), .B1(n790), .Y(n768) );
  AOI22X1TS U1300 ( .A0(\destinationAddressbuffer[3][11] ), .A1(n791), .B0(
        \destinationAddressbuffer[1][11] ), .B1(n792), .Y(n767) );
  AOI22X1TS U1301 ( .A0(\destinationAddressbuffer[7][11] ), .A1(n793), .B0(
        \destinationAddressbuffer[5][11] ), .B1(n794), .Y(n766) );
  NAND4XLTS U1302 ( .A(n769), .B(n768), .C(n767), .D(n766), .Y(n770) );
  AOI22X1TS U1303 ( .A0(destinationAddressOut[11]), .A1(n521), .B0(n819), .B1(
        n770), .Y(n771) );
  CLKBUFX2TS U1304 ( .A(dataIn_SOUTH[0]), .Y(n1501) );
  CLKBUFX2TS U1305 ( .A(dataIn_EAST[0]), .Y(n1460) );
  CLKBUFX2TS U1306 ( .A(n1460), .Y(n1108) );
  CLKBUFX2TS U1307 ( .A(n774), .Y(n844) );
  AOI22X1TS U1308 ( .A0(n1501), .A1(n784), .B0(n1108), .B1(n844), .Y(n783) );
  CLKBUFX2TS U1309 ( .A(dataIn_WEST[0]), .Y(n1499) );
  CLKBUFX2TS U1310 ( .A(n1499), .Y(n1392) );
  AOI22X1TS U1311 ( .A0(dataIn_NORTH[0]), .A1(n786), .B0(n1392), .B1(n785), 
        .Y(n782) );
  AOI22X1TS U1312 ( .A0(\dataoutbuffer[0][0] ), .A1(n788), .B0(
        \dataoutbuffer[2][0] ), .B1(n787), .Y(n778) );
  AOI22X1TS U1313 ( .A0(\dataoutbuffer[4][0] ), .A1(n790), .B0(
        \dataoutbuffer[6][0] ), .B1(n789), .Y(n777) );
  AOI22X1TS U1314 ( .A0(\dataoutbuffer[1][0] ), .A1(n792), .B0(
        \dataoutbuffer[3][0] ), .B1(n791), .Y(n776) );
  AOI22X1TS U1315 ( .A0(\dataoutbuffer[5][0] ), .A1(n794), .B0(
        \dataoutbuffer[7][0] ), .B1(n854), .Y(n775) );
  NAND4XLTS U1316 ( .A(n778), .B(n777), .C(n776), .D(n775), .Y(n779) );
  AOI22X1TS U1317 ( .A0(dataOut[0]), .A1(n780), .B0(n819), .B1(n779), .Y(n781)
         );
  CLKBUFX2TS U1318 ( .A(dataIn_SOUTH[1]), .Y(n1509) );
  CLKBUFX2TS U1319 ( .A(dataIn_EAST[1]), .Y(n1468) );
  CLKBUFX2TS U1320 ( .A(n1468), .Y(n1339) );
  AOI22X1TS U1321 ( .A0(n1509), .A1(n784), .B0(n1339), .B1(n823), .Y(n803) );
  CLKBUFX2TS U1322 ( .A(dataIn_WEST[1]), .Y(n1506) );
  CLKBUFX2TS U1323 ( .A(n1506), .Y(n1398) );
  AOI22X1TS U1324 ( .A0(dataIn_NORTH[1]), .A1(n786), .B0(n1398), .B1(n785), 
        .Y(n802) );
  AOI22X1TS U1325 ( .A0(\dataoutbuffer[0][1] ), .A1(n788), .B0(
        \dataoutbuffer[2][1] ), .B1(n787), .Y(n798) );
  AOI22X1TS U1326 ( .A0(\dataoutbuffer[4][1] ), .A1(n790), .B0(
        \dataoutbuffer[6][1] ), .B1(n789), .Y(n797) );
  AOI22X1TS U1327 ( .A0(\dataoutbuffer[1][1] ), .A1(n792), .B0(
        \dataoutbuffer[3][1] ), .B1(n791), .Y(n796) );
  AOI22X1TS U1328 ( .A0(\dataoutbuffer[5][1] ), .A1(n794), .B0(
        \dataoutbuffer[7][1] ), .B1(n793), .Y(n795) );
  NAND4XLTS U1329 ( .A(n798), .B(n797), .C(n796), .D(n795), .Y(n799) );
  AOI22X1TS U1330 ( .A0(dataOut[1]), .A1(n522), .B0(n819), .B1(n799), .Y(n801)
         );
  CLKBUFX2TS U1331 ( .A(dataIn_SOUTH[2]), .Y(n1515) );
  CLKBUFX2TS U1332 ( .A(dataIn_EAST[2]), .Y(n1474) );
  CLKBUFX2TS U1333 ( .A(n1474), .Y(n1345) );
  AOI22X1TS U1334 ( .A0(n1515), .A1(n804), .B0(n1345), .B1(n844), .Y(n822) );
  CLKBUFX2TS U1335 ( .A(n805), .Y(n847) );
  CLKBUFX2TS U1336 ( .A(dataIn_WEST[2]), .Y(n1513) );
  CLKBUFX2TS U1337 ( .A(n1513), .Y(n1403) );
  CLKBUFX2TS U1338 ( .A(n806), .Y(n846) );
  AOI22X1TS U1339 ( .A0(dataIn_NORTH[2]), .A1(n847), .B0(n1403), .B1(n846), 
        .Y(n821) );
  CLKBUFX2TS U1340 ( .A(n807), .Y(n849) );
  CLKBUFX2TS U1341 ( .A(n808), .Y(n848) );
  AOI22X1TS U1342 ( .A0(\dataoutbuffer[0][2] ), .A1(n849), .B0(
        \dataoutbuffer[2][2] ), .B1(n848), .Y(n817) );
  CLKBUFX2TS U1343 ( .A(n809), .Y(n851) );
  CLKBUFX2TS U1344 ( .A(n810), .Y(n850) );
  AOI22X1TS U1345 ( .A0(\dataoutbuffer[4][2] ), .A1(n851), .B0(
        \dataoutbuffer[6][2] ), .B1(n850), .Y(n816) );
  CLKBUFX2TS U1346 ( .A(n811), .Y(n853) );
  CLKBUFX2TS U1347 ( .A(n812), .Y(n852) );
  AOI22X1TS U1348 ( .A0(\dataoutbuffer[1][2] ), .A1(n853), .B0(
        \dataoutbuffer[3][2] ), .B1(n852), .Y(n815) );
  AOI22X1TS U1349 ( .A0(\dataoutbuffer[5][2] ), .A1(n824), .B0(
        \dataoutbuffer[7][2] ), .B1(n813), .Y(n814) );
  NAND4XLTS U1350 ( .A(n817), .B(n816), .C(n815), .D(n814), .Y(n818) );
  AOI22X1TS U1351 ( .A0(dataOut[2]), .A1(n840), .B0(n819), .B1(n818), .Y(n820)
         );
  INVX2TS U1352 ( .A(n12), .Y(n862) );
  CLKBUFX2TS U1353 ( .A(dataIn_SOUTH[3]), .Y(n1522) );
  CLKBUFX2TS U1354 ( .A(dataIn_EAST[3]), .Y(n1480) );
  CLKBUFX2TS U1355 ( .A(n1480), .Y(n1350) );
  AOI22X1TS U1356 ( .A0(n1522), .A1(n845), .B0(n1350), .B1(n823), .Y(n832) );
  CLKBUFX2TS U1357 ( .A(dataIn_WEST[3]), .Y(n1520) );
  CLKBUFX2TS U1358 ( .A(n1520), .Y(n1408) );
  AOI22X1TS U1359 ( .A0(dataIn_NORTH[3]), .A1(n847), .B0(n1408), .B1(n846), 
        .Y(n831) );
  AOI22X1TS U1360 ( .A0(\dataoutbuffer[0][3] ), .A1(n849), .B0(
        \dataoutbuffer[2][3] ), .B1(n848), .Y(n828) );
  AOI22X1TS U1361 ( .A0(\dataoutbuffer[4][3] ), .A1(n851), .B0(
        \dataoutbuffer[6][3] ), .B1(n850), .Y(n827) );
  AOI22X1TS U1362 ( .A0(\dataoutbuffer[1][3] ), .A1(n853), .B0(
        \dataoutbuffer[3][3] ), .B1(n852), .Y(n826) );
  AOI22X1TS U1363 ( .A0(\dataoutbuffer[5][3] ), .A1(n824), .B0(
        \dataoutbuffer[7][3] ), .B1(n833), .Y(n825) );
  NAND4XLTS U1364 ( .A(n828), .B(n827), .C(n826), .D(n825), .Y(n829) );
  AOI22X1TS U1365 ( .A0(dataOut[3]), .A1(n840), .B0(n839), .B1(n829), .Y(n830)
         );
  CLKBUFX2TS U1366 ( .A(dataIn_SOUTH[4]), .Y(n1531) );
  CLKBUFX2TS U1367 ( .A(dataIn_EAST[4]), .Y(n1485) );
  CLKBUFX2TS U1368 ( .A(n1485), .Y(n1355) );
  AOI22X1TS U1369 ( .A0(n1531), .A1(n845), .B0(n1355), .B1(n844), .Y(n843) );
  CLKBUFX2TS U1370 ( .A(dataIn_WEST[4]), .Y(n1527) );
  CLKBUFX2TS U1371 ( .A(n1527), .Y(n1412) );
  AOI22X1TS U1372 ( .A0(dataIn_NORTH[4]), .A1(n847), .B0(n1412), .B1(n846), 
        .Y(n842) );
  AOI22X1TS U1373 ( .A0(\dataoutbuffer[0][4] ), .A1(n849), .B0(
        \dataoutbuffer[2][4] ), .B1(n848), .Y(n837) );
  AOI22X1TS U1374 ( .A0(\dataoutbuffer[4][4] ), .A1(n851), .B0(
        \dataoutbuffer[6][4] ), .B1(n850), .Y(n836) );
  AOI22X1TS U1375 ( .A0(\dataoutbuffer[1][4] ), .A1(n853), .B0(
        \dataoutbuffer[3][4] ), .B1(n852), .Y(n835) );
  AOI22X1TS U1376 ( .A0(\dataoutbuffer[5][4] ), .A1(n855), .B0(
        \dataoutbuffer[7][4] ), .B1(n833), .Y(n834) );
  NAND4XLTS U1377 ( .A(n837), .B(n836), .C(n835), .D(n834), .Y(n838) );
  AOI22X1TS U1378 ( .A0(dataOut[4]), .A1(n840), .B0(n839), .B1(n838), .Y(n841)
         );
  CLKBUFX2TS U1379 ( .A(dataIn_SOUTH[5]), .Y(n1538) );
  CLKBUFX2TS U1380 ( .A(dataIn_EAST[5]), .Y(n1493) );
  CLKBUFX2TS U1381 ( .A(n1493), .Y(n1361) );
  AOI22X1TS U1382 ( .A0(n1538), .A1(n845), .B0(n1361), .B1(n844), .Y(n865) );
  CLKBUFX2TS U1383 ( .A(dataIn_WEST[5]), .Y(n1536) );
  CLKBUFX2TS U1384 ( .A(n1536), .Y(n1420) );
  AOI22X1TS U1385 ( .A0(dataIn_NORTH[5]), .A1(n847), .B0(n1420), .B1(n846), 
        .Y(n864) );
  AOI22X1TS U1386 ( .A0(\dataoutbuffer[0][5] ), .A1(n849), .B0(
        \dataoutbuffer[2][5] ), .B1(n848), .Y(n859) );
  AOI22X1TS U1387 ( .A0(\dataoutbuffer[4][5] ), .A1(n851), .B0(
        \dataoutbuffer[6][5] ), .B1(n850), .Y(n858) );
  AOI22X1TS U1388 ( .A0(\dataoutbuffer[1][5] ), .A1(n853), .B0(
        \dataoutbuffer[3][5] ), .B1(n852), .Y(n857) );
  AOI22X1TS U1389 ( .A0(\dataoutbuffer[5][5] ), .A1(n855), .B0(
        \dataoutbuffer[7][5] ), .B1(n854), .Y(n856) );
  NAND4XLTS U1390 ( .A(n859), .B(n858), .C(n857), .D(n856), .Y(n860) );
  AOI22X1TS U1391 ( .A0(dataOut[5]), .A1(n522), .B0(n861), .B1(n860), .Y(n863)
         );
  INVX2TS U1392 ( .A(n948), .Y(n1758) );
  AOI22X1TS U1393 ( .A0(n1758), .A1(n1635), .B0(n1655), .B1(
        \requesterAddressbuffer[7][0] ), .Y(n868) );
  CLKBUFX2TS U1394 ( .A(n1026), .Y(n918) );
  AOI22X1TS U1395 ( .A0(n76), .A1(n951), .B0(n1649), .B1(n918), .Y(n867) );
  CLKBUFX2TS U1396 ( .A(n1027), .Y(n921) );
  CLKBUFX2TS U1397 ( .A(n998), .Y(n952) );
  AOI22X1TS U1398 ( .A0(n46), .A1(n921), .B0(n869), .B1(n952), .Y(n866) );
  INVX2TS U1399 ( .A(n876), .Y(n1641) );
  INVX2TS U1400 ( .A(n1498), .Y(n1535) );
  AOI22X1TS U1401 ( .A0(n1641), .A1(n1640), .B0(n1535), .B1(
        \requesterAddressbuffer[7][1] ), .Y(n872) );
  INVX2TS U1402 ( .A(n878), .Y(n1636) );
  CLKBUFX2TS U1403 ( .A(n1032), .Y(n925) );
  AOI22X1TS U1404 ( .A0(n1528), .A1(n957), .B0(n1636), .B1(n925), .Y(n871) );
  CLKBUFX2TS U1405 ( .A(n1034), .Y(n927) );
  CLKBUFX2TS U1406 ( .A(n1005), .Y(n959) );
  AOI22X1TS U1407 ( .A0(n1660), .A1(n927), .B0(n869), .B1(n959), .Y(n870) );
  AOI22X1TS U1408 ( .A0(n34), .A1(n1648), .B0(n1535), .B1(
        \requesterAddressbuffer[7][2] ), .Y(n875) );
  CLKBUFX2TS U1409 ( .A(n1038), .Y(n931) );
  AOI22X1TS U1410 ( .A0(n1650), .A1(n964), .B0(n32), .B1(n931), .Y(n874) );
  CLKBUFX2TS U1411 ( .A(n1039), .Y(n933) );
  CLKBUFX2TS U1412 ( .A(n1012), .Y(n967) );
  AOI22X1TS U1413 ( .A0(n58), .A1(n933), .B0(n53), .B1(n967), .Y(n873) );
  INVX2TS U1414 ( .A(n876), .Y(n1657) );
  INVX2TS U1415 ( .A(n877), .Y(n1647) );
  AOI22X1TS U1416 ( .A0(n1657), .A1(n1656), .B0(n1647), .B1(
        \requesterAddressbuffer[7][3] ), .Y(n882) );
  INVX2TS U1417 ( .A(n878), .Y(n1658) );
  CLKBUFX2TS U1418 ( .A(n1046), .Y(n941) );
  AOI22X1TS U1419 ( .A0(n1528), .A1(n973), .B0(n1658), .B1(n941), .Y(n881) );
  INVX2TS U1420 ( .A(n879), .Y(n1539) );
  CLKBUFX2TS U1421 ( .A(n1048), .Y(n944) );
  CLKBUFX2TS U1422 ( .A(n1021), .Y(n974) );
  AOI22X1TS U1423 ( .A0(n1539), .A1(n944), .B0(n1530), .B1(n974), .Y(n880) );
  INVX2TS U1424 ( .A(n948), .Y(n1814) );
  AOI22X1TS U1425 ( .A0(n1814), .A1(n1664), .B0(n1685), .B1(
        \requesterAddressbuffer[6][0] ), .Y(n885) );
  INVX2TS U1426 ( .A(n1473), .Y(n1672) );
  AOI22X1TS U1427 ( .A0(n919), .A1(n1687), .B0(n918), .B1(n1672), .Y(n884) );
  AOI22X1TS U1428 ( .A0(n921), .A1(n1463), .B0(n952), .B1(n1464), .Y(n883) );
  INVX2TS U1429 ( .A(n956), .Y(n1736) );
  INVX2TS U1430 ( .A(n893), .Y(n1671) );
  INVX2TS U1431 ( .A(n1459), .Y(n1492) );
  AOI22X1TS U1432 ( .A0(n1736), .A1(n1671), .B0(n1492), .B1(
        \requesterAddressbuffer[6][1] ), .Y(n889) );
  INVX2TS U1433 ( .A(n1473), .Y(n1679) );
  AOI22X1TS U1434 ( .A0(n926), .A1(n1486), .B0(n925), .B1(n1679), .Y(n888) );
  INVX2TS U1435 ( .A(n897), .Y(n1488) );
  AOI22X1TS U1436 ( .A0(n927), .A1(n1488), .B0(n959), .B1(n93), .Y(n887) );
  INVX2TS U1437 ( .A(n963), .Y(n1742) );
  AOI22X1TS U1438 ( .A0(n1742), .A1(n1664), .B0(n1492), .B1(
        \requesterAddressbuffer[6][2] ), .Y(n892) );
  AOI22X1TS U1439 ( .A0(n932), .A1(n1461), .B0(n931), .B1(n896), .Y(n891) );
  AOI22X1TS U1440 ( .A0(n933), .A1(n98), .B0(n967), .B1(n102), .Y(n890) );
  INVX2TS U1441 ( .A(n971), .Y(n1750) );
  INVX2TS U1442 ( .A(n893), .Y(n1686) );
  INVX2TS U1443 ( .A(n894), .Y(n1678) );
  AOI22X1TS U1444 ( .A0(n1750), .A1(n1686), .B0(n1678), .B1(
        \requesterAddressbuffer[6][3] ), .Y(n900) );
  INVX2TS U1445 ( .A(n895), .Y(n1486) );
  AOI22X1TS U1446 ( .A0(n942), .A1(n1486), .B0(n941), .B1(n896), .Y(n899) );
  INVX2TS U1447 ( .A(n897), .Y(n1681) );
  AOI22X1TS U1448 ( .A0(n944), .A1(n1681), .B0(n974), .B1(n1667), .Y(n898) );
  AOI22X1TS U1449 ( .A0(n996), .A1(n1694), .B0(n1719), .B1(
        \requesterAddressbuffer[5][0] ), .Y(n904) );
  INVX2TS U1450 ( .A(n1436), .Y(n1705) );
  AOI22X1TS U1451 ( .A0(n919), .A1(n1723), .B0(n918), .B1(n1705), .Y(n903) );
  INVX2TS U1452 ( .A(n901), .Y(n1724) );
  AOI22X1TS U1453 ( .A0(n921), .A1(n1724), .B0(requesterAddressIn_NORTH[0]), 
        .B1(n1438), .Y(n902) );
  INVX2TS U1454 ( .A(n9), .Y(n1703) );
  INVX2TS U1455 ( .A(n1424), .Y(n1454) );
  AOI22X1TS U1456 ( .A0(n1640), .A1(n1703), .B0(n1454), .B1(
        \requesterAddressbuffer[5][1] ), .Y(n907) );
  INVX2TS U1457 ( .A(n1436), .Y(n1714) );
  AOI22X1TS U1458 ( .A0(n926), .A1(n1447), .B0(n925), .B1(n1714), .Y(n906) );
  AOI22X1TS U1459 ( .A0(n927), .A1(n1698), .B0(requesterAddressIn_NORTH[1]), 
        .B1(n1699), .Y(n905) );
  INVX2TS U1460 ( .A(n9), .Y(n1712) );
  AOI22X1TS U1461 ( .A0(n1648), .A1(n1712), .B0(n1454), .B1(
        \requesterAddressbuffer[5][2] ), .Y(n911) );
  AOI22X1TS U1462 ( .A0(n932), .A1(n1425), .B0(n931), .B1(n914), .Y(n910) );
  AOI22X1TS U1463 ( .A0(n933), .A1(n1426), .B0(requesterAddressIn_NORTH[2]), 
        .B1(n908), .Y(n909) );
  INVX2TS U1464 ( .A(n9), .Y(n1720) );
  INVX2TS U1465 ( .A(n912), .Y(n1711) );
  AOI22X1TS U1466 ( .A0(n1656), .A1(n1720), .B0(n1711), .B1(
        \requesterAddressbuffer[5][3] ), .Y(n917) );
  INVX2TS U1467 ( .A(n913), .Y(n1447) );
  AOI22X1TS U1468 ( .A0(n942), .A1(n1447), .B0(n941), .B1(n914), .Y(n916) );
  AOI22X1TS U1469 ( .A0(n944), .A1(n232), .B0(requesterAddressIn_NORTH[3]), 
        .B1(n1450), .Y(n915) );
  AOI22X1TS U1470 ( .A0(n996), .A1(n1728), .B0(n1748), .B1(
        \requesterAddressbuffer[4][0] ), .Y(n924) );
  INVX2TS U1471 ( .A(n1402), .Y(n1737) );
  AOI22X1TS U1472 ( .A0(n919), .A1(n1751), .B0(n918), .B1(n1737), .Y(n923) );
  AOI22X1TS U1473 ( .A0(n921), .A1(n1744), .B0(requesterAddressIn_NORTH[0]), 
        .B1(n920), .Y(n922) );
  INVX2TS U1474 ( .A(n956), .Y(n1866) );
  INVX2TS U1475 ( .A(n937), .Y(n1735) );
  INVX2TS U1476 ( .A(n1391), .Y(n1419) );
  AOI22X1TS U1477 ( .A0(n1866), .A1(n1735), .B0(n1419), .B1(
        \requesterAddressbuffer[4][1] ), .Y(n930) );
  INVX2TS U1478 ( .A(n1402), .Y(n1743) );
  AOI22X1TS U1479 ( .A0(n926), .A1(n1413), .B0(n925), .B1(n1743), .Y(n929) );
  AOI22X1TS U1480 ( .A0(n927), .A1(n1415), .B0(requesterAddressIn_NORTH[1]), 
        .B1(n1752), .Y(n928) );
  INVX2TS U1481 ( .A(n963), .Y(n1876) );
  AOI22X1TS U1482 ( .A0(n1876), .A1(n1728), .B0(n1419), .B1(
        \requesterAddressbuffer[4][2] ), .Y(n936) );
  AOI22X1TS U1483 ( .A0(n932), .A1(n1393), .B0(n931), .B1(n940), .Y(n935) );
  AOI22X1TS U1484 ( .A0(n933), .A1(n1753), .B0(requesterAddressIn_NORTH[2]), 
        .B1(n1752), .Y(n934) );
  INVX2TS U1485 ( .A(n971), .Y(n1886) );
  INVX2TS U1486 ( .A(n937), .Y(n1749) );
  INVX2TS U1487 ( .A(n938), .Y(n1741) );
  AOI22X1TS U1488 ( .A0(n1886), .A1(n1749), .B0(n1741), .B1(
        \requesterAddressbuffer[4][3] ), .Y(n947) );
  INVX2TS U1489 ( .A(n939), .Y(n1413) );
  AOI22X1TS U1490 ( .A0(n942), .A1(n1413), .B0(n941), .B1(n940), .Y(n946) );
  INVX2TS U1491 ( .A(n943), .Y(n1731) );
  AOI22X1TS U1492 ( .A0(n944), .A1(n1731), .B0(requesterAddressIn_NORTH[3]), 
        .B1(n1394), .Y(n945) );
  INVX2TS U1493 ( .A(n948), .Y(n1856) );
  AOI22X1TS U1494 ( .A0(n1856), .A1(n1757), .B0(n1780), .B1(
        \requesterAddressbuffer[3][0] ), .Y(n955) );
  INVX2TS U1495 ( .A(n949), .Y(n1373) );
  INVX2TS U1496 ( .A(n950), .Y(n1759) );
  AOI22X1TS U1497 ( .A0(n951), .A1(n1373), .B0(n997), .B1(n1759), .Y(n954) );
  INVX2TS U1498 ( .A(n965), .Y(n1775) );
  AOI22X1TS U1499 ( .A0(n999), .A1(n1775), .B0(n952), .B1(n139), .Y(n953) );
  INVX2TS U1500 ( .A(n956), .Y(n1824) );
  INVX2TS U1501 ( .A(n972), .Y(n1766) );
  INVX2TS U1502 ( .A(n1366), .Y(n1386) );
  AOI22X1TS U1503 ( .A0(n1824), .A1(n1766), .B0(n1386), .B1(
        \requesterAddressbuffer[3][1] ), .Y(n962) );
  AOI22X1TS U1504 ( .A0(n957), .A1(n141), .B0(n1004), .B1(n146), .Y(n961) );
  INVX2TS U1505 ( .A(n965), .Y(n1785) );
  AOI22X1TS U1506 ( .A0(n1006), .A1(n1785), .B0(n959), .B1(n958), .Y(n960) );
  INVX2TS U1507 ( .A(n963), .Y(n1835) );
  AOI22X1TS U1508 ( .A0(n1835), .A1(n1757), .B0(n1386), .B1(
        \requesterAddressbuffer[3][2] ), .Y(n970) );
  AOI22X1TS U1509 ( .A0(n964), .A1(n1387), .B0(n1010), .B1(n1381), .Y(n969) );
  AOI22X1TS U1510 ( .A0(n1013), .A1(n135), .B0(n967), .B1(n966), .Y(n968) );
  INVX2TS U1511 ( .A(n971), .Y(n1846) );
  INVX2TS U1512 ( .A(n972), .Y(n1781) );
  INVX2TS U1513 ( .A(n1366), .Y(n1772) );
  AOI22X1TS U1514 ( .A0(n1846), .A1(n1781), .B0(n1772), .B1(
        \requesterAddressbuffer[3][3] ), .Y(n977) );
  AOI22X1TS U1515 ( .A0(n973), .A1(n1373), .B0(n1019), .B1(n1782), .Y(n976) );
  AOI22X1TS U1516 ( .A0(n1022), .A1(n1775), .B0(n974), .B1(n1762), .Y(n975) );
  AOI22X1TS U1517 ( .A0(n1758), .A1(n1789), .B0(n1808), .B1(
        \requesterAddressbuffer[2][0] ), .Y(n980) );
  INVX2TS U1518 ( .A(n1344), .Y(n1796) );
  AOI22X1TS U1519 ( .A0(requesterAddressIn_WEST[0]), .A1(n1809), .B0(n997), 
        .B1(n1796), .Y(n979) );
  AOI22X1TS U1520 ( .A0(n999), .A1(n199), .B0(n998), .B1(n1111), .Y(n978) );
  INVX2TS U1521 ( .A(n989), .Y(n1795) );
  INVX2TS U1522 ( .A(n981), .Y(n1360) );
  AOI22X1TS U1523 ( .A0(n1866), .A1(n1795), .B0(n1360), .B1(
        \requesterAddressbuffer[2][1] ), .Y(n984) );
  INVX2TS U1524 ( .A(n1344), .Y(n1803) );
  AOI22X1TS U1525 ( .A0(requesterAddressIn_WEST[1]), .A1(n1356), .B0(n1004), 
        .B1(n1803), .Y(n983) );
  AOI22X1TS U1526 ( .A0(n1006), .A1(n1351), .B0(n1005), .B1(n1797), .Y(n982)
         );
  INVX2TS U1527 ( .A(n989), .Y(n1802) );
  AOI22X1TS U1528 ( .A0(n1876), .A1(n1802), .B0(n1360), .B1(
        \requesterAddressbuffer[2][2] ), .Y(n988) );
  AOI22X1TS U1529 ( .A0(requesterAddressIn_WEST[2]), .A1(n1109), .B0(n1010), 
        .B1(n991), .Y(n987) );
  AOI22X1TS U1530 ( .A0(n1013), .A1(n1110), .B0(n1012), .B1(n985), .Y(n986) );
  INVX2TS U1531 ( .A(n1604), .Y(n1801) );
  AOI22X1TS U1532 ( .A0(n1886), .A1(n1789), .B0(n1801), .B1(
        \requesterAddressbuffer[2][3] ), .Y(n995) );
  INVX2TS U1533 ( .A(n990), .Y(n1356) );
  AOI22X1TS U1534 ( .A0(requesterAddressIn_WEST[3]), .A1(n1356), .B0(n1019), 
        .B1(n991), .Y(n994) );
  INVX2TS U1535 ( .A(n992), .Y(n1804) );
  AOI22X1TS U1536 ( .A0(n1022), .A1(n1804), .B0(n1021), .B1(n1791), .Y(n993)
         );
  INVX2TS U1537 ( .A(n1084), .Y(n1098) );
  AOI22X1TS U1538 ( .A0(n996), .A1(n1098), .B0(n1844), .B1(
        \requesterAddressbuffer[1][0] ), .Y(n1002) );
  INVX2TS U1539 ( .A(n1089), .Y(n1826) );
  AOI22X1TS U1540 ( .A0(requesterAddressIn_WEST[0]), .A1(n1848), .B0(n997), 
        .B1(n1826), .Y(n1001) );
  AOI22X1TS U1541 ( .A0(n999), .A1(n1079), .B0(n998), .B1(n1080), .Y(n1000) );
  INVX2TS U1542 ( .A(n1084), .Y(n1834) );
  INVX2TS U1543 ( .A(n1003), .Y(n1103) );
  AOI22X1TS U1544 ( .A0(n1736), .A1(n1834), .B0(n1103), .B1(
        \requesterAddressbuffer[1][1] ), .Y(n1009) );
  INVX2TS U1545 ( .A(n1089), .Y(n1837) );
  AOI22X1TS U1546 ( .A0(requesterAddressIn_WEST[1]), .A1(n1099), .B0(n1004), 
        .B1(n1837), .Y(n1008) );
  AOI22X1TS U1547 ( .A0(n1006), .A1(n332), .B0(n1005), .B1(n1829), .Y(n1007)
         );
  AOI22X1TS U1548 ( .A0(n1742), .A1(n1845), .B0(n1103), .B1(
        \requesterAddressbuffer[1][2] ), .Y(n1016) );
  AOI22X1TS U1549 ( .A0(requesterAddressIn_WEST[2]), .A1(n1078), .B0(n1010), 
        .B1(n1018), .Y(n1015) );
  AOI22X1TS U1550 ( .A0(n1013), .A1(n1094), .B0(n1012), .B1(n1011), .Y(n1014)
         );
  INVX2TS U1551 ( .A(n1619), .Y(n1833) );
  AOI22X1TS U1552 ( .A0(n1750), .A1(n1098), .B0(n1833), .B1(
        \requesterAddressbuffer[1][3] ), .Y(n1025) );
  INVX2TS U1553 ( .A(n1017), .Y(n1099) );
  AOI22X1TS U1554 ( .A0(requesterAddressIn_WEST[3]), .A1(n1099), .B0(n1019), 
        .B1(n1018), .Y(n1024) );
  INVX2TS U1555 ( .A(n1020), .Y(n1839) );
  AOI22X1TS U1556 ( .A0(n1022), .A1(n1839), .B0(n1021), .B1(n1819), .Y(n1023)
         );
  AOI22X1TS U1557 ( .A0(readRequesterAddress[0]), .A1(n1855), .B0(n1884), .B1(
        \requesterAddressbuffer[0][0] ), .Y(n1030) );
  INVX2TS U1558 ( .A(n1061), .Y(n1867) );
  AOI22X1TS U1559 ( .A0(requesterAddressIn_WEST[0]), .A1(n1887), .B0(n1026), 
        .B1(n1867), .Y(n1029) );
  AOI22X1TS U1560 ( .A0(n1027), .A1(n1880), .B0(requesterAddressIn_NORTH[0]), 
        .B1(n1869), .Y(n1028) );
  INVX2TS U1561 ( .A(n11), .Y(n1865) );
  INVX2TS U1562 ( .A(n1031), .Y(n1074) );
  AOI22X1TS U1563 ( .A0(n1824), .A1(n1865), .B0(n1074), .B1(
        \requesterAddressbuffer[0][1] ), .Y(n1037) );
  INVX2TS U1564 ( .A(n1061), .Y(n1877) );
  AOI22X1TS U1565 ( .A0(requesterAddressIn_WEST[1]), .A1(n1069), .B0(n1032), 
        .B1(n1877), .Y(n1036) );
  AOI22X1TS U1566 ( .A0(n1034), .A1(n1070), .B0(requesterAddressIn_NORTH[1]), 
        .B1(n1033), .Y(n1035) );
  INVX2TS U1567 ( .A(n11), .Y(n1875) );
  AOI22X1TS U1568 ( .A0(n1835), .A1(n1875), .B0(n1074), .B1(
        \requesterAddressbuffer[0][2] ), .Y(n1042) );
  AOI22X1TS U1569 ( .A0(requesterAddressIn_WEST[2]), .A1(n1052), .B0(n1038), 
        .B1(n1045), .Y(n1041) );
  AOI22X1TS U1570 ( .A0(n1039), .A1(n1891), .B0(requesterAddressIn_NORTH[2]), 
        .B1(n1889), .Y(n1040) );
  INVX2TS U1571 ( .A(n11), .Y(n1885) );
  INVX2TS U1572 ( .A(n1043), .Y(n1874) );
  AOI22X1TS U1573 ( .A0(n1846), .A1(n1885), .B0(n1874), .B1(
        \requesterAddressbuffer[0][3] ), .Y(n1051) );
  INVX2TS U1574 ( .A(n1044), .Y(n1069) );
  AOI22X1TS U1575 ( .A0(requesterAddressIn_WEST[3]), .A1(n1069), .B0(n1046), 
        .B1(n1045), .Y(n1050) );
  INVX2TS U1576 ( .A(n1047), .Y(n1861) );
  AOI22X1TS U1577 ( .A0(n1048), .A1(n1861), .B0(requesterAddressIn_NORTH[3]), 
        .B1(n1053), .Y(n1049) );
  INVX2TS U1578 ( .A(n1043), .Y(n1065) );
  AOI21X1TS U1579 ( .A0(n1065), .A1(\dataoutbuffer[0][0] ), .B0(n1865), .Y(
        n1056) );
  AOI22X1TS U1580 ( .A0(n1052), .A1(n1392), .B0(n1867), .B1(n1108), .Y(n1055)
         );
  AOI22X1TS U1581 ( .A0(n415), .A1(n1501), .B0(n1053), .B1(dataIn_NORTH[0]), 
        .Y(n1054) );
  AOI21X1TS U1582 ( .A0(n1065), .A1(\dataoutbuffer[0][1] ), .B0(n1875), .Y(
        n1060) );
  AOI22X1TS U1583 ( .A0(n402), .A1(n1398), .B0(n1877), .B1(n1339), .Y(n1059)
         );
  INVX2TS U1584 ( .A(n1057), .Y(n1869) );
  AOI22X1TS U1585 ( .A0(n1880), .A1(n1509), .B0(n1869), .B1(dataIn_NORTH[1]), 
        .Y(n1058) );
  AOI21X1TS U1586 ( .A0(n1065), .A1(\dataoutbuffer[0][2] ), .B0(n1885), .Y(
        n1064) );
  AOI22X1TS U1587 ( .A0(n1069), .A1(n1403), .B0(n393), .B1(n1345), .Y(n1063)
         );
  AOI22X1TS U1588 ( .A0(n1891), .A1(n1515), .B0(n1033), .B1(dataIn_NORTH[2]), 
        .Y(n1062) );
  AOI21X1TS U1589 ( .A0(n1065), .A1(\dataoutbuffer[0][3] ), .B0(n1865), .Y(
        n1068) );
  AOI22X1TS U1590 ( .A0(n1857), .A1(n1408), .B0(n1867), .B1(n1350), .Y(n1067)
         );
  AOI22X1TS U1591 ( .A0(n415), .A1(n1522), .B0(n1859), .B1(dataIn_NORTH[3]), 
        .Y(n1066) );
  AOI21X1TS U1592 ( .A0(n1074), .A1(\dataoutbuffer[0][4] ), .B0(n1875), .Y(
        n1073) );
  AOI22X1TS U1593 ( .A0(n1069), .A1(n1412), .B0(n1877), .B1(n1355), .Y(n1072)
         );
  AOI22X1TS U1594 ( .A0(n1070), .A1(n1531), .B0(n424), .B1(dataIn_NORTH[4]), 
        .Y(n1071) );
  AOI21X1TS U1595 ( .A0(n1074), .A1(\dataoutbuffer[0][5] ), .B0(n1885), .Y(
        n1077) );
  AOI22X1TS U1596 ( .A0(n402), .A1(n1420), .B0(n393), .B1(n1361), .Y(n1076) );
  AOI22X1TS U1597 ( .A0(n1861), .A1(n1538), .B0(n1869), .B1(dataIn_NORTH[5]), 
        .Y(n1075) );
  INVX2TS U1598 ( .A(n1619), .Y(n1093) );
  AOI21X1TS U1599 ( .A0(n1093), .A1(\dataoutbuffer[1][0] ), .B0(n1098), .Y(
        n1083) );
  AOI22X1TS U1600 ( .A0(n1078), .A1(dataIn_WEST[0]), .B0(n1826), .B1(n1108), 
        .Y(n1082) );
  CLKBUFX2TS U1601 ( .A(dataIn_NORTH[0]), .Y(n1427) );
  CLKBUFX2TS U1602 ( .A(n1427), .Y(n1500) );
  CLKBUFX2TS U1603 ( .A(n1501), .Y(n1462) );
  AOI22X1TS U1604 ( .A0(n1080), .A1(n1500), .B0(n1079), .B1(n1462), .Y(n1081)
         );
  INVX2TS U1605 ( .A(n1084), .Y(n1823) );
  AOI21X1TS U1606 ( .A0(n1093), .A1(\dataoutbuffer[1][1] ), .B0(n1823), .Y(
        n1088) );
  AOI22X1TS U1607 ( .A0(n330), .A1(dataIn_WEST[1]), .B0(n1837), .B1(n1339), 
        .Y(n1087) );
  INVX2TS U1608 ( .A(n1085), .Y(n1829) );
  CLKBUFX2TS U1609 ( .A(dataIn_NORTH[1]), .Y(n1432) );
  CLKBUFX2TS U1610 ( .A(n1432), .Y(n1508) );
  CLKBUFX2TS U1611 ( .A(n1509), .Y(n1469) );
  AOI22X1TS U1612 ( .A0(n1829), .A1(n1508), .B0(n1104), .B1(n1469), .Y(n1086)
         );
  AOI21X1TS U1613 ( .A0(n1093), .A1(\dataoutbuffer[1][2] ), .B0(n1834), .Y(
        n1092) );
  AOI22X1TS U1614 ( .A0(n1099), .A1(dataIn_WEST[2]), .B0(n318), .B1(n1345), 
        .Y(n1091) );
  CLKBUFX2TS U1615 ( .A(dataIn_NORTH[2]), .Y(n1437) );
  CLKBUFX2TS U1616 ( .A(n1437), .Y(n1514) );
  CLKBUFX2TS U1617 ( .A(n1515), .Y(n1475) );
  AOI22X1TS U1618 ( .A0(n1011), .A1(n1514), .B0(n1839), .B1(n1475), .Y(n1090)
         );
  AOI21X1TS U1619 ( .A0(n1093), .A1(\dataoutbuffer[1][3] ), .B0(n1845), .Y(
        n1097) );
  AOI22X1TS U1620 ( .A0(n1816), .A1(dataIn_WEST[3]), .B0(n1826), .B1(n1350), 
        .Y(n1096) );
  CLKBUFX2TS U1621 ( .A(dataIn_NORTH[3]), .Y(n1443) );
  CLKBUFX2TS U1622 ( .A(n1443), .Y(n1521) );
  CLKBUFX2TS U1623 ( .A(n1522), .Y(n1481) );
  AOI22X1TS U1624 ( .A0(n1819), .A1(n1521), .B0(n1094), .B1(n1481), .Y(n1095)
         );
  AOI21X1TS U1625 ( .A0(n1103), .A1(\dataoutbuffer[1][4] ), .B0(n1098), .Y(
        n1102) );
  AOI22X1TS U1626 ( .A0(n1099), .A1(dataIn_WEST[4]), .B0(n1837), .B1(n1355), 
        .Y(n1101) );
  CLKBUFX2TS U1627 ( .A(dataIn_NORTH[4]), .Y(n1449) );
  CLKBUFX2TS U1628 ( .A(n1449), .Y(n1529) );
  CLKBUFX2TS U1629 ( .A(n1531), .Y(n1487) );
  AOI22X1TS U1630 ( .A0(n323), .A1(n1529), .B0(n365), .B1(n1487), .Y(n1100) );
  AOI21X1TS U1631 ( .A0(n1103), .A1(\dataoutbuffer[1][5] ), .B0(n1823), .Y(
        n1107) );
  AOI22X1TS U1632 ( .A0(n330), .A1(dataIn_WEST[5]), .B0(n318), .B1(n1361), .Y(
        n1106) );
  CLKBUFX2TS U1633 ( .A(dataIn_NORTH[5]), .Y(n1455) );
  CLKBUFX2TS U1634 ( .A(n1455), .Y(n1537) );
  CLKBUFX2TS U1635 ( .A(n1538), .Y(n1494) );
  AOI22X1TS U1636 ( .A0(n1829), .A1(n1537), .B0(n1104), .B1(n1494), .Y(n1105)
         );
  INVX2TS U1637 ( .A(n1604), .Y(n1349) );
  AOI21X1TS U1638 ( .A0(n1349), .A1(\dataoutbuffer[2][0] ), .B0(n1795), .Y(
        n1338) );
  AOI22X1TS U1639 ( .A0(n1109), .A1(dataIn_WEST[0]), .B0(n1796), .B1(n1108), 
        .Y(n1337) );
  AOI22X1TS U1640 ( .A0(n1111), .A1(n1500), .B0(n1110), .B1(dataIn_SOUTH[0]), 
        .Y(n1112) );
  AOI21X1TS U1641 ( .A0(n1349), .A1(\dataoutbuffer[2][1] ), .B0(n1802), .Y(
        n1343) );
  AOI22X1TS U1642 ( .A0(n198), .A1(dataIn_WEST[1]), .B0(n1803), .B1(n1339), 
        .Y(n1342) );
  INVX2TS U1643 ( .A(n1340), .Y(n1797) );
  AOI22X1TS U1644 ( .A0(n1797), .A1(n1508), .B0(n1362), .B1(dataIn_SOUTH[1]), 
        .Y(n1341) );
  AOI21X1TS U1645 ( .A0(n1349), .A1(\dataoutbuffer[2][2] ), .B0(n185), .Y(
        n1348) );
  AOI22X1TS U1646 ( .A0(n1356), .A1(dataIn_WEST[2]), .B0(n184), .B1(n1345), 
        .Y(n1347) );
  AOI22X1TS U1647 ( .A0(n985), .A1(n1514), .B0(n1804), .B1(dataIn_SOUTH[2]), 
        .Y(n1346) );
  AOI21X1TS U1648 ( .A0(n1349), .A1(\dataoutbuffer[2][3] ), .B0(n1795), .Y(
        n1354) );
  AOI22X1TS U1649 ( .A0(n1790), .A1(dataIn_WEST[3]), .B0(n1796), .B1(n1350), 
        .Y(n1353) );
  AOI22X1TS U1650 ( .A0(n1791), .A1(n1521), .B0(n1351), .B1(dataIn_SOUTH[3]), 
        .Y(n1352) );
  AOI21X1TS U1651 ( .A0(n1360), .A1(\dataoutbuffer[2][4] ), .B0(n1802), .Y(
        n1359) );
  AOI22X1TS U1652 ( .A0(n1356), .A1(dataIn_WEST[4]), .B0(n1803), .B1(n1355), 
        .Y(n1358) );
  AOI22X1TS U1653 ( .A0(n194), .A1(n1529), .B0(n212), .B1(dataIn_SOUTH[4]), 
        .Y(n1357) );
  AOI21X1TS U1654 ( .A0(n1360), .A1(\dataoutbuffer[2][5] ), .B0(n185), .Y(
        n1365) );
  AOI22X1TS U1655 ( .A0(n198), .A1(dataIn_WEST[5]), .B0(n184), .B1(n1361), .Y(
        n1364) );
  AOI22X1TS U1656 ( .A0(n1797), .A1(n1537), .B0(n1362), .B1(dataIn_SOUTH[5]), 
        .Y(n1363) );
  INVX2TS U1657 ( .A(n178), .Y(n1377) );
  AOI21X1TS U1658 ( .A0(n1377), .A1(\dataoutbuffer[3][0] ), .B0(n1766), .Y(
        n1369) );
  AOI22X1TS U1659 ( .A0(n1373), .A1(dataIn_WEST[0]), .B0(n1773), .B1(
        dataIn_EAST[0]), .Y(n1368) );
  AOI22X1TS U1660 ( .A0(n966), .A1(n1427), .B0(n1768), .B1(n1462), .Y(n1367)
         );
  AOI21X1TS U1661 ( .A0(n1377), .A1(\dataoutbuffer[3][1] ), .B0(n136), .Y(
        n1372) );
  AOI22X1TS U1662 ( .A0(n157), .A1(dataIn_WEST[1]), .B0(n146), .B1(
        dataIn_EAST[1]), .Y(n1371) );
  INVX2TS U1663 ( .A(n151), .Y(n1776) );
  AOI22X1TS U1664 ( .A0(n1776), .A1(n1432), .B0(n1775), .B1(n1469), .Y(n1370)
         );
  AOI21X1TS U1665 ( .A0(n1377), .A1(\dataoutbuffer[3][2] ), .B0(n1781), .Y(
        n1376) );
  AOI22X1TS U1666 ( .A0(n1373), .A1(dataIn_WEST[2]), .B0(n1759), .B1(
        dataIn_EAST[2]), .Y(n1375) );
  AOI22X1TS U1667 ( .A0(n1382), .A1(n1437), .B0(n1785), .B1(n1475), .Y(n1374)
         );
  AOI21X1TS U1668 ( .A0(n1377), .A1(\dataoutbuffer[3][3] ), .B0(n1766), .Y(
        n1380) );
  AOI22X1TS U1669 ( .A0(n1761), .A1(dataIn_WEST[3]), .B0(n1759), .B1(
        dataIn_EAST[3]), .Y(n1379) );
  AOI22X1TS U1670 ( .A0(n1762), .A1(n1443), .B0(n135), .B1(n1481), .Y(n1378)
         );
  AOI21X1TS U1671 ( .A0(n1386), .A1(\dataoutbuffer[3][4] ), .B0(n136), .Y(
        n1385) );
  AOI22X1TS U1672 ( .A0(n157), .A1(dataIn_WEST[4]), .B0(n1381), .B1(
        dataIn_EAST[4]), .Y(n1384) );
  AOI22X1TS U1673 ( .A0(n1382), .A1(n1449), .B0(n1785), .B1(n1487), .Y(n1383)
         );
  AOI21X1TS U1674 ( .A0(n1386), .A1(\dataoutbuffer[3][5] ), .B0(n1781), .Y(
        n1390) );
  AOI22X1TS U1675 ( .A0(n1387), .A1(dataIn_WEST[5]), .B0(n145), .B1(
        dataIn_EAST[5]), .Y(n1389) );
  AOI22X1TS U1676 ( .A0(n1776), .A1(n1455), .B0(n135), .B1(n1494), .Y(n1388)
         );
  INVX2TS U1677 ( .A(n938), .Y(n1407) );
  AOI21X1TS U1678 ( .A0(n1407), .A1(\dataoutbuffer[4][0] ), .B0(n1735), .Y(
        n1397) );
  AOI22X1TS U1679 ( .A0(n1393), .A1(n1392), .B0(n1737), .B1(dataIn_EAST[0]), 
        .Y(n1396) );
  AOI22X1TS U1680 ( .A0(n1731), .A1(dataIn_SOUTH[0]), .B0(n1394), .B1(n1500), 
        .Y(n1395) );
  AOI21X1TS U1681 ( .A0(n1407), .A1(\dataoutbuffer[4][1] ), .B0(n277), .Y(
        n1401) );
  AOI22X1TS U1682 ( .A0(n279), .A1(n1398), .B0(n1743), .B1(dataIn_EAST[1]), 
        .Y(n1400) );
  AOI22X1TS U1683 ( .A0(n1744), .A1(dataIn_SOUTH[1]), .B0(n1414), .B1(n1508), 
        .Y(n1399) );
  AOI21X1TS U1684 ( .A0(n1407), .A1(\dataoutbuffer[4][2] ), .B0(n1749), .Y(
        n1406) );
  AOI22X1TS U1685 ( .A0(n1413), .A1(n1403), .B0(n276), .B1(dataIn_EAST[2]), 
        .Y(n1405) );
  AOI22X1TS U1686 ( .A0(n1753), .A1(dataIn_SOUTH[2]), .B0(n1414), .B1(n1514), 
        .Y(n1404) );
  AOI21X1TS U1687 ( .A0(n1407), .A1(\dataoutbuffer[4][3] ), .B0(n1735), .Y(
        n1411) );
  AOI22X1TS U1688 ( .A0(n1729), .A1(n1408), .B0(n1737), .B1(dataIn_EAST[3]), 
        .Y(n1410) );
  AOI22X1TS U1689 ( .A0(n302), .A1(dataIn_SOUTH[3]), .B0(n1730), .B1(n1521), 
        .Y(n1409) );
  AOI21X1TS U1690 ( .A0(n1419), .A1(\dataoutbuffer[4][4] ), .B0(n277), .Y(
        n1418) );
  AOI22X1TS U1691 ( .A0(n1413), .A1(n1412), .B0(n1743), .B1(dataIn_EAST[4]), 
        .Y(n1417) );
  AOI22X1TS U1692 ( .A0(n1415), .A1(dataIn_SOUTH[4]), .B0(n1414), .B1(n1529), 
        .Y(n1416) );
  AOI21X1TS U1693 ( .A0(n1419), .A1(\dataoutbuffer[4][5] ), .B0(n1749), .Y(
        n1423) );
  AOI22X1TS U1694 ( .A0(n279), .A1(n1420), .B0(n276), .B1(dataIn_EAST[5]), .Y(
        n1422) );
  AOI22X1TS U1695 ( .A0(n1731), .A1(dataIn_SOUTH[5]), .B0(n286), .B1(n1537), 
        .Y(n1421) );
  INVX2TS U1696 ( .A(n912), .Y(n1442) );
  AOI21X1TS U1697 ( .A0(n1442), .A1(\dataoutbuffer[5][0] ), .B0(n1703), .Y(
        n1431) );
  AOI22X1TS U1698 ( .A0(n1425), .A1(n1499), .B0(n1705), .B1(n1460), .Y(n1430)
         );
  AOI22X1TS U1699 ( .A0(n1428), .A1(n1427), .B0(n1426), .B1(n1462), .Y(n1429)
         );
  AOI21X1TS U1700 ( .A0(n1442), .A1(\dataoutbuffer[5][1] ), .B0(n1712), .Y(
        n1435) );
  AOI22X1TS U1701 ( .A0(n236), .A1(n1506), .B0(n1714), .B1(n1468), .Y(n1434)
         );
  AOI22X1TS U1702 ( .A0(n1707), .A1(n1432), .B0(n1724), .B1(n1469), .Y(n1433)
         );
  AOI21X1TS U1703 ( .A0(n1442), .A1(\dataoutbuffer[5][2] ), .B0(n1720), .Y(
        n1441) );
  AOI22X1TS U1704 ( .A0(n1447), .A1(n1513), .B0(n225), .B1(n1474), .Y(n1440)
         );
  AOI22X1TS U1705 ( .A0(n1438), .A1(n1437), .B0(n1448), .B1(n1475), .Y(n1439)
         );
  AOI21X1TS U1706 ( .A0(n1442), .A1(\dataoutbuffer[5][3] ), .B0(n1703), .Y(
        n1446) );
  AOI22X1TS U1707 ( .A0(n1697), .A1(n1520), .B0(n1705), .B1(n1480), .Y(n1445)
         );
  AOI22X1TS U1708 ( .A0(n230), .A1(n1443), .B0(n1698), .B1(n1481), .Y(n1444)
         );
  AOI21X1TS U1709 ( .A0(n1454), .A1(\dataoutbuffer[5][4] ), .B0(n1712), .Y(
        n1453) );
  AOI22X1TS U1710 ( .A0(n1447), .A1(n1527), .B0(n1714), .B1(n1485), .Y(n1452)
         );
  AOI22X1TS U1711 ( .A0(n1450), .A1(n1449), .B0(n1448), .B1(n1487), .Y(n1451)
         );
  AOI21X1TS U1712 ( .A0(n1454), .A1(\dataoutbuffer[5][5] ), .B0(n1720), .Y(
        n1458) );
  AOI22X1TS U1713 ( .A0(n236), .A1(n1536), .B0(n225), .B1(n1493), .Y(n1457) );
  AOI22X1TS U1714 ( .A0(n1707), .A1(n1455), .B0(n237), .B1(n1494), .Y(n1456)
         );
  INVX2TS U1715 ( .A(n894), .Y(n1479) );
  AOI21X1TS U1716 ( .A0(n1479), .A1(\dataoutbuffer[6][0] ), .B0(n1671), .Y(
        n1467) );
  AOI22X1TS U1717 ( .A0(n1461), .A1(n1499), .B0(n1672), .B1(n1460), .Y(n1466)
         );
  AOI22X1TS U1718 ( .A0(n1464), .A1(dataIn_NORTH[0]), .B0(n1463), .B1(n1462), 
        .Y(n1465) );
  AOI21X1TS U1719 ( .A0(n1479), .A1(\dataoutbuffer[6][1] ), .B0(n88), .Y(n1472) );
  AOI22X1TS U1720 ( .A0(n90), .A1(n1506), .B0(n1679), .B1(n1468), .Y(n1471) );
  AOI22X1TS U1721 ( .A0(n1674), .A1(dataIn_NORTH[1]), .B0(n98), .B1(n1469), 
        .Y(n1470) );
  AOI21X1TS U1722 ( .A0(n1479), .A1(\dataoutbuffer[6][2] ), .B0(n1686), .Y(
        n1478) );
  AOI22X1TS U1723 ( .A0(n1486), .A1(n1513), .B0(n87), .B1(n1474), .Y(n1477) );
  AOI22X1TS U1724 ( .A0(n93), .A1(dataIn_NORTH[2]), .B0(n1488), .B1(n1475), 
        .Y(n1476) );
  AOI21X1TS U1725 ( .A0(n1479), .A1(\dataoutbuffer[6][3] ), .B0(n1671), .Y(
        n1484) );
  AOI22X1TS U1726 ( .A0(n1665), .A1(n1520), .B0(n1672), .B1(n1480), .Y(n1483)
         );
  AOI22X1TS U1727 ( .A0(n1667), .A1(dataIn_NORTH[3]), .B0(n98), .B1(n1481), 
        .Y(n1482) );
  AOI21X1TS U1728 ( .A0(n1492), .A1(\dataoutbuffer[6][4] ), .B0(n88), .Y(n1491) );
  AOI22X1TS U1729 ( .A0(n1486), .A1(n1527), .B0(n1679), .B1(n1485), .Y(n1490)
         );
  AOI22X1TS U1730 ( .A0(n102), .A1(dataIn_NORTH[4]), .B0(n1488), .B1(n1487), 
        .Y(n1489) );
  AOI21X1TS U1731 ( .A0(n1492), .A1(\dataoutbuffer[6][5] ), .B0(n1686), .Y(
        n1497) );
  AOI22X1TS U1732 ( .A0(n90), .A1(n1536), .B0(n87), .B1(n1493), .Y(n1496) );
  AOI22X1TS U1733 ( .A0(n1674), .A1(dataIn_NORTH[5]), .B0(n112), .B1(n1494), 
        .Y(n1495) );
  INVX2TS U1734 ( .A(n877), .Y(n1519) );
  AOI21X1TS U1735 ( .A0(n1519), .A1(\dataoutbuffer[7][0] ), .B0(n1641), .Y(
        n1504) );
  AOI22X1TS U1736 ( .A0(n51), .A1(n1499), .B0(n1658), .B1(dataIn_EAST[0]), .Y(
        n1503) );
  AOI22X1TS U1737 ( .A0(n1539), .A1(n1501), .B0(n72), .B1(n1500), .Y(n1502) );
  AOI21X1TS U1738 ( .A0(n1519), .A1(\dataoutbuffer[7][1] ), .B0(n34), .Y(n1512) );
  AOI22X1TS U1739 ( .A0(n67), .A1(n1506), .B0(n1636), .B1(dataIn_EAST[1]), .Y(
        n1511) );
  INVX2TS U1740 ( .A(n1507), .Y(n1651) );
  AOI22X1TS U1741 ( .A0(n63), .A1(n1509), .B0(n1651), .B1(n1508), .Y(n1510) );
  AOI21X1TS U1742 ( .A0(n1519), .A1(\dataoutbuffer[7][2] ), .B0(n1657), .Y(
        n1518) );
  AOI22X1TS U1743 ( .A0(n51), .A1(n1513), .B0(n32), .B1(dataIn_EAST[2]), .Y(
        n1517) );
  AOI22X1TS U1744 ( .A0(n1523), .A1(n1515), .B0(n1642), .B1(n1514), .Y(n1516)
         );
  AOI21X1TS U1745 ( .A0(n1519), .A1(\dataoutbuffer[7][3] ), .B0(n1641), .Y(
        n1526) );
  AOI22X1TS U1746 ( .A0(n1659), .A1(n1520), .B0(n1658), .B1(dataIn_EAST[3]), 
        .Y(n1525) );
  AOI22X1TS U1747 ( .A0(n1523), .A1(n1522), .B0(n72), .B1(n1521), .Y(n1524) );
  AOI21X1TS U1748 ( .A0(n1535), .A1(\dataoutbuffer[7][4] ), .B0(n1635), .Y(
        n1534) );
  AOI22X1TS U1749 ( .A0(n1528), .A1(n1527), .B0(n1636), .B1(dataIn_EAST[4]), 
        .Y(n1533) );
  AOI22X1TS U1750 ( .A0(n1539), .A1(n1531), .B0(n1530), .B1(n1529), .Y(n1532)
         );
  AOI21X1TS U1751 ( .A0(n1535), .A1(\dataoutbuffer[7][5] ), .B0(n1657), .Y(
        n1542) );
  AOI22X1TS U1752 ( .A0(n76), .A1(n1536), .B0(n32), .B1(dataIn_EAST[5]), .Y(
        n1541) );
  AOI22X1TS U1753 ( .A0(n1539), .A1(n1538), .B0(n1651), .B1(n1537), .Y(n1540)
         );
  CLKBUFX2TS U1754 ( .A(n1631), .Y(n1583) );
  INVX2TS U1755 ( .A(n1543), .Y(n1612) );
  AOI22X1TS U1756 ( .A0(n1545), .A1(n1566), .B0(n1565), .B1(n1544), .Y(n1547)
         );
  AOI22X1TS U1757 ( .A0(n1548), .A1(n1612), .B0(n1547), .B1(n1546), .Y(n1550)
         );
  AOI22X1TS U1758 ( .A0(n1551), .A1(n1583), .B0(n1550), .B1(n1549), .Y(n1553)
         );
  AOI32X1TS U1759 ( .A0(n1553), .A1(n1498), .A2(n1552), .B0(n1655), .B1(n1925), 
        .Y(n2052) );
  INVX2TS U1760 ( .A(n1543), .Y(n1627) );
  AOI22X1TS U1761 ( .A0(n1555), .A1(n1566), .B0(n1565), .B1(n1554), .Y(n1557)
         );
  AOI22X1TS U1762 ( .A0(n1558), .A1(n1627), .B0(n1557), .B1(n1556), .Y(n1560)
         );
  AOI22X1TS U1763 ( .A0(n1561), .A1(n1583), .B0(n1560), .B1(n1559), .Y(n1563)
         );
  AOI32X1TS U1764 ( .A0(n1563), .A1(n1459), .A2(n1562), .B0(n1685), .B1(n1926), 
        .Y(n2053) );
  AOI22X1TS U1765 ( .A0(n1567), .A1(n1566), .B0(n1565), .B1(n1564), .Y(n1569)
         );
  AOI22X1TS U1766 ( .A0(n1570), .A1(n1612), .B0(n1569), .B1(n1568), .Y(n1572)
         );
  AOI22X1TS U1767 ( .A0(n1573), .A1(n1583), .B0(n1572), .B1(n1571), .Y(n1575)
         );
  AOI32X1TS U1768 ( .A0(n1575), .A1(n1424), .A2(n1574), .B0(n1719), .B1(n1927), 
        .Y(n2054) );
  CLKBUFX2TS U1769 ( .A(n1623), .Y(n1608) );
  CLKBUFX2TS U1770 ( .A(n1622), .Y(n1607) );
  AOI22X1TS U1771 ( .A0(n1577), .A1(n1608), .B0(n1607), .B1(n1576), .Y(n1579)
         );
  AOI22X1TS U1772 ( .A0(n1580), .A1(n1627), .B0(n1579), .B1(n1578), .Y(n1582)
         );
  AOI22X1TS U1773 ( .A0(n1584), .A1(n1583), .B0(n1582), .B1(n1581), .Y(n1586)
         );
  AOI32X1TS U1774 ( .A0(n1586), .A1(n1391), .A2(n1585), .B0(n1748), .B1(n1928), 
        .Y(n2055) );
  AOI22X1TS U1775 ( .A0(n125), .A1(n1608), .B0(n1607), .B1(n26), .Y(n1588) );
  AOI22X1TS U1776 ( .A0(n1589), .A1(n1612), .B0(n1588), .B1(n1587), .Y(n1591)
         );
  AOI22X1TS U1777 ( .A0(n1592), .A1(n1631), .B0(n1591), .B1(n1590), .Y(n1594)
         );
  AOI32X1TS U1778 ( .A0(n1594), .A1(n1366), .A2(n1593), .B0(n1780), .B1(n1929), 
        .Y(n2056) );
  AOI22X1TS U1779 ( .A0(n1596), .A1(n1608), .B0(n1607), .B1(n1595), .Y(n1598)
         );
  AOI22X1TS U1780 ( .A0(n1599), .A1(n1627), .B0(n1598), .B1(n1597), .Y(n1601)
         );
  AOI22X1TS U1781 ( .A0(n1602), .A1(n1616), .B0(n1601), .B1(n1600), .Y(n1605)
         );
  AOI32X1TS U1782 ( .A0(n1605), .A1(n1604), .A2(n1603), .B0(n1808), .B1(n1930), 
        .Y(n2057) );
  AOI22X1TS U1783 ( .A0(n1609), .A1(n1608), .B0(n1607), .B1(n1606), .Y(n1611)
         );
  AOI22X1TS U1784 ( .A0(n1613), .A1(n1612), .B0(n1611), .B1(n1610), .Y(n1615)
         );
  AOI22X1TS U1785 ( .A0(n1617), .A1(n1616), .B0(n1615), .B1(n1614), .Y(n1620)
         );
  AOI32X1TS U1786 ( .A0(n1620), .A1(n1619), .A2(n1618), .B0(n1844), .B1(n1931), 
        .Y(n2058) );
  AOI22X1TS U1787 ( .A0(n1624), .A1(n1623), .B0(n1622), .B1(n1621), .Y(n1626)
         );
  AOI22X1TS U1788 ( .A0(n1628), .A1(n1627), .B0(n1626), .B1(n1625), .Y(n1630)
         );
  AOI22X1TS U1789 ( .A0(n1632), .A1(n1631), .B0(n1630), .B1(n1629), .Y(n1634)
         );
  AOI32X1TS U1790 ( .A0(n1634), .A1(n1043), .A2(n1633), .B0(n1884), .B1(n1932), 
        .Y(n2059) );
  AOI22X1TS U1791 ( .A0(n1814), .A1(n1635), .B0(n1647), .B1(
        \destinationAddressbuffer[7][0] ), .Y(n1639) );
  AOI22X1TS U1792 ( .A0(n67), .A1(n1696), .B0(n1636), .B1(n1695), .Y(n1638) );
  CLKBUFX2TS U1793 ( .A(n1666), .Y(n1818) );
  AOI22X1TS U1794 ( .A0(n1643), .A1(destinationAddressIn_SOUTH[0]), .B0(n1651), 
        .B1(n1818), .Y(n1637) );
  AOI22X1TS U1795 ( .A0(n1641), .A1(n1640), .B0(n1647), .B1(
        \destinationAddressbuffer[7][1] ), .Y(n1646) );
  AOI22X1TS U1796 ( .A0(n76), .A1(n1706), .B0(n1649), .B1(n1704), .Y(n1645) );
  CLKBUFX2TS U1797 ( .A(n1673), .Y(n1828) );
  AOI22X1TS U1798 ( .A0(n1643), .A1(destinationAddressIn_SOUTH[1]), .B0(n1642), 
        .B1(n1828), .Y(n1644) );
  AOI22X1TS U1799 ( .A0(n34), .A1(n1648), .B0(n1647), .B1(
        \destinationAddressbuffer[7][2] ), .Y(n1654) );
  AOI22X1TS U1800 ( .A0(n1650), .A1(n1715), .B0(n1649), .B1(n1713), .Y(n1653)
         );
  CLKBUFX2TS U1801 ( .A(n1680), .Y(n1840) );
  AOI22X1TS U1802 ( .A0(n58), .A1(destinationAddressIn_SOUTH[2]), .B0(n1651), 
        .B1(n1840), .Y(n1652) );
  AOI22X1TS U1803 ( .A0(n1657), .A1(n1656), .B0(n1655), .B1(
        \destinationAddressbuffer[7][3] ), .Y(n1663) );
  AOI22X1TS U1804 ( .A0(n1659), .A1(n1722), .B0(n1658), .B1(n1721), .Y(n1662)
         );
  CLKBUFX2TS U1805 ( .A(n1688), .Y(n1850) );
  AOI22X1TS U1806 ( .A0(n1660), .A1(destinationAddressIn_SOUTH[3]), .B0(n53), 
        .B1(n1850), .Y(n1661) );
  AOI22X1TS U1807 ( .A0(n1856), .A1(n1664), .B0(n1678), .B1(
        \destinationAddressbuffer[6][0] ), .Y(n1670) );
  AOI22X1TS U1808 ( .A0(n1665), .A1(n1696), .B0(n896), .B1(n1695), .Y(n1669)
         );
  CLKBUFX2TS U1809 ( .A(n1666), .Y(n1858) );
  CLKBUFX2TS U1810 ( .A(destinationAddressIn_SOUTH[0]), .Y(n1860) );
  CLKBUFX2TS U1811 ( .A(n1860), .Y(n1817) );
  AOI22X1TS U1812 ( .A0(n1667), .A1(n1858), .B0(n1689), .B1(n1817), .Y(n1668)
         );
  AOI22X1TS U1813 ( .A0(n1736), .A1(n1671), .B0(n1678), .B1(
        \destinationAddressbuffer[6][1] ), .Y(n1677) );
  AOI22X1TS U1814 ( .A0(n115), .A1(n1706), .B0(n1672), .B1(n1704), .Y(n1676)
         );
  CLKBUFX2TS U1815 ( .A(n1673), .Y(n1868) );
  CLKBUFX2TS U1816 ( .A(destinationAddressIn_SOUTH[1]), .Y(n1870) );
  CLKBUFX2TS U1817 ( .A(n1870), .Y(n1827) );
  AOI22X1TS U1818 ( .A0(n1674), .A1(n1868), .B0(n1681), .B1(n1827), .Y(n1675)
         );
  AOI22X1TS U1819 ( .A0(n1742), .A1(n88), .B0(n1678), .B1(
        \destinationAddressbuffer[6][2] ), .Y(n1684) );
  AOI22X1TS U1820 ( .A0(n1687), .A1(n1715), .B0(n1679), .B1(n1713), .Y(n1683)
         );
  CLKBUFX2TS U1821 ( .A(n1680), .Y(n1878) );
  CLKBUFX2TS U1822 ( .A(destinationAddressIn_SOUTH[2]), .Y(n1879) );
  CLKBUFX2TS U1823 ( .A(n1879), .Y(n1838) );
  AOI22X1TS U1824 ( .A0(n1690), .A1(n1878), .B0(n1681), .B1(n1838), .Y(n1682)
         );
  AOI22X1TS U1825 ( .A0(n1750), .A1(n1686), .B0(n1685), .B1(
        \destinationAddressbuffer[6][3] ), .Y(n1693) );
  AOI22X1TS U1826 ( .A0(n1687), .A1(n1722), .B0(n87), .B1(n1721), .Y(n1692) );
  CLKBUFX2TS U1827 ( .A(n1688), .Y(n1888) );
  CLKBUFX2TS U1828 ( .A(destinationAddressIn_SOUTH[3]), .Y(n1890) );
  CLKBUFX2TS U1829 ( .A(n1890), .Y(n1849) );
  AOI22X1TS U1830 ( .A0(n1690), .A1(n1888), .B0(n1689), .B1(n1849), .Y(n1691)
         );
  AOI22X1TS U1831 ( .A0(n1856), .A1(n1694), .B0(n1711), .B1(
        \destinationAddressbuffer[5][0] ), .Y(n1702) );
  AOI22X1TS U1832 ( .A0(n1697), .A1(n1696), .B0(n914), .B1(n1695), .Y(n1701)
         );
  AOI22X1TS U1833 ( .A0(n1699), .A1(n1858), .B0(n1698), .B1(
        destinationAddressIn_SOUTH[0]), .Y(n1700) );
  AOI22X1TS U1834 ( .A0(readRequesterAddress[1]), .A1(n1703), .B0(n1711), .B1(
        \destinationAddressbuffer[5][1] ), .Y(n1710) );
  AOI22X1TS U1835 ( .A0(n261), .A1(n1706), .B0(n1705), .B1(n1704), .Y(n1709)
         );
  AOI22X1TS U1836 ( .A0(n1707), .A1(n1868), .B0(n232), .B1(
        destinationAddressIn_SOUTH[1]), .Y(n1708) );
  AOI22X1TS U1837 ( .A0(readRequesterAddress[2]), .A1(n1712), .B0(n1711), .B1(
        \destinationAddressbuffer[5][2] ), .Y(n1718) );
  AOI22X1TS U1838 ( .A0(n1723), .A1(n1715), .B0(n1714), .B1(n1713), .Y(n1717)
         );
  AOI22X1TS U1839 ( .A0(n1428), .A1(n1878), .B0(n1724), .B1(
        destinationAddressIn_SOUTH[2]), .Y(n1716) );
  AOI22X1TS U1840 ( .A0(readRequesterAddress[3]), .A1(n1720), .B0(n1719), .B1(
        \destinationAddressbuffer[5][3] ), .Y(n1727) );
  AOI22X1TS U1841 ( .A0(n1723), .A1(n1722), .B0(n225), .B1(n1721), .Y(n1726)
         );
  AOI22X1TS U1842 ( .A0(n230), .A1(n1888), .B0(n1724), .B1(
        destinationAddressIn_SOUTH[3]), .Y(n1725) );
  AOI22X1TS U1843 ( .A0(n1758), .A1(n1728), .B0(n1741), .B1(
        \destinationAddressbuffer[4][0] ), .Y(n1734) );
  AOI22X1TS U1844 ( .A0(n1729), .A1(n1760), .B0(n940), .B1(
        destinationAddressIn_EAST[0]), .Y(n1733) );
  AOI22X1TS U1845 ( .A0(n1731), .A1(n1860), .B0(n1730), .B1(n1858), .Y(n1732)
         );
  AOI22X1TS U1846 ( .A0(n1736), .A1(n1735), .B0(n1741), .B1(
        \destinationAddressbuffer[4][1] ), .Y(n1740) );
  AOI22X1TS U1847 ( .A0(n309), .A1(n1767), .B0(n1737), .B1(
        destinationAddressIn_EAST[1]), .Y(n1739) );
  AOI22X1TS U1848 ( .A0(n282), .A1(n1870), .B0(n920), .B1(n1868), .Y(n1738) );
  AOI22X1TS U1849 ( .A0(n1742), .A1(n277), .B0(n1741), .B1(
        \destinationAddressbuffer[4][2] ), .Y(n1747) );
  AOI22X1TS U1850 ( .A0(n1751), .A1(n1774), .B0(n1743), .B1(
        destinationAddressIn_EAST[2]), .Y(n1746) );
  AOI22X1TS U1851 ( .A0(n1744), .A1(n1879), .B0(n1752), .B1(n1878), .Y(n1745)
         );
  AOI22X1TS U1852 ( .A0(n1750), .A1(n1749), .B0(n1748), .B1(
        \destinationAddressbuffer[4][3] ), .Y(n1756) );
  AOI22X1TS U1853 ( .A0(n1751), .A1(n1783), .B0(n276), .B1(
        destinationAddressIn_EAST[3]), .Y(n1755) );
  AOI22X1TS U1854 ( .A0(n1753), .A1(n1890), .B0(n1752), .B1(n1888), .Y(n1754)
         );
  AOI22X1TS U1855 ( .A0(n1758), .A1(n1757), .B0(n1772), .B1(
        \destinationAddressbuffer[3][0] ), .Y(n1765) );
  AOI22X1TS U1856 ( .A0(n1761), .A1(n1760), .B0(n1759), .B1(
        destinationAddressIn_EAST[0]), .Y(n1764) );
  AOI22X1TS U1857 ( .A0(n1762), .A1(n1818), .B0(n1768), .B1(n1817), .Y(n1763)
         );
  AOI22X1TS U1858 ( .A0(n1824), .A1(n1766), .B0(n1772), .B1(
        \destinationAddressbuffer[3][1] ), .Y(n1771) );
  AOI22X1TS U1859 ( .A0(n1784), .A1(n1767), .B0(n146), .B1(
        destinationAddressIn_EAST[1]), .Y(n1770) );
  AOI22X1TS U1860 ( .A0(n1776), .A1(n1828), .B0(n1768), .B1(n1827), .Y(n1769)
         );
  AOI22X1TS U1861 ( .A0(n1835), .A1(n136), .B0(n1772), .B1(
        \destinationAddressbuffer[3][2] ), .Y(n1779) );
  AOI22X1TS U1862 ( .A0(n161), .A1(n1774), .B0(n1773), .B1(
        destinationAddressIn_EAST[2]), .Y(n1778) );
  AOI22X1TS U1863 ( .A0(n1776), .A1(n1840), .B0(n1775), .B1(n1838), .Y(n1777)
         );
  AOI22X1TS U1864 ( .A0(n1846), .A1(n1781), .B0(n1780), .B1(
        \destinationAddressbuffer[3][3] ), .Y(n1788) );
  AOI22X1TS U1865 ( .A0(n1784), .A1(n1783), .B0(n1782), .B1(
        destinationAddressIn_EAST[3]), .Y(n1787) );
  AOI22X1TS U1866 ( .A0(n958), .A1(n1850), .B0(n1785), .B1(n1849), .Y(n1786)
         );
  AOI22X1TS U1867 ( .A0(n1814), .A1(n1789), .B0(n1801), .B1(
        \destinationAddressbuffer[2][0] ), .Y(n1794) );
  AOI22X1TS U1868 ( .A0(n1790), .A1(destinationAddressIn_WEST[0]), .B0(n197), 
        .B1(n1815), .Y(n1793) );
  AOI22X1TS U1869 ( .A0(n1791), .A1(n1818), .B0(n190), .B1(n1817), .Y(n1792)
         );
  AOI22X1TS U1870 ( .A0(n1866), .A1(n1795), .B0(n1801), .B1(
        \destinationAddressbuffer[2][1] ), .Y(n1800) );
  AOI22X1TS U1871 ( .A0(n209), .A1(destinationAddressIn_WEST[1]), .B0(n1796), 
        .B1(n1825), .Y(n1799) );
  AOI22X1TS U1872 ( .A0(n1797), .A1(n1828), .B0(n1804), .B1(n1827), .Y(n1798)
         );
  AOI22X1TS U1873 ( .A0(n1876), .A1(n1802), .B0(n1801), .B1(
        \destinationAddressbuffer[2][2] ), .Y(n1807) );
  AOI22X1TS U1874 ( .A0(n1809), .A1(destinationAddressIn_WEST[2]), .B0(n1803), 
        .B1(n1836), .Y(n1806) );
  AOI22X1TS U1875 ( .A0(n1810), .A1(n1840), .B0(n1804), .B1(n1838), .Y(n1805)
         );
  AOI22X1TS U1876 ( .A0(n1886), .A1(n185), .B0(n1808), .B1(
        \destinationAddressbuffer[2][3] ), .Y(n1813) );
  AOI22X1TS U1877 ( .A0(n1809), .A1(destinationAddressIn_WEST[3]), .B0(n991), 
        .B1(n1847), .Y(n1812) );
  AOI22X1TS U1878 ( .A0(n1810), .A1(n1850), .B0(n190), .B1(n1849), .Y(n1811)
         );
  AOI22X1TS U1879 ( .A0(n1814), .A1(n1823), .B0(n1833), .B1(
        \destinationAddressbuffer[1][0] ), .Y(n1822) );
  AOI22X1TS U1880 ( .A0(n1816), .A1(destinationAddressIn_WEST[0]), .B0(n1018), 
        .B1(n1815), .Y(n1821) );
  AOI22X1TS U1881 ( .A0(n1819), .A1(n1818), .B0(n325), .B1(n1817), .Y(n1820)
         );
  AOI22X1TS U1882 ( .A0(n1824), .A1(n1823), .B0(n1833), .B1(
        \destinationAddressbuffer[1][1] ), .Y(n1832) );
  AOI22X1TS U1883 ( .A0(n358), .A1(destinationAddressIn_WEST[1]), .B0(n1826), 
        .B1(n1825), .Y(n1831) );
  AOI22X1TS U1884 ( .A0(n1829), .A1(n1828), .B0(n1839), .B1(n1827), .Y(n1830)
         );
  AOI22X1TS U1885 ( .A0(n1835), .A1(n1834), .B0(n1833), .B1(
        \destinationAddressbuffer[1][2] ), .Y(n1843) );
  AOI22X1TS U1886 ( .A0(n1848), .A1(destinationAddressIn_WEST[2]), .B0(n1837), 
        .B1(n1836), .Y(n1842) );
  AOI22X1TS U1887 ( .A0(n1851), .A1(n1840), .B0(n1839), .B1(n1838), .Y(n1841)
         );
  AOI22X1TS U1888 ( .A0(n1846), .A1(n1845), .B0(n1844), .B1(
        \destinationAddressbuffer[1][3] ), .Y(n1854) );
  AOI22X1TS U1889 ( .A0(n1848), .A1(destinationAddressIn_WEST[3]), .B0(n318), 
        .B1(n1847), .Y(n1853) );
  AOI22X1TS U1890 ( .A0(n1851), .A1(n1850), .B0(n325), .B1(n1849), .Y(n1852)
         );
  AOI22X1TS U1891 ( .A0(n1856), .A1(n1855), .B0(n1874), .B1(
        \destinationAddressbuffer[0][0] ), .Y(n1864) );
  AOI22X1TS U1892 ( .A0(n1857), .A1(destinationAddressIn_WEST[0]), .B0(n1045), 
        .B1(destinationAddressIn_EAST[0]), .Y(n1863) );
  AOI22X1TS U1893 ( .A0(n1861), .A1(n1860), .B0(n1859), .B1(n1858), .Y(n1862)
         );
  AOI22X1TS U1894 ( .A0(n1866), .A1(n1865), .B0(n1874), .B1(
        \destinationAddressbuffer[0][1] ), .Y(n1873) );
  AOI22X1TS U1895 ( .A0(n422), .A1(destinationAddressIn_WEST[1]), .B0(n1867), 
        .B1(destinationAddressIn_EAST[1]), .Y(n1872) );
  AOI22X1TS U1896 ( .A0(n415), .A1(n1870), .B0(n1869), .B1(n1868), .Y(n1871)
         );
  AOI22X1TS U1897 ( .A0(n1876), .A1(n1875), .B0(n1874), .B1(
        \destinationAddressbuffer[0][2] ), .Y(n1883) );
  AOI22X1TS U1898 ( .A0(n1887), .A1(destinationAddressIn_WEST[2]), .B0(n1877), 
        .B1(destinationAddressIn_EAST[2]), .Y(n1882) );
  AOI22X1TS U1899 ( .A0(n1880), .A1(n1879), .B0(n1889), .B1(n1878), .Y(n1881)
         );
  AOI22X1TS U1900 ( .A0(n1886), .A1(n1885), .B0(n1884), .B1(
        \destinationAddressbuffer[0][3] ), .Y(n1894) );
  AOI22X1TS U1901 ( .A0(n1887), .A1(destinationAddressIn_WEST[3]), .B0(n393), 
        .B1(destinationAddressIn_EAST[3]), .Y(n1893) );
  AOI22X1TS U1902 ( .A0(n1891), .A1(n1890), .B0(n1889), .B1(n1888), .Y(n1892)
         );
endmodule


module outputPortArbiter_2 ( clk, reset, selectBit_NORTH, 
        destinationAddressIn_NORTH, requesterAddressIn_NORTH, readIn_NORTH, 
        writeIn_NORTH, dataIn_NORTH, selectBit_SOUTH, 
        destinationAddressIn_SOUTH, requesterAddressIn_SOUTH, readIn_SOUTH, 
        writeIn_SOUTH, dataIn_SOUTH, selectBit_EAST, destinationAddressIn_EAST, 
        requesterAddressIn_EAST, readIn_EAST, writeIn_EAST, dataIn_EAST, 
        selectBit_WEST, destinationAddressIn_WEST, requesterAddressIn_WEST, 
        readIn_WEST, writeIn_WEST, dataIn_WEST, readReady, 
        readRequesterAddress, cacheDataOut, destinationAddressOut, 
        requesterAddressOut, readOut, writeOut, dataOut );
  input [11:0] destinationAddressIn_NORTH;
  input [3:0] requesterAddressIn_NORTH;
  input [5:0] dataIn_NORTH;
  input [11:0] destinationAddressIn_SOUTH;
  input [3:0] requesterAddressIn_SOUTH;
  input [5:0] dataIn_SOUTH;
  input [11:0] destinationAddressIn_EAST;
  input [3:0] requesterAddressIn_EAST;
  input [5:0] dataIn_EAST;
  input [11:0] destinationAddressIn_WEST;
  input [3:0] requesterAddressIn_WEST;
  input [5:0] dataIn_WEST;
  input [3:0] readRequesterAddress;
  input [5:0] cacheDataOut;
  output [11:0] destinationAddressOut;
  output [3:0] requesterAddressOut;
  output [5:0] dataOut;
  input clk, reset, selectBit_NORTH, readIn_NORTH, writeIn_NORTH,
         selectBit_SOUTH, readIn_SOUTH, writeIn_SOUTH, selectBit_EAST,
         readIn_EAST, writeIn_EAST, selectBit_WEST, readIn_WEST, writeIn_WEST,
         readReady;
  output readOut, writeOut;
  wire   \requesterAddressbuffer[0][3] , \requesterAddressbuffer[0][2] ,
         \requesterAddressbuffer[0][1] , \requesterAddressbuffer[0][0] ,
         \requesterAddressbuffer[1][3] , \requesterAddressbuffer[1][2] ,
         \requesterAddressbuffer[1][1] , \requesterAddressbuffer[1][0] ,
         \requesterAddressbuffer[2][3] , \requesterAddressbuffer[2][2] ,
         \requesterAddressbuffer[2][1] , \requesterAddressbuffer[2][0] ,
         \requesterAddressbuffer[3][3] , \requesterAddressbuffer[3][2] ,
         \requesterAddressbuffer[3][1] , \requesterAddressbuffer[3][0] ,
         \requesterAddressbuffer[4][3] , \requesterAddressbuffer[4][2] ,
         \requesterAddressbuffer[4][1] , \requesterAddressbuffer[4][0] ,
         \requesterAddressbuffer[5][3] , \requesterAddressbuffer[5][2] ,
         \requesterAddressbuffer[5][1] , \requesterAddressbuffer[5][0] ,
         \requesterAddressbuffer[6][3] , \requesterAddressbuffer[6][2] ,
         \requesterAddressbuffer[6][1] , \requesterAddressbuffer[6][0] ,
         \requesterAddressbuffer[7][3] , \requesterAddressbuffer[7][2] ,
         \requesterAddressbuffer[7][1] , \requesterAddressbuffer[7][0] ,
         \destinationAddressbuffer[0][11] , \destinationAddressbuffer[0][10] ,
         \destinationAddressbuffer[0][9] , \destinationAddressbuffer[0][8] ,
         \destinationAddressbuffer[0][7] , \destinationAddressbuffer[0][6] ,
         \destinationAddressbuffer[0][5] , \destinationAddressbuffer[0][4] ,
         \destinationAddressbuffer[0][3] , \destinationAddressbuffer[0][2] ,
         \destinationAddressbuffer[0][1] , \destinationAddressbuffer[0][0] ,
         \destinationAddressbuffer[1][11] , \destinationAddressbuffer[1][10] ,
         \destinationAddressbuffer[1][9] , \destinationAddressbuffer[1][8] ,
         \destinationAddressbuffer[1][7] , \destinationAddressbuffer[1][6] ,
         \destinationAddressbuffer[1][5] , \destinationAddressbuffer[1][4] ,
         \destinationAddressbuffer[1][3] , \destinationAddressbuffer[1][2] ,
         \destinationAddressbuffer[1][1] , \destinationAddressbuffer[1][0] ,
         \destinationAddressbuffer[2][11] , \destinationAddressbuffer[2][10] ,
         \destinationAddressbuffer[2][9] , \destinationAddressbuffer[2][8] ,
         \destinationAddressbuffer[2][7] , \destinationAddressbuffer[2][6] ,
         \destinationAddressbuffer[2][5] , \destinationAddressbuffer[2][4] ,
         \destinationAddressbuffer[2][3] , \destinationAddressbuffer[2][2] ,
         \destinationAddressbuffer[2][1] , \destinationAddressbuffer[2][0] ,
         \destinationAddressbuffer[3][11] , \destinationAddressbuffer[3][10] ,
         \destinationAddressbuffer[3][9] , \destinationAddressbuffer[3][8] ,
         \destinationAddressbuffer[3][7] , \destinationAddressbuffer[3][6] ,
         \destinationAddressbuffer[3][5] , \destinationAddressbuffer[3][4] ,
         \destinationAddressbuffer[3][3] , \destinationAddressbuffer[3][2] ,
         \destinationAddressbuffer[3][1] , \destinationAddressbuffer[3][0] ,
         \destinationAddressbuffer[4][11] , \destinationAddressbuffer[4][10] ,
         \destinationAddressbuffer[4][9] , \destinationAddressbuffer[4][8] ,
         \destinationAddressbuffer[4][7] , \destinationAddressbuffer[4][6] ,
         \destinationAddressbuffer[4][5] , \destinationAddressbuffer[4][4] ,
         \destinationAddressbuffer[4][3] , \destinationAddressbuffer[4][2] ,
         \destinationAddressbuffer[4][1] , \destinationAddressbuffer[4][0] ,
         \destinationAddressbuffer[5][11] , \destinationAddressbuffer[5][10] ,
         \destinationAddressbuffer[5][9] , \destinationAddressbuffer[5][8] ,
         \destinationAddressbuffer[5][7] , \destinationAddressbuffer[5][6] ,
         \destinationAddressbuffer[5][5] , \destinationAddressbuffer[5][4] ,
         \destinationAddressbuffer[5][3] , \destinationAddressbuffer[5][2] ,
         \destinationAddressbuffer[5][1] , \destinationAddressbuffer[5][0] ,
         \destinationAddressbuffer[6][11] , \destinationAddressbuffer[6][10] ,
         \destinationAddressbuffer[6][9] , \destinationAddressbuffer[6][8] ,
         \destinationAddressbuffer[6][7] , \destinationAddressbuffer[6][6] ,
         \destinationAddressbuffer[6][5] , \destinationAddressbuffer[6][4] ,
         \destinationAddressbuffer[6][3] , \destinationAddressbuffer[6][2] ,
         \destinationAddressbuffer[6][1] , \destinationAddressbuffer[6][0] ,
         \destinationAddressbuffer[7][11] , \destinationAddressbuffer[7][10] ,
         \destinationAddressbuffer[7][9] , \destinationAddressbuffer[7][8] ,
         \destinationAddressbuffer[7][7] , \destinationAddressbuffer[7][6] ,
         \destinationAddressbuffer[7][5] , \destinationAddressbuffer[7][4] ,
         \destinationAddressbuffer[7][3] , \destinationAddressbuffer[7][2] ,
         \destinationAddressbuffer[7][1] , \destinationAddressbuffer[7][0] ,
         \dataoutbuffer[7][5] , \dataoutbuffer[7][4] , \dataoutbuffer[7][3] ,
         \dataoutbuffer[7][2] , \dataoutbuffer[7][1] , \dataoutbuffer[7][0] ,
         \dataoutbuffer[6][5] , \dataoutbuffer[6][4] , \dataoutbuffer[6][3] ,
         \dataoutbuffer[6][2] , \dataoutbuffer[6][1] , \dataoutbuffer[6][0] ,
         \dataoutbuffer[5][5] , \dataoutbuffer[5][4] , \dataoutbuffer[5][3] ,
         \dataoutbuffer[5][2] , \dataoutbuffer[5][1] , \dataoutbuffer[5][0] ,
         \dataoutbuffer[4][5] , \dataoutbuffer[4][4] , \dataoutbuffer[4][3] ,
         \dataoutbuffer[4][2] , \dataoutbuffer[4][1] , \dataoutbuffer[4][0] ,
         \dataoutbuffer[3][5] , \dataoutbuffer[3][4] , \dataoutbuffer[3][3] ,
         \dataoutbuffer[3][2] , \dataoutbuffer[3][1] , \dataoutbuffer[3][0] ,
         \dataoutbuffer[2][5] , \dataoutbuffer[2][4] , \dataoutbuffer[2][3] ,
         \dataoutbuffer[2][2] , \dataoutbuffer[2][1] , \dataoutbuffer[2][0] ,
         \dataoutbuffer[1][5] , \dataoutbuffer[1][4] , \dataoutbuffer[1][3] ,
         \dataoutbuffer[1][2] , \dataoutbuffer[1][1] , \dataoutbuffer[1][0] ,
         \dataoutbuffer[0][5] , \dataoutbuffer[0][4] , \dataoutbuffer[0][3] ,
         \dataoutbuffer[0][2] , \dataoutbuffer[0][1] , \dataoutbuffer[0][0] ,
         N2624, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145;
  wire   [0:7] writeOutbuffer;
  wire   [0:7] readOutbuffer;

  DFFNSRX1TS full_reg_reg ( .D(N2624), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(
        n1914) );
  DFFNSRX1TS \dataoutbuffer_reg[0][0]  ( .D(n1986), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][1]  ( .D(n1987), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][2]  ( .D(n1988), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][3]  ( .D(n1989), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][4]  ( .D(n1990), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][5]  ( .D(n1991), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][5] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[2][0]  ( .D(n1974), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[2][1]  ( .D(n1975), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[2][2]  ( .D(n1976), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[2][3]  ( .D(n1977), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][0]  ( .D(n2110), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][1]  ( .D(n2111), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][2]  ( .D(n2112), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][3]  ( .D(n2113), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][3] ) );
  DFFNSRX1TS \writeOutbuffer_reg[7]  ( .D(n2034), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[7]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][4]  ( .D(n2054), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][5]  ( .D(n2055), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][6]  ( .D(n2056), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][7]  ( .D(n2057), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][8]  ( .D(n2058), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][9]  ( .D(n2059), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][11]  ( .D(n2061), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[6]  ( .D(n2035), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[6]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][4]  ( .D(n2066), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][5]  ( .D(n2067), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][6]  ( .D(n2068), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][7]  ( .D(n2069), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][8]  ( .D(n2070), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][9]  ( .D(n2071), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][10]  ( .D(n2072), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][11]  ( .D(n2073), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[3]  ( .D(n2038), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[3]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][4]  ( .D(n2102), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][5]  ( .D(n2103), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][6]  ( .D(n2104), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][7]  ( .D(n2105), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][8]  ( .D(n2106), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][9]  ( .D(n2107), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][10]  ( .D(n2108), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][11]  ( .D(n2109), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[2]  ( .D(n2039), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[2]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][4]  ( .D(n2114), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][5]  ( .D(n2115), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][6]  ( .D(n2116), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][7]  ( .D(n2117), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][8]  ( .D(n2118), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][9]  ( .D(n2119), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][10]  ( .D(n2120), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][11]  ( .D(n2121), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][11] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][0]  ( .D(n2028), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][1]  ( .D(n2029), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][2]  ( .D(n2030), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][3]  ( .D(n2031), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][4]  ( .D(n2032), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][5]  ( .D(n2033), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][0]  ( .D(n2022), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][1]  ( .D(n2023), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][2]  ( .D(n2024), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][3]  ( .D(n2025), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][4]  ( .D(n2026), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][5]  ( .D(n2027), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][0]  ( .D(n2004), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][1]  ( .D(n2005), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][2]  ( .D(n2006), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][3]  ( .D(n2007), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][4]  ( .D(n2008), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][5]  ( .D(n2009), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][0]  ( .D(n1998), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][1]  ( .D(n1999), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][2]  ( .D(n2000), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][3]  ( .D(n2001), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][4]  ( .D(n2002), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][5]  ( .D(n2003), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][5] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[5][0]  ( .D(n1962), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[5][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[5][1]  ( .D(n1963), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[5][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[5][2]  ( .D(n1964), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[5][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[5][3]  ( .D(n1965), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[5][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][0]  ( .D(n2074), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][1]  ( .D(n2075), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][2]  ( .D(n2076), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][3]  ( .D(n2077), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[4][0]  ( .D(n1966), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[4][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[4][1]  ( .D(n1967), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[4][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[4][2]  ( .D(n1968), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[4][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[4][3]  ( .D(n1969), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[4][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][0]  ( .D(n2086), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][1]  ( .D(n2087), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][2]  ( .D(n2088), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][3]  ( .D(n2089), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[1][0]  ( .D(n1978), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[1][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[1][1]  ( .D(n1979), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[1][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[1][2]  ( .D(n1980), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[1][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[1][3]  ( .D(n1981), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[1][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][0]  ( .D(n2122), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][1]  ( .D(n2123), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][2]  ( .D(n2124), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][3]  ( .D(n2125), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[0][0]  ( .D(n1982), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[0][1]  ( .D(n1983), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[0][2]  ( .D(n1984), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[0][3]  ( .D(n1985), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][0]  ( .D(n2134), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][1]  ( .D(n2135), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][2]  ( .D(n2136), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][3]  ( .D(n2137), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][0]  ( .D(n2016), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][1]  ( .D(n2017), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][2]  ( .D(n2018), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][3]  ( .D(n2019), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][4]  ( .D(n2020), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][5]  ( .D(n2021), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][0]  ( .D(n2010), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][1]  ( .D(n2011), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][2]  ( .D(n2012), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][3]  ( .D(n2013), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][4]  ( .D(n2014), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][5]  ( .D(n2015), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][0]  ( .D(n1992), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][1]  ( .D(n1993), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][2]  ( .D(n1994), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][3]  ( .D(n1995), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][4]  ( .D(n1996), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][5]  ( .D(n1997), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][5] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[7][0]  ( .D(n1954), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[7][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[7][1]  ( .D(n1955), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[7][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[7][2]  ( .D(n1956), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[7][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[7][3]  ( .D(n1957), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[7][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][0]  ( .D(n2050), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][1]  ( .D(n2051), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][2]  ( .D(n2052), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][3]  ( .D(n2053), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[6][0]  ( .D(n1958), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[6][1]  ( .D(n1959), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[6][2]  ( .D(n1960), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[6][3]  ( .D(n1961), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][0]  ( .D(n2062), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][1]  ( .D(n2063), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][2]  ( .D(n2064), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][3]  ( .D(n2065), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[3][0]  ( .D(n1970), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[3][1]  ( .D(n1971), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[3][2]  ( .D(n1972), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[3][3]  ( .D(n1973), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][0]  ( .D(n2098), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][1]  ( .D(n2099), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][2]  ( .D(n2100), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][3]  ( .D(n2101), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][3] ) );
  DFFNSRX1TS \writeOutbuffer_reg[5]  ( .D(n2036), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[5]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][4]  ( .D(n2078), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][5]  ( .D(n2079), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][6]  ( .D(n2080), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][7]  ( .D(n2081), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][8]  ( .D(n2082), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][9]  ( .D(n2083), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][10]  ( .D(n2084), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][11]  ( .D(n2085), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[4]  ( .D(n2037), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[4]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][4]  ( .D(n2090), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][5]  ( .D(n2091), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][6]  ( .D(n2092), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][7]  ( .D(n2093), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][8]  ( .D(n2094), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][9]  ( .D(n2095), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][10]  ( .D(n2096), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][11]  ( .D(n2097), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[1]  ( .D(n2040), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[1]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][4]  ( .D(n2126), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][5]  ( .D(n2127), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][6]  ( .D(n2128), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][7]  ( .D(n2129), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][8]  ( .D(n2130), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][9]  ( .D(n2131), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][10]  ( .D(n2132), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][11]  ( .D(n2133), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[0]  ( .D(n2041), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[0]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][4]  ( .D(n2138), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][5]  ( .D(n2139), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][6]  ( .D(n2140), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][7]  ( .D(n2141), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][8]  ( .D(n2142), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][9]  ( .D(n2143), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][10]  ( .D(n2144), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][11]  ( .D(n2145), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][11] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][10]  ( .D(n2060), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][10] ) );
  DFFNSRX1TS writeOut_reg ( .D(n1931), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        writeOut) );
  DFFNSRX1TS \destinationAddressOut_reg[4]  ( .D(n1940), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[4]) );
  DFFNSRX1TS \destinationAddressOut_reg[5]  ( .D(n1941), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[5]) );
  DFFNSRX1TS \destinationAddressOut_reg[6]  ( .D(n1942), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[6]) );
  DFFNSRX1TS \destinationAddressOut_reg[7]  ( .D(n1943), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[7]) );
  DFFNSRX1TS \destinationAddressOut_reg[8]  ( .D(n1944), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[8]) );
  DFFNSRX1TS \destinationAddressOut_reg[9]  ( .D(n1945), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[9]) );
  DFFNSRX1TS \destinationAddressOut_reg[10]  ( .D(n1946), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[10]) );
  DFFNSRX1TS \destinationAddressOut_reg[11]  ( .D(n1947), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[11]) );
  DFFNSRX1TS readOut_reg ( .D(n1930), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        readOut) );
  DFFNSRX1TS \requesterAddressOut_reg[0]  ( .D(n1932), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[0]) );
  DFFNSRX1TS \requesterAddressOut_reg[1]  ( .D(n1933), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[1]) );
  DFFNSRX1TS \requesterAddressOut_reg[2]  ( .D(n1934), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[2]) );
  DFFNSRX1TS \requesterAddressOut_reg[3]  ( .D(n1935), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[3]) );
  DFFNSRX1TS \destinationAddressOut_reg[0]  ( .D(n1936), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[0]) );
  DFFNSRX1TS \destinationAddressOut_reg[1]  ( .D(n1937), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[1]) );
  DFFNSRX1TS \destinationAddressOut_reg[2]  ( .D(n1938), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[2]) );
  DFFNSRX1TS \destinationAddressOut_reg[3]  ( .D(n1939), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[3]) );
  DFFNSRX1TS \dataOut_reg[0]  ( .D(n1948), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[0]) );
  DFFNSRX1TS \dataOut_reg[1]  ( .D(n1949), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[1]) );
  DFFNSRX1TS \dataOut_reg[2]  ( .D(n1950), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[2]) );
  DFFNSRX1TS \dataOut_reg[3]  ( .D(n1951), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[3]) );
  DFFNSRX1TS \dataOut_reg[4]  ( .D(n1952), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[4]) );
  DFFNSRX1TS \dataOut_reg[5]  ( .D(n1953), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[5]) );
  DFFNSRX1TS \read_reg_reg[1]  ( .D(n1929), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1907), .QN(n1906) );
  DFFNSRX1TS \write_reg_reg[0]  ( .D(n1924), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1905), .QN(n1909) );
  DFFNSRX1TS \write_reg_reg[2]  ( .D(n1926), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1910), .QN(n1911) );
  DFFNSRX1TS \read_reg_reg[0]  ( .D(n1923), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1900), .QN(n1913) );
  DFFNSRX1TS \read_reg_reg[2]  ( .D(n1928), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1903), .QN(n1904) );
  DFFNSRX1TS empty_reg_reg ( .D(n1927), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        n1902), .QN(n1901) );
  DFFNSRX1TS \readOutbuffer_reg[7]  ( .D(n2042), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[7]), .QN(n1915) );
  DFFNSRX1TS \readOutbuffer_reg[4]  ( .D(n2045), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[4]), .QN(n1918) );
  DFFNSRX1TS \readOutbuffer_reg[6]  ( .D(n2043), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[6]), .QN(n1916) );
  DFFNSRX1TS \readOutbuffer_reg[5]  ( .D(n2044), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[5]), .QN(n1917) );
  DFFNSRX1TS \readOutbuffer_reg[3]  ( .D(n2046), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[3]), .QN(n1919) );
  DFFNSRX1TS \readOutbuffer_reg[0]  ( .D(n2049), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[0]), .QN(n1922) );
  DFFNSRX1TS \readOutbuffer_reg[2]  ( .D(n2047), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[2]), .QN(n1920) );
  DFFNSRX1TS \readOutbuffer_reg[1]  ( .D(n2048), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[1]), .QN(n1921) );
  DFFNSRX1TS \write_reg_reg[1]  ( .D(n1925), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1908), .QN(n1912) );
  CMPR32X2TS U3 ( .A(n485), .B(n484), .C(n483), .CO(n478), .S(n493) );
  CLKBUFX2TS U4 ( .A(n12), .Y(n72) );
  CMPR32X2TS U5 ( .A(n463), .B(n484), .C(n14), .CO(n15), .S(n12) );
  CMPR32X2TS U6 ( .A(n530), .B(n461), .C(n460), .CO(n452), .S(n466) );
  CMPR32X2TS U7 ( .A(n459), .B(n511), .C(n458), .CO(n462), .S(n475) );
  CMPR32X2TS U8 ( .A(selectBit_SOUTH), .B(selectBit_NORTH), .C(selectBit_EAST), 
        .CO(n463), .S(n458) );
  INVX2TS U9 ( .A(n1575), .Y(n1574) );
  OAI31X1TS U10 ( .A0(n516), .A1(n515), .A2(n537), .B0(n538), .Y(n518) );
  OR2X1TS U11 ( .A(n19), .B(n506), .Y(n8) );
  CLKBUFX2TS U12 ( .A(n18), .Y(n74) );
  ADDHXLTS U13 ( .A(n447), .B(n458), .CO(n14), .S(n13) );
  NAND2X1TS U14 ( .A(n538), .B(n520), .Y(n508) );
  INVX2TS U15 ( .A(selectBit_EAST), .Y(n510) );
  NOR2XLTS U16 ( .A(n840), .B(n519), .Y(n689) );
  NOR3XLTS U17 ( .A(n385), .B(n74), .C(n266), .Y(n1575) );
  INVX2TS U18 ( .A(n1556), .Y(n1554) );
  INVX2TS U19 ( .A(n1600), .Y(n1597) );
  INVX2TS U20 ( .A(n1616), .Y(n1613) );
  NOR3XLTS U21 ( .A(n13), .B(n174), .C(n381), .Y(n1603) );
  AOI31XLTS U22 ( .A0(n217), .A1(n1562), .A2(n214), .B0(n392), .Y(n216) );
  INVX2TS U23 ( .A(n1582), .Y(n1579) );
  NOR2XLTS U24 ( .A(n1575), .B(n275), .Y(n276) );
  NOR2XLTS U25 ( .A(n1609), .B(n326), .Y(n324) );
  CLKBUFX2TS U26 ( .A(n1087), .Y(n1082) );
  NOR2XLTS U27 ( .A(n387), .B(n1583), .Y(n271) );
  NOR2XLTS U28 ( .A(n1565), .B(n220), .Y(n219) );
  NOR2XLTS U29 ( .A(n441), .B(n1592), .Y(n126) );
  NOR2XLTS U30 ( .A(n316), .B(n1560), .Y(n78) );
  NOR2XLTS U31 ( .A(n1589), .B(n130), .Y(n131) );
  NOR2XLTS U32 ( .A(n1552), .B(n83), .Y(n84) );
  NOR3XLTS U33 ( .A(n1549), .B(n1544), .C(n30), .Y(n26) );
  NOR3XLTS U34 ( .A(n1603), .B(n1597), .C(n181), .Y(n176) );
  NOR2XLTS U35 ( .A(n1596), .B(n184), .Y(n182) );
  CLKBUFX2TS U36 ( .A(n1343), .Y(n1337) );
  NOR3XLTS U37 ( .A(n1628), .B(n1622), .C(n396), .Y(n391) );
  INVX2TS U38 ( .A(reset), .Y(n491) );
  NOR3XLTS U39 ( .A(n1571), .B(n1566), .C(n218), .Y(n1) );
  NOR2X1TS U40 ( .A(n1574), .B(n275), .Y(n279) );
  NOR2X1TS U41 ( .A(n115), .B(n128), .Y(n140) );
  NOR2X1TS U42 ( .A(n1585), .B(n128), .Y(n124) );
  NAND2BX1TS U43 ( .AN(n396), .B(n395), .Y(n397) );
  NAND2BX1TS U44 ( .AN(n181), .B(n180), .Y(n184) );
  NOR2X1TS U45 ( .A(n1543), .B(n31), .Y(n40) );
  NAND2BX1TS U46 ( .AN(n30), .B(n29), .Y(n31) );
  NOR3X1TS U47 ( .A(n1591), .B(n1586), .C(n130), .Y(n135) );
  NOR3X1TS U48 ( .A(n1616), .B(n1610), .C(n323), .Y(n318) );
  NOR2X1TS U49 ( .A(n1628), .B(n1625), .Y(n395) );
  AOI31X1TS U50 ( .A0(n123), .A1(n1585), .A2(n121), .B0(n392), .Y(n127) );
  AOI31X1TS U51 ( .A0(n29), .A1(n25), .A2(n1542), .B0(n316), .Y(n28) );
  NOR2X1TS U52 ( .A(n1591), .B(n1588), .Y(n123) );
  INVX1TS U53 ( .A(n1568), .Y(n1566) );
  NOR2X1TS U54 ( .A(n1549), .B(n1546), .Y(n29) );
  INVX1TS U55 ( .A(n1546), .Y(n1544) );
  INVX1TS U56 ( .A(n1612), .Y(n1610) );
  NOR3BX1TS U57 ( .AN(n384), .B(n383), .C(n382), .Y(n1625) );
  INVX1TS U58 ( .A(n1578), .Y(n1576) );
  NOR2X1TS U59 ( .A(n119), .B(n383), .Y(n1588) );
  NOR2X1TS U60 ( .A(n119), .B(n264), .Y(n1546) );
  NAND2BX1TS U61 ( .AN(n118), .B(n513), .Y(n383) );
  NOR3X1TS U62 ( .A(n75), .B(n74), .C(n265), .Y(n1553) );
  OAI21X1TS U63 ( .A0(selectBit_SOUTH), .A1(n19), .B0(n74), .Y(n263) );
  NOR3X1TS U64 ( .A(n313), .B(n74), .C(n265), .Y(n1596) );
  NAND3X1TS U65 ( .A(n313), .B(n213), .C(n265), .Y(n1562) );
  NOR2X1TS U66 ( .A(n213), .B(n73), .Y(n311) );
  NOR3X1TS U67 ( .A(n23), .B(n385), .C(n18), .Y(n1621) );
  NAND3X1TS U68 ( .A(n445), .B(n23), .C(n213), .Y(n1542) );
  INVX1TS U69 ( .A(n1559), .Y(n1557) );
  NOR2X1TS U70 ( .A(n387), .B(n1604), .Y(n177) );
  NOR3X1TS U71 ( .A(n313), .B(n385), .C(n8), .Y(n1609) );
  INVX1TS U72 ( .A(n1603), .Y(n1601) );
  INVX1TS U73 ( .A(n1591), .Y(n1589) );
  INVX1TS U74 ( .A(n1628), .Y(n1626) );
  NOR2X1TS U75 ( .A(n8), .B(n73), .Y(n22) );
  NOR3X1TS U76 ( .A(n174), .B(n71), .C(n381), .Y(n1591) );
  INVX1TS U77 ( .A(n1571), .Y(n1569) );
  NOR3X1TS U78 ( .A(n12), .B(n13), .C(n381), .Y(n1628) );
  INVX1TS U79 ( .A(n7), .Y(n73) );
  NOR3X1TS U80 ( .A(n12), .B(n71), .C(n262), .Y(n1571) );
  NOR3X1TS U81 ( .A(n72), .B(n71), .C(n381), .Y(n1616) );
  NOR2X1TS U82 ( .A(n840), .B(n517), .Y(n543) );
  INVX1TS U83 ( .A(n20), .Y(n120) );
  NOR2X1TS U84 ( .A(selectBit_NORTH), .B(n505), .Y(n538) );
  CLKINVX1TS U85 ( .A(n16), .Y(n17) );
  NOR2X1TS U86 ( .A(n457), .B(n504), .Y(n16) );
  NOR3X1TS U87 ( .A(n512), .B(selectBit_EAST), .C(n511), .Y(n507) );
  INVX1TS U88 ( .A(n1911), .Y(n498) );
  NAND2BX2TS U89 ( .AN(n117), .B(n459), .Y(n381) );
  INVX2TS U90 ( .A(n325), .Y(n345) );
  INVX2TS U91 ( .A(n219), .Y(n253) );
  NAND2BX1TS U92 ( .AN(n130), .B(n123), .Y(n128) );
  NAND2X1TS U93 ( .A(n127), .B(n1592), .Y(n130) );
  INVX2TS U94 ( .A(n183), .Y(n194) );
  XOR2X1TS U95 ( .A(n480), .B(n479), .Y(n495) );
  XNOR2X1TS U96 ( .A(n1910), .B(n478), .Y(n479) );
  NAND4XLTS U97 ( .A(n494), .B(n509), .C(n390), .D(n442), .Y(n1604) );
  INVX2TS U98 ( .A(n1625), .Y(n1622) );
  NAND4XLTS U99 ( .A(n494), .B(n482), .C(readReady), .D(n444), .Y(n1592) );
  NAND4XLTS U100 ( .A(n447), .B(n498), .C(readReady), .D(n314), .Y(n1572) );
  NAND4XLTS U101 ( .A(n445), .B(n498), .C(n509), .D(n390), .Y(n1560) );
  NOR3XLTS U102 ( .A(n13), .B(n174), .C(n262), .Y(n1559) );
  NAND4XLTS U103 ( .A(n269), .B(n514), .C(n390), .D(n314), .Y(n1583) );
  NOR3XLTS U104 ( .A(n72), .B(n116), .C(n262), .Y(n1582) );
  CLKAND2X2TS U105 ( .A(n523), .B(n521), .Y(n551) );
  INVX2TS U106 ( .A(n1422), .Y(n1451) );
  CLKAND2X2TS U107 ( .A(n477), .B(n475), .Y(n481) );
  NOR2XLTS U108 ( .A(reset), .B(n24), .Y(n496) );
  INVX2TS U109 ( .A(selectBit_NORTH), .Y(n504) );
  AO21X1TS U110 ( .A0(n457), .A1(n504), .B0(n315), .Y(n19) );
  NOR3BXLTS U111 ( .AN(n514), .B(selectBit_WEST), .C(n513), .Y(n537) );
  NAND3XLTS U112 ( .A(n505), .B(n507), .C(n504), .Y(n517) );
  NAND3XLTS U113 ( .A(selectBit_NORTH), .B(n507), .C(n506), .Y(n519) );
  NOR2XLTS U114 ( .A(n1582), .B(n1578), .Y(n273) );
  NOR2XLTS U115 ( .A(n1616), .B(n1612), .Y(n322) );
  NOR2XLTS U116 ( .A(n1571), .B(n1568), .Y(n217) );
  NOR2XLTS U117 ( .A(n1559), .B(n1556), .Y(n80) );
  NOR2XLTS U118 ( .A(n1603), .B(n1600), .Y(n180) );
  XOR2XLTS U119 ( .A(n452), .B(n454), .Y(n472) );
  OAI21XLTS U120 ( .A0(n455), .A1(n1906), .B0(n454), .Y(n456) );
  NAND3XLTS U121 ( .A(n315), .B(n451), .C(n389), .Y(n214) );
  INVX2TS U122 ( .A(n265), .Y(n385) );
  XOR2X1TS U123 ( .A(n498), .B(n15), .Y(n117) );
  NAND2BXLTS U124 ( .AN(n274), .B(n273), .Y(n275) );
  NAND2BXLTS U125 ( .AN(n81), .B(n80), .Y(n83) );
  CLKAND2X2TS U126 ( .A(n477), .B(n476), .Y(n483) );
  NOR2XLTS U127 ( .A(n267), .B(reset), .Y(n497) );
  NAND4XLTS U128 ( .A(n1905), .B(readReady), .C(n442), .D(n389), .Y(n1617) );
  INVX2TS U129 ( .A(n1609), .Y(n1607) );
  NOR3XLTS U130 ( .A(n312), .B(n311), .C(n383), .Y(n1612) );
  INVX2TS U131 ( .A(n1596), .Y(n1594) );
  NAND4XLTS U132 ( .A(n509), .B(n390), .C(n389), .D(n442), .Y(n1629) );
  INVX2TS U133 ( .A(n1621), .Y(n1620) );
  INVX2TS U134 ( .A(n1588), .Y(n1586) );
  NOR3XLTS U135 ( .A(n312), .B(n311), .C(n264), .Y(n1568) );
  INVX2TS U136 ( .A(n1553), .Y(n1552) );
  NOR3BXLTS U137 ( .AN(n384), .B(n264), .C(n263), .Y(n1578) );
  NAND4XLTS U138 ( .A(n72), .B(n116), .C(n117), .D(selectBit_WEST), .Y(n1547)
         );
  NAND4XLTS U139 ( .A(n482), .B(n484), .C(n269), .D(n514), .Y(n1550) );
  INVX2TS U140 ( .A(n1542), .Y(n1543) );
  INVX2TS U141 ( .A(n1422), .Y(n257) );
  INVX2TS U142 ( .A(destinationAddressIn_SOUTH[11]), .Y(n154) );
  INVX2TS U143 ( .A(destinationAddressIn_SOUTH[10]), .Y(n162) );
  INVX2TS U144 ( .A(destinationAddressIn_SOUTH[9]), .Y(n168) );
  INVX2TS U145 ( .A(destinationAddressIn_SOUTH[8]), .Y(n158) );
  AO22XLTS U146 ( .A0(n498), .A1(n497), .B0(n496), .B1(n495), .Y(n1926) );
  AO22XLTS U147 ( .A0(n1905), .A1(n497), .B0(n496), .B1(n492), .Y(n1924) );
  AO22XLTS U148 ( .A0(n494), .A1(n497), .B0(n496), .B1(n493), .Y(n1925) );
  OAI21XLTS U149 ( .A0(n267), .A1(n449), .B0(n491), .Y(n1927) );
  NAND4XLTS U150 ( .A(n866), .B(n865), .C(n864), .D(n863), .Y(n1953) );
  NAND4XLTS U151 ( .A(n844), .B(n843), .C(n842), .D(n863), .Y(n1952) );
  NAND4XLTS U152 ( .A(n833), .B(n832), .C(n831), .D(n863), .Y(n1951) );
  NAND4XLTS U153 ( .A(n823), .B(n822), .C(n821), .D(n863), .Y(n1950) );
  NAND4XLTS U154 ( .A(n804), .B(n803), .C(n802), .D(n801), .Y(n1949) );
  NAND4XLTS U155 ( .A(n784), .B(n783), .C(n782), .D(n801), .Y(n1948) );
  NAND4XLTS U156 ( .A(n655), .B(n654), .C(n653), .D(n652), .Y(n1939) );
  NAND4XLTS U157 ( .A(n644), .B(n643), .C(n642), .D(n641), .Y(n1938) );
  NAND4XLTS U158 ( .A(n626), .B(n625), .C(n624), .D(n623), .Y(n1937) );
  NAND4XLTS U159 ( .A(n611), .B(n610), .C(n609), .D(n608), .Y(n1936) );
  NAND4XLTS U160 ( .A(n599), .B(n598), .C(n597), .D(n652), .Y(n1935) );
  NAND4XLTS U161 ( .A(n588), .B(n587), .C(n586), .D(n641), .Y(n1934) );
  NAND4XLTS U162 ( .A(n579), .B(n578), .C(n577), .D(n623), .Y(n1933) );
  NAND4XLTS U163 ( .A(n562), .B(n561), .C(n560), .D(n608), .Y(n1932) );
  NAND4XLTS U164 ( .A(n541), .B(n540), .C(n539), .D(n801), .Y(n1930) );
  NAND3XLTS U165 ( .A(n774), .B(n773), .C(n772), .Y(n1947) );
  NAND3XLTS U166 ( .A(n760), .B(n759), .C(n758), .Y(n1946) );
  NAND3XLTS U167 ( .A(n744), .B(n743), .C(n742), .Y(n1945) );
  NAND3XLTS U168 ( .A(n726), .B(n725), .C(n724), .Y(n1944) );
  NAND3XLTS U169 ( .A(n712), .B(n711), .C(n710), .Y(n1943) );
  NAND3XLTS U170 ( .A(n701), .B(n700), .C(n699), .Y(n1942) );
  NAND3XLTS U171 ( .A(n687), .B(n686), .C(n685), .Y(n1941) );
  NAND3XLTS U172 ( .A(n666), .B(n665), .C(n664), .Y(n1940) );
  NAND3XLTS U173 ( .A(n554), .B(n553), .C(n552), .Y(n1931) );
  NAND3XLTS U174 ( .A(n1781), .B(n1780), .C(n1779), .Y(n2101) );
  NAND3XLTS U175 ( .A(n1772), .B(n1771), .C(n1770), .Y(n2100) );
  NAND3XLTS U176 ( .A(n1764), .B(n1763), .C(n1762), .Y(n2099) );
  NAND3XLTS U177 ( .A(n1756), .B(n1755), .C(n1754), .Y(n2098) );
  NAND3XLTS U178 ( .A(n977), .B(n976), .C(n975), .Y(n1973) );
  NAND3XLTS U179 ( .A(n970), .B(n969), .C(n968), .Y(n1972) );
  NAND3XLTS U180 ( .A(n962), .B(n961), .C(n960), .Y(n1971) );
  NAND3XLTS U181 ( .A(n955), .B(n954), .C(n953), .Y(n1970) );
  NAND3XLTS U182 ( .A(n1686), .B(n1685), .C(n1684), .Y(n2065) );
  NAND3XLTS U183 ( .A(n1679), .B(n1678), .C(n1677), .Y(n2064) );
  NAND3XLTS U184 ( .A(n1672), .B(n1671), .C(n1670), .Y(n2063) );
  NAND3XLTS U185 ( .A(n1667), .B(n1666), .C(n1665), .Y(n2062) );
  NAND3XLTS U186 ( .A(n902), .B(n901), .C(n900), .Y(n1961) );
  NAND3XLTS U187 ( .A(n894), .B(n893), .C(n892), .Y(n1960) );
  NAND3XLTS U188 ( .A(n890), .B(n889), .C(n888), .Y(n1959) );
  NAND3XLTS U189 ( .A(n886), .B(n885), .C(n884), .Y(n1958) );
  NAND3XLTS U190 ( .A(n1661), .B(n1660), .C(n1659), .Y(n2053) );
  NAND3XLTS U191 ( .A(n1651), .B(n1650), .C(n1649), .Y(n2052) );
  NAND3XLTS U192 ( .A(n1641), .B(n1640), .C(n1639), .Y(n2051) );
  NAND3XLTS U193 ( .A(n1634), .B(n1633), .C(n1632), .Y(n2050) );
  NAND3XLTS U194 ( .A(n883), .B(n882), .C(n881), .Y(n1957) );
  NAND3XLTS U195 ( .A(n878), .B(n877), .C(n876), .Y(n1956) );
  NAND3XLTS U196 ( .A(n875), .B(n874), .C(n873), .Y(n1955) );
  NAND3XLTS U197 ( .A(n870), .B(n869), .C(n868), .Y(n1954) );
  NAND3XLTS U198 ( .A(n1105), .B(n1104), .C(n1103), .Y(n1997) );
  NAND3XLTS U199 ( .A(n1101), .B(n1100), .C(n1099), .Y(n1996) );
  NAND3XLTS U200 ( .A(n1094), .B(n1093), .C(n1092), .Y(n1995) );
  NAND3XLTS U201 ( .A(n1090), .B(n1089), .C(n1088), .Y(n1994) );
  NAND3XLTS U202 ( .A(n1085), .B(n1084), .C(n1083), .Y(n1993) );
  NAND3XLTS U203 ( .A(n1080), .B(n1079), .C(n1078), .Y(n1992) );
  NAND3XLTS U204 ( .A(n1421), .B(n1420), .C(n1419), .Y(n2015) );
  NAND3XLTS U205 ( .A(n1416), .B(n1415), .C(n1414), .Y(n2014) );
  NAND3XLTS U206 ( .A(n1410), .B(n1409), .C(n1408), .Y(n2013) );
  NAND3XLTS U207 ( .A(n1405), .B(n1404), .C(n1403), .Y(n2012) );
  NAND3XLTS U208 ( .A(n1400), .B(n1399), .C(n1398), .Y(n2011) );
  NAND3XLTS U209 ( .A(n1396), .B(n1395), .C(n1394), .Y(n2010) );
  NAND3XLTS U210 ( .A(n1455), .B(n1454), .C(n1453), .Y(n2021) );
  NAND3XLTS U211 ( .A(n1450), .B(n1449), .C(n1448), .Y(n2020) );
  NAND3XLTS U212 ( .A(n1444), .B(n1443), .C(n1442), .Y(n2019) );
  NAND3XLTS U213 ( .A(n1439), .B(n1438), .C(n1437), .Y(n2018) );
  NAND3XLTS U214 ( .A(n1433), .B(n1432), .C(n1431), .Y(n2017) );
  NAND3XLTS U215 ( .A(n1429), .B(n1428), .C(n1427), .Y(n2016) );
  NAND3XLTS U216 ( .A(n1884), .B(n1883), .C(n1882), .Y(n2137) );
  NAND3XLTS U217 ( .A(n1873), .B(n1872), .C(n1871), .Y(n2136) );
  NAND3XLTS U218 ( .A(n1863), .B(n1862), .C(n1861), .Y(n2135) );
  NAND3XLTS U219 ( .A(n1855), .B(n1854), .C(n1853), .Y(n2134) );
  NAND3XLTS U220 ( .A(n1049), .B(n1048), .C(n1047), .Y(n1985) );
  NAND3XLTS U221 ( .A(n1040), .B(n1039), .C(n1038), .Y(n1984) );
  NAND3XLTS U222 ( .A(n1035), .B(n1034), .C(n1033), .Y(n1983) );
  NAND3XLTS U223 ( .A(n1030), .B(n1029), .C(n1028), .Y(n1982) );
  NAND3XLTS U224 ( .A(n1845), .B(n1844), .C(n1843), .Y(n2125) );
  NAND3XLTS U225 ( .A(n1834), .B(n1833), .C(n1832), .Y(n2124) );
  NAND3XLTS U226 ( .A(n1824), .B(n1823), .C(n1822), .Y(n2123) );
  NAND3XLTS U227 ( .A(n1815), .B(n1814), .C(n1813), .Y(n2122) );
  NAND3XLTS U228 ( .A(n1025), .B(n1024), .C(n1023), .Y(n1981) );
  NAND3XLTS U229 ( .A(n1016), .B(n1015), .C(n1014), .Y(n1980) );
  NAND3XLTS U230 ( .A(n1010), .B(n1009), .C(n1008), .Y(n1979) );
  NAND3XLTS U231 ( .A(n1003), .B(n1002), .C(n1001), .Y(n1978) );
  NAND3XLTS U232 ( .A(n1748), .B(n1747), .C(n1746), .Y(n2089) );
  NAND3XLTS U233 ( .A(n1739), .B(n1738), .C(n1737), .Y(n2088) );
  NAND3XLTS U234 ( .A(n1732), .B(n1731), .C(n1730), .Y(n2087) );
  NAND3XLTS U235 ( .A(n1724), .B(n1723), .C(n1722), .Y(n2086) );
  NAND3XLTS U236 ( .A(n948), .B(n947), .C(n946), .Y(n1969) );
  NAND3XLTS U237 ( .A(n940), .B(n939), .C(n938), .Y(n1968) );
  NAND3XLTS U238 ( .A(n935), .B(n934), .C(n933), .Y(n1967) );
  NAND3XLTS U239 ( .A(n927), .B(n926), .C(n925), .Y(n1966) );
  NAND3XLTS U240 ( .A(n1719), .B(n1718), .C(n1717), .Y(n2077) );
  NAND3XLTS U241 ( .A(n1710), .B(n1709), .C(n1708), .Y(n2076) );
  NAND3XLTS U242 ( .A(n1703), .B(n1702), .C(n1701), .Y(n2075) );
  NAND3XLTS U243 ( .A(n1695), .B(n1694), .C(n1693), .Y(n2074) );
  NAND3XLTS U244 ( .A(n920), .B(n919), .C(n918), .Y(n1965) );
  NAND3XLTS U245 ( .A(n914), .B(n913), .C(n912), .Y(n1964) );
  NAND3XLTS U246 ( .A(n910), .B(n909), .C(n908), .Y(n1963) );
  NAND3XLTS U247 ( .A(n906), .B(n905), .C(n904), .Y(n1962) );
  NAND3XLTS U248 ( .A(n1363), .B(n1362), .C(n1361), .Y(n2003) );
  NAND3XLTS U249 ( .A(n1358), .B(n1357), .C(n1356), .Y(n2002) );
  NAND3XLTS U250 ( .A(n1351), .B(n1350), .C(n1349), .Y(n2001) );
  NAND3XLTS U251 ( .A(n1346), .B(n1345), .C(n1344), .Y(n2000) );
  NAND3XLTS U252 ( .A(n1340), .B(n1339), .C(n1338), .Y(n1999) );
  NAND3XLTS U253 ( .A(n1111), .B(n1110), .C(n1109), .Y(n1998) );
  NAND3XLTS U254 ( .A(n1389), .B(n1388), .C(n1387), .Y(n2009) );
  NAND3XLTS U255 ( .A(n1384), .B(n1383), .C(n1382), .Y(n2008) );
  NAND3XLTS U256 ( .A(n1380), .B(n1379), .C(n1378), .Y(n2007) );
  NAND3XLTS U257 ( .A(n1376), .B(n1375), .C(n1374), .Y(n2006) );
  NAND3XLTS U258 ( .A(n1372), .B(n1371), .C(n1370), .Y(n2005) );
  NAND3XLTS U259 ( .A(n1368), .B(n1367), .C(n1366), .Y(n2004) );
  NAND3XLTS U260 ( .A(n1494), .B(n1493), .C(n1492), .Y(n2027) );
  NAND3XLTS U261 ( .A(n1488), .B(n1487), .C(n1486), .Y(n2026) );
  NAND3XLTS U262 ( .A(n1481), .B(n1480), .C(n1479), .Y(n2025) );
  NAND3XLTS U263 ( .A(n1475), .B(n1474), .C(n1473), .Y(n2024) );
  NAND3XLTS U264 ( .A(n1469), .B(n1468), .C(n1467), .Y(n2023) );
  NAND3XLTS U265 ( .A(n1464), .B(n1463), .C(n1462), .Y(n2022) );
  NAND3XLTS U266 ( .A(n1541), .B(n1540), .C(n1539), .Y(n2033) );
  NAND3XLTS U267 ( .A(n1533), .B(n1532), .C(n1531), .Y(n2032) );
  NAND3XLTS U268 ( .A(n1524), .B(n1523), .C(n1522), .Y(n2031) );
  NAND3XLTS U269 ( .A(n1517), .B(n1516), .C(n1515), .Y(n2030) );
  NAND3XLTS U270 ( .A(n1510), .B(n1509), .C(n1508), .Y(n2029) );
  NAND3XLTS U271 ( .A(n1502), .B(n1501), .C(n1500), .Y(n2028) );
  NAND3XLTS U272 ( .A(n1805), .B(n1804), .C(n1803), .Y(n2113) );
  NAND3XLTS U273 ( .A(n1799), .B(n1798), .C(n1797), .Y(n2112) );
  NAND3XLTS U274 ( .A(n1793), .B(n1792), .C(n1791), .Y(n2111) );
  NAND3XLTS U275 ( .A(n1788), .B(n1787), .C(n1786), .Y(n2110) );
  NAND3XLTS U276 ( .A(n995), .B(n994), .C(n993), .Y(n1977) );
  NAND3XLTS U277 ( .A(n988), .B(n987), .C(n986), .Y(n1976) );
  NAND3XLTS U278 ( .A(n985), .B(n984), .C(n983), .Y(n1975) );
  NAND3XLTS U279 ( .A(n981), .B(n980), .C(n979), .Y(n1974) );
  NAND3XLTS U280 ( .A(n1075), .B(n1074), .C(n1073), .Y(n1991) );
  NAND3XLTS U281 ( .A(n1071), .B(n1070), .C(n1069), .Y(n1990) );
  NAND3XLTS U282 ( .A(n1065), .B(n1064), .C(n1063), .Y(n1989) );
  NAND3XLTS U283 ( .A(n1061), .B(n1060), .C(n1059), .Y(n1988) );
  NAND3XLTS U284 ( .A(n1057), .B(n1056), .C(n1055), .Y(n1987) );
  NAND3XLTS U285 ( .A(n1054), .B(n1053), .C(n1052), .Y(n1986) );
  AOI211XLTS U286 ( .A0(n489), .A1(n525), .B0(n488), .C0(n487), .Y(n490) );
  XOR2XLTS U287 ( .A(n524), .B(n492), .Y(n488) );
  OR2X1TS U288 ( .A(n272), .B(n1720), .Y(n1390) );
  OR2X1TS U289 ( .A(n393), .B(n1846), .Y(n1031) );
  OR2X1TS U290 ( .A(n178), .B(n1782), .Y(n982) );
  OR2X1TS U291 ( .A(n127), .B(n1749), .Y(n1364) );
  OR2X1TS U292 ( .A(n79), .B(n1662), .Y(n1456) );
  OR2X1TS U293 ( .A(n28), .B(n1654), .Y(n1495) );
  NOR2XLTS U294 ( .A(n24), .B(n1572), .Y(n215) );
  OR2X1TS U295 ( .A(n1620), .B(n397), .Y(n2) );
  OR2X1TS U296 ( .A(n1594), .B(n184), .Y(n3) );
  OR2X1TS U297 ( .A(n1607), .B(n326), .Y(n4) );
  OR2X1TS U298 ( .A(n1621), .B(n397), .Y(n5) );
  OR2X1TS U299 ( .A(n1553), .B(n83), .Y(n6) );
  OA21XLTS U300 ( .A0(n315), .A1(n455), .B0(n20), .Y(n7) );
  CLKBUFX2TS U301 ( .A(n182), .Y(n183) );
  CLKBUFX2TS U302 ( .A(n324), .Y(n325) );
  NOR3XLTS U303 ( .A(n1559), .B(n1554), .C(n81), .Y(n77) );
  NOR3XLTS U304 ( .A(n1582), .B(n1576), .C(n274), .Y(n270) );
  OR2X1TS U305 ( .A(n392), .B(n1629), .Y(n9) );
  AND3X1TS U306 ( .A(n538), .B(n1902), .C(n537), .Y(n10) );
  INVX2TS U307 ( .A(destinationAddressIn_EAST[7]), .Y(n63) );
  INVX2TS U308 ( .A(destinationAddressIn_EAST[6]), .Y(n66) );
  INVX2TS U309 ( .A(destinationAddressIn_EAST[5]), .Y(n57) );
  INVX2TS U310 ( .A(destinationAddressIn_EAST[4]), .Y(n53) );
  INVX2TS U311 ( .A(destinationAddressIn_EAST[9]), .Y(n34) );
  INVX2TS U312 ( .A(destinationAddressIn_EAST[11]), .Y(n39) );
  INVX2TS U313 ( .A(destinationAddressIn_EAST[8]), .Y(n43) );
  INVX2TS U314 ( .A(destinationAddressIn_EAST[10]), .Y(n27) );
  INVX2TS U315 ( .A(writeIn_EAST), .Y(n47) );
  CLKBUFX2TS U316 ( .A(n1906), .Y(n11) );
  INVX2TS U332 ( .A(n1912), .Y(n484) );
  INVX2TS U333 ( .A(n1909), .Y(n447) );
  INVX2TS U334 ( .A(n13), .Y(n71) );
  INVX2TS U335 ( .A(n71), .Y(n116) );
  INVX2TS U336 ( .A(selectBit_WEST), .Y(n453) );
  INVX2TS U337 ( .A(n1547), .Y(n1549) );
  INVX2TS U338 ( .A(n1905), .Y(n457) );
  INVX2TS U339 ( .A(n17), .Y(n315) );
  INVX2TS U340 ( .A(selectBit_SOUTH), .Y(n506) );
  INVX2TS U341 ( .A(n8), .Y(n213) );
  INVX2TS U342 ( .A(n1912), .Y(n455) );
  NAND2X1TS U343 ( .A(n16), .B(n455), .Y(n20) );
  NAND2X1TS U344 ( .A(selectBit_SOUTH), .B(n19), .Y(n18) );
  NAND2X1TS U345 ( .A(n311), .B(n263), .Y(n119) );
  INVX2TS U346 ( .A(n1911), .Y(n269) );
  INVX2TS U347 ( .A(n1910), .Y(n450) );
  AOI22X1TS U348 ( .A0(n269), .A1(n20), .B0(n120), .B1(n450), .Y(n75) );
  NAND2X1TS U349 ( .A(n22), .B(n75), .Y(n21) );
  INVX2TS U350 ( .A(n21), .Y(n115) );
  OAI21XLTS U351 ( .A0(n22), .A1(n75), .B0(n21), .Y(n118) );
  NAND2X1TS U352 ( .A(selectBit_EAST), .B(n118), .Y(n264) );
  NAND2X1TS U353 ( .A(n269), .B(n120), .Y(n25) );
  INVX2TS U354 ( .A(n1912), .Y(n445) );
  CLKBUFX2TS U355 ( .A(n75), .Y(n266) );
  INVX2TS U356 ( .A(n266), .Y(n23) );
  INVX2TS U357 ( .A(n506), .Y(n505) );
  INVX2TS U358 ( .A(n453), .Y(n512) );
  INVX2TS U359 ( .A(readReady), .Y(n122) );
  INVX2TS U360 ( .A(n122), .Y(n511) );
  NAND2X1TS U361 ( .A(n538), .B(n507), .Y(n523) );
  NAND2X1TS U362 ( .A(n523), .B(n1914), .Y(n24) );
  INVX2TS U363 ( .A(n24), .Y(n125) );
  INVX2TS U364 ( .A(n125), .Y(n316) );
  INVX2TS U365 ( .A(n1909), .Y(n482) );
  INVX2TS U366 ( .A(n122), .Y(n514) );
  NAND2X1TS U367 ( .A(n28), .B(n1550), .Y(n30) );
  INVX2TS U368 ( .A(n26), .Y(n880) );
  INVX2TS U369 ( .A(n880), .Y(n1645) );
  CLKBUFX2TS U370 ( .A(n1645), .Y(n38) );
  INVX2TS U371 ( .A(n38), .Y(n62) );
  INVX2TS U372 ( .A(destinationAddressIn_EAST[10]), .Y(n223) );
  INVX2TS U373 ( .A(n125), .Y(n387) );
  INVX2TS U374 ( .A(n387), .Y(n267) );
  OR2X1TS U375 ( .A(n1550), .B(n316), .Y(n1503) );
  INVX2TS U376 ( .A(n1503), .Y(n1654) );
  INVX2TS U377 ( .A(n1495), .Y(n44) );
  OR2X1TS U378 ( .A(n1547), .B(n30), .Y(n48) );
  INVX2TS U379 ( .A(n48), .Y(n1646) );
  CLKBUFX2TS U380 ( .A(destinationAddressIn_WEST[10]), .Y(n412) );
  CLKBUFX2TS U381 ( .A(n412), .Y(n745) );
  AOI22X1TS U382 ( .A0(n44), .A1(\destinationAddressbuffer[7][10] ), .B0(n1646), .B1(n745), .Y(n33) );
  OR2X1TS U383 ( .A(n1542), .B(n31), .Y(n54) );
  INVX2TS U384 ( .A(n54), .Y(n872) );
  INVX2TS U385 ( .A(n162), .Y(n748) );
  INVX2TS U386 ( .A(n40), .Y(n59) );
  INVX2TS U387 ( .A(n59), .Y(n1647) );
  CLKBUFX2TS U388 ( .A(destinationAddressIn_NORTH[10]), .Y(n749) );
  CLKBUFX2TS U389 ( .A(n749), .Y(n339) );
  AOI22X1TS U390 ( .A0(n872), .A1(n748), .B0(n1647), .B1(n339), .Y(n32) );
  OAI211XLTS U391 ( .A0(n62), .A1(n223), .B0(n33), .C0(n32), .Y(n2060) );
  INVX2TS U392 ( .A(destinationAddressIn_EAST[9]), .Y(n226) );
  INVX2TS U393 ( .A(n48), .Y(n1527) );
  CLKBUFX2TS U394 ( .A(destinationAddressIn_WEST[9]), .Y(n394) );
  CLKBUFX2TS U395 ( .A(n394), .Y(n728) );
  AOI22X1TS U396 ( .A0(n44), .A1(\destinationAddressbuffer[7][9] ), .B0(n49), 
        .B1(n728), .Y(n37) );
  INVX2TS U397 ( .A(n54), .Y(n1530) );
  INVX2TS U398 ( .A(n1530), .Y(n1505) );
  INVX2TS U399 ( .A(n1505), .Y(n1638) );
  INVX2TS U400 ( .A(n168), .Y(n729) );
  INVX2TS U401 ( .A(n59), .Y(n35) );
  CLKBUFX2TS U402 ( .A(destinationAddressIn_NORTH[9]), .Y(n731) );
  CLKBUFX2TS U403 ( .A(n731), .Y(n333) );
  AOI22X1TS U404 ( .A0(n1638), .A1(n729), .B0(n871), .B1(n333), .Y(n36) );
  OAI211XLTS U405 ( .A0(n62), .A1(n226), .B0(n37), .C0(n36), .Y(n2059) );
  INVX2TS U406 ( .A(n38), .Y(n70) );
  INVX2TS U407 ( .A(destinationAddressIn_EAST[11]), .Y(n238) );
  CLKBUFX2TS U408 ( .A(destinationAddressIn_WEST[11]), .Y(n401) );
  CLKBUFX2TS U409 ( .A(n401), .Y(n761) );
  AOI22X1TS U410 ( .A0(n44), .A1(\destinationAddressbuffer[7][11] ), .B0(n58), 
        .B1(n761), .Y(n42) );
  INVX2TS U411 ( .A(n154), .Y(n764) );
  INVX2TS U412 ( .A(n40), .Y(n1497) );
  INVX2TS U413 ( .A(n1497), .Y(n871) );
  CLKBUFX2TS U414 ( .A(destinationAddressIn_NORTH[11]), .Y(n765) );
  CLKBUFX2TS U415 ( .A(n765), .Y(n348) );
  AOI22X1TS U416 ( .A0(n1530), .A1(n764), .B0(n871), .B1(n348), .Y(n41) );
  OAI211XLTS U417 ( .A0(n70), .A1(n238), .B0(n42), .C0(n41), .Y(n2061) );
  INVX2TS U418 ( .A(destinationAddressIn_EAST[8]), .Y(n232) );
  INVX2TS U419 ( .A(n48), .Y(n1656) );
  CLKBUFX2TS U420 ( .A(destinationAddressIn_WEST[8]), .Y(n407) );
  CLKBUFX2TS U421 ( .A(n407), .Y(n713) );
  AOI22X1TS U422 ( .A0(n44), .A1(\destinationAddressbuffer[7][8] ), .B0(n1656), 
        .B1(n713), .Y(n46) );
  INVX2TS U423 ( .A(n158), .Y(n714) );
  CLKBUFX2TS U424 ( .A(destinationAddressIn_NORTH[8]), .Y(n715) );
  CLKBUFX2TS U425 ( .A(n715), .Y(n328) );
  AOI22X1TS U426 ( .A0(n872), .A1(n714), .B0(n871), .B1(n328), .Y(n45) );
  OAI211XLTS U427 ( .A0(n62), .A1(n232), .B0(n46), .C0(n45), .Y(n2058) );
  INVX2TS U428 ( .A(writeIn_EAST), .Y(n243) );
  CLKBUFX2TS U429 ( .A(n1495), .Y(n879) );
  INVX2TS U430 ( .A(n879), .Y(n1652) );
  INVX2TS U431 ( .A(n48), .Y(n49) );
  INVX2TS U432 ( .A(n49), .Y(n867) );
  INVX2TS U433 ( .A(n867), .Y(n58) );
  CLKBUFX2TS U434 ( .A(writeIn_WEST), .Y(n420) );
  CLKBUFX2TS U435 ( .A(n420), .Y(n542) );
  AOI22X1TS U436 ( .A0(n1652), .A1(writeOutbuffer[7]), .B0(n58), .B1(n542), 
        .Y(n52) );
  INVX2TS U437 ( .A(n54), .Y(n50) );
  INVX2TS U438 ( .A(writeIn_SOUTH), .Y(n172) );
  INVX2TS U439 ( .A(n172), .Y(n544) );
  INVX2TS U440 ( .A(n59), .Y(n1657) );
  CLKBUFX2TS U441 ( .A(writeIn_NORTH), .Y(n545) );
  CLKBUFX2TS U442 ( .A(n545), .Y(n354) );
  AOI22X1TS U443 ( .A0(n50), .A1(n544), .B0(n1657), .B1(n354), .Y(n51) );
  OAI211XLTS U444 ( .A0(n70), .A1(n243), .B0(n52), .C0(n51), .Y(n2034) );
  INVX2TS U445 ( .A(destinationAddressIn_EAST[4]), .Y(n260) );
  INVX2TS U446 ( .A(n879), .Y(n67) );
  AOI22X1TS U447 ( .A0(n67), .A1(\destinationAddressbuffer[7][4] ), .B0(n1646), 
        .B1(destinationAddressIn_WEST[4]), .Y(n56) );
  INVX2TS U448 ( .A(n54), .Y(n1658) );
  INVX2TS U449 ( .A(destinationAddressIn_SOUTH[4]), .Y(n150) );
  INVX2TS U450 ( .A(n150), .Y(n658) );
  AOI22X1TS U451 ( .A0(n1658), .A1(n658), .B0(n1657), .B1(
        destinationAddressIn_NORTH[4]), .Y(n55) );
  OAI211XLTS U452 ( .A0(n70), .A1(n260), .B0(n56), .C0(n55), .Y(n2054) );
  INVX2TS U453 ( .A(destinationAddressIn_EAST[5]), .Y(n247) );
  AOI22X1TS U454 ( .A0(n67), .A1(\destinationAddressbuffer[7][5] ), .B0(n58), 
        .B1(destinationAddressIn_WEST[5]), .Y(n61) );
  INVX2TS U455 ( .A(destinationAddressIn_SOUTH[5]), .Y(n144) );
  INVX2TS U456 ( .A(n144), .Y(n670) );
  INVX2TS U457 ( .A(n59), .Y(n1537) );
  AOI22X1TS U458 ( .A0(n50), .A1(n670), .B0(n1537), .B1(
        destinationAddressIn_NORTH[5]), .Y(n60) );
  OAI211XLTS U459 ( .A0(n62), .A1(n247), .B0(n61), .C0(n60), .Y(n2055) );
  INVX2TS U460 ( .A(destinationAddressIn_EAST[7]), .Y(n256) );
  AOI22X1TS U461 ( .A0(n67), .A1(\destinationAddressbuffer[7][7] ), .B0(n1656), 
        .B1(destinationAddressIn_WEST[7]), .Y(n65) );
  INVX2TS U462 ( .A(destinationAddressIn_SOUTH[7]), .Y(n138) );
  INVX2TS U463 ( .A(n138), .Y(n703) );
  AOI22X1TS U464 ( .A0(n1658), .A1(n703), .B0(n1647), .B1(
        destinationAddressIn_NORTH[7]), .Y(n64) );
  OAI211XLTS U465 ( .A0(n880), .A1(n256), .B0(n65), .C0(n64), .Y(n2057) );
  INVX2TS U466 ( .A(destinationAddressIn_EAST[6]), .Y(n251) );
  AOI22X1TS U467 ( .A0(n67), .A1(\destinationAddressbuffer[7][6] ), .B0(n1527), 
        .B1(destinationAddressIn_WEST[6]), .Y(n69) );
  INVX2TS U468 ( .A(destinationAddressIn_SOUTH[6]), .Y(n134) );
  INVX2TS U469 ( .A(n134), .Y(n690) );
  AOI22X1TS U470 ( .A0(n1638), .A1(n690), .B0(n1637), .B1(
        destinationAddressIn_NORTH[6]), .Y(n68) );
  OAI211XLTS U471 ( .A0(n70), .A1(n251), .B0(n69), .C0(n68), .Y(n2056) );
  INVX2TS U472 ( .A(n72), .Y(n174) );
  NAND2X1TS U473 ( .A(n117), .B(n459), .Y(n262) );
  AOI21X1TS U474 ( .A0(n213), .A1(n73), .B0(n311), .Y(n384) );
  NOR3XLTS U475 ( .A(n384), .B(n264), .C(n263), .Y(n1556) );
  NOR2XLTS U476 ( .A(n447), .B(n504), .Y(n386) );
  INVX2TS U477 ( .A(n7), .Y(n265) );
  AOI31XLTS U478 ( .A0(n451), .A1(n445), .A2(n386), .B0(n1553), .Y(n76) );
  INVX2TS U479 ( .A(n125), .Y(n392) );
  AOI21X1TS U480 ( .A0(n80), .A1(n76), .B0(n392), .Y(n79) );
  INVX2TS U481 ( .A(n122), .Y(n509) );
  INVX2TS U482 ( .A(n1905), .Y(n390) );
  NAND2X1TS U483 ( .A(n79), .B(n1560), .Y(n81) );
  INVX2TS U484 ( .A(n77), .Y(n1470) );
  INVX2TS U485 ( .A(n1470), .Y(n898) );
  CLKBUFX2TS U486 ( .A(n898), .Y(n90) );
  INVX2TS U487 ( .A(n90), .Y(n107) );
  INVX2TS U488 ( .A(n78), .Y(n895) );
  INVX2TS U489 ( .A(n895), .Y(n1662) );
  CLKBUFX2TS U490 ( .A(n1456), .Y(n896) );
  INVX2TS U491 ( .A(n896), .Y(n94) );
  OR2X1TS U492 ( .A(n1557), .B(n81), .Y(n98) );
  INVX2TS U493 ( .A(n98), .Y(n1663) );
  AOI22X1TS U494 ( .A0(n94), .A1(\destinationAddressbuffer[6][10] ), .B0(n1663), .B1(n745), .Y(n86) );
  INVX2TS U495 ( .A(n6), .Y(n82) );
  INVX2TS U496 ( .A(n82), .Y(n887) );
  INVX2TS U497 ( .A(n887), .Y(n87) );
  CLKBUFX2TS U498 ( .A(n749), .Y(n414) );
  INVX2TS U499 ( .A(n84), .Y(n95) );
  INVX2TS U500 ( .A(n162), .Y(n338) );
  AOI22X1TS U501 ( .A0(n87), .A1(n414), .B0(n104), .B1(n338), .Y(n85) );
  OAI211XLTS U502 ( .A0(n107), .A1(n223), .B0(n86), .C0(n85), .Y(n2072) );
  INVX2TS U503 ( .A(n98), .Y(n1681) );
  AOI22X1TS U504 ( .A0(n94), .A1(\destinationAddressbuffer[6][11] ), .B0(n108), 
        .B1(n761), .Y(n89) );
  CLKBUFX2TS U505 ( .A(n765), .Y(n403) );
  INVX2TS U506 ( .A(n154), .Y(n347) );
  AOI22X1TS U507 ( .A0(n87), .A1(n403), .B0(n84), .B1(n347), .Y(n88) );
  OAI211XLTS U508 ( .A0(n107), .A1(n238), .B0(n89), .C0(n88), .Y(n2073) );
  INVX2TS U509 ( .A(n90), .Y(n114) );
  AOI22X1TS U510 ( .A0(n94), .A1(\destinationAddressbuffer[6][9] ), .B0(n99), 
        .B1(n728), .Y(n93) );
  INVX2TS U511 ( .A(n887), .Y(n891) );
  CLKBUFX2TS U512 ( .A(n731), .Y(n398) );
  INVX2TS U513 ( .A(n95), .Y(n1460) );
  INVX2TS U514 ( .A(n95), .Y(n91) );
  INVX2TS U515 ( .A(n168), .Y(n332) );
  AOI22X1TS U516 ( .A0(n891), .A1(n398), .B0(n91), .B1(n332), .Y(n92) );
  OAI211XLTS U517 ( .A0(n114), .A1(n226), .B0(n93), .C0(n92), .Y(n2071) );
  INVX2TS U518 ( .A(n98), .Y(n1458) );
  AOI22X1TS U519 ( .A0(n94), .A1(\destinationAddressbuffer[6][8] ), .B0(n1458), 
        .B1(n713), .Y(n97) );
  INVX2TS U520 ( .A(n6), .Y(n1683) );
  CLKBUFX2TS U521 ( .A(n715), .Y(n409) );
  INVX2TS U522 ( .A(n84), .Y(n899) );
  INVX2TS U523 ( .A(n899), .Y(n104) );
  INVX2TS U524 ( .A(n158), .Y(n327) );
  AOI22X1TS U525 ( .A0(n1683), .A1(n409), .B0(n104), .B1(n327), .Y(n96) );
  OAI211XLTS U526 ( .A0(n107), .A1(n232), .B0(n97), .C0(n96), .Y(n2070) );
  INVX2TS U527 ( .A(n896), .Y(n1680) );
  INVX2TS U528 ( .A(n98), .Y(n99) );
  INVX2TS U529 ( .A(n99), .Y(n897) );
  INVX2TS U530 ( .A(n897), .Y(n108) );
  AOI22X1TS U531 ( .A0(n1680), .A1(writeOutbuffer[6]), .B0(n108), .B1(n542), 
        .Y(n101) );
  INVX2TS U532 ( .A(n6), .Y(n1664) );
  CLKBUFX2TS U533 ( .A(n545), .Y(n421) );
  INVX2TS U534 ( .A(n172), .Y(n352) );
  AOI22X1TS U535 ( .A0(n1664), .A1(n421), .B0(n1676), .B1(n352), .Y(n100) );
  OAI211XLTS U536 ( .A0(n114), .A1(n243), .B0(n101), .C0(n100), .Y(n2035) );
  INVX2TS U537 ( .A(n1456), .Y(n111) );
  AOI22X1TS U538 ( .A0(n111), .A1(\destinationAddressbuffer[6][4] ), .B0(n1663), .B1(destinationAddressIn_WEST[4]), .Y(n103) );
  CLKBUFX2TS U539 ( .A(destinationAddressIn_NORTH[4]), .Y(n360) );
  CLKBUFX2TS U540 ( .A(n360), .Y(n438) );
  INVX2TS U541 ( .A(n150), .Y(n359) );
  AOI22X1TS U542 ( .A0(n1683), .A1(n438), .B0(n84), .B1(n359), .Y(n102) );
  OAI211XLTS U543 ( .A0(n114), .A1(n260), .B0(n103), .C0(n102), .Y(n2066) );
  AOI22X1TS U544 ( .A0(n111), .A1(\destinationAddressbuffer[6][6] ), .B0(n1681), .B1(destinationAddressIn_WEST[6]), .Y(n106) );
  CLKBUFX2TS U545 ( .A(destinationAddressIn_NORTH[6]), .Y(n365) );
  CLKBUFX2TS U546 ( .A(n365), .Y(n427) );
  INVX2TS U547 ( .A(n134), .Y(n364) );
  AOI22X1TS U548 ( .A0(n891), .A1(n427), .B0(n104), .B1(n364), .Y(n105) );
  OAI211XLTS U549 ( .A0(n107), .A1(n251), .B0(n106), .C0(n105), .Y(n2068) );
  AOI22X1TS U550 ( .A0(n111), .A1(\destinationAddressbuffer[6][5] ), .B0(n108), 
        .B1(destinationAddressIn_WEST[5]), .Y(n110) );
  INVX2TS U551 ( .A(n6), .Y(n1461) );
  CLKBUFX2TS U552 ( .A(destinationAddressIn_NORTH[5]), .Y(n371) );
  CLKBUFX2TS U553 ( .A(n371), .Y(n433) );
  INVX2TS U554 ( .A(n95), .Y(n1682) );
  INVX2TS U555 ( .A(n144), .Y(n370) );
  AOI22X1TS U556 ( .A0(n1461), .A1(n433), .B0(n1682), .B1(n370), .Y(n109) );
  OAI211XLTS U557 ( .A0(n1470), .A1(n247), .B0(n110), .C0(n109), .Y(n2067) );
  AOI22X1TS U558 ( .A0(n111), .A1(\destinationAddressbuffer[6][7] ), .B0(n1458), .B1(destinationAddressIn_WEST[7]), .Y(n113) );
  CLKBUFX2TS U559 ( .A(destinationAddressIn_NORTH[7]), .Y(n377) );
  CLKBUFX2TS U560 ( .A(n377), .Y(n424) );
  INVX2TS U561 ( .A(n138), .Y(n376) );
  AOI22X1TS U562 ( .A0(n1461), .A1(n424), .B0(n1460), .B1(n376), .Y(n112) );
  OAI211XLTS U563 ( .A0(n114), .A1(n256), .B0(n113), .C0(n112), .Y(n2069) );
  INVX2TS U564 ( .A(n115), .Y(n1585) );
  INVX2TS U565 ( .A(n510), .Y(n513) );
  INVX2TS U566 ( .A(n1910), .Y(n444) );
  NAND2X1TS U567 ( .A(n120), .B(n444), .Y(n121) );
  INVX2TS U568 ( .A(n1912), .Y(n494) );
  INVX2TS U569 ( .A(n124), .Y(n965) );
  INVX2TS U570 ( .A(n965), .Y(n1760) );
  CLKBUFX2TS U571 ( .A(n1760), .Y(n139) );
  INVX2TS U572 ( .A(n139), .Y(n163) );
  INVX2TS U573 ( .A(n125), .Y(n441) );
  INVX2TS U574 ( .A(n126), .Y(n972) );
  INVX2TS U575 ( .A(n972), .Y(n1749) );
  CLKBUFX2TS U576 ( .A(n1364), .Y(n169) );
  INVX2TS U577 ( .A(n169), .Y(n146) );
  INVX2TS U578 ( .A(n135), .Y(n957) );
  INVX2TS U579 ( .A(n957), .Y(n164) );
  AOI22X1TS U580 ( .A0(n146), .A1(\destinationAddressbuffer[3][6] ), .B0(n164), 
        .B1(destinationAddressIn_EAST[6]), .Y(n133) );
  INVX2TS U581 ( .A(n140), .Y(n159) );
  INVX2TS U582 ( .A(n159), .Y(n129) );
  INVX2TS U583 ( .A(n131), .Y(n147) );
  INVX2TS U584 ( .A(n147), .Y(n1752) );
  CLKBUFX2TS U585 ( .A(destinationAddressIn_WEST[6]), .Y(n688) );
  CLKBUFX2TS U586 ( .A(n688), .Y(n363) );
  AOI22X1TS U587 ( .A0(n129), .A1(n365), .B0(n1752), .B1(n363), .Y(n132) );
  OAI211XLTS U588 ( .A0(n163), .A1(n134), .B0(n133), .C0(n132), .Y(n2104) );
  INVX2TS U589 ( .A(n135), .Y(n155) );
  INVX2TS U590 ( .A(n155), .Y(n1774) );
  AOI22X1TS U591 ( .A0(n146), .A1(\destinationAddressbuffer[3][7] ), .B0(n1774), .B1(destinationAddressIn_EAST[7]), .Y(n137) );
  INVX2TS U592 ( .A(n147), .Y(n1776) );
  CLKBUFX2TS U593 ( .A(destinationAddressIn_WEST[7]), .Y(n702) );
  CLKBUFX2TS U594 ( .A(n702), .Y(n374) );
  AOI22X1TS U595 ( .A0(n129), .A1(n377), .B0(n1776), .B1(n374), .Y(n136) );
  OAI211XLTS U596 ( .A0(n163), .A1(n138), .B0(n137), .C0(n136), .Y(n2105) );
  INVX2TS U597 ( .A(n139), .Y(n173) );
  INVX2TS U598 ( .A(n155), .Y(n1767) );
  AOI22X1TS U599 ( .A0(n146), .A1(\destinationAddressbuffer[3][5] ), .B0(n1767), .B1(destinationAddressIn_EAST[5]), .Y(n143) );
  INVX2TS U600 ( .A(n140), .Y(n1369) );
  INVX2TS U601 ( .A(n1369), .Y(n966) );
  INVX2TS U602 ( .A(n147), .Y(n141) );
  INVX2TS U603 ( .A(n141), .Y(n950) );
  INVX2TS U604 ( .A(n950), .Y(n151) );
  CLKBUFX2TS U605 ( .A(destinationAddressIn_WEST[5]), .Y(n668) );
  CLKBUFX2TS U606 ( .A(n668), .Y(n369) );
  AOI22X1TS U607 ( .A0(n966), .A1(n371), .B0(n151), .B1(n369), .Y(n142) );
  OAI211XLTS U608 ( .A0(n173), .A1(n144), .B0(n143), .C0(n142), .Y(n2103) );
  INVX2TS U609 ( .A(n155), .Y(n145) );
  AOI22X1TS U610 ( .A0(n146), .A1(\destinationAddressbuffer[3][4] ), .B0(n164), 
        .B1(destinationAddressIn_EAST[4]), .Y(n149) );
  INVX2TS U611 ( .A(n159), .Y(n1778) );
  INVX2TS U612 ( .A(n147), .Y(n1386) );
  CLKBUFX2TS U613 ( .A(destinationAddressIn_WEST[4]), .Y(n656) );
  CLKBUFX2TS U614 ( .A(n656), .Y(n357) );
  AOI22X1TS U615 ( .A0(n1778), .A1(n360), .B0(n1386), .B1(n357), .Y(n148) );
  OAI211XLTS U616 ( .A0(n163), .A1(n150), .B0(n149), .C0(n148), .Y(n2102) );
  INVX2TS U617 ( .A(n169), .Y(n165) );
  AOI22X1TS U618 ( .A0(n165), .A1(\destinationAddressbuffer[3][11] ), .B0(
        n1767), .B1(destinationAddressIn_EAST[11]), .Y(n153) );
  CLKBUFX2TS U619 ( .A(n401), .Y(n343) );
  AOI22X1TS U620 ( .A0(n1778), .A1(n348), .B0(n151), .B1(n343), .Y(n152) );
  OAI211XLTS U621 ( .A0(n173), .A1(n154), .B0(n153), .C0(n152), .Y(n2109) );
  INVX2TS U622 ( .A(n155), .Y(n1381) );
  AOI22X1TS U623 ( .A0(n165), .A1(\destinationAddressbuffer[3][8] ), .B0(n1381), .B1(destinationAddressIn_EAST[8]), .Y(n157) );
  INVX2TS U624 ( .A(n159), .Y(n1753) );
  CLKBUFX2TS U625 ( .A(n407), .Y(n321) );
  AOI22X1TS U626 ( .A0(n1753), .A1(n328), .B0(n1752), .B1(n321), .Y(n156) );
  OAI211XLTS U627 ( .A0(n173), .A1(n158), .B0(n157), .C0(n156), .Y(n2106) );
  AOI22X1TS U628 ( .A0(n165), .A1(\destinationAddressbuffer[3][10] ), .B0(
        n1381), .B1(destinationAddressIn_EAST[10]), .Y(n161) );
  INVX2TS U629 ( .A(n159), .Y(n1365) );
  CLKBUFX2TS U630 ( .A(n412), .Y(n337) );
  AOI22X1TS U631 ( .A0(n1365), .A1(n339), .B0(n1386), .B1(n337), .Y(n160) );
  OAI211XLTS U632 ( .A0(n163), .A1(n162), .B0(n161), .C0(n160), .Y(n2108) );
  AOI22X1TS U633 ( .A0(n165), .A1(\destinationAddressbuffer[3][9] ), .B0(n164), 
        .B1(destinationAddressIn_EAST[9]), .Y(n167) );
  CLKBUFX2TS U634 ( .A(n394), .Y(n331) );
  AOI22X1TS U635 ( .A0(n966), .A1(n333), .B0(n131), .B1(n331), .Y(n166) );
  OAI211XLTS U636 ( .A0(n965), .A1(n168), .B0(n167), .C0(n166), .Y(n2107) );
  INVX2TS U637 ( .A(n169), .Y(n1773) );
  AOI22X1TS U638 ( .A0(n1773), .A1(writeOutbuffer[3]), .B0(n1774), .B1(
        writeIn_EAST), .Y(n171) );
  CLKBUFX2TS U639 ( .A(n420), .Y(n351) );
  AOI22X1TS U640 ( .A0(n1365), .A1(n354), .B0(n1776), .B1(n351), .Y(n170) );
  OAI211XLTS U641 ( .A0(n173), .A1(n172), .B0(n171), .C0(n170), .Y(n2038) );
  INVX2TS U642 ( .A(n263), .Y(n312) );
  INVX2TS U643 ( .A(n312), .Y(n382) );
  NOR3XLTS U644 ( .A(n384), .B(n382), .C(n383), .Y(n1600) );
  INVX2TS U645 ( .A(n266), .Y(n313) );
  AOI31XLTS U646 ( .A0(n494), .A1(n386), .A2(n450), .B0(n1596), .Y(n175) );
  AOI21X1TS U647 ( .A0(n180), .A1(n175), .B0(n441), .Y(n178) );
  INVX2TS U648 ( .A(n1910), .Y(n442) );
  NAND2X1TS U649 ( .A(n178), .B(n1604), .Y(n181) );
  INVX2TS U650 ( .A(n176), .Y(n1341) );
  INVX2TS U651 ( .A(n1341), .Y(n991) );
  CLKBUFX2TS U652 ( .A(n991), .Y(n189) );
  INVX2TS U653 ( .A(n189), .Y(n205) );
  INVX2TS U654 ( .A(n177), .Y(n989) );
  INVX2TS U655 ( .A(n989), .Y(n1782) );
  INVX2TS U656 ( .A(n982), .Y(n193) );
  OR2X1TS U657 ( .A(n1601), .B(n181), .Y(n192) );
  INVX2TS U658 ( .A(n192), .Y(n179) );
  INVX2TS U659 ( .A(n179), .Y(n990) );
  INVX2TS U660 ( .A(n990), .Y(n208) );
  AOI22X1TS U661 ( .A0(n193), .A1(\destinationAddressbuffer[2][8] ), .B0(n208), 
        .B1(n321), .Y(n186) );
  INVX2TS U662 ( .A(n194), .Y(n1355) );
  INVX2TS U663 ( .A(n3), .Y(n1108) );
  AOI22X1TS U664 ( .A0(n1355), .A1(n328), .B0(n1108), .B1(n327), .Y(n185) );
  OAI211XLTS U665 ( .A0(n205), .A1(n232), .B0(n186), .C0(n185), .Y(n2118) );
  INVX2TS U666 ( .A(n192), .Y(n1801) );
  AOI22X1TS U667 ( .A0(n193), .A1(\destinationAddressbuffer[2][9] ), .B0(n1801), .B1(n331), .Y(n188) );
  INVX2TS U668 ( .A(n194), .Y(n992) );
  INVX2TS U669 ( .A(n3), .Y(n1784) );
  AOI22X1TS U670 ( .A0(n992), .A1(n333), .B0(n1784), .B1(n332), .Y(n187) );
  OAI211XLTS U671 ( .A0(n205), .A1(n226), .B0(n188), .C0(n187), .Y(n2119) );
  INVX2TS U672 ( .A(n189), .Y(n212) );
  INVX2TS U673 ( .A(n192), .Y(n1107) );
  AOI22X1TS U674 ( .A0(n193), .A1(\destinationAddressbuffer[2][10] ), .B0(
        n1107), .B1(n337), .Y(n191) );
  INVX2TS U675 ( .A(n194), .Y(n1343) );
  INVX2TS U676 ( .A(n3), .Y(n1354) );
  AOI22X1TS U677 ( .A0(n1337), .A1(n339), .B0(n1354), .B1(n338), .Y(n190) );
  OAI211XLTS U678 ( .A0(n212), .A1(n223), .B0(n191), .C0(n190), .Y(n2120) );
  INVX2TS U679 ( .A(n192), .Y(n1783) );
  AOI22X1TS U680 ( .A0(n193), .A1(\destinationAddressbuffer[2][11] ), .B0(
        n1783), .B1(n343), .Y(n197) );
  INVX2TS U681 ( .A(n194), .Y(n1785) );
  INVX2TS U682 ( .A(n3), .Y(n195) );
  INVX2TS U683 ( .A(n195), .Y(n978) );
  INVX2TS U684 ( .A(n978), .Y(n198) );
  AOI22X1TS U685 ( .A0(n1785), .A1(n348), .B0(n198), .B1(n347), .Y(n196) );
  OAI211XLTS U686 ( .A0(n205), .A1(n238), .B0(n197), .C0(n196), .Y(n2121) );
  CLKBUFX2TS U687 ( .A(n982), .Y(n1605) );
  INVX2TS U688 ( .A(n1605), .Y(n1800) );
  AOI22X1TS U689 ( .A0(n1800), .A1(writeOutbuffer[2]), .B0(n208), .B1(n351), 
        .Y(n200) );
  AOI22X1TS U690 ( .A0(n1355), .A1(n354), .B0(n198), .B1(n352), .Y(n199) );
  OAI211XLTS U691 ( .A0(n212), .A1(n243), .B0(n200), .C0(n199), .Y(n2039) );
  INVX2TS U692 ( .A(n982), .Y(n209) );
  AOI22X1TS U693 ( .A0(n209), .A1(\destinationAddressbuffer[2][6] ), .B0(n179), 
        .B1(n363), .Y(n202) );
  AOI22X1TS U694 ( .A0(n1343), .A1(destinationAddressIn_NORTH[6]), .B0(n195), 
        .B1(n364), .Y(n201) );
  OAI211XLTS U695 ( .A0(n212), .A1(n251), .B0(n202), .C0(n201), .Y(n2116) );
  AOI22X1TS U696 ( .A0(n209), .A1(\destinationAddressbuffer[2][5] ), .B0(n1107), .B1(n369), .Y(n204) );
  AOI22X1TS U697 ( .A0(n1337), .A1(destinationAddressIn_NORTH[5]), .B0(n198), 
        .B1(n370), .Y(n203) );
  OAI211XLTS U698 ( .A0(n205), .A1(n247), .B0(n204), .C0(n203), .Y(n2115) );
  AOI22X1TS U699 ( .A0(n209), .A1(\destinationAddressbuffer[2][7] ), .B0(n1783), .B1(n374), .Y(n207) );
  AOI22X1TS U700 ( .A0(n992), .A1(destinationAddressIn_NORTH[7]), .B0(n1108), 
        .B1(n376), .Y(n206) );
  OAI211XLTS U701 ( .A0(n1341), .A1(n256), .B0(n207), .C0(n206), .Y(n2117) );
  AOI22X1TS U702 ( .A0(n209), .A1(\destinationAddressbuffer[2][4] ), .B0(n208), 
        .B1(n357), .Y(n211) );
  AOI22X1TS U703 ( .A0(n992), .A1(destinationAddressIn_NORTH[4]), .B0(n1354), 
        .B1(n359), .Y(n210) );
  OAI211XLTS U704 ( .A0(n212), .A1(n260), .B0(n211), .C0(n210), .Y(n2114) );
  INVX2TS U705 ( .A(n1908), .Y(n389) );
  INVX2TS U706 ( .A(n1908), .Y(n314) );
  NAND2X1TS U707 ( .A(n216), .B(n1572), .Y(n218) );
  INVX2TS U708 ( .A(n1), .Y(n1434) );
  INVX2TS U709 ( .A(n1434), .Y(n917) );
  CLKBUFX2TS U710 ( .A(n917), .Y(n227) );
  INVX2TS U711 ( .A(n227), .Y(n252) );
  INVX2TS U712 ( .A(n215), .Y(n915) );
  INVX2TS U713 ( .A(n915), .Y(n1687) );
  OR2X1TS U714 ( .A(n216), .B(n1687), .Y(n1422) );
  CLKBUFX2TS U715 ( .A(n1422), .Y(n916) );
  INVX2TS U716 ( .A(n916), .Y(n234) );
  OR2X1TS U717 ( .A(n1569), .B(n218), .Y(n233) );
  INVX2TS U718 ( .A(n233), .Y(n1423) );
  AOI22X1TS U719 ( .A0(n234), .A1(\destinationAddressbuffer[5][10] ), .B0(
        n1423), .B1(n745), .Y(n222) );
  INVX2TS U720 ( .A(n1562), .Y(n1565) );
  NAND2BX1TS U721 ( .AN(n218), .B(n217), .Y(n220) );
  INVX2TS U722 ( .A(n253), .Y(n1692) );
  INVX2TS U723 ( .A(n1692), .Y(n244) );
  INVX2TS U724 ( .A(n244), .Y(n911) );
  OR2X1TS U725 ( .A(n1562), .B(n220), .Y(n240) );
  INVX2TS U726 ( .A(n240), .Y(n1445) );
  AOI22X1TS U727 ( .A0(n911), .A1(n414), .B0(n1445), .B1(n338), .Y(n221) );
  OAI211XLTS U728 ( .A0(n252), .A1(n223), .B0(n222), .C0(n221), .Y(n2084) );
  INVX2TS U729 ( .A(n233), .Y(n1715) );
  INVX2TS U730 ( .A(n1715), .Y(n907) );
  INVX2TS U731 ( .A(n907), .Y(n248) );
  AOI22X1TS U732 ( .A0(n234), .A1(\destinationAddressbuffer[5][9] ), .B0(n248), 
        .B1(n728), .Y(n225) );
  INVX2TS U733 ( .A(n253), .Y(n1426) );
  INVX2TS U734 ( .A(n240), .Y(n1691) );
  AOI22X1TS U735 ( .A0(n1426), .A1(n398), .B0(n1691), .B1(n332), .Y(n224) );
  OAI211XLTS U736 ( .A0(n252), .A1(n226), .B0(n225), .C0(n224), .Y(n2083) );
  INVX2TS U737 ( .A(n227), .Y(n261) );
  INVX2TS U738 ( .A(n233), .Y(n228) );
  AOI22X1TS U739 ( .A0(n234), .A1(\destinationAddressbuffer[5][8] ), .B0(n228), 
        .B1(n713), .Y(n231) );
  INVX2TS U740 ( .A(n240), .Y(n229) );
  INVX2TS U741 ( .A(n229), .Y(n903) );
  INVX2TS U742 ( .A(n903), .Y(n235) );
  AOI22X1TS U743 ( .A0(n1436), .A1(n409), .B0(n235), .B1(n327), .Y(n230) );
  OAI211XLTS U744 ( .A0(n261), .A1(n232), .B0(n231), .C0(n230), .Y(n2082) );
  INVX2TS U745 ( .A(n233), .Y(n1690) );
  AOI22X1TS U746 ( .A0(n234), .A1(\destinationAddressbuffer[5][11] ), .B0(
        n1690), .B1(n761), .Y(n237) );
  INVX2TS U747 ( .A(n253), .Y(n1447) );
  AOI22X1TS U748 ( .A0(n1447), .A1(n403), .B0(n235), .B1(n347), .Y(n236) );
  OAI211XLTS U749 ( .A0(n252), .A1(n238), .B0(n237), .C0(n236), .Y(n2085) );
  INVX2TS U750 ( .A(n916), .Y(n1711) );
  INVX2TS U751 ( .A(n907), .Y(n239) );
  AOI22X1TS U752 ( .A0(n1711), .A1(writeOutbuffer[5]), .B0(n239), .B1(n542), 
        .Y(n242) );
  INVX2TS U753 ( .A(n240), .Y(n1424) );
  AOI22X1TS U754 ( .A0(n1426), .A1(n421), .B0(n1424), .B1(n352), .Y(n241) );
  OAI211XLTS U755 ( .A0(n261), .A1(n243), .B0(n242), .C0(n241), .Y(n2036) );
  AOI22X1TS U756 ( .A0(n257), .A1(\destinationAddressbuffer[5][5] ), .B0(n1423), .B1(n668), .Y(n246) );
  INVX2TS U757 ( .A(n244), .Y(n1700) );
  AOI22X1TS U758 ( .A0(n1700), .A1(n433), .B0(n1445), .B1(n370), .Y(n245) );
  OAI211XLTS U759 ( .A0(n261), .A1(n247), .B0(n246), .C0(n245), .Y(n2079) );
  AOI22X1TS U760 ( .A0(n257), .A1(\destinationAddressbuffer[5][6] ), .B0(n248), 
        .B1(n688), .Y(n250) );
  AOI22X1TS U761 ( .A0(n1692), .A1(n427), .B0(n229), .B1(n364), .Y(n249) );
  OAI211XLTS U762 ( .A0(n252), .A1(n251), .B0(n250), .C0(n249), .Y(n2080) );
  AOI22X1TS U763 ( .A0(n257), .A1(\destinationAddressbuffer[5][7] ), .B0(n1690), .B1(n702), .Y(n255) );
  INVX2TS U764 ( .A(n253), .Y(n1436) );
  AOI22X1TS U765 ( .A0(n1436), .A1(n424), .B0(n1424), .B1(n376), .Y(n254) );
  OAI211XLTS U766 ( .A0(n1434), .A1(n256), .B0(n255), .C0(n254), .Y(n2081) );
  AOI22X1TS U767 ( .A0(n257), .A1(\destinationAddressbuffer[5][4] ), .B0(n228), 
        .B1(n656), .Y(n259) );
  AOI22X1TS U768 ( .A0(n1447), .A1(n438), .B0(n235), .B1(n359), .Y(n258) );
  OAI211XLTS U769 ( .A0(n261), .A1(n260), .B0(n259), .C0(n258), .Y(n2078) );
  AOI31XLTS U770 ( .A0(n451), .A1(n386), .A2(n314), .B0(n1575), .Y(n268) );
  AOI21X1TS U771 ( .A0(n273), .A1(n268), .B0(n441), .Y(n272) );
  NAND2X1TS U772 ( .A(n272), .B(n1583), .Y(n274) );
  INVX2TS U773 ( .A(n270), .Y(n1401) );
  INVX2TS U774 ( .A(n1401), .Y(n943) );
  CLKBUFX2TS U775 ( .A(n943), .Y(n282) );
  INVX2TS U776 ( .A(n282), .Y(n302) );
  INVX2TS U777 ( .A(n271), .Y(n941) );
  INVX2TS U778 ( .A(n941), .Y(n1720) );
  CLKBUFX2TS U779 ( .A(n1390), .Y(n942) );
  INVX2TS U780 ( .A(n942), .Y(n288) );
  OR2X1TS U781 ( .A(n1579), .B(n274), .Y(n287) );
  INVX2TS U782 ( .A(n287), .Y(n1392) );
  AOI22X1TS U783 ( .A0(n288), .A1(\destinationAddressbuffer[4][10] ), .B0(
        n1392), .B1(n337), .Y(n278) );
  INVX2TS U784 ( .A(n279), .Y(n1393) );
  INVX2TS U785 ( .A(n1393), .Y(n308) );
  INVX2TS U786 ( .A(n276), .Y(n294) );
  INVX2TS U787 ( .A(n276), .Y(n923) );
  INVX2TS U788 ( .A(n923), .Y(n289) );
  AOI22X1TS U789 ( .A0(n308), .A1(n748), .B0(n289), .B1(n414), .Y(n277) );
  OAI211XLTS U790 ( .A0(n302), .A1(n27), .B0(n278), .C0(n277), .Y(n2096) );
  INVX2TS U791 ( .A(n282), .Y(n306) );
  INVX2TS U792 ( .A(n287), .Y(n1743) );
  INVX2TS U793 ( .A(n1743), .Y(n928) );
  INVX2TS U794 ( .A(n928), .Y(n303) );
  AOI22X1TS U795 ( .A0(n288), .A1(\destinationAddressbuffer[4][9] ), .B0(n303), 
        .B1(n331), .Y(n281) );
  INVX2TS U796 ( .A(n279), .Y(n293) );
  INVX2TS U797 ( .A(n293), .Y(n1745) );
  INVX2TS U798 ( .A(n294), .Y(n1744) );
  INVX2TS U799 ( .A(n294), .Y(n931) );
  AOI22X1TS U800 ( .A0(n1745), .A1(n729), .B0(n931), .B1(n398), .Y(n280) );
  OAI211XLTS U801 ( .A0(n306), .A1(n34), .B0(n281), .C0(n280), .Y(n2095) );
  INVX2TS U802 ( .A(n287), .Y(n283) );
  AOI22X1TS U803 ( .A0(n288), .A1(\destinationAddressbuffer[4][8] ), .B0(n283), 
        .B1(n321), .Y(n286) );
  INVX2TS U804 ( .A(n293), .Y(n284) );
  AOI22X1TS U805 ( .A0(n284), .A1(n714), .B0(n289), .B1(n409), .Y(n285) );
  OAI211XLTS U806 ( .A0(n302), .A1(n43), .B0(n286), .C0(n285), .Y(n2094) );
  INVX2TS U807 ( .A(n287), .Y(n1721) );
  AOI22X1TS U808 ( .A0(n288), .A1(\destinationAddressbuffer[4][11] ), .B0(
        n1721), .B1(n343), .Y(n291) );
  INVX2TS U809 ( .A(n293), .Y(n1736) );
  AOI22X1TS U810 ( .A0(n1736), .A1(n764), .B0(n289), .B1(n403), .Y(n290) );
  OAI211XLTS U811 ( .A0(n302), .A1(n39), .B0(n291), .C0(n290), .Y(n2097) );
  INVX2TS U812 ( .A(n942), .Y(n1740) );
  INVX2TS U813 ( .A(n928), .Y(n292) );
  AOI22X1TS U814 ( .A0(n1740), .A1(writeOutbuffer[4]), .B0(n292), .B1(n351), 
        .Y(n296) );
  INVX2TS U815 ( .A(n293), .Y(n1413) );
  AOI22X1TS U816 ( .A0(n1413), .A1(n544), .B0(n276), .B1(n421), .Y(n295) );
  OAI211XLTS U817 ( .A0(n306), .A1(n47), .B0(n296), .C0(n295), .Y(n2037) );
  INVX2TS U818 ( .A(n1390), .Y(n307) );
  AOI22X1TS U819 ( .A0(n307), .A1(\destinationAddressbuffer[4][5] ), .B0(n1392), .B1(n369), .Y(n299) );
  INVX2TS U820 ( .A(n294), .Y(n297) );
  AOI22X1TS U821 ( .A0(n1413), .A1(n670), .B0(n297), .B1(n433), .Y(n298) );
  OAI211XLTS U822 ( .A0(n306), .A1(n57), .B0(n299), .C0(n298), .Y(n2091) );
  AOI22X1TS U823 ( .A0(n307), .A1(\destinationAddressbuffer[4][4] ), .B0(n283), 
        .B1(n357), .Y(n301) );
  AOI22X1TS U824 ( .A0(n308), .A1(n658), .B0(n297), .B1(n438), .Y(n300) );
  OAI211XLTS U825 ( .A0(n302), .A1(n53), .B0(n301), .C0(n300), .Y(n2090) );
  AOI22X1TS U826 ( .A0(n307), .A1(\destinationAddressbuffer[4][6] ), .B0(n303), 
        .B1(n363), .Y(n305) );
  AOI22X1TS U827 ( .A0(n284), .A1(n690), .B0(n931), .B1(n427), .Y(n304) );
  OAI211XLTS U828 ( .A0(n306), .A1(n66), .B0(n305), .C0(n304), .Y(n2092) );
  AOI22X1TS U829 ( .A0(n307), .A1(\destinationAddressbuffer[4][7] ), .B0(n1721), .B1(n374), .Y(n310) );
  AOI22X1TS U830 ( .A0(n308), .A1(n703), .B0(n276), .B1(n424), .Y(n309) );
  OAI211XLTS U831 ( .A0(n1401), .A1(n63), .B0(n310), .C0(n309), .Y(n2093) );
  AOI31XLTS U832 ( .A0(n315), .A1(n314), .A2(n450), .B0(n1609), .Y(n317) );
  AOI21X1TS U833 ( .A0(n322), .A1(n317), .B0(n316), .Y(n319) );
  NAND2X1TS U834 ( .A(n319), .B(n1617), .Y(n323) );
  INVX2TS U835 ( .A(n318), .Y(n1086) );
  INVX2TS U836 ( .A(n1086), .Y(n1018) );
  CLKBUFX2TS U837 ( .A(n1018), .Y(n336) );
  INVX2TS U838 ( .A(n336), .Y(n368) );
  OR2X1TS U839 ( .A(n441), .B(n1617), .Y(n1081) );
  INVX2TS U840 ( .A(n1081), .Y(n1836) );
  OR2X1TS U841 ( .A(n319), .B(n1836), .Y(n1004) );
  INVX2TS U842 ( .A(n1004), .Y(n344) );
  OR2X1TS U843 ( .A(n1613), .B(n323), .Y(n342) );
  INVX2TS U844 ( .A(n342), .Y(n320) );
  INVX2TS U845 ( .A(n320), .Y(n1017) );
  INVX2TS U846 ( .A(n1017), .Y(n358) );
  AOI22X1TS U847 ( .A0(n344), .A1(\destinationAddressbuffer[1][8] ), .B0(n358), 
        .B1(n321), .Y(n330) );
  NAND2BX1TS U848 ( .AN(n323), .B(n322), .Y(n326) );
  INVX2TS U849 ( .A(n345), .Y(n1098) );
  INVX2TS U850 ( .A(n4), .Y(n1077) );
  AOI22X1TS U851 ( .A0(n1098), .A1(n328), .B0(n1077), .B1(n327), .Y(n329) );
  OAI211XLTS U852 ( .A0(n368), .A1(n43), .B0(n330), .C0(n329), .Y(n2130) );
  INVX2TS U853 ( .A(n342), .Y(n1839) );
  AOI22X1TS U854 ( .A0(n344), .A1(\destinationAddressbuffer[1][9] ), .B0(n1839), .B1(n331), .Y(n335) );
  INVX2TS U855 ( .A(n345), .Y(n1020) );
  INVX2TS U856 ( .A(n4), .Y(n1810) );
  AOI22X1TS U857 ( .A0(n1020), .A1(n333), .B0(n1810), .B1(n332), .Y(n334) );
  OAI211XLTS U858 ( .A0(n368), .A1(n34), .B0(n335), .C0(n334), .Y(n2131) );
  INVX2TS U859 ( .A(n336), .Y(n380) );
  INVX2TS U860 ( .A(n342), .Y(n1076) );
  AOI22X1TS U861 ( .A0(n344), .A1(\destinationAddressbuffer[1][10] ), .B0(
        n1076), .B1(n337), .Y(n341) );
  INVX2TS U862 ( .A(n345), .Y(n1087) );
  INVX2TS U863 ( .A(n4), .Y(n1097) );
  AOI22X1TS U864 ( .A0(n1082), .A1(n339), .B0(n1097), .B1(n338), .Y(n340) );
  OAI211XLTS U865 ( .A0(n380), .A1(n27), .B0(n341), .C0(n340), .Y(n2132) );
  INVX2TS U866 ( .A(n342), .Y(n1808) );
  AOI22X1TS U867 ( .A0(n344), .A1(\destinationAddressbuffer[1][11] ), .B0(
        n1808), .B1(n343), .Y(n350) );
  INVX2TS U868 ( .A(n345), .Y(n1812) );
  INVX2TS U869 ( .A(n4), .Y(n346) );
  INVX2TS U870 ( .A(n346), .Y(n998) );
  INVX2TS U871 ( .A(n998), .Y(n353) );
  AOI22X1TS U872 ( .A0(n1812), .A1(n348), .B0(n353), .B1(n347), .Y(n349) );
  OAI211XLTS U873 ( .A0(n368), .A1(n39), .B0(n350), .C0(n349), .Y(n2133) );
  CLKBUFX2TS U874 ( .A(n1004), .Y(n1618) );
  INVX2TS U875 ( .A(n1618), .Y(n1835) );
  AOI22X1TS U876 ( .A0(n1835), .A1(writeOutbuffer[1]), .B0(n358), .B1(n351), 
        .Y(n356) );
  AOI22X1TS U877 ( .A0(n1098), .A1(n354), .B0(n353), .B1(n352), .Y(n355) );
  OAI211XLTS U878 ( .A0(n380), .A1(n47), .B0(n356), .C0(n355), .Y(n2040) );
  INVX2TS U879 ( .A(n1004), .Y(n375) );
  AOI22X1TS U880 ( .A0(n375), .A1(\destinationAddressbuffer[1][4] ), .B0(n358), 
        .B1(n357), .Y(n362) );
  AOI22X1TS U881 ( .A0(n1098), .A1(n360), .B0(n1097), .B1(n359), .Y(n361) );
  OAI211XLTS U882 ( .A0(n380), .A1(n53), .B0(n362), .C0(n361), .Y(n2126) );
  AOI22X1TS U883 ( .A0(n375), .A1(\destinationAddressbuffer[1][6] ), .B0(n320), 
        .B1(n363), .Y(n367) );
  AOI22X1TS U884 ( .A0(n1087), .A1(n365), .B0(n346), .B1(n364), .Y(n366) );
  OAI211XLTS U885 ( .A0(n368), .A1(n66), .B0(n367), .C0(n366), .Y(n2128) );
  AOI22X1TS U886 ( .A0(n375), .A1(\destinationAddressbuffer[1][5] ), .B0(n1076), .B1(n369), .Y(n373) );
  AOI22X1TS U887 ( .A0(n1082), .A1(n371), .B0(n353), .B1(n370), .Y(n372) );
  OAI211XLTS U888 ( .A0(n1086), .A1(n57), .B0(n373), .C0(n372), .Y(n2127) );
  AOI22X1TS U889 ( .A0(n375), .A1(\destinationAddressbuffer[1][7] ), .B0(n1808), .B1(n374), .Y(n379) );
  AOI22X1TS U890 ( .A0(n1020), .A1(n377), .B0(n1077), .B1(n376), .Y(n378) );
  OAI211XLTS U891 ( .A0(n380), .A1(n63), .B0(n379), .C0(n378), .Y(n2129) );
  AOI31XLTS U892 ( .A0(n386), .A1(n389), .A2(n444), .B0(n1621), .Y(n388) );
  AOI21X1TS U893 ( .A0(n395), .A1(n388), .B0(n387), .Y(n393) );
  NAND2X1TS U894 ( .A(n393), .B(n1629), .Y(n396) );
  INVX2TS U895 ( .A(n391), .Y(n1058) );
  INVX2TS U896 ( .A(n1058), .Y(n1043) );
  CLKBUFX2TS U897 ( .A(n1043), .Y(n406) );
  INVX2TS U898 ( .A(n406), .Y(n431) );
  INVX2TS U899 ( .A(n9), .Y(n1846) );
  CLKBUFX2TS U900 ( .A(n1031), .Y(n1041) );
  INVX2TS U901 ( .A(n1041), .Y(n413) );
  OR2X1TS U902 ( .A(n1626), .B(n396), .Y(n418) );
  INVX2TS U903 ( .A(n418), .Y(n1877) );
  AOI22X1TS U904 ( .A0(n413), .A1(\destinationAddressbuffer[0][9] ), .B0(n419), 
        .B1(n394), .Y(n400) );
  INVX2TS U905 ( .A(n2), .Y(n1881) );
  INVX2TS U906 ( .A(n5), .Y(n1879) );
  AOI22X1TS U907 ( .A0(n1881), .A1(n729), .B0(n1879), .B1(n398), .Y(n399) );
  OAI211XLTS U908 ( .A0(n431), .A1(n34), .B0(n400), .C0(n399), .Y(n2143) );
  INVX2TS U909 ( .A(n406), .Y(n436) );
  AOI22X1TS U910 ( .A0(n413), .A1(\destinationAddressbuffer[0][11] ), .B0(n432), .B1(n401), .Y(n405) );
  INVX2TS U911 ( .A(n2), .Y(n1870) );
  INVX2TS U912 ( .A(n5), .Y(n402) );
  INVX2TS U913 ( .A(n402), .Y(n1027) );
  INVX2TS U914 ( .A(n1027), .Y(n415) );
  AOI22X1TS U915 ( .A0(n1870), .A1(n764), .B0(n415), .B1(n403), .Y(n404) );
  OAI211XLTS U916 ( .A0(n436), .A1(n39), .B0(n405), .C0(n404), .Y(n2145) );
  INVX2TS U917 ( .A(n418), .Y(n1050) );
  AOI22X1TS U918 ( .A0(n413), .A1(\destinationAddressbuffer[0][8] ), .B0(n1050), .B1(n407), .Y(n411) );
  INVX2TS U919 ( .A(n2), .Y(n408) );
  INVX2TS U920 ( .A(n408), .Y(n1045) );
  INVX2TS U921 ( .A(n1045), .Y(n428) );
  INVX2TS U922 ( .A(n5), .Y(n1850) );
  AOI22X1TS U923 ( .A0(n428), .A1(n714), .B0(n1850), .B1(n409), .Y(n410) );
  OAI211XLTS U924 ( .A0(n431), .A1(n43), .B0(n411), .C0(n410), .Y(n2142) );
  INVX2TS U925 ( .A(n418), .Y(n1848) );
  AOI22X1TS U926 ( .A0(n413), .A1(\destinationAddressbuffer[0][10] ), .B0(
        n1848), .B1(n412), .Y(n417) );
  AOI22X1TS U927 ( .A0(n408), .A1(n748), .B0(n415), .B1(n414), .Y(n416) );
  OAI211XLTS U928 ( .A0(n431), .A1(n27), .B0(n417), .C0(n416), .Y(n2144) );
  INVX2TS U929 ( .A(n1031), .Y(n1874) );
  INVX2TS U930 ( .A(n418), .Y(n419) );
  INVX2TS U931 ( .A(n419), .Y(n1042) );
  INVX2TS U932 ( .A(n1042), .Y(n432) );
  AOI22X1TS U933 ( .A0(n1874), .A1(writeOutbuffer[0]), .B0(n432), .B1(n420), 
        .Y(n423) );
  INVX2TS U934 ( .A(n2), .Y(n1068) );
  INVX2TS U935 ( .A(n5), .Y(n1051) );
  AOI22X1TS U936 ( .A0(n1068), .A1(n544), .B0(n1051), .B1(n421), .Y(n422) );
  OAI211XLTS U937 ( .A0(n436), .A1(n47), .B0(n423), .C0(n422), .Y(n2041) );
  INVX2TS U938 ( .A(n1031), .Y(n437) );
  AOI22X1TS U939 ( .A0(n437), .A1(\destinationAddressbuffer[0][7] ), .B0(n1050), .B1(destinationAddressIn_WEST[7]), .Y(n426) );
  AOI22X1TS U940 ( .A0(n408), .A1(n703), .B0(n1051), .B1(n424), .Y(n425) );
  OAI211XLTS U941 ( .A0(n436), .A1(n63), .B0(n426), .C0(n425), .Y(n2141) );
  AOI22X1TS U942 ( .A0(n437), .A1(\destinationAddressbuffer[0][6] ), .B0(n1877), .B1(destinationAddressIn_WEST[6]), .Y(n430) );
  AOI22X1TS U943 ( .A0(n428), .A1(n690), .B0(n402), .B1(n427), .Y(n429) );
  OAI211XLTS U944 ( .A0(n431), .A1(n66), .B0(n430), .C0(n429), .Y(n2140) );
  AOI22X1TS U945 ( .A0(n437), .A1(\destinationAddressbuffer[0][5] ), .B0(n432), 
        .B1(destinationAddressIn_WEST[5]), .Y(n435) );
  AOI22X1TS U946 ( .A0(n1068), .A1(n670), .B0(n415), .B1(n433), .Y(n434) );
  OAI211XLTS U947 ( .A0(n436), .A1(n57), .B0(n435), .C0(n434), .Y(n2139) );
  AOI22X1TS U948 ( .A0(n437), .A1(\destinationAddressbuffer[0][4] ), .B0(n1848), .B1(destinationAddressIn_WEST[4]), .Y(n440) );
  AOI22X1TS U949 ( .A0(n408), .A1(n658), .B0(n1850), .B1(n438), .Y(n439) );
  OAI211XLTS U950 ( .A0(n1058), .A1(n53), .B0(n440), .C0(n439), .Y(n2138) );
  INVX2TS U951 ( .A(n1913), .Y(n527) );
  INVX2TS U952 ( .A(n1913), .Y(n524) );
  INVX2TS U953 ( .A(n1906), .Y(n530) );
  NAND2X1TS U954 ( .A(n524), .B(n530), .Y(n528) );
  OAI21XLTS U955 ( .A0(n527), .A1(n1907), .B0(n528), .Y(n502) );
  INVX2TS U956 ( .A(n1903), .Y(n531) );
  INVX2TS U957 ( .A(n1903), .Y(n526) );
  NOR2XLTS U958 ( .A(n528), .B(n526), .Y(n834) );
  CLKBUFX2TS U959 ( .A(n834), .Y(n794) );
  CLKBUFX2TS U960 ( .A(n794), .Y(n814) );
  AOI21X1TS U961 ( .A0(n528), .A1(n531), .B0(n814), .Y(n499) );
  OAI22X1TS U962 ( .A0(n484), .A1(n502), .B0(n442), .B1(n499), .Y(n443) );
  AOI221XLTS U963 ( .A0(n502), .A1(n445), .B0(n444), .B1(n499), .C0(n443), .Y(
        n448) );
  INVX2TS U964 ( .A(n1900), .Y(n446) );
  NAND2X1TS U965 ( .A(n447), .B(n446), .Y(n460) );
  OAI21XLTS U966 ( .A0(n482), .A1(n1913), .B0(n460), .Y(n464) );
  AOI21X1TS U967 ( .A0(n448), .A1(n464), .B0(n1902), .Y(n449) );
  NAND2X1TS U968 ( .A(n491), .B(n1902), .Y(n503) );
  INVX2TS U969 ( .A(n1908), .Y(n461) );
  INVX2TS U970 ( .A(n1911), .Y(n451) );
  INVX2TS U971 ( .A(n1904), .Y(n529) );
  AOI22X1TS U972 ( .A0(n451), .A1(n526), .B0(n529), .B1(n450), .Y(n454) );
  INVX2TS U973 ( .A(n453), .Y(n459) );
  INVX2TS U974 ( .A(n474), .Y(n471) );
  AOI21X1TS U975 ( .A0(n527), .A1(n457), .B0(n456), .Y(n470) );
  ADDHXLTS U976 ( .A(n463), .B(n462), .CO(n474), .S(n476) );
  INVX2TS U977 ( .A(n476), .Y(n465) );
  AOI21X1TS U978 ( .A0(n466), .A1(n465), .B0(n464), .Y(n468) );
  OAI22X1TS U979 ( .A0(n466), .A1(n465), .B0(n472), .B1(n471), .Y(n467) );
  AOI21X1TS U980 ( .A0(n475), .A1(n468), .B0(n467), .Y(n469) );
  AOI211X1TS U981 ( .A0(n472), .A1(n471), .B0(n470), .C0(n469), .Y(n473) );
  INVX2TS U982 ( .A(n473), .Y(n477) );
  NAND2X1TS U983 ( .A(n477), .B(n474), .Y(n480) );
  INVX2TS U984 ( .A(n495), .Y(n489) );
  INVX2TS U985 ( .A(n1904), .Y(n525) );
  ADDHXLTS U986 ( .A(n482), .B(n481), .CO(n485), .S(n492) );
  XNOR2X1TS U987 ( .A(n1907), .B(n493), .Y(n486) );
  OAI21X1TS U988 ( .A0(n489), .A1(n525), .B0(n486), .Y(n487) );
  OAI2BB2XLTS U989 ( .B0(n1914), .B1(n503), .A0N(n496), .A1N(n490), .Y(N2624)
         );
  CLKBUFX2TS U990 ( .A(n1901), .Y(n640) );
  CLKBUFX2TS U991 ( .A(n640), .Y(n607) );
  NAND2X1TS U992 ( .A(n491), .B(n607), .Y(n501) );
  AOI22X1TS U993 ( .A0(n1900), .A1(n503), .B0(n501), .B1(n446), .Y(n1923) );
  INVX2TS U994 ( .A(n499), .Y(n500) );
  OAI22X1TS U995 ( .A0(n531), .A1(n503), .B0(n500), .B1(n501), .Y(n1928) );
  OAI22X1TS U996 ( .A0(n11), .A1(n503), .B0(n502), .B1(n501), .Y(n1929) );
  CLKBUFX2TS U997 ( .A(readIn_SOUTH), .Y(n1564) );
  CLKBUFX2TS U998 ( .A(n1901), .Y(n840) );
  CLKBUFX2TS U999 ( .A(n543), .Y(n846) );
  CLKBUFX2TS U1000 ( .A(readIn_WEST), .Y(n1581) );
  CLKBUFX2TS U1001 ( .A(n1581), .Y(n1615) );
  INVX2TS U1002 ( .A(n1901), .Y(n520) );
  NOR4XLTS U1003 ( .A(n514), .B(n513), .C(n453), .D(n508), .Y(n613) );
  CLKBUFX2TS U1004 ( .A(n613), .Y(n627) );
  CLKBUFX2TS U1005 ( .A(n627), .Y(n807) );
  CLKBUFX2TS U1006 ( .A(n807), .Y(n564) );
  AOI22X1TS U1007 ( .A0(n1564), .A1(n846), .B0(n1615), .B1(n564), .Y(n541) );
  CLKBUFX2TS U1008 ( .A(readIn_NORTH), .Y(n1595) );
  CLKBUFX2TS U1009 ( .A(n1595), .Y(n1563) );
  CLKBUFX2TS U1010 ( .A(n689), .Y(n563) );
  NOR4XLTS U1011 ( .A(n512), .B(n511), .C(n510), .D(n508), .Y(n589) );
  CLKBUFX2TS U1012 ( .A(n589), .Y(n600) );
  CLKBUFX2TS U1013 ( .A(n600), .Y(n775) );
  CLKBUFX2TS U1014 ( .A(n775), .Y(n824) );
  AOI22X1TS U1015 ( .A0(n1563), .A1(n563), .B0(readIn_EAST), .B1(n824), .Y(
        n540) );
  NOR3XLTS U1016 ( .A(n513), .B(n509), .C(n453), .Y(n516) );
  NOR3XLTS U1017 ( .A(n512), .B(n511), .C(n510), .Y(n515) );
  NAND4XLTS U1018 ( .A(n520), .B(n519), .C(n518), .D(n517), .Y(n732) );
  INVX2TS U1019 ( .A(n732), .Y(n521) );
  INVX2TS U1020 ( .A(n521), .Y(n580) );
  INVX2TS U1021 ( .A(n580), .Y(n522) );
  NOR3XLTS U1022 ( .A(n524), .B(n525), .C(n1906), .Y(n716) );
  CLKBUFX2TS U1023 ( .A(n716), .Y(n628) );
  CLKBUFX2TS U1024 ( .A(n628), .Y(n566) );
  NOR3XLTS U1025 ( .A(n527), .B(n1907), .C(n525), .Y(n691) );
  CLKBUFX2TS U1026 ( .A(n691), .Y(n629) );
  CLKBUFX2TS U1027 ( .A(n629), .Y(n565) );
  AOI22X1TS U1028 ( .A0(readOutbuffer[2]), .A1(n566), .B0(readOutbuffer[0]), 
        .B1(n565), .Y(n535) );
  NOR3XLTS U1029 ( .A(n524), .B(n11), .C(n526), .Y(n717) );
  CLKBUFX2TS U1030 ( .A(n717), .Y(n630) );
  CLKBUFX2TS U1031 ( .A(n630), .Y(n568) );
  NOR3XLTS U1032 ( .A(n527), .B(n530), .C(n531), .Y(n692) );
  CLKBUFX2TS U1033 ( .A(n692), .Y(n631) );
  CLKBUFX2TS U1034 ( .A(n631), .Y(n567) );
  AOI22X1TS U1035 ( .A0(readOutbuffer[6]), .A1(n568), .B0(readOutbuffer[4]), 
        .B1(n567), .Y(n534) );
  NOR2XLTS U1036 ( .A(n529), .B(n528), .Y(n718) );
  CLKBUFX2TS U1037 ( .A(n718), .Y(n632) );
  CLKBUFX2TS U1038 ( .A(n632), .Y(n570) );
  NOR3XLTS U1039 ( .A(n530), .B(n529), .C(n1913), .Y(n693) );
  CLKBUFX2TS U1040 ( .A(n693), .Y(n633) );
  CLKBUFX2TS U1041 ( .A(n633), .Y(n569) );
  AOI22X1TS U1042 ( .A0(readOutbuffer[3]), .A1(n570), .B0(readOutbuffer[1]), 
        .B1(n569), .Y(n533) );
  CLKBUFX2TS U1043 ( .A(n834), .Y(n855) );
  NOR3XLTS U1044 ( .A(n1907), .B(n446), .C(n531), .Y(n856) );
  CLKBUFX2TS U1045 ( .A(n856), .Y(n634) );
  CLKBUFX2TS U1046 ( .A(n634), .Y(n571) );
  AOI22X1TS U1047 ( .A0(readOutbuffer[7]), .A1(n855), .B0(readOutbuffer[5]), 
        .B1(n571), .Y(n532) );
  NAND4XLTS U1048 ( .A(n535), .B(n534), .C(n533), .D(n532), .Y(n536) );
  AOI22X1TS U1049 ( .A0(readOut), .A1(n551), .B0(n607), .B1(n536), .Y(n539) );
  INVX2TS U1050 ( .A(n10), .Y(n801) );
  CLKBUFX2TS U1051 ( .A(n775), .Y(n746) );
  AOI22X1TS U1052 ( .A0(writeIn_EAST), .A1(n746), .B0(n542), .B1(n564), .Y(
        n554) );
  CLKBUFX2TS U1053 ( .A(n543), .Y(n669) );
  CLKBUFX2TS U1054 ( .A(n669), .Y(n763) );
  AOI22X1TS U1055 ( .A0(n545), .A1(n563), .B0(n544), .B1(n763), .Y(n553) );
  AOI22X1TS U1056 ( .A0(writeOutbuffer[2]), .A1(n566), .B0(writeOutbuffer[0]), 
        .B1(n565), .Y(n549) );
  AOI22X1TS U1057 ( .A0(writeOutbuffer[6]), .A1(n568), .B0(writeOutbuffer[4]), 
        .B1(n567), .Y(n548) );
  AOI22X1TS U1058 ( .A0(writeOutbuffer[3]), .A1(n570), .B0(writeOutbuffer[1]), 
        .B1(n569), .Y(n547) );
  AOI22X1TS U1059 ( .A0(writeOutbuffer[7]), .A1(n855), .B0(writeOutbuffer[5]), 
        .B1(n571), .Y(n546) );
  NAND4XLTS U1060 ( .A(n549), .B(n548), .C(n547), .D(n546), .Y(n550) );
  AOI22X1TS U1061 ( .A0(writeOut), .A1(n551), .B0(n607), .B1(n550), .Y(n552)
         );
  CLKBUFX2TS U1062 ( .A(requesterAddressIn_NORTH[0]), .Y(n999) );
  CLKBUFX2TS U1063 ( .A(requesterAddressIn_EAST[0]), .Y(n1026) );
  CLKBUFX2TS U1064 ( .A(n1026), .Y(n997) );
  AOI22X1TS U1065 ( .A0(n999), .A1(n563), .B0(n997), .B1(n600), .Y(n562) );
  CLKBUFX2TS U1066 ( .A(requesterAddressIn_SOUTH[0]), .Y(n1000) );
  CLKBUFX2TS U1067 ( .A(n669), .Y(n657) );
  CLKBUFX2TS U1068 ( .A(requesterAddressIn_WEST[0]), .Y(n922) );
  CLKBUFX2TS U1069 ( .A(n922), .Y(n951) );
  AOI22X1TS U1070 ( .A0(n1000), .A1(n657), .B0(n951), .B1(n564), .Y(n561) );
  INVX2TS U1071 ( .A(n732), .Y(n684) );
  CLKBUFX2TS U1072 ( .A(n640), .Y(n595) );
  AOI22X1TS U1073 ( .A0(\requesterAddressbuffer[2][0] ), .A1(n566), .B0(
        \requesterAddressbuffer[0][0] ), .B1(n565), .Y(n558) );
  AOI22X1TS U1074 ( .A0(\requesterAddressbuffer[6][0] ), .A1(n568), .B0(
        \requesterAddressbuffer[4][0] ), .B1(n567), .Y(n557) );
  AOI22X1TS U1075 ( .A0(\requesterAddressbuffer[3][0] ), .A1(n570), .B0(
        \requesterAddressbuffer[1][0] ), .B1(n569), .Y(n556) );
  CLKBUFX2TS U1076 ( .A(n794), .Y(n750) );
  CLKBUFX2TS U1077 ( .A(n750), .Y(n601) );
  AOI22X1TS U1078 ( .A0(\requesterAddressbuffer[7][0] ), .A1(n601), .B0(
        \requesterAddressbuffer[5][0] ), .B1(n571), .Y(n555) );
  NAND4XLTS U1079 ( .A(n558), .B(n557), .C(n556), .D(n555), .Y(n559) );
  AOI22X1TS U1080 ( .A0(requesterAddressOut[0]), .A1(n684), .B0(n595), .B1(
        n559), .Y(n560) );
  INVX2TS U1081 ( .A(readRequesterAddress[0]), .Y(n949) );
  INVX2TS U1082 ( .A(n949), .Y(n996) );
  INVX2TS U1083 ( .A(n801), .Y(n596) );
  NAND2X1TS U1084 ( .A(n996), .B(n596), .Y(n608) );
  CLKBUFX2TS U1085 ( .A(requesterAddressIn_NORTH[1]), .Y(n1006) );
  CLKBUFX2TS U1086 ( .A(requesterAddressIn_EAST[1]), .Y(n1032) );
  CLKBUFX2TS U1087 ( .A(n1032), .Y(n1005) );
  AOI22X1TS U1088 ( .A0(n1006), .A1(n563), .B0(n1005), .B1(n589), .Y(n579) );
  CLKBUFX2TS U1089 ( .A(requesterAddressIn_SOUTH[1]), .Y(n1007) );
  CLKBUFX2TS U1090 ( .A(n543), .Y(n805) );
  CLKBUFX2TS U1091 ( .A(requesterAddressIn_WEST[1]), .Y(n930) );
  CLKBUFX2TS U1092 ( .A(n930), .Y(n958) );
  AOI22X1TS U1093 ( .A0(n1007), .A1(n805), .B0(n958), .B1(n564), .Y(n578) );
  INVX2TS U1094 ( .A(n732), .Y(n781) );
  AOI22X1TS U1095 ( .A0(\requesterAddressbuffer[2][1] ), .A1(n566), .B0(
        \requesterAddressbuffer[0][1] ), .B1(n565), .Y(n575) );
  AOI22X1TS U1096 ( .A0(\requesterAddressbuffer[6][1] ), .A1(n568), .B0(
        \requesterAddressbuffer[4][1] ), .B1(n567), .Y(n574) );
  AOI22X1TS U1097 ( .A0(\requesterAddressbuffer[3][1] ), .A1(n570), .B0(
        \requesterAddressbuffer[1][1] ), .B1(n569), .Y(n573) );
  AOI22X1TS U1098 ( .A0(\requesterAddressbuffer[7][1] ), .A1(n601), .B0(
        \requesterAddressbuffer[5][1] ), .B1(n571), .Y(n572) );
  NAND4XLTS U1099 ( .A(n575), .B(n574), .C(n573), .D(n572), .Y(n576) );
  AOI22X1TS U1100 ( .A0(requesterAddressOut[1]), .A1(n781), .B0(n595), .B1(
        n576), .Y(n577) );
  INVX2TS U1101 ( .A(readRequesterAddress[1]), .Y(n956) );
  INVX2TS U1102 ( .A(n956), .Y(n1635) );
  NAND2X1TS U1103 ( .A(n1635), .B(n596), .Y(n623) );
  CLKBUFX2TS U1104 ( .A(requesterAddressIn_NORTH[2]), .Y(n1012) );
  CLKBUFX2TS U1105 ( .A(n689), .Y(n612) );
  CLKBUFX2TS U1106 ( .A(requesterAddressIn_EAST[2]), .Y(n1036) );
  CLKBUFX2TS U1107 ( .A(n1036), .Y(n1011) );
  AOI22X1TS U1108 ( .A0(n1012), .A1(n612), .B0(n1011), .B1(n589), .Y(n588) );
  CLKBUFX2TS U1109 ( .A(requesterAddressIn_SOUTH[2]), .Y(n1013) );
  CLKBUFX2TS U1110 ( .A(requesterAddressIn_WEST[2]), .Y(n937) );
  CLKBUFX2TS U1111 ( .A(n937), .Y(n964) );
  AOI22X1TS U1112 ( .A0(n1013), .A1(n657), .B0(n964), .B1(n627), .Y(n587) );
  INVX2TS U1113 ( .A(n580), .Y(n757) );
  CLKBUFX2TS U1114 ( .A(n628), .Y(n614) );
  AOI22X1TS U1115 ( .A0(\requesterAddressbuffer[2][2] ), .A1(n614), .B0(
        \requesterAddressbuffer[0][2] ), .B1(n691), .Y(n584) );
  CLKBUFX2TS U1116 ( .A(n630), .Y(n615) );
  AOI22X1TS U1117 ( .A0(\requesterAddressbuffer[6][2] ), .A1(n615), .B0(
        \requesterAddressbuffer[4][2] ), .B1(n692), .Y(n583) );
  CLKBUFX2TS U1118 ( .A(n632), .Y(n616) );
  AOI22X1TS U1119 ( .A0(\requesterAddressbuffer[3][2] ), .A1(n616), .B0(
        \requesterAddressbuffer[1][2] ), .B1(n693), .Y(n582) );
  CLKBUFX2TS U1120 ( .A(n634), .Y(n617) );
  AOI22X1TS U1121 ( .A0(\requesterAddressbuffer[7][2] ), .A1(n601), .B0(
        \requesterAddressbuffer[5][2] ), .B1(n617), .Y(n581) );
  NAND4XLTS U1122 ( .A(n584), .B(n583), .C(n582), .D(n581), .Y(n585) );
  AOI22X1TS U1123 ( .A0(requesterAddressOut[2]), .A1(n757), .B0(n595), .B1(
        n585), .Y(n586) );
  INVX2TS U1124 ( .A(readRequesterAddress[2]), .Y(n963) );
  INVX2TS U1125 ( .A(n963), .Y(n1643) );
  NAND2X1TS U1126 ( .A(n1643), .B(n596), .Y(n641) );
  CLKBUFX2TS U1127 ( .A(requesterAddressIn_NORTH[3]), .Y(n1021) );
  CLKBUFX2TS U1128 ( .A(requesterAddressIn_EAST[3]), .Y(n1044) );
  CLKBUFX2TS U1129 ( .A(n1044), .Y(n1019) );
  AOI22X1TS U1130 ( .A0(n1021), .A1(n612), .B0(n1019), .B1(n589), .Y(n599) );
  CLKBUFX2TS U1131 ( .A(requesterAddressIn_SOUTH[3]), .Y(n1022) );
  CLKBUFX2TS U1132 ( .A(requesterAddressIn_WEST[3]), .Y(n945) );
  CLKBUFX2TS U1133 ( .A(n945), .Y(n973) );
  AOI22X1TS U1134 ( .A0(n1022), .A1(n805), .B0(n973), .B1(n613), .Y(n598) );
  AOI22X1TS U1135 ( .A0(\requesterAddressbuffer[2][3] ), .A1(n614), .B0(
        \requesterAddressbuffer[0][3] ), .B1(n691), .Y(n593) );
  AOI22X1TS U1136 ( .A0(\requesterAddressbuffer[6][3] ), .A1(n615), .B0(
        \requesterAddressbuffer[4][3] ), .B1(n692), .Y(n592) );
  AOI22X1TS U1137 ( .A0(\requesterAddressbuffer[3][3] ), .A1(n616), .B0(
        \requesterAddressbuffer[1][3] ), .B1(n693), .Y(n591) );
  CLKBUFX2TS U1138 ( .A(n750), .Y(n646) );
  AOI22X1TS U1139 ( .A0(\requesterAddressbuffer[7][3] ), .A1(n646), .B0(
        \requesterAddressbuffer[5][3] ), .B1(n617), .Y(n590) );
  NAND4XLTS U1140 ( .A(n593), .B(n592), .C(n591), .D(n590), .Y(n594) );
  AOI22X1TS U1141 ( .A0(requesterAddressOut[3]), .A1(n522), .B0(n595), .B1(
        n594), .Y(n597) );
  INVX2TS U1142 ( .A(readRequesterAddress[3]), .Y(n971) );
  INVX2TS U1143 ( .A(n971), .Y(n1653) );
  NAND2X1TS U1144 ( .A(n1653), .B(n596), .Y(n652) );
  CLKBUFX2TS U1145 ( .A(destinationAddressIn_EAST[0]), .Y(n1807) );
  CLKBUFX2TS U1146 ( .A(n1807), .Y(n1688) );
  CLKBUFX2TS U1147 ( .A(n600), .Y(n645) );
  AOI22X1TS U1148 ( .A0(destinationAddressIn_NORTH[0]), .A1(n612), .B0(n1688), 
        .B1(n645), .Y(n611) );
  CLKBUFX2TS U1149 ( .A(destinationAddressIn_WEST[0]), .Y(n1689) );
  CLKBUFX2TS U1150 ( .A(n1689), .Y(n1751) );
  AOI22X1TS U1151 ( .A0(destinationAddressIn_SOUTH[0]), .A1(n657), .B0(n1751), 
        .B1(n613), .Y(n610) );
  AOI22X1TS U1152 ( .A0(\destinationAddressbuffer[2][0] ), .A1(n614), .B0(
        \destinationAddressbuffer[0][0] ), .B1(n629), .Y(n605) );
  AOI22X1TS U1153 ( .A0(\destinationAddressbuffer[6][0] ), .A1(n615), .B0(
        \destinationAddressbuffer[4][0] ), .B1(n631), .Y(n604) );
  AOI22X1TS U1154 ( .A0(\destinationAddressbuffer[3][0] ), .A1(n616), .B0(
        \destinationAddressbuffer[1][0] ), .B1(n633), .Y(n603) );
  AOI22X1TS U1155 ( .A0(\destinationAddressbuffer[7][0] ), .A1(n601), .B0(
        \destinationAddressbuffer[5][0] ), .B1(n617), .Y(n602) );
  NAND4XLTS U1156 ( .A(n605), .B(n604), .C(n603), .D(n602), .Y(n606) );
  AOI22X1TS U1157 ( .A0(destinationAddressOut[0]), .A1(n684), .B0(n607), .B1(
        n606), .Y(n609) );
  CLKBUFX2TS U1158 ( .A(destinationAddressIn_EAST[1]), .Y(n1818) );
  CLKBUFX2TS U1159 ( .A(n1818), .Y(n1697) );
  AOI22X1TS U1160 ( .A0(destinationAddressIn_NORTH[1]), .A1(n612), .B0(n1697), 
        .B1(n645), .Y(n626) );
  CLKBUFX2TS U1161 ( .A(destinationAddressIn_WEST[1]), .Y(n1699) );
  CLKBUFX2TS U1162 ( .A(n1699), .Y(n1759) );
  AOI22X1TS U1163 ( .A0(destinationAddressIn_SOUTH[1]), .A1(n805), .B0(n1759), 
        .B1(n613), .Y(n625) );
  AOI22X1TS U1164 ( .A0(\destinationAddressbuffer[2][1] ), .A1(n614), .B0(
        \destinationAddressbuffer[0][1] ), .B1(n629), .Y(n621) );
  AOI22X1TS U1165 ( .A0(\destinationAddressbuffer[6][1] ), .A1(n615), .B0(
        \destinationAddressbuffer[4][1] ), .B1(n631), .Y(n620) );
  AOI22X1TS U1166 ( .A0(\destinationAddressbuffer[3][1] ), .A1(n616), .B0(
        \destinationAddressbuffer[1][1] ), .B1(n633), .Y(n619) );
  AOI22X1TS U1167 ( .A0(\destinationAddressbuffer[7][1] ), .A1(n646), .B0(
        \destinationAddressbuffer[5][1] ), .B1(n617), .Y(n618) );
  NAND4XLTS U1168 ( .A(n621), .B(n620), .C(n619), .D(n618), .Y(n622) );
  AOI22X1TS U1169 ( .A0(destinationAddressOut[1]), .A1(n684), .B0(n640), .B1(
        n622), .Y(n624) );
  CLKBUFX2TS U1170 ( .A(n689), .Y(n671) );
  CLKBUFX2TS U1171 ( .A(destinationAddressIn_EAST[2]), .Y(n1828) );
  CLKBUFX2TS U1172 ( .A(n1828), .Y(n1705) );
  AOI22X1TS U1173 ( .A0(destinationAddressIn_NORTH[2]), .A1(n671), .B0(n1705), 
        .B1(n645), .Y(n644) );
  CLKBUFX2TS U1174 ( .A(n543), .Y(n785) );
  CLKBUFX2TS U1175 ( .A(destinationAddressIn_WEST[2]), .Y(n1707) );
  CLKBUFX2TS U1176 ( .A(n1707), .Y(n1768) );
  CLKBUFX2TS U1177 ( .A(n627), .Y(n667) );
  AOI22X1TS U1178 ( .A0(destinationAddressIn_SOUTH[2]), .A1(n785), .B0(n1768), 
        .B1(n667), .Y(n643) );
  CLKBUFX2TS U1179 ( .A(n628), .Y(n673) );
  CLKBUFX2TS U1180 ( .A(n629), .Y(n672) );
  AOI22X1TS U1181 ( .A0(\destinationAddressbuffer[2][2] ), .A1(n673), .B0(
        \destinationAddressbuffer[0][2] ), .B1(n672), .Y(n638) );
  CLKBUFX2TS U1182 ( .A(n630), .Y(n675) );
  CLKBUFX2TS U1183 ( .A(n631), .Y(n674) );
  AOI22X1TS U1184 ( .A0(\destinationAddressbuffer[6][2] ), .A1(n675), .B0(
        \destinationAddressbuffer[4][2] ), .B1(n674), .Y(n637) );
  CLKBUFX2TS U1185 ( .A(n632), .Y(n677) );
  CLKBUFX2TS U1186 ( .A(n633), .Y(n676) );
  AOI22X1TS U1187 ( .A0(\destinationAddressbuffer[3][2] ), .A1(n677), .B0(
        \destinationAddressbuffer[1][2] ), .B1(n676), .Y(n636) );
  CLKBUFX2TS U1188 ( .A(n634), .Y(n678) );
  AOI22X1TS U1189 ( .A0(\destinationAddressbuffer[7][2] ), .A1(n646), .B0(
        \destinationAddressbuffer[5][2] ), .B1(n678), .Y(n635) );
  NAND4XLTS U1190 ( .A(n638), .B(n637), .C(n636), .D(n635), .Y(n639) );
  AOI22X1TS U1191 ( .A0(destinationAddressOut[2]), .A1(n522), .B0(n640), .B1(
        n639), .Y(n642) );
  CLKBUFX2TS U1192 ( .A(destinationAddressIn_EAST[3]), .Y(n1838) );
  CLKBUFX2TS U1193 ( .A(n1838), .Y(n1713) );
  AOI22X1TS U1194 ( .A0(destinationAddressIn_NORTH[3]), .A1(n671), .B0(n1713), 
        .B1(n645), .Y(n655) );
  CLKBUFX2TS U1195 ( .A(destinationAddressIn_WEST[3]), .Y(n1714) );
  CLKBUFX2TS U1196 ( .A(n1714), .Y(n1775) );
  AOI22X1TS U1197 ( .A0(destinationAddressIn_SOUTH[3]), .A1(n785), .B0(n1775), 
        .B1(n667), .Y(n654) );
  AOI22X1TS U1198 ( .A0(\destinationAddressbuffer[2][3] ), .A1(n673), .B0(
        \destinationAddressbuffer[0][3] ), .B1(n672), .Y(n650) );
  AOI22X1TS U1199 ( .A0(\destinationAddressbuffer[6][3] ), .A1(n675), .B0(
        \destinationAddressbuffer[4][3] ), .B1(n674), .Y(n649) );
  AOI22X1TS U1200 ( .A0(\destinationAddressbuffer[3][3] ), .A1(n677), .B0(
        \destinationAddressbuffer[1][3] ), .B1(n676), .Y(n648) );
  AOI22X1TS U1201 ( .A0(\destinationAddressbuffer[7][3] ), .A1(n646), .B0(
        \destinationAddressbuffer[5][3] ), .B1(n678), .Y(n647) );
  NAND4XLTS U1202 ( .A(n650), .B(n649), .C(n648), .D(n647), .Y(n651) );
  AOI22X1TS U1203 ( .A0(destinationAddressOut[3]), .A1(n757), .B0(n1901), .B1(
        n651), .Y(n653) );
  AOI22X1TS U1204 ( .A0(destinationAddressIn_EAST[4]), .A1(n746), .B0(n656), 
        .B1(n667), .Y(n666) );
  AOI22X1TS U1205 ( .A0(destinationAddressIn_NORTH[4]), .A1(n671), .B0(n658), 
        .B1(n657), .Y(n665) );
  INVX2TS U1206 ( .A(n1902), .Y(n766) );
  CLKBUFX2TS U1207 ( .A(n766), .Y(n862) );
  AOI22X1TS U1208 ( .A0(\destinationAddressbuffer[2][4] ), .A1(n673), .B0(
        \destinationAddressbuffer[0][4] ), .B1(n672), .Y(n662) );
  AOI22X1TS U1209 ( .A0(\destinationAddressbuffer[6][4] ), .A1(n675), .B0(
        \destinationAddressbuffer[4][4] ), .B1(n674), .Y(n661) );
  AOI22X1TS U1210 ( .A0(\destinationAddressbuffer[3][4] ), .A1(n677), .B0(
        \destinationAddressbuffer[1][4] ), .B1(n676), .Y(n660) );
  CLKBUFX2TS U1211 ( .A(n750), .Y(n704) );
  AOI22X1TS U1212 ( .A0(\destinationAddressbuffer[7][4] ), .A1(n704), .B0(
        \destinationAddressbuffer[5][4] ), .B1(n678), .Y(n659) );
  NAND4XLTS U1213 ( .A(n662), .B(n661), .C(n660), .D(n659), .Y(n663) );
  AOI22X1TS U1214 ( .A0(destinationAddressOut[4]), .A1(n781), .B0(n862), .B1(
        n663), .Y(n664) );
  CLKBUFX2TS U1215 ( .A(n775), .Y(n762) );
  AOI22X1TS U1216 ( .A0(destinationAddressIn_EAST[5]), .A1(n762), .B0(n668), 
        .B1(n667), .Y(n687) );
  CLKBUFX2TS U1217 ( .A(n669), .Y(n747) );
  AOI22X1TS U1218 ( .A0(destinationAddressIn_NORTH[5]), .A1(n671), .B0(n670), 
        .B1(n747), .Y(n686) );
  AOI22X1TS U1219 ( .A0(\destinationAddressbuffer[2][5] ), .A1(n673), .B0(
        \destinationAddressbuffer[0][5] ), .B1(n672), .Y(n682) );
  AOI22X1TS U1220 ( .A0(\destinationAddressbuffer[6][5] ), .A1(n675), .B0(
        \destinationAddressbuffer[4][5] ), .B1(n674), .Y(n681) );
  AOI22X1TS U1221 ( .A0(\destinationAddressbuffer[3][5] ), .A1(n677), .B0(
        \destinationAddressbuffer[1][5] ), .B1(n676), .Y(n680) );
  AOI22X1TS U1222 ( .A0(\destinationAddressbuffer[7][5] ), .A1(n704), .B0(
        \destinationAddressbuffer[5][5] ), .B1(n678), .Y(n679) );
  NAND4XLTS U1223 ( .A(n682), .B(n681), .C(n680), .D(n679), .Y(n683) );
  AOI22X1TS U1224 ( .A0(destinationAddressOut[5]), .A1(n684), .B0(n862), .B1(
        n683), .Y(n685) );
  CLKBUFX2TS U1225 ( .A(n807), .Y(n727) );
  AOI22X1TS U1226 ( .A0(destinationAddressIn_EAST[6]), .A1(n762), .B0(n688), 
        .B1(n727), .Y(n701) );
  CLKBUFX2TS U1227 ( .A(n689), .Y(n806) );
  CLKBUFX2TS U1228 ( .A(n806), .Y(n730) );
  AOI22X1TS U1229 ( .A0(destinationAddressIn_NORTH[6]), .A1(n730), .B0(n690), 
        .B1(n747), .Y(n700) );
  CLKBUFX2TS U1230 ( .A(n691), .Y(n808) );
  CLKBUFX2TS U1231 ( .A(n808), .Y(n733) );
  AOI22X1TS U1232 ( .A0(\destinationAddressbuffer[2][6] ), .A1(n716), .B0(
        \destinationAddressbuffer[0][6] ), .B1(n733), .Y(n697) );
  CLKBUFX2TS U1233 ( .A(n692), .Y(n810) );
  CLKBUFX2TS U1234 ( .A(n810), .Y(n734) );
  AOI22X1TS U1235 ( .A0(\destinationAddressbuffer[6][6] ), .A1(n717), .B0(
        \destinationAddressbuffer[4][6] ), .B1(n734), .Y(n696) );
  CLKBUFX2TS U1236 ( .A(n693), .Y(n812) );
  CLKBUFX2TS U1237 ( .A(n812), .Y(n735) );
  AOI22X1TS U1238 ( .A0(\destinationAddressbuffer[3][6] ), .A1(n718), .B0(
        \destinationAddressbuffer[1][6] ), .B1(n735), .Y(n695) );
  CLKBUFX2TS U1239 ( .A(n856), .Y(n825) );
  CLKBUFX2TS U1240 ( .A(n825), .Y(n736) );
  AOI22X1TS U1241 ( .A0(\destinationAddressbuffer[7][6] ), .A1(n704), .B0(
        \destinationAddressbuffer[5][6] ), .B1(n736), .Y(n694) );
  NAND4XLTS U1242 ( .A(n697), .B(n696), .C(n695), .D(n694), .Y(n698) );
  AOI22X1TS U1243 ( .A0(destinationAddressOut[6]), .A1(n781), .B0(n862), .B1(
        n698), .Y(n699) );
  AOI22X1TS U1244 ( .A0(destinationAddressIn_EAST[7]), .A1(n824), .B0(n702), 
        .B1(n727), .Y(n712) );
  AOI22X1TS U1245 ( .A0(destinationAddressIn_NORTH[7]), .A1(n730), .B0(n703), 
        .B1(n763), .Y(n711) );
  CLKBUFX2TS U1246 ( .A(n766), .Y(n756) );
  AOI22X1TS U1247 ( .A0(\destinationAddressbuffer[2][7] ), .A1(n716), .B0(
        \destinationAddressbuffer[0][7] ), .B1(n733), .Y(n708) );
  AOI22X1TS U1248 ( .A0(\destinationAddressbuffer[6][7] ), .A1(n717), .B0(
        \destinationAddressbuffer[4][7] ), .B1(n734), .Y(n707) );
  AOI22X1TS U1249 ( .A0(\destinationAddressbuffer[3][7] ), .A1(n718), .B0(
        \destinationAddressbuffer[1][7] ), .B1(n735), .Y(n706) );
  AOI22X1TS U1250 ( .A0(\destinationAddressbuffer[7][7] ), .A1(n704), .B0(
        \destinationAddressbuffer[5][7] ), .B1(n736), .Y(n705) );
  NAND4XLTS U1251 ( .A(n708), .B(n707), .C(n706), .D(n705), .Y(n709) );
  AOI22X1TS U1252 ( .A0(destinationAddressOut[7]), .A1(n521), .B0(n756), .B1(
        n709), .Y(n710) );
  AOI22X1TS U1253 ( .A0(destinationAddressIn_EAST[8]), .A1(n746), .B0(n713), 
        .B1(n727), .Y(n726) );
  AOI22X1TS U1254 ( .A0(n715), .A1(n730), .B0(n714), .B1(n747), .Y(n725) );
  CLKBUFX2TS U1255 ( .A(n716), .Y(n809) );
  AOI22X1TS U1256 ( .A0(\destinationAddressbuffer[2][8] ), .A1(n809), .B0(
        \destinationAddressbuffer[0][8] ), .B1(n733), .Y(n722) );
  CLKBUFX2TS U1257 ( .A(n717), .Y(n811) );
  AOI22X1TS U1258 ( .A0(\destinationAddressbuffer[6][8] ), .A1(n811), .B0(
        \destinationAddressbuffer[4][8] ), .B1(n734), .Y(n721) );
  CLKBUFX2TS U1259 ( .A(n718), .Y(n813) );
  AOI22X1TS U1260 ( .A0(\destinationAddressbuffer[3][8] ), .A1(n813), .B0(
        \destinationAddressbuffer[1][8] ), .B1(n735), .Y(n720) );
  AOI22X1TS U1261 ( .A0(\destinationAddressbuffer[7][8] ), .A1(n814), .B0(
        \destinationAddressbuffer[5][8] ), .B1(n736), .Y(n719) );
  NAND4XLTS U1262 ( .A(n722), .B(n721), .C(n720), .D(n719), .Y(n723) );
  AOI22X1TS U1263 ( .A0(destinationAddressOut[8]), .A1(n757), .B0(n756), .B1(
        n723), .Y(n724) );
  AOI22X1TS U1264 ( .A0(destinationAddressIn_EAST[9]), .A1(n762), .B0(n728), 
        .B1(n727), .Y(n744) );
  AOI22X1TS U1265 ( .A0(n731), .A1(n730), .B0(n729), .B1(n763), .Y(n743) );
  INVX2TS U1266 ( .A(n732), .Y(n841) );
  AOI22X1TS U1267 ( .A0(\destinationAddressbuffer[2][9] ), .A1(n809), .B0(
        \destinationAddressbuffer[0][9] ), .B1(n733), .Y(n740) );
  AOI22X1TS U1268 ( .A0(\destinationAddressbuffer[6][9] ), .A1(n811), .B0(
        \destinationAddressbuffer[4][9] ), .B1(n734), .Y(n739) );
  AOI22X1TS U1269 ( .A0(\destinationAddressbuffer[3][9] ), .A1(n813), .B0(
        \destinationAddressbuffer[1][9] ), .B1(n735), .Y(n738) );
  AOI22X1TS U1270 ( .A0(\destinationAddressbuffer[7][9] ), .A1(n814), .B0(
        \destinationAddressbuffer[5][9] ), .B1(n736), .Y(n737) );
  NAND4XLTS U1271 ( .A(n740), .B(n739), .C(n738), .D(n737), .Y(n741) );
  AOI22X1TS U1272 ( .A0(destinationAddressOut[9]), .A1(n841), .B0(n756), .B1(
        n741), .Y(n742) );
  CLKBUFX2TS U1273 ( .A(n807), .Y(n786) );
  AOI22X1TS U1274 ( .A0(destinationAddressIn_EAST[10]), .A1(n746), .B0(n745), 
        .B1(n786), .Y(n760) );
  CLKBUFX2TS U1275 ( .A(n806), .Y(n787) );
  AOI22X1TS U1276 ( .A0(n749), .A1(n787), .B0(n748), .B1(n747), .Y(n759) );
  CLKBUFX2TS U1277 ( .A(n809), .Y(n788) );
  CLKBUFX2TS U1278 ( .A(n808), .Y(n789) );
  AOI22X1TS U1279 ( .A0(\destinationAddressbuffer[2][10] ), .A1(n788), .B0(
        \destinationAddressbuffer[0][10] ), .B1(n789), .Y(n754) );
  CLKBUFX2TS U1280 ( .A(n811), .Y(n790) );
  CLKBUFX2TS U1281 ( .A(n810), .Y(n791) );
  AOI22X1TS U1282 ( .A0(\destinationAddressbuffer[6][10] ), .A1(n790), .B0(
        \destinationAddressbuffer[4][10] ), .B1(n791), .Y(n753) );
  CLKBUFX2TS U1283 ( .A(n813), .Y(n792) );
  CLKBUFX2TS U1284 ( .A(n812), .Y(n793) );
  AOI22X1TS U1285 ( .A0(\destinationAddressbuffer[3][10] ), .A1(n792), .B0(
        \destinationAddressbuffer[1][10] ), .B1(n793), .Y(n752) );
  CLKBUFX2TS U1286 ( .A(n825), .Y(n795) );
  AOI22X1TS U1287 ( .A0(\destinationAddressbuffer[7][10] ), .A1(n750), .B0(
        \destinationAddressbuffer[5][10] ), .B1(n795), .Y(n751) );
  NAND4XLTS U1288 ( .A(n754), .B(n753), .C(n752), .D(n751), .Y(n755) );
  AOI22X1TS U1289 ( .A0(destinationAddressOut[10]), .A1(n757), .B0(n756), .B1(
        n755), .Y(n758) );
  AOI22X1TS U1290 ( .A0(destinationAddressIn_EAST[11]), .A1(n762), .B0(n761), 
        .B1(n786), .Y(n774) );
  AOI22X1TS U1291 ( .A0(n765), .A1(n787), .B0(n764), .B1(n763), .Y(n773) );
  CLKBUFX2TS U1292 ( .A(n766), .Y(n820) );
  AOI22X1TS U1293 ( .A0(\destinationAddressbuffer[2][11] ), .A1(n788), .B0(
        \destinationAddressbuffer[0][11] ), .B1(n789), .Y(n770) );
  AOI22X1TS U1294 ( .A0(\destinationAddressbuffer[6][11] ), .A1(n790), .B0(
        \destinationAddressbuffer[4][11] ), .B1(n791), .Y(n769) );
  AOI22X1TS U1295 ( .A0(\destinationAddressbuffer[3][11] ), .A1(n792), .B0(
        \destinationAddressbuffer[1][11] ), .B1(n793), .Y(n768) );
  AOI22X1TS U1296 ( .A0(\destinationAddressbuffer[7][11] ), .A1(n794), .B0(
        \destinationAddressbuffer[5][11] ), .B1(n795), .Y(n767) );
  NAND4XLTS U1297 ( .A(n770), .B(n769), .C(n768), .D(n767), .Y(n771) );
  AOI22X1TS U1298 ( .A0(destinationAddressOut[11]), .A1(n521), .B0(n820), .B1(
        n771), .Y(n772) );
  CLKBUFX2TS U1299 ( .A(dataIn_EAST[0]), .Y(n1457) );
  CLKBUFX2TS U1300 ( .A(n1457), .Y(n1106) );
  CLKBUFX2TS U1301 ( .A(n775), .Y(n845) );
  AOI22X1TS U1302 ( .A0(dataIn_SOUTH[0]), .A1(n785), .B0(n1106), .B1(n845), 
        .Y(n784) );
  CLKBUFX2TS U1303 ( .A(dataIn_WEST[0]), .Y(n1496) );
  CLKBUFX2TS U1304 ( .A(n1496), .Y(n1391) );
  AOI22X1TS U1305 ( .A0(dataIn_NORTH[0]), .A1(n787), .B0(n1391), .B1(n786), 
        .Y(n783) );
  AOI22X1TS U1306 ( .A0(\dataoutbuffer[0][0] ), .A1(n789), .B0(
        \dataoutbuffer[2][0] ), .B1(n788), .Y(n779) );
  AOI22X1TS U1307 ( .A0(\dataoutbuffer[4][0] ), .A1(n791), .B0(
        \dataoutbuffer[6][0] ), .B1(n790), .Y(n778) );
  AOI22X1TS U1308 ( .A0(\dataoutbuffer[1][0] ), .A1(n793), .B0(
        \dataoutbuffer[3][0] ), .B1(n792), .Y(n777) );
  AOI22X1TS U1309 ( .A0(\dataoutbuffer[5][0] ), .A1(n795), .B0(
        \dataoutbuffer[7][0] ), .B1(n855), .Y(n776) );
  NAND4XLTS U1310 ( .A(n779), .B(n778), .C(n777), .D(n776), .Y(n780) );
  AOI22X1TS U1311 ( .A0(dataOut[0]), .A1(n781), .B0(n820), .B1(n780), .Y(n782)
         );
  CLKBUFX2TS U1312 ( .A(dataIn_EAST[1]), .Y(n1465) );
  CLKBUFX2TS U1313 ( .A(n1465), .Y(n1112) );
  AOI22X1TS U1314 ( .A0(dataIn_SOUTH[1]), .A1(n785), .B0(n1112), .B1(n824), 
        .Y(n804) );
  CLKBUFX2TS U1315 ( .A(dataIn_WEST[1]), .Y(n1504) );
  CLKBUFX2TS U1316 ( .A(n1504), .Y(n1397) );
  AOI22X1TS U1317 ( .A0(dataIn_NORTH[1]), .A1(n787), .B0(n1397), .B1(n786), 
        .Y(n803) );
  AOI22X1TS U1318 ( .A0(\dataoutbuffer[0][1] ), .A1(n789), .B0(
        \dataoutbuffer[2][1] ), .B1(n788), .Y(n799) );
  AOI22X1TS U1319 ( .A0(\dataoutbuffer[4][1] ), .A1(n791), .B0(
        \dataoutbuffer[6][1] ), .B1(n790), .Y(n798) );
  AOI22X1TS U1320 ( .A0(\dataoutbuffer[1][1] ), .A1(n793), .B0(
        \dataoutbuffer[3][1] ), .B1(n792), .Y(n797) );
  AOI22X1TS U1321 ( .A0(\dataoutbuffer[5][1] ), .A1(n795), .B0(
        \dataoutbuffer[7][1] ), .B1(n794), .Y(n796) );
  NAND4XLTS U1322 ( .A(n799), .B(n798), .C(n797), .D(n796), .Y(n800) );
  AOI22X1TS U1323 ( .A0(dataOut[1]), .A1(n522), .B0(n820), .B1(n800), .Y(n802)
         );
  CLKBUFX2TS U1324 ( .A(dataIn_EAST[2]), .Y(n1471) );
  CLKBUFX2TS U1325 ( .A(n1471), .Y(n1342) );
  AOI22X1TS U1326 ( .A0(dataIn_SOUTH[2]), .A1(n805), .B0(n1342), .B1(n845), 
        .Y(n823) );
  CLKBUFX2TS U1327 ( .A(n806), .Y(n848) );
  CLKBUFX2TS U1328 ( .A(dataIn_WEST[2]), .Y(n1511) );
  CLKBUFX2TS U1329 ( .A(n1511), .Y(n1402) );
  CLKBUFX2TS U1330 ( .A(n807), .Y(n847) );
  AOI22X1TS U1331 ( .A0(dataIn_NORTH[2]), .A1(n848), .B0(n1402), .B1(n847), 
        .Y(n822) );
  CLKBUFX2TS U1332 ( .A(n808), .Y(n850) );
  CLKBUFX2TS U1333 ( .A(n809), .Y(n849) );
  AOI22X1TS U1334 ( .A0(\dataoutbuffer[0][2] ), .A1(n850), .B0(
        \dataoutbuffer[2][2] ), .B1(n849), .Y(n818) );
  CLKBUFX2TS U1335 ( .A(n810), .Y(n852) );
  CLKBUFX2TS U1336 ( .A(n811), .Y(n851) );
  AOI22X1TS U1337 ( .A0(\dataoutbuffer[4][2] ), .A1(n852), .B0(
        \dataoutbuffer[6][2] ), .B1(n851), .Y(n817) );
  CLKBUFX2TS U1338 ( .A(n812), .Y(n854) );
  CLKBUFX2TS U1339 ( .A(n813), .Y(n853) );
  AOI22X1TS U1340 ( .A0(\dataoutbuffer[1][2] ), .A1(n854), .B0(
        \dataoutbuffer[3][2] ), .B1(n853), .Y(n816) );
  AOI22X1TS U1341 ( .A0(\dataoutbuffer[5][2] ), .A1(n825), .B0(
        \dataoutbuffer[7][2] ), .B1(n814), .Y(n815) );
  NAND4XLTS U1342 ( .A(n818), .B(n817), .C(n816), .D(n815), .Y(n819) );
  AOI22X1TS U1343 ( .A0(dataOut[2]), .A1(n841), .B0(n820), .B1(n819), .Y(n821)
         );
  INVX2TS U1344 ( .A(n10), .Y(n863) );
  CLKBUFX2TS U1345 ( .A(dataIn_EAST[3]), .Y(n1477) );
  CLKBUFX2TS U1346 ( .A(n1477), .Y(n1348) );
  AOI22X1TS U1347 ( .A0(dataIn_SOUTH[3]), .A1(n846), .B0(n1348), .B1(n824), 
        .Y(n833) );
  CLKBUFX2TS U1348 ( .A(dataIn_WEST[3]), .Y(n1519) );
  CLKBUFX2TS U1349 ( .A(n1519), .Y(n1407) );
  AOI22X1TS U1350 ( .A0(dataIn_NORTH[3]), .A1(n848), .B0(n1407), .B1(n847), 
        .Y(n832) );
  AOI22X1TS U1351 ( .A0(\dataoutbuffer[0][3] ), .A1(n850), .B0(
        \dataoutbuffer[2][3] ), .B1(n849), .Y(n829) );
  AOI22X1TS U1352 ( .A0(\dataoutbuffer[4][3] ), .A1(n852), .B0(
        \dataoutbuffer[6][3] ), .B1(n851), .Y(n828) );
  AOI22X1TS U1353 ( .A0(\dataoutbuffer[1][3] ), .A1(n854), .B0(
        \dataoutbuffer[3][3] ), .B1(n853), .Y(n827) );
  AOI22X1TS U1354 ( .A0(\dataoutbuffer[5][3] ), .A1(n825), .B0(
        \dataoutbuffer[7][3] ), .B1(n834), .Y(n826) );
  NAND4XLTS U1355 ( .A(n829), .B(n828), .C(n827), .D(n826), .Y(n830) );
  AOI22X1TS U1356 ( .A0(dataOut[3]), .A1(n841), .B0(n840), .B1(n830), .Y(n831)
         );
  CLKBUFX2TS U1357 ( .A(dataIn_EAST[4]), .Y(n1482) );
  CLKBUFX2TS U1358 ( .A(n1482), .Y(n1352) );
  AOI22X1TS U1359 ( .A0(dataIn_SOUTH[4]), .A1(n846), .B0(n1352), .B1(n845), 
        .Y(n844) );
  CLKBUFX2TS U1360 ( .A(dataIn_WEST[4]), .Y(n1526) );
  CLKBUFX2TS U1361 ( .A(n1526), .Y(n1411) );
  AOI22X1TS U1362 ( .A0(dataIn_NORTH[4]), .A1(n848), .B0(n1411), .B1(n847), 
        .Y(n843) );
  AOI22X1TS U1363 ( .A0(\dataoutbuffer[0][4] ), .A1(n850), .B0(
        \dataoutbuffer[2][4] ), .B1(n849), .Y(n838) );
  AOI22X1TS U1364 ( .A0(\dataoutbuffer[4][4] ), .A1(n852), .B0(
        \dataoutbuffer[6][4] ), .B1(n851), .Y(n837) );
  AOI22X1TS U1365 ( .A0(\dataoutbuffer[1][4] ), .A1(n854), .B0(
        \dataoutbuffer[3][4] ), .B1(n853), .Y(n836) );
  AOI22X1TS U1366 ( .A0(\dataoutbuffer[5][4] ), .A1(n856), .B0(
        \dataoutbuffer[7][4] ), .B1(n834), .Y(n835) );
  NAND4XLTS U1367 ( .A(n838), .B(n837), .C(n836), .D(n835), .Y(n839) );
  AOI22X1TS U1368 ( .A0(dataOut[4]), .A1(n841), .B0(n840), .B1(n839), .Y(n842)
         );
  CLKBUFX2TS U1369 ( .A(dataIn_EAST[5]), .Y(n1490) );
  CLKBUFX2TS U1370 ( .A(n1490), .Y(n1360) );
  AOI22X1TS U1371 ( .A0(dataIn_SOUTH[5]), .A1(n846), .B0(n1360), .B1(n845), 
        .Y(n866) );
  CLKBUFX2TS U1372 ( .A(dataIn_WEST[5]), .Y(n1535) );
  CLKBUFX2TS U1373 ( .A(n1535), .Y(n1418) );
  AOI22X1TS U1374 ( .A0(dataIn_NORTH[5]), .A1(n848), .B0(n1418), .B1(n847), 
        .Y(n865) );
  AOI22X1TS U1375 ( .A0(\dataoutbuffer[0][5] ), .A1(n850), .B0(
        \dataoutbuffer[2][5] ), .B1(n849), .Y(n860) );
  AOI22X1TS U1376 ( .A0(\dataoutbuffer[4][5] ), .A1(n852), .B0(
        \dataoutbuffer[6][5] ), .B1(n851), .Y(n859) );
  AOI22X1TS U1377 ( .A0(\dataoutbuffer[1][5] ), .A1(n854), .B0(
        \dataoutbuffer[3][5] ), .B1(n853), .Y(n858) );
  AOI22X1TS U1378 ( .A0(\dataoutbuffer[5][5] ), .A1(n856), .B0(
        \dataoutbuffer[7][5] ), .B1(n855), .Y(n857) );
  NAND4XLTS U1379 ( .A(n860), .B(n859), .C(n858), .D(n857), .Y(n861) );
  AOI22X1TS U1380 ( .A0(dataOut[5]), .A1(n522), .B0(n862), .B1(n861), .Y(n864)
         );
  INVX2TS U1381 ( .A(n949), .Y(n1750) );
  INVX2TS U1382 ( .A(n1503), .Y(n1525) );
  AOI22X1TS U1383 ( .A0(n1750), .A1(n1525), .B0(n1652), .B1(
        \requesterAddressbuffer[7][0] ), .Y(n870) );
  INVX2TS U1384 ( .A(n867), .Y(n1512) );
  CLKBUFX2TS U1385 ( .A(n1026), .Y(n921) );
  AOI22X1TS U1386 ( .A0(n1512), .A1(n951), .B0(n1645), .B1(n921), .Y(n869) );
  CLKBUFX2TS U1387 ( .A(requesterAddressIn_SOUTH[0]), .Y(n924) );
  CLKBUFX2TS U1388 ( .A(n999), .Y(n952) );
  AOI22X1TS U1389 ( .A0(n872), .A1(n924), .B0(n1537), .B1(n952), .Y(n868) );
  INVX2TS U1390 ( .A(n1503), .Y(n1644) );
  INVX2TS U1391 ( .A(n1495), .Y(n1534) );
  AOI22X1TS U1392 ( .A0(n1644), .A1(n1635), .B0(n1534), .B1(
        \requesterAddressbuffer[7][1] ), .Y(n875) );
  INVX2TS U1393 ( .A(n880), .Y(n1631) );
  CLKBUFX2TS U1394 ( .A(n1032), .Y(n929) );
  AOI22X1TS U1395 ( .A0(n1527), .A1(n958), .B0(n1631), .B1(n929), .Y(n874) );
  CLKBUFX2TS U1396 ( .A(requesterAddressIn_SOUTH[1]), .Y(n932) );
  CLKBUFX2TS U1397 ( .A(n1006), .Y(n959) );
  AOI22X1TS U1398 ( .A0(n872), .A1(n932), .B0(n871), .B1(n959), .Y(n873) );
  AOI22X1TS U1399 ( .A0(n1654), .A1(n1643), .B0(n1534), .B1(
        \requesterAddressbuffer[7][2] ), .Y(n878) );
  CLKBUFX2TS U1400 ( .A(n1036), .Y(n936) );
  AOI22X1TS U1401 ( .A0(n1646), .A1(n964), .B0(n26), .B1(n936), .Y(n877) );
  CLKBUFX2TS U1402 ( .A(requesterAddressIn_SOUTH[2]), .Y(n1037) );
  CLKBUFX2TS U1403 ( .A(n1012), .Y(n967) );
  AOI22X1TS U1404 ( .A0(n50), .A1(n1037), .B0(n1537), .B1(n967), .Y(n876) );
  INVX2TS U1405 ( .A(n879), .Y(n1642) );
  AOI22X1TS U1406 ( .A0(n1525), .A1(n1653), .B0(n1642), .B1(
        \requesterAddressbuffer[7][3] ), .Y(n883) );
  INVX2TS U1407 ( .A(n880), .Y(n1655) );
  CLKBUFX2TS U1408 ( .A(n1044), .Y(n944) );
  AOI22X1TS U1409 ( .A0(n1527), .A1(n973), .B0(n1655), .B1(n944), .Y(n882) );
  CLKBUFX2TS U1410 ( .A(requesterAddressIn_SOUTH[3]), .Y(n1046) );
  CLKBUFX2TS U1411 ( .A(n1021), .Y(n974) );
  AOI22X1TS U1412 ( .A0(n1530), .A1(n1046), .B0(n35), .B1(n974), .Y(n881) );
  INVX2TS U1413 ( .A(n949), .Y(n1806) );
  AOI22X1TS U1414 ( .A0(n1806), .A1(n1662), .B0(n1680), .B1(
        \requesterAddressbuffer[6][0] ), .Y(n886) );
  INVX2TS U1415 ( .A(n1470), .Y(n1669) );
  AOI22X1TS U1416 ( .A0(n922), .A1(n1681), .B0(n921), .B1(n1669), .Y(n885) );
  AOI22X1TS U1417 ( .A0(n924), .A1(n1460), .B0(n952), .B1(n1461), .Y(n884) );
  INVX2TS U1418 ( .A(n956), .Y(n1726) );
  INVX2TS U1419 ( .A(n895), .Y(n1668) );
  INVX2TS U1420 ( .A(n1456), .Y(n1489) );
  AOI22X1TS U1421 ( .A0(n1726), .A1(n1668), .B0(n1489), .B1(
        \requesterAddressbuffer[6][1] ), .Y(n890) );
  INVX2TS U1422 ( .A(n1470), .Y(n1675) );
  AOI22X1TS U1423 ( .A0(n930), .A1(n1483), .B0(n929), .B1(n1675), .Y(n889) );
  INVX2TS U1424 ( .A(n899), .Y(n1485) );
  AOI22X1TS U1425 ( .A0(n932), .A1(n1485), .B0(n959), .B1(n87), .Y(n888) );
  INVX2TS U1426 ( .A(n963), .Y(n1734) );
  INVX2TS U1427 ( .A(n895), .Y(n1674) );
  AOI22X1TS U1428 ( .A0(n1734), .A1(n1674), .B0(n1489), .B1(
        \requesterAddressbuffer[6][2] ), .Y(n894) );
  AOI22X1TS U1429 ( .A0(n937), .A1(n1458), .B0(n936), .B1(n898), .Y(n893) );
  AOI22X1TS U1430 ( .A0(requesterAddressIn_SOUTH[2]), .A1(n91), .B0(n967), 
        .B1(n891), .Y(n892) );
  INVX2TS U1431 ( .A(n971), .Y(n1742) );
  INVX2TS U1432 ( .A(n896), .Y(n1673) );
  AOI22X1TS U1433 ( .A0(n1742), .A1(n1662), .B0(n1673), .B1(
        \requesterAddressbuffer[6][3] ), .Y(n902) );
  INVX2TS U1434 ( .A(n897), .Y(n1483) );
  AOI22X1TS U1435 ( .A0(n945), .A1(n1483), .B0(n944), .B1(n898), .Y(n901) );
  INVX2TS U1436 ( .A(n899), .Y(n1676) );
  AOI22X1TS U1437 ( .A0(requesterAddressIn_SOUTH[3]), .A1(n1676), .B0(n974), 
        .B1(n1664), .Y(n900) );
  AOI22X1TS U1438 ( .A0(n996), .A1(n1687), .B0(n1711), .B1(
        \requesterAddressbuffer[5][0] ), .Y(n906) );
  INVX2TS U1439 ( .A(n1434), .Y(n1698) );
  AOI22X1TS U1440 ( .A0(n922), .A1(n1715), .B0(n921), .B1(n1698), .Y(n905) );
  INVX2TS U1441 ( .A(n903), .Y(n1716) );
  AOI22X1TS U1442 ( .A0(n924), .A1(n1716), .B0(requesterAddressIn_NORTH[0]), 
        .B1(n1436), .Y(n904) );
  INVX2TS U1443 ( .A(n915), .Y(n1696) );
  AOI22X1TS U1444 ( .A0(n1635), .A1(n1696), .B0(n1451), .B1(
        \requesterAddressbuffer[5][1] ), .Y(n910) );
  INVX2TS U1445 ( .A(n1434), .Y(n1706) );
  AOI22X1TS U1446 ( .A0(n930), .A1(n248), .B0(n929), .B1(n1706), .Y(n909) );
  AOI22X1TS U1447 ( .A0(n932), .A1(n1691), .B0(requesterAddressIn_NORTH[1]), 
        .B1(n1692), .Y(n908) );
  AOI22X1TS U1448 ( .A0(n1643), .A1(n1687), .B0(n1451), .B1(
        \requesterAddressbuffer[5][2] ), .Y(n914) );
  AOI22X1TS U1449 ( .A0(n937), .A1(n1423), .B0(n936), .B1(n917), .Y(n913) );
  AOI22X1TS U1450 ( .A0(n1037), .A1(n1424), .B0(requesterAddressIn_NORTH[2]), 
        .B1(n911), .Y(n912) );
  INVX2TS U1451 ( .A(n915), .Y(n1712) );
  INVX2TS U1452 ( .A(n916), .Y(n1704) );
  AOI22X1TS U1453 ( .A0(n1653), .A1(n1712), .B0(n1704), .B1(
        \requesterAddressbuffer[5][3] ), .Y(n920) );
  AOI22X1TS U1454 ( .A0(n945), .A1(n239), .B0(n944), .B1(n917), .Y(n919) );
  AOI22X1TS U1455 ( .A0(n1046), .A1(n229), .B0(requesterAddressIn_NORTH[3]), 
        .B1(n1447), .Y(n918) );
  AOI22X1TS U1456 ( .A0(n996), .A1(n1720), .B0(n1740), .B1(
        \requesterAddressbuffer[4][0] ), .Y(n927) );
  INVX2TS U1457 ( .A(n1401), .Y(n1727) );
  AOI22X1TS U1458 ( .A0(n922), .A1(n1743), .B0(n921), .B1(n1727), .Y(n926) );
  INVX2TS U1459 ( .A(n923), .Y(n1412) );
  AOI22X1TS U1460 ( .A0(n924), .A1(n1736), .B0(requesterAddressIn_NORTH[0]), 
        .B1(n1412), .Y(n925) );
  INVX2TS U1461 ( .A(n956), .Y(n1857) );
  INVX2TS U1462 ( .A(n941), .Y(n1725) );
  INVX2TS U1463 ( .A(n1390), .Y(n1417) );
  AOI22X1TS U1464 ( .A0(n1857), .A1(n1725), .B0(n1417), .B1(
        \requesterAddressbuffer[4][1] ), .Y(n935) );
  INVX2TS U1465 ( .A(n1401), .Y(n1735) );
  AOI22X1TS U1466 ( .A0(n930), .A1(n303), .B0(n929), .B1(n1735), .Y(n934) );
  AOI22X1TS U1467 ( .A0(n932), .A1(n1413), .B0(requesterAddressIn_NORTH[1]), 
        .B1(n931), .Y(n933) );
  INVX2TS U1468 ( .A(n963), .Y(n1866) );
  AOI22X1TS U1469 ( .A0(n1866), .A1(n1720), .B0(n1417), .B1(
        \requesterAddressbuffer[4][2] ), .Y(n940) );
  AOI22X1TS U1470 ( .A0(n937), .A1(n1392), .B0(n936), .B1(n943), .Y(n939) );
  AOI22X1TS U1471 ( .A0(n1037), .A1(n1745), .B0(requesterAddressIn_NORTH[2]), 
        .B1(n1744), .Y(n938) );
  INVX2TS U1472 ( .A(n971), .Y(n1876) );
  INVX2TS U1473 ( .A(n941), .Y(n1741) );
  INVX2TS U1474 ( .A(n942), .Y(n1733) );
  AOI22X1TS U1475 ( .A0(n1876), .A1(n1741), .B0(n1733), .B1(
        \requesterAddressbuffer[4][3] ), .Y(n948) );
  AOI22X1TS U1476 ( .A0(n945), .A1(n292), .B0(n944), .B1(n943), .Y(n947) );
  AOI22X1TS U1477 ( .A0(n1046), .A1(n1729), .B0(requesterAddressIn_NORTH[3]), 
        .B1(n1412), .Y(n946) );
  INVX2TS U1478 ( .A(n949), .Y(n1847) );
  AOI22X1TS U1479 ( .A0(n1847), .A1(n1749), .B0(n1773), .B1(
        \requesterAddressbuffer[3][0] ), .Y(n955) );
  INVX2TS U1480 ( .A(n950), .Y(n1373) );
  AOI22X1TS U1481 ( .A0(n951), .A1(n1373), .B0(n997), .B1(n145), .Y(n954) );
  INVX2TS U1482 ( .A(n965), .Y(n1769) );
  AOI22X1TS U1483 ( .A0(n1000), .A1(n1769), .B0(n952), .B1(n1761), .Y(n953) );
  INVX2TS U1484 ( .A(n956), .Y(n1817) );
  INVX2TS U1485 ( .A(n972), .Y(n1757) );
  INVX2TS U1486 ( .A(n1364), .Y(n1385) );
  AOI22X1TS U1487 ( .A0(n1817), .A1(n1757), .B0(n1385), .B1(
        \requesterAddressbuffer[3][1] ), .Y(n962) );
  INVX2TS U1488 ( .A(n957), .Y(n1758) );
  AOI22X1TS U1489 ( .A0(n958), .A1(n131), .B0(n1005), .B1(n1758), .Y(n961) );
  INVX2TS U1490 ( .A(n965), .Y(n1777) );
  AOI22X1TS U1491 ( .A0(n1007), .A1(n1777), .B0(n959), .B1(n1365), .Y(n960) );
  INVX2TS U1492 ( .A(n963), .Y(n1827) );
  INVX2TS U1493 ( .A(n972), .Y(n1766) );
  AOI22X1TS U1494 ( .A0(n1827), .A1(n1766), .B0(n1385), .B1(
        \requesterAddressbuffer[3][2] ), .Y(n970) );
  AOI22X1TS U1495 ( .A0(n964), .A1(n1386), .B0(n1011), .B1(n1381), .Y(n969) );
  AOI22X1TS U1496 ( .A0(n1013), .A1(n124), .B0(n967), .B1(n966), .Y(n968) );
  INVX2TS U1497 ( .A(n971), .Y(n1837) );
  INVX2TS U1498 ( .A(n1364), .Y(n1765) );
  AOI22X1TS U1499 ( .A0(n1837), .A1(n1749), .B0(n1765), .B1(
        \requesterAddressbuffer[3][3] ), .Y(n977) );
  AOI22X1TS U1500 ( .A0(n973), .A1(n1373), .B0(n1019), .B1(n1774), .Y(n976) );
  AOI22X1TS U1501 ( .A0(n1022), .A1(n1769), .B0(n974), .B1(n1753), .Y(n975) );
  AOI22X1TS U1502 ( .A0(n1750), .A1(n1782), .B0(n1800), .B1(
        \requesterAddressbuffer[2][0] ), .Y(n981) );
  INVX2TS U1503 ( .A(n1341), .Y(n1790) );
  AOI22X1TS U1504 ( .A0(requesterAddressIn_WEST[0]), .A1(n1801), .B0(n997), 
        .B1(n1790), .Y(n980) );
  INVX2TS U1505 ( .A(n978), .Y(n1802) );
  AOI22X1TS U1506 ( .A0(n1000), .A1(n1802), .B0(n999), .B1(n1785), .Y(n979) );
  INVX2TS U1507 ( .A(n989), .Y(n1789) );
  INVX2TS U1508 ( .A(n982), .Y(n1359) );
  AOI22X1TS U1509 ( .A0(n1857), .A1(n1789), .B0(n1359), .B1(
        \requesterAddressbuffer[2][1] ), .Y(n985) );
  INVX2TS U1510 ( .A(n1341), .Y(n1796) );
  AOI22X1TS U1511 ( .A0(requesterAddressIn_WEST[1]), .A1(n1353), .B0(n1005), 
        .B1(n1796), .Y(n984) );
  AOI22X1TS U1512 ( .A0(n1007), .A1(n1784), .B0(n1006), .B1(n1343), .Y(n983)
         );
  INVX2TS U1513 ( .A(n989), .Y(n1795) );
  AOI22X1TS U1514 ( .A0(n1866), .A1(n1795), .B0(n1359), .B1(
        \requesterAddressbuffer[2][2] ), .Y(n988) );
  AOI22X1TS U1515 ( .A0(requesterAddressIn_WEST[2]), .A1(n1107), .B0(n1011), 
        .B1(n991), .Y(n987) );
  AOI22X1TS U1516 ( .A0(n1013), .A1(n1108), .B0(n1012), .B1(n1337), .Y(n986)
         );
  INVX2TS U1517 ( .A(n1605), .Y(n1794) );
  AOI22X1TS U1518 ( .A0(n1876), .A1(n1782), .B0(n1794), .B1(
        \requesterAddressbuffer[2][3] ), .Y(n995) );
  INVX2TS U1519 ( .A(n990), .Y(n1353) );
  AOI22X1TS U1520 ( .A0(requesterAddressIn_WEST[3]), .A1(n1353), .B0(n1019), 
        .B1(n991), .Y(n994) );
  AOI22X1TS U1521 ( .A0(n1022), .A1(n195), .B0(n1021), .B1(n992), .Y(n993) );
  INVX2TS U1522 ( .A(n1081), .Y(n1095) );
  AOI22X1TS U1523 ( .A0(n996), .A1(n1095), .B0(n1835), .B1(
        \requesterAddressbuffer[1][0] ), .Y(n1003) );
  INVX2TS U1524 ( .A(n1086), .Y(n1819) );
  AOI22X1TS U1525 ( .A0(requesterAddressIn_WEST[0]), .A1(n1839), .B0(n997), 
        .B1(n1819), .Y(n1002) );
  INVX2TS U1526 ( .A(n998), .Y(n1841) );
  AOI22X1TS U1527 ( .A0(n1000), .A1(n1841), .B0(n999), .B1(n1812), .Y(n1001)
         );
  INVX2TS U1528 ( .A(n1081), .Y(n1826) );
  INVX2TS U1529 ( .A(n1004), .Y(n1102) );
  AOI22X1TS U1530 ( .A0(n1726), .A1(n1826), .B0(n1102), .B1(
        \requesterAddressbuffer[1][1] ), .Y(n1010) );
  INVX2TS U1531 ( .A(n1086), .Y(n1829) );
  AOI22X1TS U1532 ( .A0(requesterAddressIn_WEST[1]), .A1(n1096), .B0(n1005), 
        .B1(n1829), .Y(n1009) );
  AOI22X1TS U1533 ( .A0(n1007), .A1(n1810), .B0(n1006), .B1(n1087), .Y(n1008)
         );
  AOI22X1TS U1534 ( .A0(n1734), .A1(n1836), .B0(n1102), .B1(
        \requesterAddressbuffer[1][2] ), .Y(n1016) );
  AOI22X1TS U1535 ( .A0(requesterAddressIn_WEST[2]), .A1(n1076), .B0(n1011), 
        .B1(n1018), .Y(n1015) );
  AOI22X1TS U1536 ( .A0(n1013), .A1(n1077), .B0(n1012), .B1(n1082), .Y(n1014)
         );
  INVX2TS U1537 ( .A(n1618), .Y(n1825) );
  AOI22X1TS U1538 ( .A0(n1742), .A1(n1095), .B0(n1825), .B1(
        \requesterAddressbuffer[1][3] ), .Y(n1025) );
  INVX2TS U1539 ( .A(n1017), .Y(n1096) );
  AOI22X1TS U1540 ( .A0(requesterAddressIn_WEST[3]), .A1(n1096), .B0(n1019), 
        .B1(n1018), .Y(n1024) );
  AOI22X1TS U1541 ( .A0(n1022), .A1(n346), .B0(n1021), .B1(n1020), .Y(n1023)
         );
  AOI22X1TS U1542 ( .A0(readRequesterAddress[0]), .A1(n1846), .B0(n1874), .B1(
        \requesterAddressbuffer[0][0] ), .Y(n1030) );
  INVX2TS U1543 ( .A(n1058), .Y(n1858) );
  AOI22X1TS U1544 ( .A0(requesterAddressIn_WEST[0]), .A1(n1877), .B0(n1026), 
        .B1(n1858), .Y(n1029) );
  INVX2TS U1545 ( .A(n1027), .Y(n1067) );
  AOI22X1TS U1546 ( .A0(requesterAddressIn_SOUTH[0]), .A1(n1870), .B0(
        requesterAddressIn_NORTH[0]), .B1(n1067), .Y(n1028) );
  INVX2TS U1547 ( .A(n9), .Y(n1856) );
  INVX2TS U1548 ( .A(n1031), .Y(n1072) );
  AOI22X1TS U1549 ( .A0(n1817), .A1(n1856), .B0(n1072), .B1(
        \requesterAddressbuffer[0][1] ), .Y(n1035) );
  INVX2TS U1550 ( .A(n1058), .Y(n1867) );
  AOI22X1TS U1551 ( .A0(requesterAddressIn_WEST[1]), .A1(n1066), .B0(n1032), 
        .B1(n1867), .Y(n1034) );
  AOI22X1TS U1552 ( .A0(requesterAddressIn_SOUTH[1]), .A1(n1068), .B0(
        requesterAddressIn_NORTH[1]), .B1(n1067), .Y(n1033) );
  INVX2TS U1553 ( .A(n9), .Y(n1865) );
  AOI22X1TS U1554 ( .A0(n1827), .A1(n1865), .B0(n1072), .B1(
        \requesterAddressbuffer[0][2] ), .Y(n1040) );
  AOI22X1TS U1555 ( .A0(requesterAddressIn_WEST[2]), .A1(n1050), .B0(n1036), 
        .B1(n1043), .Y(n1039) );
  AOI22X1TS U1556 ( .A0(n1037), .A1(n1881), .B0(requesterAddressIn_NORTH[2]), 
        .B1(n1879), .Y(n1038) );
  INVX2TS U1557 ( .A(n9), .Y(n1875) );
  INVX2TS U1558 ( .A(n1041), .Y(n1864) );
  AOI22X1TS U1559 ( .A0(n1837), .A1(n1875), .B0(n1864), .B1(
        \requesterAddressbuffer[0][3] ), .Y(n1049) );
  INVX2TS U1560 ( .A(n1042), .Y(n1066) );
  AOI22X1TS U1561 ( .A0(requesterAddressIn_WEST[3]), .A1(n1066), .B0(n1044), 
        .B1(n1043), .Y(n1048) );
  INVX2TS U1562 ( .A(n1045), .Y(n1852) );
  AOI22X1TS U1563 ( .A0(n1046), .A1(n1852), .B0(requesterAddressIn_NORTH[3]), 
        .B1(n1051), .Y(n1047) );
  INVX2TS U1564 ( .A(n1041), .Y(n1062) );
  AOI21X1TS U1565 ( .A0(n1062), .A1(\dataoutbuffer[0][0] ), .B0(n1856), .Y(
        n1054) );
  AOI22X1TS U1566 ( .A0(n1050), .A1(n1391), .B0(n1858), .B1(n1106), .Y(n1053)
         );
  CLKBUFX2TS U1567 ( .A(dataIn_SOUTH[0]), .Y(n1499) );
  AOI22X1TS U1568 ( .A0(n1852), .A1(n1499), .B0(n1051), .B1(dataIn_NORTH[0]), 
        .Y(n1052) );
  AOI21X1TS U1569 ( .A0(n1062), .A1(\dataoutbuffer[0][1] ), .B0(n1865), .Y(
        n1057) );
  AOI22X1TS U1570 ( .A0(n419), .A1(n1397), .B0(n1867), .B1(n1112), .Y(n1056)
         );
  CLKBUFX2TS U1571 ( .A(dataIn_SOUTH[1]), .Y(n1507) );
  AOI22X1TS U1572 ( .A0(n1870), .A1(n1507), .B0(n402), .B1(dataIn_NORTH[1]), 
        .Y(n1055) );
  AOI21X1TS U1573 ( .A0(n1062), .A1(\dataoutbuffer[0][2] ), .B0(n1875), .Y(
        n1061) );
  AOI22X1TS U1574 ( .A0(n1066), .A1(n1402), .B0(n391), .B1(n1342), .Y(n1060)
         );
  CLKBUFX2TS U1575 ( .A(dataIn_SOUTH[2]), .Y(n1514) );
  AOI22X1TS U1576 ( .A0(n1881), .A1(n1514), .B0(n1067), .B1(dataIn_NORTH[2]), 
        .Y(n1059) );
  AOI21X1TS U1577 ( .A0(n1062), .A1(\dataoutbuffer[0][3] ), .B0(n1856), .Y(
        n1065) );
  AOI22X1TS U1578 ( .A0(n1848), .A1(n1407), .B0(n1858), .B1(n1348), .Y(n1064)
         );
  CLKBUFX2TS U1579 ( .A(dataIn_SOUTH[3]), .Y(n1521) );
  AOI22X1TS U1580 ( .A0(n428), .A1(n1521), .B0(n1850), .B1(dataIn_NORTH[3]), 
        .Y(n1063) );
  AOI21X1TS U1581 ( .A0(n1072), .A1(\dataoutbuffer[0][4] ), .B0(n1865), .Y(
        n1071) );
  AOI22X1TS U1582 ( .A0(n1066), .A1(n1411), .B0(n1867), .B1(n1352), .Y(n1070)
         );
  CLKBUFX2TS U1583 ( .A(dataIn_SOUTH[4]), .Y(n1529) );
  AOI22X1TS U1584 ( .A0(n1068), .A1(n1529), .B0(n1067), .B1(dataIn_NORTH[4]), 
        .Y(n1069) );
  AOI21X1TS U1585 ( .A0(n1072), .A1(\dataoutbuffer[0][5] ), .B0(n1875), .Y(
        n1075) );
  AOI22X1TS U1586 ( .A0(n419), .A1(n1418), .B0(n391), .B1(n1360), .Y(n1074) );
  CLKBUFX2TS U1587 ( .A(dataIn_SOUTH[5]), .Y(n1538) );
  AOI22X1TS U1588 ( .A0(n1852), .A1(n1538), .B0(n402), .B1(dataIn_NORTH[5]), 
        .Y(n1073) );
  INVX2TS U1589 ( .A(n1618), .Y(n1091) );
  AOI21X1TS U1590 ( .A0(n1091), .A1(\dataoutbuffer[1][0] ), .B0(n1095), .Y(
        n1080) );
  AOI22X1TS U1591 ( .A0(n1076), .A1(dataIn_WEST[0]), .B0(n1819), .B1(n1106), 
        .Y(n1079) );
  CLKBUFX2TS U1592 ( .A(dataIn_NORTH[0]), .Y(n1425) );
  CLKBUFX2TS U1593 ( .A(n1425), .Y(n1498) );
  CLKBUFX2TS U1594 ( .A(n1499), .Y(n1459) );
  AOI22X1TS U1595 ( .A0(n1082), .A1(n1498), .B0(n1077), .B1(n1459), .Y(n1078)
         );
  INVX2TS U1596 ( .A(n1081), .Y(n1816) );
  AOI21X1TS U1597 ( .A0(n1091), .A1(\dataoutbuffer[1][1] ), .B0(n1816), .Y(
        n1085) );
  AOI22X1TS U1598 ( .A0(n320), .A1(dataIn_WEST[1]), .B0(n1829), .B1(n1112), 
        .Y(n1084) );
  CLKBUFX2TS U1599 ( .A(dataIn_NORTH[1]), .Y(n1430) );
  CLKBUFX2TS U1600 ( .A(n1430), .Y(n1506) );
  CLKBUFX2TS U1601 ( .A(n1507), .Y(n1466) );
  AOI22X1TS U1602 ( .A0(n325), .A1(n1506), .B0(n353), .B1(n1466), .Y(n1083) );
  AOI21X1TS U1603 ( .A0(n1091), .A1(\dataoutbuffer[1][2] ), .B0(n1826), .Y(
        n1090) );
  AOI22X1TS U1604 ( .A0(n1096), .A1(dataIn_WEST[2]), .B0(n318), .B1(n1342), 
        .Y(n1089) );
  CLKBUFX2TS U1605 ( .A(dataIn_NORTH[2]), .Y(n1435) );
  CLKBUFX2TS U1606 ( .A(n1435), .Y(n1513) );
  CLKBUFX2TS U1607 ( .A(n1514), .Y(n1472) );
  AOI22X1TS U1608 ( .A0(n1087), .A1(n1513), .B0(n1097), .B1(n1472), .Y(n1088)
         );
  AOI21X1TS U1609 ( .A0(n1091), .A1(\dataoutbuffer[1][3] ), .B0(n1836), .Y(
        n1094) );
  AOI22X1TS U1610 ( .A0(n1808), .A1(dataIn_WEST[3]), .B0(n1819), .B1(n1348), 
        .Y(n1093) );
  CLKBUFX2TS U1611 ( .A(dataIn_NORTH[3]), .Y(n1441) );
  CLKBUFX2TS U1612 ( .A(n1441), .Y(n1520) );
  CLKBUFX2TS U1613 ( .A(n1521), .Y(n1478) );
  AOI22X1TS U1614 ( .A0(n325), .A1(n1520), .B0(n1810), .B1(n1478), .Y(n1092)
         );
  AOI21X1TS U1615 ( .A0(n1102), .A1(\dataoutbuffer[1][4] ), .B0(n1095), .Y(
        n1101) );
  AOI22X1TS U1616 ( .A0(n1096), .A1(dataIn_WEST[4]), .B0(n1829), .B1(n1352), 
        .Y(n1100) );
  CLKBUFX2TS U1617 ( .A(dataIn_NORTH[4]), .Y(n1446) );
  CLKBUFX2TS U1618 ( .A(n1446), .Y(n1528) );
  CLKBUFX2TS U1619 ( .A(n1529), .Y(n1484) );
  AOI22X1TS U1620 ( .A0(n1098), .A1(n1528), .B0(n1097), .B1(n1484), .Y(n1099)
         );
  AOI21X1TS U1621 ( .A0(n1102), .A1(\dataoutbuffer[1][5] ), .B0(n1816), .Y(
        n1105) );
  AOI22X1TS U1622 ( .A0(n320), .A1(dataIn_WEST[5]), .B0(n318), .B1(n1360), .Y(
        n1104) );
  CLKBUFX2TS U1623 ( .A(dataIn_NORTH[5]), .Y(n1452) );
  CLKBUFX2TS U1624 ( .A(n1452), .Y(n1536) );
  CLKBUFX2TS U1625 ( .A(n1538), .Y(n1491) );
  AOI22X1TS U1626 ( .A0(n324), .A1(n1536), .B0(n346), .B1(n1491), .Y(n1103) );
  INVX2TS U1627 ( .A(n1605), .Y(n1347) );
  AOI21X1TS U1628 ( .A0(n1347), .A1(\dataoutbuffer[2][0] ), .B0(n1789), .Y(
        n1111) );
  AOI22X1TS U1629 ( .A0(n1107), .A1(dataIn_WEST[0]), .B0(n1790), .B1(n1106), 
        .Y(n1110) );
  AOI22X1TS U1630 ( .A0(n1337), .A1(n1498), .B0(n1108), .B1(dataIn_SOUTH[0]), 
        .Y(n1109) );
  AOI21X1TS U1631 ( .A0(n1347), .A1(\dataoutbuffer[2][1] ), .B0(n1795), .Y(
        n1340) );
  AOI22X1TS U1632 ( .A0(n179), .A1(dataIn_WEST[1]), .B0(n1796), .B1(n1112), 
        .Y(n1339) );
  AOI22X1TS U1633 ( .A0(n182), .A1(n1506), .B0(n198), .B1(dataIn_SOUTH[1]), 
        .Y(n1338) );
  AOI21X1TS U1634 ( .A0(n1347), .A1(\dataoutbuffer[2][2] ), .B0(n177), .Y(
        n1346) );
  AOI22X1TS U1635 ( .A0(n1353), .A1(dataIn_WEST[2]), .B0(n176), .B1(n1342), 
        .Y(n1345) );
  AOI22X1TS U1636 ( .A0(n1343), .A1(n1513), .B0(n1354), .B1(dataIn_SOUTH[2]), 
        .Y(n1344) );
  AOI21X1TS U1637 ( .A0(n1347), .A1(\dataoutbuffer[2][3] ), .B0(n1789), .Y(
        n1351) );
  AOI22X1TS U1638 ( .A0(n1783), .A1(dataIn_WEST[3]), .B0(n1790), .B1(n1348), 
        .Y(n1350) );
  AOI22X1TS U1639 ( .A0(n183), .A1(n1520), .B0(n1784), .B1(dataIn_SOUTH[3]), 
        .Y(n1349) );
  AOI21X1TS U1640 ( .A0(n1359), .A1(\dataoutbuffer[2][4] ), .B0(n1795), .Y(
        n1358) );
  AOI22X1TS U1641 ( .A0(n1353), .A1(dataIn_WEST[4]), .B0(n1796), .B1(n1352), 
        .Y(n1357) );
  AOI22X1TS U1642 ( .A0(n1355), .A1(n1528), .B0(n1354), .B1(dataIn_SOUTH[4]), 
        .Y(n1356) );
  AOI21X1TS U1643 ( .A0(n1359), .A1(\dataoutbuffer[2][5] ), .B0(n177), .Y(
        n1363) );
  AOI22X1TS U1644 ( .A0(n179), .A1(dataIn_WEST[5]), .B0(n176), .B1(n1360), .Y(
        n1362) );
  AOI22X1TS U1645 ( .A0(n182), .A1(n1536), .B0(n195), .B1(dataIn_SOUTH[5]), 
        .Y(n1361) );
  INVX2TS U1646 ( .A(n169), .Y(n1377) );
  AOI21X1TS U1647 ( .A0(n1377), .A1(\dataoutbuffer[3][0] ), .B0(n1757), .Y(
        n1368) );
  AOI22X1TS U1648 ( .A0(n1373), .A1(dataIn_WEST[0]), .B0(n1767), .B1(
        dataIn_EAST[0]), .Y(n1367) );
  AOI22X1TS U1649 ( .A0(n1365), .A1(n1425), .B0(n1760), .B1(n1459), .Y(n1366)
         );
  AOI21X1TS U1650 ( .A0(n1377), .A1(\dataoutbuffer[3][1] ), .B0(n1766), .Y(
        n1372) );
  AOI22X1TS U1651 ( .A0(n141), .A1(dataIn_WEST[1]), .B0(n1758), .B1(
        dataIn_EAST[1]), .Y(n1371) );
  INVX2TS U1652 ( .A(n1369), .Y(n1761) );
  AOI22X1TS U1653 ( .A0(n1761), .A1(n1430), .B0(n1769), .B1(n1466), .Y(n1370)
         );
  AOI21X1TS U1654 ( .A0(n1377), .A1(\dataoutbuffer[3][2] ), .B0(n126), .Y(
        n1376) );
  AOI22X1TS U1655 ( .A0(n1373), .A1(dataIn_WEST[2]), .B0(n164), .B1(
        dataIn_EAST[2]), .Y(n1375) );
  AOI22X1TS U1656 ( .A0(n966), .A1(n1435), .B0(n1777), .B1(n1472), .Y(n1374)
         );
  AOI21X1TS U1657 ( .A0(n1377), .A1(\dataoutbuffer[3][3] ), .B0(n1757), .Y(
        n1380) );
  AOI22X1TS U1658 ( .A0(n1752), .A1(dataIn_WEST[3]), .B0(n145), .B1(
        dataIn_EAST[3]), .Y(n1379) );
  AOI22X1TS U1659 ( .A0(n1753), .A1(n1441), .B0(n124), .B1(n1478), .Y(n1378)
         );
  AOI21X1TS U1660 ( .A0(n1385), .A1(\dataoutbuffer[3][4] ), .B0(n1766), .Y(
        n1384) );
  AOI22X1TS U1661 ( .A0(n141), .A1(dataIn_WEST[4]), .B0(n1381), .B1(
        dataIn_EAST[4]), .Y(n1383) );
  AOI22X1TS U1662 ( .A0(n129), .A1(n1446), .B0(n1777), .B1(n1484), .Y(n1382)
         );
  AOI21X1TS U1663 ( .A0(n1385), .A1(\dataoutbuffer[3][5] ), .B0(n126), .Y(
        n1389) );
  AOI22X1TS U1664 ( .A0(n1386), .A1(dataIn_WEST[5]), .B0(n1758), .B1(
        dataIn_EAST[5]), .Y(n1388) );
  AOI22X1TS U1665 ( .A0(n1761), .A1(n1452), .B0(n124), .B1(n1491), .Y(n1387)
         );
  INVX2TS U1666 ( .A(n942), .Y(n1406) );
  AOI21X1TS U1667 ( .A0(n1406), .A1(\dataoutbuffer[4][0] ), .B0(n1725), .Y(
        n1396) );
  AOI22X1TS U1668 ( .A0(n1392), .A1(n1391), .B0(n1727), .B1(dataIn_EAST[0]), 
        .Y(n1395) );
  INVX2TS U1669 ( .A(n1393), .Y(n1729) );
  AOI22X1TS U1670 ( .A0(n1729), .A1(dataIn_SOUTH[0]), .B0(n297), .B1(n1498), 
        .Y(n1394) );
  AOI21X1TS U1671 ( .A0(n1406), .A1(\dataoutbuffer[4][1] ), .B0(n271), .Y(
        n1400) );
  AOI22X1TS U1672 ( .A0(n303), .A1(n1397), .B0(n1735), .B1(dataIn_EAST[1]), 
        .Y(n1399) );
  INVX2TS U1673 ( .A(n294), .Y(n1728) );
  AOI22X1TS U1674 ( .A0(n1736), .A1(dataIn_SOUTH[1]), .B0(n1728), .B1(n1506), 
        .Y(n1398) );
  AOI21X1TS U1675 ( .A0(n1406), .A1(\dataoutbuffer[4][2] ), .B0(n1741), .Y(
        n1405) );
  AOI22X1TS U1676 ( .A0(n283), .A1(n1402), .B0(n270), .B1(dataIn_EAST[2]), .Y(
        n1404) );
  AOI22X1TS U1677 ( .A0(n1745), .A1(dataIn_SOUTH[2]), .B0(n1412), .B1(n1513), 
        .Y(n1403) );
  AOI21X1TS U1678 ( .A0(n1406), .A1(\dataoutbuffer[4][3] ), .B0(n1725), .Y(
        n1410) );
  AOI22X1TS U1679 ( .A0(n1721), .A1(n1407), .B0(n1727), .B1(dataIn_EAST[3]), 
        .Y(n1409) );
  AOI22X1TS U1680 ( .A0(n1729), .A1(dataIn_SOUTH[3]), .B0(n289), .B1(n1520), 
        .Y(n1408) );
  AOI21X1TS U1681 ( .A0(n1417), .A1(\dataoutbuffer[4][4] ), .B0(n271), .Y(
        n1416) );
  AOI22X1TS U1682 ( .A0(n283), .A1(n1411), .B0(n1735), .B1(dataIn_EAST[4]), 
        .Y(n1415) );
  AOI22X1TS U1683 ( .A0(n1413), .A1(dataIn_SOUTH[4]), .B0(n1412), .B1(n1528), 
        .Y(n1414) );
  AOI21X1TS U1684 ( .A0(n1417), .A1(\dataoutbuffer[4][5] ), .B0(n1741), .Y(
        n1421) );
  AOI22X1TS U1685 ( .A0(n292), .A1(n1418), .B0(n270), .B1(dataIn_EAST[5]), .Y(
        n1420) );
  AOI22X1TS U1686 ( .A0(n284), .A1(dataIn_SOUTH[5]), .B0(n1728), .B1(n1536), 
        .Y(n1419) );
  INVX2TS U1687 ( .A(n916), .Y(n1440) );
  AOI21X1TS U1688 ( .A0(n1440), .A1(\dataoutbuffer[5][0] ), .B0(n1696), .Y(
        n1429) );
  AOI22X1TS U1689 ( .A0(n1423), .A1(n1496), .B0(n1698), .B1(n1457), .Y(n1428)
         );
  AOI22X1TS U1690 ( .A0(n1426), .A1(n1425), .B0(n1424), .B1(n1459), .Y(n1427)
         );
  AOI21X1TS U1691 ( .A0(n1440), .A1(\dataoutbuffer[5][1] ), .B0(n215), .Y(
        n1433) );
  AOI22X1TS U1692 ( .A0(n248), .A1(n1504), .B0(n1706), .B1(n1465), .Y(n1432)
         );
  AOI22X1TS U1693 ( .A0(n1700), .A1(n1430), .B0(n1716), .B1(n1466), .Y(n1431)
         );
  AOI21X1TS U1694 ( .A0(n1440), .A1(\dataoutbuffer[5][2] ), .B0(n1712), .Y(
        n1439) );
  AOI22X1TS U1695 ( .A0(n228), .A1(n1511), .B0(n1), .B1(n1471), .Y(n1438) );
  AOI22X1TS U1696 ( .A0(n1436), .A1(n1435), .B0(n1445), .B1(n1472), .Y(n1437)
         );
  AOI21X1TS U1697 ( .A0(n1440), .A1(\dataoutbuffer[5][3] ), .B0(n1696), .Y(
        n1444) );
  AOI22X1TS U1698 ( .A0(n1690), .A1(n1519), .B0(n1698), .B1(n1477), .Y(n1443)
         );
  AOI22X1TS U1699 ( .A0(n219), .A1(n1441), .B0(n1691), .B1(n1478), .Y(n1442)
         );
  AOI21X1TS U1700 ( .A0(n1451), .A1(\dataoutbuffer[5][4] ), .B0(n215), .Y(
        n1450) );
  AOI22X1TS U1701 ( .A0(n228), .A1(n1526), .B0(n1706), .B1(n1482), .Y(n1449)
         );
  AOI22X1TS U1702 ( .A0(n1447), .A1(n1446), .B0(n1445), .B1(n1484), .Y(n1448)
         );
  AOI21X1TS U1703 ( .A0(n1451), .A1(\dataoutbuffer[5][5] ), .B0(n1712), .Y(
        n1455) );
  AOI22X1TS U1704 ( .A0(n239), .A1(n1535), .B0(n1), .B1(n1490), .Y(n1454) );
  AOI22X1TS U1705 ( .A0(n1700), .A1(n1452), .B0(n235), .B1(n1491), .Y(n1453)
         );
  INVX2TS U1706 ( .A(n896), .Y(n1476) );
  AOI21X1TS U1707 ( .A0(n1476), .A1(\dataoutbuffer[6][0] ), .B0(n1668), .Y(
        n1464) );
  AOI22X1TS U1708 ( .A0(n1458), .A1(n1496), .B0(n1669), .B1(n1457), .Y(n1463)
         );
  AOI22X1TS U1709 ( .A0(n1461), .A1(dataIn_NORTH[0]), .B0(n1460), .B1(n1459), 
        .Y(n1462) );
  AOI21X1TS U1710 ( .A0(n1476), .A1(\dataoutbuffer[6][1] ), .B0(n1674), .Y(
        n1469) );
  AOI22X1TS U1711 ( .A0(n99), .A1(n1504), .B0(n1675), .B1(n1465), .Y(n1468) );
  AOI22X1TS U1712 ( .A0(n891), .A1(dataIn_NORTH[1]), .B0(n91), .B1(n1466), .Y(
        n1467) );
  AOI21X1TS U1713 ( .A0(n1476), .A1(\dataoutbuffer[6][2] ), .B0(n78), .Y(n1475) );
  AOI22X1TS U1714 ( .A0(n1483), .A1(n1511), .B0(n77), .B1(n1471), .Y(n1474) );
  AOI22X1TS U1715 ( .A0(n82), .A1(dataIn_NORTH[2]), .B0(n1485), .B1(n1472), 
        .Y(n1473) );
  AOI21X1TS U1716 ( .A0(n1476), .A1(\dataoutbuffer[6][3] ), .B0(n1668), .Y(
        n1481) );
  AOI22X1TS U1717 ( .A0(n1663), .A1(n1519), .B0(n1669), .B1(n1477), .Y(n1480)
         );
  AOI22X1TS U1718 ( .A0(n1664), .A1(dataIn_NORTH[3]), .B0(n91), .B1(n1478), 
        .Y(n1479) );
  AOI21X1TS U1719 ( .A0(n1489), .A1(\dataoutbuffer[6][4] ), .B0(n1674), .Y(
        n1488) );
  AOI22X1TS U1720 ( .A0(n1483), .A1(n1526), .B0(n1675), .B1(n1482), .Y(n1487)
         );
  AOI22X1TS U1721 ( .A0(n82), .A1(dataIn_NORTH[4]), .B0(n1485), .B1(n1484), 
        .Y(n1486) );
  AOI21X1TS U1722 ( .A0(n1489), .A1(\dataoutbuffer[6][5] ), .B0(n78), .Y(n1494) );
  AOI22X1TS U1723 ( .A0(n99), .A1(n1535), .B0(n77), .B1(n1490), .Y(n1493) );
  AOI22X1TS U1724 ( .A0(n87), .A1(dataIn_NORTH[5]), .B0(n104), .B1(n1491), .Y(
        n1492) );
  INVX2TS U1725 ( .A(n879), .Y(n1518) );
  AOI21X1TS U1726 ( .A0(n1518), .A1(\dataoutbuffer[7][0] ), .B0(n1525), .Y(
        n1502) );
  AOI22X1TS U1727 ( .A0(n1512), .A1(n1496), .B0(n1655), .B1(dataIn_EAST[0]), 
        .Y(n1501) );
  INVX2TS U1728 ( .A(n1497), .Y(n1637) );
  AOI22X1TS U1729 ( .A0(n50), .A1(n1499), .B0(n1637), .B1(n1498), .Y(n1500) );
  INVX2TS U1730 ( .A(n1503), .Y(n1636) );
  AOI21X1TS U1731 ( .A0(n1518), .A1(\dataoutbuffer[7][1] ), .B0(n1636), .Y(
        n1510) );
  AOI22X1TS U1732 ( .A0(n49), .A1(n1504), .B0(n1631), .B1(dataIn_EAST[1]), .Y(
        n1509) );
  INVX2TS U1733 ( .A(n1505), .Y(n1648) );
  AOI22X1TS U1734 ( .A0(n1648), .A1(n1507), .B0(n1647), .B1(n1506), .Y(n1508)
         );
  AOI21X1TS U1735 ( .A0(n1518), .A1(\dataoutbuffer[7][2] ), .B0(n1644), .Y(
        n1517) );
  AOI22X1TS U1736 ( .A0(n1512), .A1(n1511), .B0(n26), .B1(dataIn_EAST[2]), .Y(
        n1516) );
  AOI22X1TS U1737 ( .A0(n1638), .A1(n1514), .B0(n35), .B1(n1513), .Y(n1515) );
  AOI21X1TS U1738 ( .A0(n1518), .A1(\dataoutbuffer[7][3] ), .B0(n1654), .Y(
        n1524) );
  AOI22X1TS U1739 ( .A0(n1656), .A1(n1519), .B0(n1655), .B1(dataIn_EAST[3]), 
        .Y(n1523) );
  AOI22X1TS U1740 ( .A0(n1658), .A1(n1521), .B0(n1637), .B1(n1520), .Y(n1522)
         );
  AOI21X1TS U1741 ( .A0(n1534), .A1(\dataoutbuffer[7][4] ), .B0(n1525), .Y(
        n1533) );
  AOI22X1TS U1742 ( .A0(n1527), .A1(n1526), .B0(n1631), .B1(dataIn_EAST[4]), 
        .Y(n1532) );
  AOI22X1TS U1743 ( .A0(n1530), .A1(n1529), .B0(n1657), .B1(n1528), .Y(n1531)
         );
  AOI21X1TS U1744 ( .A0(n1534), .A1(\dataoutbuffer[7][5] ), .B0(n1636), .Y(
        n1541) );
  AOI22X1TS U1745 ( .A0(n49), .A1(n1535), .B0(n26), .B1(dataIn_EAST[5]), .Y(
        n1540) );
  AOI22X1TS U1746 ( .A0(n1648), .A1(n1538), .B0(n1537), .B1(n1536), .Y(n1539)
         );
  INVX2TS U1747 ( .A(readIn_EAST), .Y(n1624) );
  AOI22X1TS U1748 ( .A0(n1543), .A1(n1564), .B0(n1563), .B1(n1542), .Y(n1545)
         );
  AOI22X1TS U1749 ( .A0(n1546), .A1(n1624), .B0(n1545), .B1(n1544), .Y(n1548)
         );
  AOI22X1TS U1750 ( .A0(n1549), .A1(n1615), .B0(n1548), .B1(n1547), .Y(n1551)
         );
  AOI32X1TS U1751 ( .A0(n1551), .A1(n1495), .A2(n1550), .B0(n1652), .B1(n1915), 
        .Y(n2042) );
  INVX2TS U1752 ( .A(readIn_EAST), .Y(n1599) );
  AOI22X1TS U1753 ( .A0(n1553), .A1(n1564), .B0(n1563), .B1(n1552), .Y(n1555)
         );
  AOI22X1TS U1754 ( .A0(n1556), .A1(n1599), .B0(n1555), .B1(n1554), .Y(n1558)
         );
  AOI22X1TS U1755 ( .A0(n1559), .A1(n1581), .B0(n1558), .B1(n1557), .Y(n1561)
         );
  AOI32X1TS U1756 ( .A0(n1561), .A1(n1456), .A2(n1560), .B0(n1680), .B1(n1916), 
        .Y(n2043) );
  AOI22X1TS U1757 ( .A0(n1565), .A1(n1564), .B0(n1563), .B1(n1562), .Y(n1567)
         );
  AOI22X1TS U1758 ( .A0(n1568), .A1(n1599), .B0(n1567), .B1(n1566), .Y(n1570)
         );
  AOI22X1TS U1759 ( .A0(n1571), .A1(n1581), .B0(n1570), .B1(n1569), .Y(n1573)
         );
  AOI32X1TS U1760 ( .A0(n1573), .A1(n1422), .A2(n1572), .B0(n1711), .B1(n1917), 
        .Y(n2044) );
  CLKBUFX2TS U1761 ( .A(readIn_SOUTH), .Y(n1608) );
  AOI22X1TS U1762 ( .A0(n1575), .A1(n1608), .B0(n1595), .B1(n1574), .Y(n1577)
         );
  AOI22X1TS U1763 ( .A0(n1578), .A1(n1624), .B0(n1577), .B1(n1576), .Y(n1580)
         );
  AOI22X1TS U1764 ( .A0(n1582), .A1(n1581), .B0(n1580), .B1(n1579), .Y(n1584)
         );
  AOI32X1TS U1765 ( .A0(n1584), .A1(n1390), .A2(n1583), .B0(n1740), .B1(n1918), 
        .Y(n2045) );
  AOI22X1TS U1766 ( .A0(n115), .A1(n1608), .B0(readIn_NORTH), .B1(n1585), .Y(
        n1587) );
  AOI22X1TS U1767 ( .A0(n1588), .A1(n1599), .B0(n1587), .B1(n1586), .Y(n1590)
         );
  AOI22X1TS U1768 ( .A0(n1591), .A1(readIn_WEST), .B0(n1590), .B1(n1589), .Y(
        n1593) );
  AOI32X1TS U1769 ( .A0(n1593), .A1(n1364), .A2(n1592), .B0(n1773), .B1(n1919), 
        .Y(n2046) );
  AOI22X1TS U1770 ( .A0(n1596), .A1(n1608), .B0(n1595), .B1(n1594), .Y(n1598)
         );
  AOI22X1TS U1771 ( .A0(n1600), .A1(n1599), .B0(n1598), .B1(n1597), .Y(n1602)
         );
  AOI22X1TS U1772 ( .A0(n1603), .A1(readIn_WEST), .B0(n1602), .B1(n1601), .Y(
        n1606) );
  AOI32X1TS U1773 ( .A0(n1606), .A1(n1605), .A2(n1604), .B0(n1800), .B1(n1920), 
        .Y(n2047) );
  AOI22X1TS U1774 ( .A0(n1609), .A1(n1608), .B0(readIn_NORTH), .B1(n1607), .Y(
        n1611) );
  AOI22X1TS U1775 ( .A0(n1612), .A1(n1624), .B0(n1611), .B1(n1610), .Y(n1614)
         );
  AOI22X1TS U1776 ( .A0(n1616), .A1(n1615), .B0(n1614), .B1(n1613), .Y(n1619)
         );
  AOI32X1TS U1777 ( .A0(n1619), .A1(n1618), .A2(n1617), .B0(n1835), .B1(n1921), 
        .Y(n2048) );
  AOI22X1TS U1778 ( .A0(n1621), .A1(readIn_SOUTH), .B0(readIn_NORTH), .B1(
        n1620), .Y(n1623) );
  AOI22X1TS U1779 ( .A0(n1625), .A1(n1624), .B0(n1623), .B1(n1622), .Y(n1627)
         );
  AOI22X1TS U1780 ( .A0(n1628), .A1(readIn_WEST), .B0(n1627), .B1(n1626), .Y(
        n1630) );
  AOI32X1TS U1781 ( .A0(n1630), .A1(n1041), .A2(n1629), .B0(n1874), .B1(n1922), 
        .Y(n2049) );
  AOI22X1TS U1782 ( .A0(n1806), .A1(n1636), .B0(n1642), .B1(
        \destinationAddressbuffer[7][0] ), .Y(n1634) );
  AOI22X1TS U1783 ( .A0(n1512), .A1(n1689), .B0(n1631), .B1(n1688), .Y(n1633)
         );
  CLKBUFX2TS U1784 ( .A(destinationAddressIn_NORTH[0]), .Y(n1811) );
  AOI22X1TS U1785 ( .A0(n1648), .A1(destinationAddressIn_SOUTH[0]), .B0(n35), 
        .B1(n1811), .Y(n1632) );
  AOI22X1TS U1786 ( .A0(n1636), .A1(n1635), .B0(n1642), .B1(
        \destinationAddressbuffer[7][1] ), .Y(n1641) );
  AOI22X1TS U1787 ( .A0(n58), .A1(n1699), .B0(n1645), .B1(n1697), .Y(n1640) );
  CLKBUFX2TS U1788 ( .A(destinationAddressIn_NORTH[1]), .Y(n1821) );
  AOI22X1TS U1789 ( .A0(n1638), .A1(destinationAddressIn_SOUTH[1]), .B0(n1637), 
        .B1(n1821), .Y(n1639) );
  AOI22X1TS U1790 ( .A0(n1644), .A1(n1643), .B0(n1642), .B1(
        \destinationAddressbuffer[7][2] ), .Y(n1651) );
  AOI22X1TS U1791 ( .A0(n1646), .A1(n1707), .B0(n1645), .B1(n1705), .Y(n1650)
         );
  CLKBUFX2TS U1792 ( .A(destinationAddressIn_NORTH[2]), .Y(n1831) );
  AOI22X1TS U1793 ( .A0(n1648), .A1(destinationAddressIn_SOUTH[2]), .B0(n1647), 
        .B1(n1831), .Y(n1649) );
  AOI22X1TS U1794 ( .A0(n1654), .A1(n1653), .B0(n1652), .B1(
        \destinationAddressbuffer[7][3] ), .Y(n1661) );
  AOI22X1TS U1795 ( .A0(n1656), .A1(n1714), .B0(n1655), .B1(n1713), .Y(n1660)
         );
  CLKBUFX2TS U1796 ( .A(destinationAddressIn_NORTH[3]), .Y(n1842) );
  AOI22X1TS U1797 ( .A0(n1658), .A1(destinationAddressIn_SOUTH[3]), .B0(n1657), 
        .B1(n1842), .Y(n1659) );
  AOI22X1TS U1798 ( .A0(n1847), .A1(n1662), .B0(n1673), .B1(
        \destinationAddressbuffer[6][0] ), .Y(n1667) );
  AOI22X1TS U1799 ( .A0(n1663), .A1(n1689), .B0(n898), .B1(n1688), .Y(n1666)
         );
  CLKBUFX2TS U1800 ( .A(destinationAddressIn_NORTH[0]), .Y(n1849) );
  CLKBUFX2TS U1801 ( .A(destinationAddressIn_SOUTH[0]), .Y(n1851) );
  CLKBUFX2TS U1802 ( .A(n1851), .Y(n1809) );
  AOI22X1TS U1803 ( .A0(n1664), .A1(n1849), .B0(n1682), .B1(n1809), .Y(n1665)
         );
  AOI22X1TS U1804 ( .A0(n1726), .A1(n1668), .B0(n1673), .B1(
        \destinationAddressbuffer[6][1] ), .Y(n1672) );
  AOI22X1TS U1805 ( .A0(n108), .A1(n1699), .B0(n1669), .B1(n1697), .Y(n1671)
         );
  CLKBUFX2TS U1806 ( .A(destinationAddressIn_NORTH[1]), .Y(n1859) );
  CLKBUFX2TS U1807 ( .A(destinationAddressIn_SOUTH[1]), .Y(n1860) );
  CLKBUFX2TS U1808 ( .A(n1860), .Y(n1820) );
  AOI22X1TS U1809 ( .A0(n82), .A1(n1859), .B0(n1676), .B1(n1820), .Y(n1670) );
  AOI22X1TS U1810 ( .A0(n1734), .A1(n1674), .B0(n1673), .B1(
        \destinationAddressbuffer[6][2] ), .Y(n1679) );
  AOI22X1TS U1811 ( .A0(n1681), .A1(n1707), .B0(n1675), .B1(n1705), .Y(n1678)
         );
  CLKBUFX2TS U1812 ( .A(destinationAddressIn_NORTH[2]), .Y(n1868) );
  CLKBUFX2TS U1813 ( .A(destinationAddressIn_SOUTH[2]), .Y(n1869) );
  CLKBUFX2TS U1814 ( .A(n1869), .Y(n1830) );
  AOI22X1TS U1815 ( .A0(n1683), .A1(n1868), .B0(n1676), .B1(n1830), .Y(n1677)
         );
  AOI22X1TS U1816 ( .A0(n1742), .A1(n78), .B0(n1680), .B1(
        \destinationAddressbuffer[6][3] ), .Y(n1686) );
  AOI22X1TS U1817 ( .A0(n1681), .A1(n1714), .B0(n77), .B1(n1713), .Y(n1685) );
  CLKBUFX2TS U1818 ( .A(destinationAddressIn_NORTH[3]), .Y(n1878) );
  CLKBUFX2TS U1819 ( .A(destinationAddressIn_SOUTH[3]), .Y(n1880) );
  CLKBUFX2TS U1820 ( .A(n1880), .Y(n1840) );
  AOI22X1TS U1821 ( .A0(n1683), .A1(n1878), .B0(n1682), .B1(n1840), .Y(n1684)
         );
  AOI22X1TS U1822 ( .A0(n1847), .A1(n1687), .B0(n1704), .B1(
        \destinationAddressbuffer[5][0] ), .Y(n1695) );
  AOI22X1TS U1823 ( .A0(n1690), .A1(n1689), .B0(n917), .B1(n1688), .Y(n1694)
         );
  AOI22X1TS U1824 ( .A0(n1692), .A1(n1849), .B0(n1691), .B1(
        destinationAddressIn_SOUTH[0]), .Y(n1693) );
  AOI22X1TS U1825 ( .A0(readRequesterAddress[1]), .A1(n1696), .B0(n1704), .B1(
        \destinationAddressbuffer[5][1] ), .Y(n1703) );
  AOI22X1TS U1826 ( .A0(n239), .A1(n1699), .B0(n1698), .B1(n1697), .Y(n1702)
         );
  AOI22X1TS U1827 ( .A0(n1700), .A1(n1859), .B0(n229), .B1(
        destinationAddressIn_SOUTH[1]), .Y(n1701) );
  AOI22X1TS U1828 ( .A0(readRequesterAddress[2]), .A1(n215), .B0(n1704), .B1(
        \destinationAddressbuffer[5][2] ), .Y(n1710) );
  AOI22X1TS U1829 ( .A0(n1715), .A1(n1707), .B0(n1706), .B1(n1705), .Y(n1709)
         );
  AOI22X1TS U1830 ( .A0(n1426), .A1(n1868), .B0(n1716), .B1(
        destinationAddressIn_SOUTH[2]), .Y(n1708) );
  AOI22X1TS U1831 ( .A0(readRequesterAddress[3]), .A1(n1712), .B0(n1711), .B1(
        \destinationAddressbuffer[5][3] ), .Y(n1719) );
  AOI22X1TS U1832 ( .A0(n1715), .A1(n1714), .B0(n1), .B1(n1713), .Y(n1718) );
  AOI22X1TS U1833 ( .A0(n219), .A1(n1878), .B0(n1716), .B1(
        destinationAddressIn_SOUTH[3]), .Y(n1717) );
  AOI22X1TS U1834 ( .A0(n1750), .A1(n1720), .B0(n1733), .B1(
        \destinationAddressbuffer[4][0] ), .Y(n1724) );
  AOI22X1TS U1835 ( .A0(n1721), .A1(n1751), .B0(n943), .B1(
        destinationAddressIn_EAST[0]), .Y(n1723) );
  AOI22X1TS U1836 ( .A0(n308), .A1(n1851), .B0(n1728), .B1(n1849), .Y(n1722)
         );
  AOI22X1TS U1837 ( .A0(n1726), .A1(n1725), .B0(n1733), .B1(
        \destinationAddressbuffer[4][1] ), .Y(n1732) );
  AOI22X1TS U1838 ( .A0(n292), .A1(n1759), .B0(n1727), .B1(
        destinationAddressIn_EAST[1]), .Y(n1731) );
  AOI22X1TS U1839 ( .A0(n1729), .A1(n1860), .B0(n1728), .B1(n1859), .Y(n1730)
         );
  AOI22X1TS U1840 ( .A0(n1734), .A1(n271), .B0(n1733), .B1(
        \destinationAddressbuffer[4][2] ), .Y(n1739) );
  AOI22X1TS U1841 ( .A0(n1743), .A1(n1768), .B0(n1735), .B1(
        destinationAddressIn_EAST[2]), .Y(n1738) );
  AOI22X1TS U1842 ( .A0(n1736), .A1(n1869), .B0(n1744), .B1(n1868), .Y(n1737)
         );
  AOI22X1TS U1843 ( .A0(n1742), .A1(n1741), .B0(n1740), .B1(
        \destinationAddressbuffer[4][3] ), .Y(n1748) );
  AOI22X1TS U1844 ( .A0(n1743), .A1(n1775), .B0(n270), .B1(
        destinationAddressIn_EAST[3]), .Y(n1747) );
  AOI22X1TS U1845 ( .A0(n1745), .A1(n1880), .B0(n1744), .B1(n1878), .Y(n1746)
         );
  AOI22X1TS U1846 ( .A0(n1750), .A1(n1749), .B0(n1765), .B1(
        \destinationAddressbuffer[3][0] ), .Y(n1756) );
  AOI22X1TS U1847 ( .A0(n1752), .A1(n1751), .B0(n145), .B1(
        destinationAddressIn_EAST[0]), .Y(n1755) );
  AOI22X1TS U1848 ( .A0(n1753), .A1(n1811), .B0(n1760), .B1(n1809), .Y(n1754)
         );
  AOI22X1TS U1849 ( .A0(n1817), .A1(n1757), .B0(n1765), .B1(
        \destinationAddressbuffer[3][1] ), .Y(n1764) );
  AOI22X1TS U1850 ( .A0(n1776), .A1(n1759), .B0(n1758), .B1(
        destinationAddressIn_EAST[1]), .Y(n1763) );
  AOI22X1TS U1851 ( .A0(n1761), .A1(n1821), .B0(n1760), .B1(n1820), .Y(n1762)
         );
  AOI22X1TS U1852 ( .A0(n1827), .A1(n1766), .B0(n1765), .B1(
        \destinationAddressbuffer[3][2] ), .Y(n1772) );
  AOI22X1TS U1853 ( .A0(n151), .A1(n1768), .B0(n1767), .B1(
        destinationAddressIn_EAST[2]), .Y(n1771) );
  AOI22X1TS U1854 ( .A0(n1778), .A1(n1831), .B0(n1769), .B1(n1830), .Y(n1770)
         );
  AOI22X1TS U1855 ( .A0(n1837), .A1(n126), .B0(n1773), .B1(
        \destinationAddressbuffer[3][3] ), .Y(n1781) );
  AOI22X1TS U1856 ( .A0(n1776), .A1(n1775), .B0(n1774), .B1(
        destinationAddressIn_EAST[3]), .Y(n1780) );
  AOI22X1TS U1857 ( .A0(n1778), .A1(n1842), .B0(n1777), .B1(n1840), .Y(n1779)
         );
  AOI22X1TS U1858 ( .A0(n1806), .A1(n1782), .B0(n1794), .B1(
        \destinationAddressbuffer[2][0] ), .Y(n1788) );
  AOI22X1TS U1859 ( .A0(n1783), .A1(destinationAddressIn_WEST[0]), .B0(n991), 
        .B1(n1807), .Y(n1787) );
  AOI22X1TS U1860 ( .A0(n1785), .A1(n1811), .B0(n1784), .B1(n1809), .Y(n1786)
         );
  AOI22X1TS U1861 ( .A0(n1857), .A1(n1789), .B0(n1794), .B1(
        \destinationAddressbuffer[2][1] ), .Y(n1793) );
  AOI22X1TS U1862 ( .A0(n208), .A1(destinationAddressIn_WEST[1]), .B0(n1790), 
        .B1(n1818), .Y(n1792) );
  AOI22X1TS U1863 ( .A0(n182), .A1(n1821), .B0(n1802), .B1(n1820), .Y(n1791)
         );
  AOI22X1TS U1864 ( .A0(n1866), .A1(n1795), .B0(n1794), .B1(
        \destinationAddressbuffer[2][2] ), .Y(n1799) );
  AOI22X1TS U1865 ( .A0(n1801), .A1(destinationAddressIn_WEST[2]), .B0(n1796), 
        .B1(n1828), .Y(n1798) );
  AOI22X1TS U1866 ( .A0(n1355), .A1(n1831), .B0(n1802), .B1(n1830), .Y(n1797)
         );
  AOI22X1TS U1867 ( .A0(n1876), .A1(n177), .B0(n1800), .B1(
        \destinationAddressbuffer[2][3] ), .Y(n1805) );
  AOI22X1TS U1868 ( .A0(n1801), .A1(destinationAddressIn_WEST[3]), .B0(n176), 
        .B1(n1838), .Y(n1804) );
  AOI22X1TS U1869 ( .A0(n1785), .A1(n1842), .B0(n1802), .B1(n1840), .Y(n1803)
         );
  AOI22X1TS U1870 ( .A0(n1806), .A1(n1816), .B0(n1825), .B1(
        \destinationAddressbuffer[1][0] ), .Y(n1815) );
  AOI22X1TS U1871 ( .A0(n1808), .A1(destinationAddressIn_WEST[0]), .B0(n336), 
        .B1(n1807), .Y(n1814) );
  AOI22X1TS U1872 ( .A0(n1812), .A1(n1811), .B0(n1810), .B1(n1809), .Y(n1813)
         );
  AOI22X1TS U1873 ( .A0(n1817), .A1(n1816), .B0(n1825), .B1(
        \destinationAddressbuffer[1][1] ), .Y(n1824) );
  AOI22X1TS U1874 ( .A0(n358), .A1(destinationAddressIn_WEST[1]), .B0(n1819), 
        .B1(n1818), .Y(n1823) );
  AOI22X1TS U1875 ( .A0(n325), .A1(n1821), .B0(n1841), .B1(n1820), .Y(n1822)
         );
  AOI22X1TS U1876 ( .A0(n1827), .A1(n1826), .B0(n1825), .B1(
        \destinationAddressbuffer[1][2] ), .Y(n1834) );
  AOI22X1TS U1877 ( .A0(n1839), .A1(destinationAddressIn_WEST[2]), .B0(n1829), 
        .B1(n1828), .Y(n1833) );
  AOI22X1TS U1878 ( .A0(n1020), .A1(n1831), .B0(n1841), .B1(n1830), .Y(n1832)
         );
  AOI22X1TS U1879 ( .A0(n1837), .A1(n1836), .B0(n1835), .B1(
        \destinationAddressbuffer[1][3] ), .Y(n1845) );
  AOI22X1TS U1880 ( .A0(n1839), .A1(destinationAddressIn_WEST[3]), .B0(n1018), 
        .B1(n1838), .Y(n1844) );
  AOI22X1TS U1881 ( .A0(n1812), .A1(n1842), .B0(n1841), .B1(n1840), .Y(n1843)
         );
  AOI22X1TS U1882 ( .A0(n1847), .A1(n1846), .B0(n1864), .B1(
        \destinationAddressbuffer[0][0] ), .Y(n1855) );
  AOI22X1TS U1883 ( .A0(n1848), .A1(destinationAddressIn_WEST[0]), .B0(n1043), 
        .B1(destinationAddressIn_EAST[0]), .Y(n1854) );
  AOI22X1TS U1884 ( .A0(n1852), .A1(n1851), .B0(n1850), .B1(n1849), .Y(n1853)
         );
  AOI22X1TS U1885 ( .A0(n1857), .A1(n1856), .B0(n1864), .B1(
        \destinationAddressbuffer[0][1] ), .Y(n1863) );
  AOI22X1TS U1886 ( .A0(n432), .A1(destinationAddressIn_WEST[1]), .B0(n1858), 
        .B1(destinationAddressIn_EAST[1]), .Y(n1862) );
  AOI22X1TS U1887 ( .A0(n428), .A1(n1860), .B0(n415), .B1(n1859), .Y(n1861) );
  AOI22X1TS U1888 ( .A0(n1866), .A1(n1865), .B0(n1864), .B1(
        \destinationAddressbuffer[0][2] ), .Y(n1873) );
  AOI22X1TS U1889 ( .A0(n1877), .A1(destinationAddressIn_WEST[2]), .B0(n1867), 
        .B1(destinationAddressIn_EAST[2]), .Y(n1872) );
  AOI22X1TS U1890 ( .A0(n1870), .A1(n1869), .B0(n1879), .B1(n1868), .Y(n1871)
         );
  AOI22X1TS U1891 ( .A0(n1876), .A1(n1875), .B0(n1874), .B1(
        \destinationAddressbuffer[0][3] ), .Y(n1884) );
  AOI22X1TS U1892 ( .A0(n1877), .A1(destinationAddressIn_WEST[3]), .B0(n391), 
        .B1(destinationAddressIn_EAST[3]), .Y(n1883) );
  AOI22X1TS U1893 ( .A0(n1881), .A1(n1880), .B0(n1879), .B1(n1878), .Y(n1882)
         );
endmodule


module outputPortArbiter_3 ( clk, reset, selectBit_NORTH, 
        destinationAddressIn_NORTH, requesterAddressIn_NORTH, readIn_NORTH, 
        writeIn_NORTH, dataIn_NORTH, selectBit_SOUTH, 
        destinationAddressIn_SOUTH, requesterAddressIn_SOUTH, readIn_SOUTH, 
        writeIn_SOUTH, dataIn_SOUTH, selectBit_EAST, destinationAddressIn_EAST, 
        requesterAddressIn_EAST, readIn_EAST, writeIn_EAST, dataIn_EAST, 
        selectBit_WEST, destinationAddressIn_WEST, requesterAddressIn_WEST, 
        readIn_WEST, writeIn_WEST, dataIn_WEST, readReady, 
        readRequesterAddress, cacheDataOut, destinationAddressOut, 
        requesterAddressOut, readOut, writeOut, dataOut );
  input [11:0] destinationAddressIn_NORTH;
  input [3:0] requesterAddressIn_NORTH;
  input [5:0] dataIn_NORTH;
  input [11:0] destinationAddressIn_SOUTH;
  input [3:0] requesterAddressIn_SOUTH;
  input [5:0] dataIn_SOUTH;
  input [11:0] destinationAddressIn_EAST;
  input [3:0] requesterAddressIn_EAST;
  input [5:0] dataIn_EAST;
  input [11:0] destinationAddressIn_WEST;
  input [3:0] requesterAddressIn_WEST;
  input [5:0] dataIn_WEST;
  input [3:0] readRequesterAddress;
  input [5:0] cacheDataOut;
  output [11:0] destinationAddressOut;
  output [3:0] requesterAddressOut;
  output [5:0] dataOut;
  input clk, reset, selectBit_NORTH, readIn_NORTH, writeIn_NORTH,
         selectBit_SOUTH, readIn_SOUTH, writeIn_SOUTH, selectBit_EAST,
         readIn_EAST, writeIn_EAST, selectBit_WEST, readIn_WEST, writeIn_WEST,
         readReady;
  output readOut, writeOut;
  wire   \requesterAddressbuffer[0][3] , \requesterAddressbuffer[0][2] ,
         \requesterAddressbuffer[0][1] , \requesterAddressbuffer[0][0] ,
         \requesterAddressbuffer[1][3] , \requesterAddressbuffer[1][2] ,
         \requesterAddressbuffer[1][1] , \requesterAddressbuffer[1][0] ,
         \requesterAddressbuffer[2][3] , \requesterAddressbuffer[2][2] ,
         \requesterAddressbuffer[2][1] , \requesterAddressbuffer[2][0] ,
         \requesterAddressbuffer[3][3] , \requesterAddressbuffer[3][2] ,
         \requesterAddressbuffer[3][1] , \requesterAddressbuffer[3][0] ,
         \requesterAddressbuffer[4][3] , \requesterAddressbuffer[4][2] ,
         \requesterAddressbuffer[4][1] , \requesterAddressbuffer[4][0] ,
         \requesterAddressbuffer[5][3] , \requesterAddressbuffer[5][2] ,
         \requesterAddressbuffer[5][1] , \requesterAddressbuffer[5][0] ,
         \requesterAddressbuffer[6][3] , \requesterAddressbuffer[6][2] ,
         \requesterAddressbuffer[6][1] , \requesterAddressbuffer[6][0] ,
         \requesterAddressbuffer[7][3] , \requesterAddressbuffer[7][2] ,
         \requesterAddressbuffer[7][1] , \requesterAddressbuffer[7][0] ,
         \destinationAddressbuffer[0][11] , \destinationAddressbuffer[0][10] ,
         \destinationAddressbuffer[0][9] , \destinationAddressbuffer[0][8] ,
         \destinationAddressbuffer[0][7] , \destinationAddressbuffer[0][6] ,
         \destinationAddressbuffer[0][5] , \destinationAddressbuffer[0][4] ,
         \destinationAddressbuffer[0][3] , \destinationAddressbuffer[0][2] ,
         \destinationAddressbuffer[0][1] , \destinationAddressbuffer[0][0] ,
         \destinationAddressbuffer[1][11] , \destinationAddressbuffer[1][10] ,
         \destinationAddressbuffer[1][9] , \destinationAddressbuffer[1][8] ,
         \destinationAddressbuffer[1][7] , \destinationAddressbuffer[1][6] ,
         \destinationAddressbuffer[1][5] , \destinationAddressbuffer[1][4] ,
         \destinationAddressbuffer[1][3] , \destinationAddressbuffer[1][2] ,
         \destinationAddressbuffer[1][1] , \destinationAddressbuffer[1][0] ,
         \destinationAddressbuffer[2][11] , \destinationAddressbuffer[2][10] ,
         \destinationAddressbuffer[2][9] , \destinationAddressbuffer[2][8] ,
         \destinationAddressbuffer[2][7] , \destinationAddressbuffer[2][6] ,
         \destinationAddressbuffer[2][5] , \destinationAddressbuffer[2][4] ,
         \destinationAddressbuffer[2][3] , \destinationAddressbuffer[2][2] ,
         \destinationAddressbuffer[2][1] , \destinationAddressbuffer[2][0] ,
         \destinationAddressbuffer[3][11] , \destinationAddressbuffer[3][10] ,
         \destinationAddressbuffer[3][9] , \destinationAddressbuffer[3][8] ,
         \destinationAddressbuffer[3][7] , \destinationAddressbuffer[3][6] ,
         \destinationAddressbuffer[3][5] , \destinationAddressbuffer[3][4] ,
         \destinationAddressbuffer[3][3] , \destinationAddressbuffer[3][2] ,
         \destinationAddressbuffer[3][1] , \destinationAddressbuffer[3][0] ,
         \destinationAddressbuffer[4][11] , \destinationAddressbuffer[4][10] ,
         \destinationAddressbuffer[4][9] , \destinationAddressbuffer[4][8] ,
         \destinationAddressbuffer[4][7] , \destinationAddressbuffer[4][6] ,
         \destinationAddressbuffer[4][5] , \destinationAddressbuffer[4][4] ,
         \destinationAddressbuffer[4][3] , \destinationAddressbuffer[4][2] ,
         \destinationAddressbuffer[4][1] , \destinationAddressbuffer[4][0] ,
         \destinationAddressbuffer[5][11] , \destinationAddressbuffer[5][10] ,
         \destinationAddressbuffer[5][9] , \destinationAddressbuffer[5][8] ,
         \destinationAddressbuffer[5][7] , \destinationAddressbuffer[5][6] ,
         \destinationAddressbuffer[5][5] , \destinationAddressbuffer[5][4] ,
         \destinationAddressbuffer[5][3] , \destinationAddressbuffer[5][2] ,
         \destinationAddressbuffer[5][1] , \destinationAddressbuffer[5][0] ,
         \destinationAddressbuffer[6][11] , \destinationAddressbuffer[6][10] ,
         \destinationAddressbuffer[6][9] , \destinationAddressbuffer[6][8] ,
         \destinationAddressbuffer[6][7] , \destinationAddressbuffer[6][6] ,
         \destinationAddressbuffer[6][5] , \destinationAddressbuffer[6][4] ,
         \destinationAddressbuffer[6][3] , \destinationAddressbuffer[6][2] ,
         \destinationAddressbuffer[6][1] , \destinationAddressbuffer[6][0] ,
         \destinationAddressbuffer[7][11] , \destinationAddressbuffer[7][10] ,
         \destinationAddressbuffer[7][9] , \destinationAddressbuffer[7][8] ,
         \destinationAddressbuffer[7][7] , \destinationAddressbuffer[7][6] ,
         \destinationAddressbuffer[7][5] , \destinationAddressbuffer[7][4] ,
         \destinationAddressbuffer[7][3] , \destinationAddressbuffer[7][2] ,
         \destinationAddressbuffer[7][1] , \destinationAddressbuffer[7][0] ,
         \dataoutbuffer[7][5] , \dataoutbuffer[7][4] , \dataoutbuffer[7][3] ,
         \dataoutbuffer[7][2] , \dataoutbuffer[7][1] , \dataoutbuffer[7][0] ,
         \dataoutbuffer[6][5] , \dataoutbuffer[6][4] , \dataoutbuffer[6][3] ,
         \dataoutbuffer[6][2] , \dataoutbuffer[6][1] , \dataoutbuffer[6][0] ,
         \dataoutbuffer[5][5] , \dataoutbuffer[5][4] , \dataoutbuffer[5][3] ,
         \dataoutbuffer[5][2] , \dataoutbuffer[5][1] , \dataoutbuffer[5][0] ,
         \dataoutbuffer[4][5] , \dataoutbuffer[4][4] , \dataoutbuffer[4][3] ,
         \dataoutbuffer[4][2] , \dataoutbuffer[4][1] , \dataoutbuffer[4][0] ,
         \dataoutbuffer[3][5] , \dataoutbuffer[3][4] , \dataoutbuffer[3][3] ,
         \dataoutbuffer[3][2] , \dataoutbuffer[3][1] , \dataoutbuffer[3][0] ,
         \dataoutbuffer[2][5] , \dataoutbuffer[2][4] , \dataoutbuffer[2][3] ,
         \dataoutbuffer[2][2] , \dataoutbuffer[2][1] , \dataoutbuffer[2][0] ,
         \dataoutbuffer[1][5] , \dataoutbuffer[1][4] , \dataoutbuffer[1][3] ,
         \dataoutbuffer[1][2] , \dataoutbuffer[1][1] , \dataoutbuffer[1][0] ,
         \dataoutbuffer[0][5] , \dataoutbuffer[0][4] , \dataoutbuffer[0][3] ,
         \dataoutbuffer[0][2] , \dataoutbuffer[0][1] , \dataoutbuffer[0][0] ,
         N2624, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151;
  wire   [0:7] writeOutbuffer;
  wire   [0:7] readOutbuffer;

  DFFNSRX1TS full_reg_reg ( .D(N2624), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(
        n1920) );
  DFFNSRX1TS \dataoutbuffer_reg[0][0]  ( .D(n1992), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][1]  ( .D(n1993), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][2]  ( .D(n1994), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][3]  ( .D(n1995), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][4]  ( .D(n1996), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][5]  ( .D(n1997), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][5] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[2][0]  ( .D(n1980), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[2][1]  ( .D(n1981), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[2][2]  ( .D(n1982), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[2][3]  ( .D(n1983), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][0]  ( .D(n2116), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][1]  ( .D(n2117), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][2]  ( .D(n2118), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][3]  ( .D(n2119), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][3] ) );
  DFFNSRX1TS \writeOutbuffer_reg[7]  ( .D(n2040), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[7]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][4]  ( .D(n2060), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][5]  ( .D(n2061), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][6]  ( .D(n2062), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][7]  ( .D(n2063), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][8]  ( .D(n2064), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][9]  ( .D(n2065), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][11]  ( .D(n2067), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[6]  ( .D(n2041), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[6]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][4]  ( .D(n2072), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][5]  ( .D(n2073), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][6]  ( .D(n2074), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][7]  ( .D(n2075), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][8]  ( .D(n2076), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][9]  ( .D(n2077), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][10]  ( .D(n2078), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][11]  ( .D(n2079), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[3]  ( .D(n2044), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[3]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][4]  ( .D(n2108), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][5]  ( .D(n2109), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][6]  ( .D(n2110), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][7]  ( .D(n2111), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][8]  ( .D(n2112), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][9]  ( .D(n2113), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][10]  ( .D(n2114), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][11]  ( .D(n2115), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[2]  ( .D(n2045), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[2]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][4]  ( .D(n2120), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][5]  ( .D(n2121), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][6]  ( .D(n2122), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][7]  ( .D(n2123), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][8]  ( .D(n2124), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][9]  ( .D(n2125), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][10]  ( .D(n2126), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][11]  ( .D(n2127), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][11] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][0]  ( .D(n2034), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][1]  ( .D(n2035), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][2]  ( .D(n2036), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][3]  ( .D(n2037), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][4]  ( .D(n2038), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][5]  ( .D(n2039), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][0]  ( .D(n2028), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][1]  ( .D(n2029), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][2]  ( .D(n2030), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][3]  ( .D(n2031), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][4]  ( .D(n2032), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][5]  ( .D(n2033), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][0]  ( .D(n2010), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][1]  ( .D(n2011), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][2]  ( .D(n2012), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][3]  ( .D(n2013), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][4]  ( .D(n2014), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][5]  ( .D(n2015), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][0]  ( .D(n2004), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][1]  ( .D(n2005), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][2]  ( .D(n2006), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][3]  ( .D(n2007), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][4]  ( .D(n2008), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][5]  ( .D(n2009), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][5] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[5][0]  ( .D(n1968), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[5][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[5][1]  ( .D(n1969), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[5][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[5][2]  ( .D(n1970), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[5][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[5][3]  ( .D(n1971), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[5][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][0]  ( .D(n2080), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][1]  ( .D(n2081), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][2]  ( .D(n2082), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][3]  ( .D(n2083), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[4][0]  ( .D(n1972), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[4][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[4][1]  ( .D(n1973), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[4][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[4][2]  ( .D(n1974), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[4][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[4][3]  ( .D(n1975), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[4][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][0]  ( .D(n2092), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][1]  ( .D(n2093), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][2]  ( .D(n2094), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][3]  ( .D(n2095), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[1][0]  ( .D(n1984), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[1][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[1][1]  ( .D(n1985), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[1][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[1][2]  ( .D(n1986), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[1][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[1][3]  ( .D(n1987), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[1][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][0]  ( .D(n2128), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][1]  ( .D(n2129), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][2]  ( .D(n2130), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][3]  ( .D(n2131), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[0][0]  ( .D(n1988), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[0][1]  ( .D(n1989), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[0][2]  ( .D(n1990), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[0][3]  ( .D(n1991), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][0]  ( .D(n2140), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][1]  ( .D(n2141), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][2]  ( .D(n2142), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][3]  ( .D(n2143), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][0]  ( .D(n2022), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][1]  ( .D(n2023), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][2]  ( .D(n2024), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][3]  ( .D(n2025), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][4]  ( .D(n2026), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][5]  ( .D(n2027), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][0]  ( .D(n2016), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][1]  ( .D(n2017), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][2]  ( .D(n2018), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][3]  ( .D(n2019), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][4]  ( .D(n2020), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][5]  ( .D(n2021), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][0]  ( .D(n1998), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][1]  ( .D(n1999), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][2]  ( .D(n2000), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][3]  ( .D(n2001), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][4]  ( .D(n2002), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][5]  ( .D(n2003), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][5] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[7][0]  ( .D(n1960), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[7][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[7][1]  ( .D(n1961), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[7][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[7][2]  ( .D(n1962), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[7][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[7][3]  ( .D(n1963), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[7][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][0]  ( .D(n2056), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][1]  ( .D(n2057), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][2]  ( .D(n2058), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][3]  ( .D(n2059), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[6][0]  ( .D(n1964), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[6][1]  ( .D(n1965), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[6][2]  ( .D(n1966), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[6][3]  ( .D(n1967), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][0]  ( .D(n2068), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][1]  ( .D(n2069), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][2]  ( .D(n2070), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][3]  ( .D(n2071), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[3][0]  ( .D(n1976), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[3][1]  ( .D(n1977), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[3][2]  ( .D(n1978), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[3][3]  ( .D(n1979), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][0]  ( .D(n2104), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][1]  ( .D(n2105), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][2]  ( .D(n2106), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][3]  ( .D(n2107), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][3] ) );
  DFFNSRX1TS \writeOutbuffer_reg[5]  ( .D(n2042), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[5]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][4]  ( .D(n2084), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][5]  ( .D(n2085), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][6]  ( .D(n2086), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][7]  ( .D(n2087), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][8]  ( .D(n2088), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][9]  ( .D(n2089), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][10]  ( .D(n2090), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][11]  ( .D(n2091), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[4]  ( .D(n2043), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[4]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][4]  ( .D(n2096), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][5]  ( .D(n2097), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][6]  ( .D(n2098), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][7]  ( .D(n2099), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][8]  ( .D(n2100), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][9]  ( .D(n2101), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][10]  ( .D(n2102), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][11]  ( .D(n2103), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[1]  ( .D(n2046), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[1]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][4]  ( .D(n2132), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][5]  ( .D(n2133), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][6]  ( .D(n2134), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][7]  ( .D(n2135), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][8]  ( .D(n2136), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][9]  ( .D(n2137), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][10]  ( .D(n2138), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][11]  ( .D(n2139), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[0]  ( .D(n2047), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[0]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][4]  ( .D(n2144), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][5]  ( .D(n2145), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][6]  ( .D(n2146), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][7]  ( .D(n2147), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][8]  ( .D(n2148), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][9]  ( .D(n2149), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][10]  ( .D(n2150), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][11]  ( .D(n2151), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][11] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][10]  ( .D(n2066), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][10] ) );
  DFFNSRX1TS writeOut_reg ( .D(n1937), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        writeOut) );
  DFFNSRX1TS \destinationAddressOut_reg[4]  ( .D(n1946), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[4]) );
  DFFNSRX1TS \destinationAddressOut_reg[5]  ( .D(n1947), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[5]) );
  DFFNSRX1TS \destinationAddressOut_reg[6]  ( .D(n1948), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[6]) );
  DFFNSRX1TS \destinationAddressOut_reg[7]  ( .D(n1949), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[7]) );
  DFFNSRX1TS \destinationAddressOut_reg[8]  ( .D(n1950), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[8]) );
  DFFNSRX1TS \destinationAddressOut_reg[9]  ( .D(n1951), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[9]) );
  DFFNSRX1TS \destinationAddressOut_reg[10]  ( .D(n1952), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[10]) );
  DFFNSRX1TS \destinationAddressOut_reg[11]  ( .D(n1953), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[11]) );
  DFFNSRX1TS readOut_reg ( .D(n1936), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        readOut) );
  DFFNSRX1TS \requesterAddressOut_reg[0]  ( .D(n1938), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[0]) );
  DFFNSRX1TS \requesterAddressOut_reg[1]  ( .D(n1939), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[1]) );
  DFFNSRX1TS \requesterAddressOut_reg[2]  ( .D(n1940), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[2]) );
  DFFNSRX1TS \requesterAddressOut_reg[3]  ( .D(n1941), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[3]) );
  DFFNSRX1TS \destinationAddressOut_reg[0]  ( .D(n1942), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[0]) );
  DFFNSRX1TS \destinationAddressOut_reg[1]  ( .D(n1943), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[1]) );
  DFFNSRX1TS \destinationAddressOut_reg[2]  ( .D(n1944), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[2]) );
  DFFNSRX1TS \destinationAddressOut_reg[3]  ( .D(n1945), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[3]) );
  DFFNSRX1TS \dataOut_reg[0]  ( .D(n1954), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[0]) );
  DFFNSRX1TS \dataOut_reg[1]  ( .D(n1955), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[1]) );
  DFFNSRX1TS \dataOut_reg[2]  ( .D(n1956), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[2]) );
  DFFNSRX1TS \dataOut_reg[3]  ( .D(n1957), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[3]) );
  DFFNSRX1TS \dataOut_reg[4]  ( .D(n1958), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[4]) );
  DFFNSRX1TS \dataOut_reg[5]  ( .D(n1959), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[5]) );
  DFFNSRX1TS \read_reg_reg[1]  ( .D(n1935), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1913), .QN(n1912) );
  DFFNSRX1TS \write_reg_reg[0]  ( .D(n1930), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1911), .QN(n1915) );
  DFFNSRX1TS \write_reg_reg[2]  ( .D(n1932), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1916), .QN(n1917) );
  DFFNSRX1TS \read_reg_reg[0]  ( .D(n1929), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1906), .QN(n1918) );
  DFFNSRX1TS \read_reg_reg[2]  ( .D(n1934), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1909), .QN(n1910) );
  DFFNSRX1TS empty_reg_reg ( .D(n1933), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        n1908), .QN(n1907) );
  DFFNSRX1TS \readOutbuffer_reg[7]  ( .D(n2048), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[7]), .QN(n1921) );
  DFFNSRX1TS \readOutbuffer_reg[4]  ( .D(n2051), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[4]), .QN(n1924) );
  DFFNSRX1TS \readOutbuffer_reg[6]  ( .D(n2049), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[6]), .QN(n1922) );
  DFFNSRX1TS \readOutbuffer_reg[5]  ( .D(n2050), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[5]), .QN(n1923) );
  DFFNSRX1TS \readOutbuffer_reg[0]  ( .D(n2055), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[0]), .QN(n1928) );
  DFFNSRX1TS \readOutbuffer_reg[3]  ( .D(n2052), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[3]), .QN(n1925) );
  DFFNSRX1TS \readOutbuffer_reg[2]  ( .D(n2053), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[2]), .QN(n1926) );
  DFFNSRX1TS \readOutbuffer_reg[1]  ( .D(n2054), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[1]), .QN(n1927) );
  DFFNSRX1TS \write_reg_reg[1]  ( .D(n1931), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1914), .QN(n1919) );
  CLKBUFX2TS U3 ( .A(n14), .Y(n72) );
  CMPR32X2TS U4 ( .A(n454), .B(n475), .C(n16), .CO(n17), .S(n14) );
  CMPR32X2TS U5 ( .A(n531), .B(n452), .C(n455), .CO(n445), .S(n458) );
  CLKBUFX2TS U6 ( .A(n20), .Y(n74) );
  CMPR32X2TS U7 ( .A(n451), .B(n513), .C(n450), .CO(n453), .S(n467) );
  CMPR32X2TS U8 ( .A(selectBit_SOUTH), .B(selectBit_NORTH), .C(selectBit_EAST), 
        .CO(n454), .S(n450) );
  NOR2XLTS U9 ( .A(n9), .B(n73), .Y(n27) );
  OR2X1TS U10 ( .A(n449), .B(n505), .Y(n2) );
  OR2X1TS U11 ( .A(n21), .B(n507), .Y(n9) );
  INVX2TS U12 ( .A(n22), .Y(n120) );
  OAI31X1TS U13 ( .A0(n517), .A1(n516), .A2(n538), .B0(n539), .Y(n519) );
  NOR3XLTS U14 ( .A(n28), .B(n75), .C(n9), .Y(n1610) );
  NOR2XLTS U15 ( .A(n1598), .B(n179), .Y(n188) );
  NOR2XLTS U16 ( .A(n1593), .B(n1590), .Y(n124) );
  ADDHXLTS U17 ( .A(n493), .B(n450), .CO(n16), .S(n15) );
  NOR2XLTS U18 ( .A(n1551), .B(n1548), .Y(n34) );
  NAND2X1TS U19 ( .A(n539), .B(n521), .Y(n509) );
  NOR2XLTS U20 ( .A(selectBit_NORTH), .B(selectBit_SOUTH), .Y(n539) );
  NOR2XLTS U21 ( .A(n841), .B(n520), .Y(n690) );
  INVX2TS U22 ( .A(n1580), .Y(n1578) );
  INVX2TS U23 ( .A(n1558), .Y(n1556) );
  INVX2TS U24 ( .A(n1601), .Y(n1599) );
  INVX2TS U25 ( .A(n1628), .Y(n1625) );
  INVX2TS U26 ( .A(n1618), .Y(n1615) );
  INVX2TS U27 ( .A(n1561), .Y(n1559) );
  AOI31XLTS U28 ( .A0(n34), .A1(n30), .A2(n1544), .B0(n218), .Y(n33) );
  NOR2XLTS U29 ( .A(n1544), .B(n36), .Y(n39) );
  NOR2XLTS U30 ( .A(n1608), .B(n315), .Y(n316) );
  NOR3XLTS U31 ( .A(n1584), .B(n1578), .C(n271), .Y(n267) );
  NOR2XLTS U32 ( .A(n441), .B(n1585), .Y(n268) );
  NOR2XLTS U33 ( .A(n1567), .B(n223), .Y(n222) );
  NOR2XLTS U34 ( .A(n482), .B(n1562), .Y(n78) );
  NOR2XLTS U35 ( .A(n1552), .B(n218), .Y(n32) );
  NOR2XLTS U36 ( .A(n1587), .B(n129), .Y(n125) );
  NOR3XLTS U37 ( .A(n1561), .B(n1556), .C(n82), .Y(n77) );
  NOR3XLTS U38 ( .A(n1551), .B(n1546), .C(n35), .Y(n31) );
  NOR2XLTS U39 ( .A(n306), .B(n1605), .Y(n175) );
  NOR2XLTS U40 ( .A(n1596), .B(n179), .Y(n180) );
  NOR2X1TS U41 ( .A(n1610), .B(n315), .Y(n322) );
  NOR2X1TS U42 ( .A(n1554), .B(n83), .Y(n84) );
  INVX2TS U43 ( .A(n77), .Y(n1472) );
  INVX1TS U44 ( .A(n139), .Y(n954) );
  NOR3X1TS U45 ( .A(n1573), .B(n1568), .C(n221), .Y(n216) );
  NAND2BXLTS U46 ( .AN(n271), .B(n270), .Y(n272) );
  NAND2BXLTS U47 ( .AN(n82), .B(n81), .Y(n83) );
  NAND2BXLTS U48 ( .AN(n387), .B(n386), .Y(n388) );
  AOI31X1TS U49 ( .A0(n220), .A1(n1564), .A2(n215), .B0(n482), .Y(n219) );
  INVX1TS U50 ( .A(n1548), .Y(n1546) );
  INVX1TS U51 ( .A(n1614), .Y(n1611) );
  INVX1TS U52 ( .A(n1570), .Y(n1568) );
  NOR2X1TS U53 ( .A(n119), .B(n264), .Y(n1548) );
  NOR2X1TS U54 ( .A(n119), .B(n376), .Y(n1590) );
  NAND2BX1TS U55 ( .AN(n118), .B(n515), .Y(n376) );
  ADDFX1TS U56 ( .A(n476), .B(n475), .CI(n474), .CO(n470), .S(n494) );
  NOR3X1TS U57 ( .A(n28), .B(n74), .C(n19), .Y(n1598) );
  NAND3X1TS U58 ( .A(n475), .B(n28), .C(n214), .Y(n1544) );
  OAI21X1TS U59 ( .A0(n27), .A1(n25), .B0(n26), .Y(n118) );
  NAND3X1TS U60 ( .A(n28), .B(n214), .C(n19), .Y(n1564) );
  INVX1TS U61 ( .A(n1555), .Y(n1554) );
  INVX1TS U62 ( .A(n1604), .Y(n1602) );
  INVX1TS U63 ( .A(n1593), .Y(n1591) );
  NOR3X1TS U64 ( .A(n24), .B(n75), .C(n74), .Y(n1624) );
  NOR2X1TS U65 ( .A(n214), .B(n73), .Y(n303) );
  INVX1TS U66 ( .A(n1577), .Y(n1576) );
  OAI21X1TS U67 ( .A0(n506), .A1(n21), .B0(n74), .Y(n213) );
  INVX1TS U68 ( .A(n1631), .Y(n1629) );
  NOR3X1TS U69 ( .A(n116), .B(n172), .C(n263), .Y(n1561) );
  NOR3X1TS U70 ( .A(n172), .B(n71), .C(n374), .Y(n1593) );
  NAND2BX1TS U71 ( .AN(n117), .B(n451), .Y(n374) );
  OAI21X1TS U72 ( .A0(n305), .A1(n495), .B0(n22), .Y(n19) );
  NOR2X1TS U73 ( .A(n841), .B(n518), .Y(n544) );
  NOR3X1TS U74 ( .A(n514), .B(selectBit_EAST), .C(n513), .Y(n508) );
  INVX1TS U75 ( .A(selectBit_EAST), .Y(n512) );
  CLKBUFX2TS U76 ( .A(readIn_EAST), .Y(n1543) );
  INVX1TS U77 ( .A(n1917), .Y(n499) );
  CLKINVX1TS U78 ( .A(n465), .Y(n469) );
  XOR2X1TS U79 ( .A(n472), .B(n471), .Y(n496) );
  INVX2TS U80 ( .A(selectBit_NORTH), .Y(n505) );
  NOR2XLTS U81 ( .A(n1631), .B(n1628), .Y(n386) );
  NOR2XLTS U82 ( .A(n1584), .B(n1580), .Y(n270) );
  NOR2XLTS U83 ( .A(n1618), .B(n1614), .Y(n312) );
  NOR2XLTS U84 ( .A(n1604), .B(n1601), .Y(n177) );
  NAND2BX1TS U85 ( .AN(n313), .B(n312), .Y(n315) );
  INVX2TS U86 ( .A(n222), .Y(n246) );
  NAND2BX1TS U87 ( .AN(n178), .B(n177), .Y(n179) );
  CLKAND2X2TS U88 ( .A(n469), .B(n468), .Y(n474) );
  NOR3X1TS U89 ( .A(n72), .B(n71), .C(n374), .Y(n1618) );
  INVX2TS U90 ( .A(n1610), .Y(n1608) );
  NAND4XLTS U91 ( .A(n495), .B(n510), .C(n382), .D(n483), .Y(n1605) );
  NOR3X1TS U92 ( .A(n15), .B(n172), .C(n374), .Y(n1604) );
  INVX2TS U93 ( .A(n1598), .Y(n1596) );
  NAND4XLTS U94 ( .A(n484), .B(n1911), .C(n510), .D(n486), .Y(n1594) );
  NOR3X1TS U95 ( .A(n72), .B(n15), .C(n374), .Y(n1631) );
  NOR3X1TS U96 ( .A(n14), .B(n71), .C(n263), .Y(n1573) );
  NAND4XLTS U97 ( .A(n487), .B(n499), .C(n513), .D(n382), .Y(n1562) );
  NAND4XLTS U98 ( .A(n266), .B(n511), .C(n382), .D(n308), .Y(n1585) );
  NOR3X1TS U99 ( .A(n72), .B(n15), .C(n263), .Y(n1584) );
  NAND4XLTS U100 ( .A(n1911), .B(n484), .C(n499), .D(n511), .Y(n1552) );
  CLKAND2X2TS U101 ( .A(n524), .B(n522), .Y(n552) );
  AO21X1TS U102 ( .A0(n449), .A1(n505), .B0(n305), .Y(n21) );
  NOR3BXLTS U103 ( .AN(readReady), .B(selectBit_WEST), .C(n515), .Y(n538) );
  NAND3XLTS U104 ( .A(n506), .B(n508), .C(n505), .Y(n518) );
  NAND3XLTS U105 ( .A(selectBit_NORTH), .B(n508), .C(n507), .Y(n520) );
  AOI21X1TS U106 ( .A0(n312), .A1(n307), .B0(n306), .Y(n310) );
  NOR2XLTS U107 ( .A(n1573), .B(n1570), .Y(n220) );
  NAND2X1TS U108 ( .A(n127), .B(n1594), .Y(n130) );
  NOR2XLTS U109 ( .A(n1561), .B(n1558), .Y(n81) );
  AOI21X1TS U110 ( .A0(n177), .A1(n173), .B0(n218), .Y(n176) );
  AOI21X1TS U111 ( .A0(n386), .A1(n380), .B0(n306), .Y(n384) );
  XOR2XLTS U112 ( .A(n445), .B(n447), .Y(n464) );
  OAI21XLTS U113 ( .A0(n487), .A1(n1912), .B0(n447), .Y(n448) );
  NAND3XLTS U114 ( .A(n305), .B(n266), .C(n381), .Y(n215) );
  AOI21X1TS U115 ( .A0(n270), .A1(n265), .B0(n482), .Y(n269) );
  XOR2X1TS U116 ( .A(n499), .B(n17), .Y(n117) );
  NOR2XLTS U117 ( .A(n379), .B(reset), .Y(n498) );
  NAND4XLTS U118 ( .A(n493), .B(n510), .C(n443), .D(n308), .Y(n1619) );
  NOR3XLTS U119 ( .A(n304), .B(n303), .C(n376), .Y(n1614) );
  INVX2TS U120 ( .A(n1590), .Y(n1588) );
  NAND4XLTS U121 ( .A(n511), .B(n382), .C(n381), .D(n486), .Y(n1632) );
  INVX2TS U122 ( .A(n1624), .Y(n1622) );
  NOR3BXLTS U123 ( .AN(n377), .B(n376), .C(n375), .Y(n1628) );
  NAND4XLTS U124 ( .A(n493), .B(n266), .C(readReady), .D(n308), .Y(n1574) );
  INVX2TS U125 ( .A(n1573), .Y(n1571) );
  NOR3XLTS U126 ( .A(n304), .B(n303), .C(n264), .Y(n1570) );
  NOR3XLTS U127 ( .A(n75), .B(n20), .C(n23), .Y(n1577) );
  INVX2TS U128 ( .A(n1584), .Y(n1581) );
  NOR3BXLTS U129 ( .AN(n377), .B(n264), .C(n375), .Y(n1580) );
  NAND4XLTS U130 ( .A(n14), .B(n116), .C(n117), .D(selectBit_WEST), .Y(n1549)
         );
  INVX2TS U131 ( .A(n1544), .Y(n1545) );
  INVX2TS U132 ( .A(destinationAddressIn_SOUTH[11]), .Y(n152) );
  INVX2TS U133 ( .A(destinationAddressIn_SOUTH[10]), .Y(n160) );
  INVX2TS U134 ( .A(destinationAddressIn_SOUTH[9]), .Y(n166) );
  INVX2TS U135 ( .A(destinationAddressIn_SOUTH[8]), .Y(n156) );
  CLKAND2X2TS U136 ( .A(n469), .B(n467), .Y(n473) );
  NOR2XLTS U137 ( .A(reset), .B(n441), .Y(n497) );
  AO22XLTS U138 ( .A0(n499), .A1(n498), .B0(n497), .B1(n496), .Y(n1932) );
  AO22XLTS U139 ( .A0(n493), .A1(n498), .B0(n497), .B1(n492), .Y(n1930) );
  AO22XLTS U140 ( .A0(n495), .A1(n498), .B0(n497), .B1(n494), .Y(n1931) );
  OAI21XLTS U141 ( .A0(n379), .A1(n490), .B0(n491), .Y(n1933) );
  NAND4XLTS U142 ( .A(n867), .B(n866), .C(n865), .D(n864), .Y(n1959) );
  NAND4XLTS U143 ( .A(n845), .B(n844), .C(n843), .D(n864), .Y(n1958) );
  NAND4XLTS U144 ( .A(n834), .B(n833), .C(n832), .D(n864), .Y(n1957) );
  NAND4XLTS U145 ( .A(n824), .B(n823), .C(n822), .D(n864), .Y(n1956) );
  NAND4XLTS U146 ( .A(n805), .B(n804), .C(n803), .D(n802), .Y(n1955) );
  NAND4XLTS U147 ( .A(n785), .B(n784), .C(n783), .D(n802), .Y(n1954) );
  NAND4XLTS U148 ( .A(n656), .B(n655), .C(n654), .D(n653), .Y(n1945) );
  NAND4XLTS U149 ( .A(n645), .B(n644), .C(n643), .D(n642), .Y(n1944) );
  NAND4XLTS U150 ( .A(n627), .B(n626), .C(n625), .D(n624), .Y(n1943) );
  NAND4XLTS U151 ( .A(n612), .B(n611), .C(n610), .D(n609), .Y(n1942) );
  NAND4XLTS U152 ( .A(n600), .B(n599), .C(n598), .D(n653), .Y(n1941) );
  NAND4XLTS U153 ( .A(n589), .B(n588), .C(n587), .D(n642), .Y(n1940) );
  NAND4XLTS U154 ( .A(n580), .B(n579), .C(n578), .D(n624), .Y(n1939) );
  NAND4XLTS U155 ( .A(n563), .B(n562), .C(n561), .D(n609), .Y(n1938) );
  NAND4XLTS U156 ( .A(n542), .B(n541), .C(n540), .D(n802), .Y(n1936) );
  NAND3XLTS U157 ( .A(n775), .B(n774), .C(n773), .Y(n1953) );
  NAND3XLTS U158 ( .A(n761), .B(n760), .C(n759), .Y(n1952) );
  NAND3XLTS U159 ( .A(n745), .B(n744), .C(n743), .Y(n1951) );
  NAND3XLTS U160 ( .A(n727), .B(n726), .C(n725), .Y(n1950) );
  NAND3XLTS U161 ( .A(n713), .B(n712), .C(n711), .Y(n1949) );
  NAND3XLTS U162 ( .A(n702), .B(n701), .C(n700), .Y(n1948) );
  NAND3XLTS U163 ( .A(n688), .B(n687), .C(n686), .Y(n1947) );
  NAND3XLTS U164 ( .A(n667), .B(n666), .C(n665), .Y(n1946) );
  NAND3XLTS U165 ( .A(n555), .B(n554), .C(n553), .Y(n1937) );
  NAND3XLTS U166 ( .A(n1785), .B(n1784), .C(n1783), .Y(n2107) );
  NAND3XLTS U167 ( .A(n1775), .B(n1774), .C(n1773), .Y(n2106) );
  NAND3XLTS U168 ( .A(n1768), .B(n1767), .C(n1766), .Y(n2105) );
  NAND3XLTS U169 ( .A(n1761), .B(n1760), .C(n1759), .Y(n2104) );
  NAND3XLTS U170 ( .A(n977), .B(n976), .C(n975), .Y(n1979) );
  NAND3XLTS U171 ( .A(n969), .B(n968), .C(n967), .Y(n1978) );
  NAND3XLTS U172 ( .A(n961), .B(n960), .C(n959), .Y(n1977) );
  NAND3XLTS U173 ( .A(n952), .B(n951), .C(n950), .Y(n1976) );
  NAND3XLTS U174 ( .A(n1690), .B(n1689), .C(n1688), .Y(n2071) );
  NAND3XLTS U175 ( .A(n1681), .B(n1680), .C(n1679), .Y(n2070) );
  NAND3XLTS U176 ( .A(n1674), .B(n1673), .C(n1672), .Y(n2069) );
  NAND3XLTS U177 ( .A(n1668), .B(n1667), .C(n1666), .Y(n2068) );
  NAND3XLTS U178 ( .A(n903), .B(n902), .C(n901), .Y(n1967) );
  NAND3XLTS U179 ( .A(n895), .B(n894), .C(n893), .Y(n1966) );
  NAND3XLTS U180 ( .A(n892), .B(n891), .C(n890), .Y(n1965) );
  NAND3XLTS U181 ( .A(n888), .B(n887), .C(n886), .Y(n1964) );
  NAND3XLTS U182 ( .A(n1661), .B(n1660), .C(n1659), .Y(n2059) );
  NAND3XLTS U183 ( .A(n1651), .B(n1650), .C(n1649), .Y(n2058) );
  NAND3XLTS U184 ( .A(n1644), .B(n1643), .C(n1642), .Y(n2057) );
  NAND3XLTS U185 ( .A(n1638), .B(n1637), .C(n1636), .Y(n2056) );
  NAND3XLTS U186 ( .A(n885), .B(n884), .C(n883), .Y(n1963) );
  NAND3XLTS U187 ( .A(n879), .B(n878), .C(n877), .Y(n1962) );
  NAND3XLTS U188 ( .A(n874), .B(n873), .C(n872), .Y(n1961) );
  NAND3XLTS U189 ( .A(n870), .B(n869), .C(n868), .Y(n1960) );
  NAND3XLTS U190 ( .A(n1107), .B(n1106), .C(n1105), .Y(n2003) );
  NAND3XLTS U191 ( .A(n1102), .B(n1101), .C(n1100), .Y(n2002) );
  NAND3XLTS U192 ( .A(n1097), .B(n1096), .C(n1095), .Y(n2001) );
  NAND3XLTS U193 ( .A(n1092), .B(n1091), .C(n1090), .Y(n2000) );
  NAND3XLTS U194 ( .A(n1088), .B(n1087), .C(n1086), .Y(n1999) );
  NAND3XLTS U195 ( .A(n1083), .B(n1082), .C(n1081), .Y(n1998) );
  NAND3XLTS U196 ( .A(n1422), .B(n1421), .C(n1420), .Y(n2021) );
  NAND3XLTS U197 ( .A(n1417), .B(n1416), .C(n1415), .Y(n2020) );
  NAND3XLTS U198 ( .A(n1410), .B(n1409), .C(n1408), .Y(n2019) );
  NAND3XLTS U199 ( .A(n1405), .B(n1404), .C(n1403), .Y(n2018) );
  NAND3XLTS U200 ( .A(n1400), .B(n1399), .C(n1398), .Y(n2017) );
  NAND3XLTS U201 ( .A(n1396), .B(n1395), .C(n1394), .Y(n2016) );
  NAND3XLTS U202 ( .A(n1457), .B(n1456), .C(n1455), .Y(n2027) );
  NAND3XLTS U203 ( .A(n1452), .B(n1451), .C(n1450), .Y(n2026) );
  NAND3XLTS U204 ( .A(n1445), .B(n1444), .C(n1443), .Y(n2025) );
  NAND3XLTS U205 ( .A(n1440), .B(n1439), .C(n1438), .Y(n2024) );
  NAND3XLTS U206 ( .A(n1434), .B(n1433), .C(n1432), .Y(n2023) );
  NAND3XLTS U207 ( .A(n1430), .B(n1429), .C(n1428), .Y(n2022) );
  NAND3XLTS U208 ( .A(n1890), .B(n1889), .C(n1888), .Y(n2143) );
  NAND3XLTS U209 ( .A(n1879), .B(n1878), .C(n1877), .Y(n2142) );
  NAND3XLTS U210 ( .A(n1869), .B(n1868), .C(n1867), .Y(n2141) );
  NAND3XLTS U211 ( .A(n1861), .B(n1860), .C(n1859), .Y(n2140) );
  NAND3XLTS U212 ( .A(n1051), .B(n1050), .C(n1049), .Y(n1991) );
  NAND3XLTS U213 ( .A(n1042), .B(n1041), .C(n1040), .Y(n1990) );
  NAND3XLTS U214 ( .A(n1037), .B(n1036), .C(n1035), .Y(n1989) );
  NAND3XLTS U215 ( .A(n1031), .B(n1030), .C(n1029), .Y(n1988) );
  NAND3XLTS U216 ( .A(n1851), .B(n1850), .C(n1849), .Y(n2131) );
  NAND3XLTS U217 ( .A(n1840), .B(n1839), .C(n1838), .Y(n2130) );
  NAND3XLTS U218 ( .A(n1829), .B(n1828), .C(n1827), .Y(n2129) );
  NAND3XLTS U219 ( .A(n1819), .B(n1818), .C(n1817), .Y(n2128) );
  NAND3XLTS U220 ( .A(n1025), .B(n1024), .C(n1023), .Y(n1987) );
  NAND3XLTS U221 ( .A(n1016), .B(n1015), .C(n1014), .Y(n1986) );
  NAND3XLTS U222 ( .A(n1009), .B(n1008), .C(n1007), .Y(n1985) );
  NAND3XLTS U223 ( .A(n1002), .B(n1001), .C(n1000), .Y(n1984) );
  NAND3XLTS U224 ( .A(n1753), .B(n1752), .C(n1751), .Y(n2095) );
  NAND3XLTS U225 ( .A(n1744), .B(n1743), .C(n1742), .Y(n2094) );
  NAND3XLTS U226 ( .A(n1737), .B(n1736), .C(n1735), .Y(n2093) );
  NAND3XLTS U227 ( .A(n1731), .B(n1730), .C(n1729), .Y(n2092) );
  NAND3XLTS U228 ( .A(n946), .B(n945), .C(n944), .Y(n1975) );
  NAND3XLTS U229 ( .A(n936), .B(n935), .C(n934), .Y(n1974) );
  NAND3XLTS U230 ( .A(n931), .B(n930), .C(n929), .Y(n1973) );
  NAND3XLTS U231 ( .A(n926), .B(n925), .C(n924), .Y(n1972) );
  NAND3XLTS U232 ( .A(n1724), .B(n1723), .C(n1722), .Y(n2083) );
  NAND3XLTS U233 ( .A(n1715), .B(n1714), .C(n1713), .Y(n2082) );
  NAND3XLTS U234 ( .A(n1707), .B(n1706), .C(n1705), .Y(n2081) );
  NAND3XLTS U235 ( .A(n1699), .B(n1698), .C(n1697), .Y(n2080) );
  NAND3XLTS U236 ( .A(n920), .B(n919), .C(n918), .Y(n1971) );
  NAND3XLTS U237 ( .A(n914), .B(n913), .C(n912), .Y(n1970) );
  NAND3XLTS U238 ( .A(n910), .B(n909), .C(n908), .Y(n1969) );
  NAND3XLTS U239 ( .A(n907), .B(n906), .C(n905), .Y(n1968) );
  NAND3XLTS U240 ( .A(n1365), .B(n1364), .C(n1363), .Y(n2009) );
  NAND3XLTS U241 ( .A(n1359), .B(n1358), .C(n1357), .Y(n2008) );
  NAND3XLTS U242 ( .A(n1354), .B(n1353), .C(n1352), .Y(n2007) );
  NAND3XLTS U243 ( .A(n1348), .B(n1347), .C(n1346), .Y(n2006) );
  NAND3XLTS U244 ( .A(n1343), .B(n1342), .C(n1341), .Y(n2005) );
  NAND3XLTS U245 ( .A(n1338), .B(n1337), .C(n1112), .Y(n2004) );
  NAND3XLTS U246 ( .A(n1389), .B(n1388), .C(n1387), .Y(n2015) );
  NAND3XLTS U247 ( .A(n1384), .B(n1383), .C(n1382), .Y(n2014) );
  NAND3XLTS U248 ( .A(n1380), .B(n1379), .C(n1378), .Y(n2013) );
  NAND3XLTS U249 ( .A(n1376), .B(n1375), .C(n1374), .Y(n2012) );
  NAND3XLTS U250 ( .A(n1373), .B(n1372), .C(n1371), .Y(n2011) );
  NAND3XLTS U251 ( .A(n1370), .B(n1369), .C(n1368), .Y(n2010) );
  NAND3XLTS U252 ( .A(n1497), .B(n1496), .C(n1495), .Y(n2033) );
  NAND3XLTS U253 ( .A(n1491), .B(n1490), .C(n1489), .Y(n2032) );
  NAND3XLTS U254 ( .A(n1483), .B(n1482), .C(n1481), .Y(n2031) );
  NAND3XLTS U255 ( .A(n1477), .B(n1476), .C(n1475), .Y(n2030) );
  NAND3XLTS U256 ( .A(n1471), .B(n1470), .C(n1469), .Y(n2029) );
  NAND3XLTS U257 ( .A(n1466), .B(n1465), .C(n1464), .Y(n2028) );
  NAND3XLTS U258 ( .A(n1542), .B(n1541), .C(n1540), .Y(n2039) );
  NAND3XLTS U259 ( .A(n1535), .B(n1534), .C(n1533), .Y(n2038) );
  NAND3XLTS U260 ( .A(n1528), .B(n1527), .C(n1526), .Y(n2037) );
  NAND3XLTS U261 ( .A(n1520), .B(n1519), .C(n1518), .Y(n2036) );
  NAND3XLTS U262 ( .A(n1511), .B(n1510), .C(n1509), .Y(n2035) );
  NAND3XLTS U263 ( .A(n1504), .B(n1503), .C(n1502), .Y(n2034) );
  NAND3XLTS U264 ( .A(n1810), .B(n1809), .C(n1808), .Y(n2119) );
  NAND3XLTS U265 ( .A(n1804), .B(n1803), .C(n1802), .Y(n2118) );
  NAND3XLTS U266 ( .A(n1797), .B(n1796), .C(n1795), .Y(n2117) );
  NAND3XLTS U267 ( .A(n1791), .B(n1790), .C(n1789), .Y(n2116) );
  NAND3XLTS U268 ( .A(n995), .B(n994), .C(n993), .Y(n1983) );
  NAND3XLTS U269 ( .A(n988), .B(n987), .C(n986), .Y(n1982) );
  NAND3XLTS U270 ( .A(n984), .B(n983), .C(n982), .Y(n1981) );
  NAND3XLTS U271 ( .A(n980), .B(n979), .C(n978), .Y(n1980) );
  NAND3XLTS U272 ( .A(n1077), .B(n1076), .C(n1075), .Y(n1997) );
  NAND3XLTS U273 ( .A(n1073), .B(n1072), .C(n1071), .Y(n1996) );
  NAND3XLTS U274 ( .A(n1067), .B(n1066), .C(n1065), .Y(n1995) );
  NAND3XLTS U275 ( .A(n1063), .B(n1062), .C(n1061), .Y(n1994) );
  NAND3XLTS U276 ( .A(n1059), .B(n1058), .C(n1057), .Y(n1993) );
  NAND3XLTS U277 ( .A(n1056), .B(n1055), .C(n1054), .Y(n1992) );
  OAI2BB2XLTS U278 ( .B0(n1920), .B1(n504), .A0N(n497), .A1N(n481), .Y(N2624)
         );
  AOI211XLTS U279 ( .A0(n480), .A1(n526), .B0(n479), .C0(n478), .Y(n481) );
  XOR2XLTS U280 ( .A(n525), .B(n492), .Y(n479) );
  OAI21XLTS U281 ( .A0(n480), .A1(n526), .B0(n477), .Y(n478) );
  OR2X1TS U282 ( .A(n176), .B(n1786), .Y(n981) );
  OR2X1TS U283 ( .A(n127), .B(n1754), .Y(n1366) );
  OR2X1TS U284 ( .A(n384), .B(n1852), .Y(n1032) );
  OR2X1TS U285 ( .A(n269), .B(n1725), .Y(n1390) );
  OR2X1TS U286 ( .A(n79), .B(n1662), .Y(n1458) );
  OR2X1TS U287 ( .A(n33), .B(n1634), .Y(n1498) );
  NAND2X1TS U288 ( .A(n27), .B(n25), .Y(n26) );
  NAND2X1TS U289 ( .A(n524), .B(n1920), .Y(n29) );
  OR2X1TS U290 ( .A(n1576), .B(n272), .Y(n3) );
  OR2X1TS U291 ( .A(n1622), .B(n388), .Y(n4) );
  OR2X1TS U292 ( .A(n1555), .B(n83), .Y(n5) );
  OR2X1TS U293 ( .A(n1591), .B(n130), .Y(n6) );
  OR2X1TS U294 ( .A(n1624), .B(n388), .Y(n7) );
  OR2X1TS U295 ( .A(n1577), .B(n272), .Y(n8) );
  OR2X1TS U296 ( .A(n218), .B(n1574), .Y(n10) );
  NOR3XLTS U297 ( .A(n1604), .B(n1599), .C(n178), .Y(n174) );
  NOR3XLTS U298 ( .A(n1618), .B(n1611), .C(n313), .Y(n309) );
  NOR3XLTS U299 ( .A(n1631), .B(n1625), .C(n387), .Y(n383) );
  OR2X1TS U300 ( .A(n219), .B(n1691), .Y(n1423) );
  INVX2TS U301 ( .A(n25), .Y(n28) );
  OR2X1TS U302 ( .A(n29), .B(n1632), .Y(n11) );
  NOR2XLTS U303 ( .A(n29), .B(n1594), .Y(n126) );
  AND3X1TS U304 ( .A(n539), .B(n1908), .C(n538), .Y(n12) );
  CLKBUFX2TS U305 ( .A(n1912), .Y(n13) );
  INVX2TS U321 ( .A(n1919), .Y(n475) );
  INVX2TS U322 ( .A(n1915), .Y(n493) );
  INVX2TS U323 ( .A(n15), .Y(n71) );
  INVX2TS U324 ( .A(n71), .Y(n116) );
  INVX2TS U325 ( .A(selectBit_WEST), .Y(n446) );
  INVX2TS U326 ( .A(n1549), .Y(n1551) );
  INVX2TS U327 ( .A(n1911), .Y(n449) );
  INVX2TS U328 ( .A(n2), .Y(n305) );
  INVX2TS U329 ( .A(selectBit_SOUTH), .Y(n507) );
  INVX2TS U330 ( .A(n9), .Y(n214) );
  INVX2TS U331 ( .A(n1919), .Y(n495) );
  INVX2TS U332 ( .A(n2), .Y(n18) );
  INVX2TS U333 ( .A(n1919), .Y(n484) );
  NAND2X1TS U334 ( .A(n18), .B(n484), .Y(n22) );
  INVX2TS U335 ( .A(n19), .Y(n75) );
  INVX2TS U336 ( .A(n75), .Y(n73) );
  INVX2TS U337 ( .A(n507), .Y(n506) );
  NAND2X1TS U338 ( .A(selectBit_SOUTH), .B(n21), .Y(n20) );
  NAND2X1TS U339 ( .A(n303), .B(n213), .Y(n119) );
  INVX2TS U340 ( .A(n1917), .Y(n266) );
  INVX2TS U341 ( .A(n1916), .Y(n443) );
  AOI22X1TS U342 ( .A0(n266), .A1(n22), .B0(n120), .B1(n443), .Y(n23) );
  INVX2TS U343 ( .A(n23), .Y(n24) );
  INVX2TS U344 ( .A(n24), .Y(n25) );
  INVX2TS U345 ( .A(n26), .Y(n115) );
  NAND2X1TS U346 ( .A(selectBit_EAST), .B(n118), .Y(n264) );
  NAND2X1TS U347 ( .A(n444), .B(n120), .Y(n30) );
  INVX2TS U348 ( .A(n446), .Y(n514) );
  INVX2TS U349 ( .A(readReady), .Y(n123) );
  INVX2TS U350 ( .A(n123), .Y(n513) );
  NAND2X1TS U351 ( .A(n539), .B(n508), .Y(n524) );
  INVX2TS U352 ( .A(n29), .Y(n121) );
  INVX2TS U353 ( .A(n121), .Y(n218) );
  INVX2TS U354 ( .A(n123), .Y(n511) );
  NAND2X1TS U355 ( .A(n33), .B(n1552), .Y(n35) );
  INVX2TS U356 ( .A(n31), .Y(n1512) );
  INVX2TS U357 ( .A(n1512), .Y(n875) );
  CLKBUFX2TS U358 ( .A(n875), .Y(n42) );
  INVX2TS U359 ( .A(n42), .Y(n60) );
  INVX2TS U360 ( .A(destinationAddressIn_EAST[8]), .Y(n234) );
  INVX2TS U361 ( .A(n121), .Y(n482) );
  INVX2TS U362 ( .A(n482), .Y(n379) );
  INVX2TS U363 ( .A(n32), .Y(n880) );
  INVX2TS U364 ( .A(n880), .Y(n1634) );
  INVX2TS U365 ( .A(n1498), .Y(n48) );
  OR2X1TS U366 ( .A(n1549), .B(n35), .Y(n46) );
  INVX2TS U367 ( .A(n46), .Y(n1523) );
  CLKBUFX2TS U368 ( .A(destinationAddressIn_WEST[8]), .Y(n400) );
  CLKBUFX2TS U369 ( .A(n400), .Y(n714) );
  AOI22X1TS U370 ( .A0(n48), .A1(\destinationAddressbuffer[7][8] ), .B0(n1523), 
        .B1(n714), .Y(n38) );
  NAND2BX1TS U371 ( .AN(n35), .B(n34), .Y(n36) );
  INVX2TS U372 ( .A(n156), .Y(n715) );
  OR2X1TS U373 ( .A(n1545), .B(n36), .Y(n55) );
  INVX2TS U374 ( .A(n55), .Y(n1531) );
  CLKBUFX2TS U375 ( .A(destinationAddressIn_NORTH[8]), .Y(n716) );
  CLKBUFX2TS U376 ( .A(n716), .Y(n332) );
  AOI22X1TS U377 ( .A0(n43), .A1(n715), .B0(n1531), .B1(n332), .Y(n37) );
  OAI211XLTS U378 ( .A0(n60), .A1(n234), .B0(n38), .C0(n37), .Y(n2064) );
  INVX2TS U379 ( .A(n42), .Y(n65) );
  INVX2TS U380 ( .A(destinationAddressIn_EAST[10]), .Y(n217) );
  INVX2TS U381 ( .A(n46), .Y(n1656) );
  CLKBUFX2TS U382 ( .A(destinationAddressIn_WEST[10]), .Y(n385) );
  CLKBUFX2TS U383 ( .A(n385), .Y(n746) );
  AOI22X1TS U384 ( .A0(n48), .A1(\destinationAddressbuffer[7][10] ), .B0(n1656), .B1(n746), .Y(n41) );
  INVX2TS U385 ( .A(n39), .Y(n62) );
  INVX2TS U386 ( .A(n62), .Y(n1648) );
  INVX2TS U387 ( .A(n160), .Y(n749) );
  INVX2TS U388 ( .A(n55), .Y(n871) );
  CLKBUFX2TS U389 ( .A(destinationAddressIn_NORTH[10]), .Y(n750) );
  CLKBUFX2TS U390 ( .A(n750), .Y(n318) );
  AOI22X1TS U391 ( .A0(n1648), .A1(n749), .B0(n871), .B1(n318), .Y(n40) );
  OAI211XLTS U392 ( .A0(n65), .A1(n217), .B0(n41), .C0(n40), .Y(n2066) );
  INVX2TS U393 ( .A(destinationAddressIn_EAST[9]), .Y(n226) );
  INVX2TS U394 ( .A(n46), .Y(n1647) );
  INVX2TS U395 ( .A(n1647), .Y(n1505) );
  INVX2TS U396 ( .A(n1505), .Y(n61) );
  CLKBUFX2TS U397 ( .A(destinationAddressIn_WEST[9]), .Y(n394) );
  CLKBUFX2TS U398 ( .A(n394), .Y(n729) );
  AOI22X1TS U399 ( .A0(n48), .A1(\destinationAddressbuffer[7][9] ), .B0(n61), 
        .B1(n729), .Y(n45) );
  INVX2TS U400 ( .A(n62), .Y(n43) );
  INVX2TS U401 ( .A(n43), .Y(n882) );
  INVX2TS U402 ( .A(n882), .Y(n68) );
  INVX2TS U403 ( .A(n166), .Y(n730) );
  CLKBUFX2TS U404 ( .A(destinationAddressIn_NORTH[9]), .Y(n732) );
  CLKBUFX2TS U405 ( .A(n732), .Y(n324) );
  AOI22X1TS U406 ( .A0(n68), .A1(n730), .B0(n49), .B1(n324), .Y(n44) );
  OAI211XLTS U407 ( .A0(n60), .A1(n226), .B0(n45), .C0(n44), .Y(n2065) );
  INVX2TS U408 ( .A(destinationAddressIn_EAST[11]), .Y(n230) );
  INVX2TS U409 ( .A(n46), .Y(n47) );
  CLKBUFX2TS U410 ( .A(destinationAddressIn_WEST[11]), .Y(n406) );
  CLKBUFX2TS U411 ( .A(n406), .Y(n762) );
  AOI22X1TS U412 ( .A0(n48), .A1(\destinationAddressbuffer[7][11] ), .B0(n47), 
        .B1(n762), .Y(n51) );
  INVX2TS U413 ( .A(n152), .Y(n765) );
  INVX2TS U414 ( .A(n55), .Y(n49) );
  INVX2TS U415 ( .A(n49), .Y(n876) );
  INVX2TS U416 ( .A(n876), .Y(n67) );
  CLKBUFX2TS U417 ( .A(destinationAddressIn_NORTH[11]), .Y(n766) );
  CLKBUFX2TS U418 ( .A(n766), .Y(n340) );
  AOI22X1TS U419 ( .A0(n43), .A1(n765), .B0(n67), .B1(n340), .Y(n50) );
  OAI211XLTS U420 ( .A0(n60), .A1(n230), .B0(n51), .C0(n50), .Y(n2067) );
  INVX2TS U421 ( .A(writeIn_EAST), .Y(n241) );
  CLKBUFX2TS U422 ( .A(n1498), .Y(n881) );
  INVX2TS U423 ( .A(n881), .Y(n1652) );
  INVX2TS U424 ( .A(n1505), .Y(n52) );
  CLKBUFX2TS U425 ( .A(writeIn_WEST), .Y(n415) );
  CLKBUFX2TS U426 ( .A(n415), .Y(n543) );
  AOI22X1TS U427 ( .A0(n1652), .A1(writeOutbuffer[7]), .B0(n52), .B1(n543), 
        .Y(n54) );
  INVX2TS U428 ( .A(n62), .Y(n1658) );
  INVX2TS U429 ( .A(writeIn_SOUTH), .Y(n171) );
  INVX2TS U430 ( .A(n171), .Y(n545) );
  CLKBUFX2TS U431 ( .A(writeIn_NORTH), .Y(n546) );
  CLKBUFX2TS U432 ( .A(n546), .Y(n345) );
  AOI22X1TS U433 ( .A0(n1658), .A1(n545), .B0(n871), .B1(n345), .Y(n53) );
  OAI211XLTS U434 ( .A0(n65), .A1(n241), .B0(n54), .C0(n53), .Y(n2040) );
  INVX2TS U435 ( .A(destinationAddressIn_EAST[4]), .Y(n249) );
  INVX2TS U436 ( .A(n881), .Y(n66) );
  AOI22X1TS U437 ( .A0(n66), .A1(\destinationAddressbuffer[7][4] ), .B0(n1656), 
        .B1(destinationAddressIn_WEST[4]), .Y(n57) );
  INVX2TS U438 ( .A(destinationAddressIn_SOUTH[4]), .Y(n133) );
  INVX2TS U439 ( .A(n133), .Y(n659) );
  INVX2TS U440 ( .A(n55), .Y(n1657) );
  AOI22X1TS U441 ( .A0(n1648), .A1(n659), .B0(n1657), .B1(
        destinationAddressIn_NORTH[4]), .Y(n56) );
  OAI211XLTS U442 ( .A0(n65), .A1(n249), .B0(n57), .C0(n56), .Y(n2060) );
  INVX2TS U443 ( .A(destinationAddressIn_EAST[7]), .Y(n245) );
  AOI22X1TS U444 ( .A0(n66), .A1(\destinationAddressbuffer[7][7] ), .B0(n1523), 
        .B1(destinationAddressIn_WEST[7]), .Y(n59) );
  INVX2TS U445 ( .A(destinationAddressIn_SOUTH[7]), .Y(n149) );
  INVX2TS U446 ( .A(n149), .Y(n704) );
  AOI22X1TS U447 ( .A0(n1658), .A1(n704), .B0(n1657), .B1(
        destinationAddressIn_NORTH[7]), .Y(n58) );
  OAI211XLTS U448 ( .A0(n60), .A1(n245), .B0(n59), .C0(n58), .Y(n2063) );
  INVX2TS U449 ( .A(destinationAddressIn_EAST[6]), .Y(n254) );
  AOI22X1TS U450 ( .A0(n66), .A1(\destinationAddressbuffer[7][6] ), .B0(n61), 
        .B1(destinationAddressIn_WEST[6]), .Y(n64) );
  INVX2TS U451 ( .A(n62), .Y(n1517) );
  INVX2TS U452 ( .A(destinationAddressIn_SOUTH[6]), .Y(n144) );
  INVX2TS U453 ( .A(n144), .Y(n691) );
  AOI22X1TS U454 ( .A0(n1517), .A1(n691), .B0(n67), .B1(
        destinationAddressIn_NORTH[6]), .Y(n63) );
  OAI211XLTS U455 ( .A0(n65), .A1(n254), .B0(n64), .C0(n63), .Y(n2062) );
  INVX2TS U456 ( .A(destinationAddressIn_EAST[5]), .Y(n258) );
  AOI22X1TS U457 ( .A0(n66), .A1(\destinationAddressbuffer[7][5] ), .B0(n47), 
        .B1(destinationAddressIn_WEST[5]), .Y(n70) );
  INVX2TS U458 ( .A(destinationAddressIn_SOUTH[5]), .Y(n137) );
  INVX2TS U459 ( .A(n137), .Y(n671) );
  AOI22X1TS U460 ( .A0(n68), .A1(n671), .B0(n67), .B1(
        destinationAddressIn_NORTH[5]), .Y(n69) );
  OAI211XLTS U461 ( .A0(n1512), .A1(n258), .B0(n70), .C0(n69), .Y(n2061) );
  INVX2TS U462 ( .A(n72), .Y(n172) );
  NAND2X1TS U463 ( .A(n117), .B(n451), .Y(n263) );
  AOI21X1TS U464 ( .A0(n214), .A1(n73), .B0(n303), .Y(n377) );
  NOR3XLTS U465 ( .A(n377), .B(n264), .C(n213), .Y(n1558) );
  INVX2TS U466 ( .A(n1919), .Y(n487) );
  NOR2XLTS U467 ( .A(n456), .B(n505), .Y(n378) );
  NOR3XLTS U468 ( .A(n23), .B(n74), .C(n73), .Y(n1555) );
  AOI31XLTS U469 ( .A0(n444), .A1(n487), .A2(n378), .B0(n1555), .Y(n76) );
  INVX2TS U470 ( .A(n121), .Y(n441) );
  AOI21X1TS U471 ( .A0(n81), .A1(n76), .B0(n441), .Y(n79) );
  INVX2TS U472 ( .A(n1911), .Y(n382) );
  NAND2X1TS U473 ( .A(n79), .B(n1562), .Y(n82) );
  INVX2TS U474 ( .A(n1472), .Y(n899) );
  CLKBUFX2TS U475 ( .A(n899), .Y(n89) );
  INVX2TS U476 ( .A(n89), .Y(n104) );
  INVX2TS U477 ( .A(n78), .Y(n896) );
  INVX2TS U478 ( .A(n896), .Y(n1662) );
  CLKBUFX2TS U479 ( .A(n1458), .Y(n897) );
  INVX2TS U480 ( .A(n897), .Y(n93) );
  OR2X1TS U481 ( .A(n1559), .B(n82), .Y(n92) );
  INVX2TS U482 ( .A(n92), .Y(n80) );
  INVX2TS U483 ( .A(n80), .Y(n898) );
  INVX2TS U484 ( .A(n898), .Y(n109) );
  AOI22X1TS U485 ( .A0(n93), .A1(\destinationAddressbuffer[6][11] ), .B0(n109), 
        .B1(n762), .Y(n86) );
  INVX2TS U486 ( .A(n5), .Y(n1687) );
  CLKBUFX2TS U487 ( .A(n766), .Y(n408) );
  INVX2TS U488 ( .A(n84), .Y(n96) );
  INVX2TS U489 ( .A(n96), .Y(n1462) );
  INVX2TS U490 ( .A(n152), .Y(n339) );
  AOI22X1TS U491 ( .A0(n1687), .A1(n408), .B0(n1462), .B1(n339), .Y(n85) );
  OAI211XLTS U492 ( .A0(n104), .A1(n230), .B0(n86), .C0(n85), .Y(n2079) );
  INVX2TS U493 ( .A(n92), .Y(n1663) );
  AOI22X1TS U494 ( .A0(n93), .A1(\destinationAddressbuffer[6][10] ), .B0(n1663), .B1(n746), .Y(n88) );
  INVX2TS U495 ( .A(n5), .Y(n1463) );
  CLKBUFX2TS U496 ( .A(n750), .Y(n390) );
  INVX2TS U497 ( .A(n84), .Y(n900) );
  INVX2TS U498 ( .A(n900), .Y(n105) );
  INVX2TS U499 ( .A(n160), .Y(n317) );
  AOI22X1TS U500 ( .A0(n1463), .A1(n390), .B0(n105), .B1(n317), .Y(n87) );
  OAI211XLTS U501 ( .A0(n104), .A1(n217), .B0(n88), .C0(n87), .Y(n2078) );
  INVX2TS U502 ( .A(n89), .Y(n114) );
  INVX2TS U503 ( .A(n92), .Y(n1684) );
  AOI22X1TS U504 ( .A0(n93), .A1(\destinationAddressbuffer[6][9] ), .B0(n80), 
        .B1(n729), .Y(n91) );
  CLKBUFX2TS U505 ( .A(n732), .Y(n395) );
  INVX2TS U506 ( .A(n900), .Y(n1686) );
  INVX2TS U507 ( .A(n166), .Y(n323) );
  AOI22X1TS U508 ( .A0(n106), .A1(n395), .B0(n1686), .B1(n323), .Y(n90) );
  OAI211XLTS U509 ( .A0(n114), .A1(n226), .B0(n91), .C0(n90), .Y(n2077) );
  INVX2TS U510 ( .A(n92), .Y(n1460) );
  AOI22X1TS U511 ( .A0(n93), .A1(\destinationAddressbuffer[6][8] ), .B0(n1460), 
        .B1(n714), .Y(n95) );
  INVX2TS U512 ( .A(n5), .Y(n1665) );
  CLKBUFX2TS U513 ( .A(n716), .Y(n402) );
  INVX2TS U514 ( .A(n156), .Y(n331) );
  AOI22X1TS U515 ( .A0(n1665), .A1(n402), .B0(n105), .B1(n331), .Y(n94) );
  OAI211XLTS U516 ( .A0(n104), .A1(n234), .B0(n95), .C0(n94), .Y(n2076) );
  INVX2TS U517 ( .A(n897), .Y(n1682) );
  AOI22X1TS U518 ( .A0(n1682), .A1(writeOutbuffer[6]), .B0(n109), .B1(n543), 
        .Y(n98) );
  CLKBUFX2TS U519 ( .A(n546), .Y(n416) );
  INVX2TS U520 ( .A(n171), .Y(n344) );
  AOI22X1TS U521 ( .A0(n1463), .A1(n416), .B0(n84), .B1(n344), .Y(n97) );
  OAI211XLTS U522 ( .A0(n114), .A1(n241), .B0(n98), .C0(n97), .Y(n2041) );
  INVX2TS U523 ( .A(n1458), .Y(n110) );
  AOI22X1TS U524 ( .A0(n110), .A1(\destinationAddressbuffer[6][7] ), .B0(n1460), .B1(destinationAddressIn_WEST[7]), .Y(n101) );
  INVX2TS U525 ( .A(n5), .Y(n99) );
  INVX2TS U526 ( .A(n99), .Y(n889) );
  INVX2TS U527 ( .A(n889), .Y(n106) );
  CLKBUFX2TS U528 ( .A(destinationAddressIn_NORTH[7]), .Y(n357) );
  CLKBUFX2TS U529 ( .A(n357), .Y(n424) );
  INVX2TS U530 ( .A(n149), .Y(n356) );
  AOI22X1TS U531 ( .A0(n106), .A1(n424), .B0(n84), .B1(n356), .Y(n100) );
  OAI211XLTS U532 ( .A0(n114), .A1(n245), .B0(n101), .C0(n100), .Y(n2075) );
  AOI22X1TS U533 ( .A0(n110), .A1(\destinationAddressbuffer[6][6] ), .B0(n1684), .B1(destinationAddressIn_WEST[6]), .Y(n103) );
  CLKBUFX2TS U534 ( .A(destinationAddressIn_NORTH[6]), .Y(n351) );
  CLKBUFX2TS U535 ( .A(n351), .Y(n435) );
  INVX2TS U536 ( .A(n144), .Y(n349) );
  AOI22X1TS U537 ( .A0(n106), .A1(n435), .B0(n1678), .B1(n349), .Y(n102) );
  OAI211XLTS U538 ( .A0(n104), .A1(n254), .B0(n103), .C0(n102), .Y(n2074) );
  AOI22X1TS U539 ( .A0(n110), .A1(\destinationAddressbuffer[6][4] ), .B0(n1663), .B1(destinationAddressIn_WEST[4]), .Y(n108) );
  CLKBUFX2TS U540 ( .A(destinationAddressIn_NORTH[4]), .Y(n364) );
  CLKBUFX2TS U541 ( .A(n364), .Y(n420) );
  INVX2TS U542 ( .A(n133), .Y(n363) );
  AOI22X1TS U543 ( .A0(n106), .A1(n420), .B0(n105), .B1(n363), .Y(n107) );
  OAI211XLTS U544 ( .A0(n1472), .A1(n249), .B0(n108), .C0(n107), .Y(n2072) );
  AOI22X1TS U545 ( .A0(n110), .A1(\destinationAddressbuffer[6][5] ), .B0(n109), 
        .B1(destinationAddressIn_WEST[5]), .Y(n113) );
  CLKBUFX2TS U546 ( .A(destinationAddressIn_NORTH[5]), .Y(n370) );
  CLKBUFX2TS U547 ( .A(n370), .Y(n430) );
  INVX2TS U548 ( .A(n96), .Y(n111) );
  INVX2TS U549 ( .A(n137), .Y(n369) );
  AOI22X1TS U550 ( .A0(n1687), .A1(n430), .B0(n111), .B1(n369), .Y(n112) );
  OAI211XLTS U551 ( .A0(n114), .A1(n258), .B0(n113), .C0(n112), .Y(n2073) );
  INVX2TS U552 ( .A(n115), .Y(n1587) );
  INVX2TS U553 ( .A(n512), .Y(n515) );
  INVX2TS U554 ( .A(n1916), .Y(n483) );
  NAND2X1TS U555 ( .A(n120), .B(n483), .Y(n122) );
  INVX2TS U556 ( .A(n121), .Y(n306) );
  AOI31X1TS U557 ( .A0(n124), .A1(n1587), .A2(n122), .B0(n306), .Y(n127) );
  INVX2TS U558 ( .A(n123), .Y(n510) );
  INVX2TS U559 ( .A(n1916), .Y(n486) );
  NAND2BX1TS U560 ( .AN(n130), .B(n124), .Y(n129) );
  INVX2TS U561 ( .A(n125), .Y(n964) );
  INVX2TS U562 ( .A(n964), .Y(n1765) );
  CLKBUFX2TS U563 ( .A(n1765), .Y(n138) );
  INVX2TS U564 ( .A(n138), .Y(n161) );
  INVX2TS U565 ( .A(n126), .Y(n971) );
  INVX2TS U566 ( .A(n971), .Y(n1754) );
  CLKBUFX2TS U567 ( .A(n1366), .Y(n168) );
  INVX2TS U568 ( .A(n168), .Y(n145) );
  NOR3XLTS U569 ( .A(n1593), .B(n1588), .C(n130), .Y(n139) );
  INVX2TS U570 ( .A(n139), .Y(n153) );
  INVX2TS U571 ( .A(n153), .Y(n128) );
  AOI22X1TS U572 ( .A0(n145), .A1(\destinationAddressbuffer[3][4] ), .B0(n162), 
        .B1(destinationAddressIn_EAST[4]), .Y(n132) );
  OR2X1TS U573 ( .A(n115), .B(n129), .Y(n157) );
  INVX2TS U574 ( .A(n157), .Y(n1782) );
  INVX2TS U575 ( .A(n6), .Y(n1386) );
  CLKBUFX2TS U576 ( .A(destinationAddressIn_WEST[4]), .Y(n657) );
  CLKBUFX2TS U577 ( .A(n657), .Y(n361) );
  AOI22X1TS U578 ( .A0(n1782), .A1(n364), .B0(n1386), .B1(n361), .Y(n131) );
  OAI211XLTS U579 ( .A0(n161), .A1(n133), .B0(n132), .C0(n131), .Y(n2108) );
  INVX2TS U580 ( .A(n138), .Y(n167) );
  INVX2TS U581 ( .A(n153), .Y(n1770) );
  AOI22X1TS U582 ( .A0(n145), .A1(\destinationAddressbuffer[3][5] ), .B0(n1770), .B1(destinationAddressIn_EAST[5]), .Y(n136) );
  INVX2TS U583 ( .A(n146), .Y(n965) );
  INVX2TS U584 ( .A(n6), .Y(n134) );
  CLKBUFX2TS U585 ( .A(destinationAddressIn_WEST[5]), .Y(n669) );
  CLKBUFX2TS U586 ( .A(n669), .Y(n367) );
  AOI22X1TS U587 ( .A0(n965), .A1(n370), .B0(n134), .B1(n367), .Y(n135) );
  OAI211XLTS U588 ( .A0(n167), .A1(n137), .B0(n136), .C0(n135), .Y(n2109) );
  INVX2TS U589 ( .A(n954), .Y(n162) );
  AOI22X1TS U590 ( .A0(n145), .A1(\destinationAddressbuffer[3][6] ), .B0(n162), 
        .B1(destinationAddressIn_EAST[6]), .Y(n143) );
  INVX2TS U591 ( .A(n157), .Y(n140) );
  INVX2TS U592 ( .A(n140), .Y(n146) );
  INVX2TS U593 ( .A(n146), .Y(n957) );
  INVX2TS U594 ( .A(n6), .Y(n1757) );
  INVX2TS U595 ( .A(n1757), .Y(n972) );
  INVX2TS U596 ( .A(n972), .Y(n141) );
  CLKBUFX2TS U597 ( .A(destinationAddressIn_WEST[6]), .Y(n689) );
  CLKBUFX2TS U598 ( .A(n689), .Y(n348) );
  AOI22X1TS U599 ( .A0(n957), .A1(n351), .B0(n141), .B1(n348), .Y(n142) );
  OAI211XLTS U600 ( .A0(n161), .A1(n144), .B0(n143), .C0(n142), .Y(n2110) );
  INVX2TS U601 ( .A(n153), .Y(n1778) );
  AOI22X1TS U602 ( .A0(n145), .A1(\destinationAddressbuffer[3][7] ), .B0(n1778), .B1(destinationAddressIn_EAST[7]), .Y(n148) );
  INVX2TS U603 ( .A(n6), .Y(n1780) );
  CLKBUFX2TS U604 ( .A(destinationAddressIn_WEST[7]), .Y(n703) );
  CLKBUFX2TS U605 ( .A(n703), .Y(n354) );
  AOI22X1TS U606 ( .A0(n965), .A1(n357), .B0(n1780), .B1(n354), .Y(n147) );
  OAI211XLTS U607 ( .A0(n161), .A1(n149), .B0(n148), .C0(n147), .Y(n2111) );
  INVX2TS U608 ( .A(n168), .Y(n163) );
  AOI22X1TS U609 ( .A0(n163), .A1(\destinationAddressbuffer[3][11] ), .B0(
        n1770), .B1(destinationAddressIn_EAST[11]), .Y(n151) );
  CLKBUFX2TS U610 ( .A(n406), .Y(n336) );
  AOI22X1TS U611 ( .A0(n1782), .A1(n340), .B0(n134), .B1(n336), .Y(n150) );
  OAI211XLTS U612 ( .A0(n167), .A1(n152), .B0(n151), .C0(n150), .Y(n2115) );
  INVX2TS U613 ( .A(n153), .Y(n1381) );
  AOI22X1TS U614 ( .A0(n163), .A1(\destinationAddressbuffer[3][8] ), .B0(n1381), .B1(destinationAddressIn_EAST[8]), .Y(n155) );
  INVX2TS U615 ( .A(n157), .Y(n1758) );
  CLKBUFX2TS U616 ( .A(n400), .Y(n329) );
  AOI22X1TS U617 ( .A0(n1758), .A1(n332), .B0(n1757), .B1(n329), .Y(n154) );
  OAI211XLTS U618 ( .A0(n964), .A1(n156), .B0(n155), .C0(n154), .Y(n2112) );
  AOI22X1TS U619 ( .A0(n163), .A1(\destinationAddressbuffer[3][10] ), .B0(
        n1381), .B1(destinationAddressIn_EAST[10]), .Y(n159) );
  INVX2TS U620 ( .A(n157), .Y(n1367) );
  CLKBUFX2TS U621 ( .A(n385), .Y(n311) );
  AOI22X1TS U622 ( .A0(n1367), .A1(n318), .B0(n1386), .B1(n311), .Y(n158) );
  OAI211XLTS U623 ( .A0(n161), .A1(n160), .B0(n159), .C0(n158), .Y(n2114) );
  AOI22X1TS U624 ( .A0(n163), .A1(\destinationAddressbuffer[3][9] ), .B0(n162), 
        .B1(destinationAddressIn_EAST[9]), .Y(n165) );
  INVX2TS U625 ( .A(n972), .Y(n955) );
  CLKBUFX2TS U626 ( .A(n394), .Y(n321) );
  AOI22X1TS U627 ( .A0(n965), .A1(n324), .B0(n955), .B1(n321), .Y(n164) );
  OAI211XLTS U628 ( .A0(n167), .A1(n166), .B0(n165), .C0(n164), .Y(n2113) );
  INVX2TS U629 ( .A(n168), .Y(n1776) );
  AOI22X1TS U630 ( .A0(n1776), .A1(writeOutbuffer[3]), .B0(n1778), .B1(
        writeIn_EAST), .Y(n170) );
  CLKBUFX2TS U631 ( .A(n415), .Y(n343) );
  AOI22X1TS U632 ( .A0(n1367), .A1(n345), .B0(n1780), .B1(n343), .Y(n169) );
  OAI211XLTS U633 ( .A0(n167), .A1(n171), .B0(n170), .C0(n169), .Y(n2044) );
  NOR3XLTS U634 ( .A(n377), .B(n213), .C(n376), .Y(n1601) );
  AOI31XLTS U635 ( .A0(n495), .A1(n378), .A2(n443), .B0(n1598), .Y(n173) );
  NAND2X1TS U636 ( .A(n176), .B(n1605), .Y(n178) );
  INVX2TS U637 ( .A(n174), .Y(n1344) );
  INVX2TS U638 ( .A(n1344), .Y(n991) );
  CLKBUFX2TS U639 ( .A(n991), .Y(n187) );
  INVX2TS U640 ( .A(n187), .Y(n205) );
  INVX2TS U641 ( .A(n175), .Y(n989) );
  INVX2TS U642 ( .A(n989), .Y(n1786) );
  INVX2TS U643 ( .A(n981), .Y(n192) );
  OR2X1TS U644 ( .A(n1602), .B(n178), .Y(n191) );
  INVX2TS U645 ( .A(n191), .Y(n1787) );
  AOI22X1TS U646 ( .A0(n192), .A1(\destinationAddressbuffer[2][10] ), .B0(
        n1787), .B1(n311), .Y(n183) );
  INVX2TS U647 ( .A(n188), .Y(n201) );
  INVX2TS U648 ( .A(n201), .Y(n1111) );
  INVX2TS U649 ( .A(n180), .Y(n195) );
  INVX2TS U650 ( .A(n195), .Y(n181) );
  INVX2TS U651 ( .A(n181), .Y(n992) );
  INVX2TS U652 ( .A(n992), .Y(n206) );
  AOI22X1TS U653 ( .A0(n1111), .A1(n318), .B0(n206), .B1(n317), .Y(n182) );
  OAI211XLTS U654 ( .A0(n205), .A1(n217), .B0(n183), .C0(n182), .Y(n2126) );
  INVX2TS U655 ( .A(n191), .Y(n184) );
  INVX2TS U656 ( .A(n184), .Y(n990) );
  INVX2TS U657 ( .A(n990), .Y(n198) );
  AOI22X1TS U658 ( .A0(n192), .A1(\destinationAddressbuffer[2][11] ), .B0(n198), .B1(n336), .Y(n186) );
  INVX2TS U659 ( .A(n201), .Y(n1807) );
  INVX2TS U660 ( .A(n195), .Y(n1110) );
  AOI22X1TS U661 ( .A0(n1807), .A1(n340), .B0(n1110), .B1(n339), .Y(n185) );
  OAI211XLTS U662 ( .A0(n205), .A1(n230), .B0(n186), .C0(n185), .Y(n2127) );
  INVX2TS U663 ( .A(n187), .Y(n212) );
  INVX2TS U664 ( .A(n191), .Y(n1806) );
  AOI22X1TS U665 ( .A0(n192), .A1(\destinationAddressbuffer[2][9] ), .B0(n1806), .B1(n321), .Y(n190) );
  INVX2TS U666 ( .A(n188), .Y(n1340) );
  INVX2TS U667 ( .A(n1340), .Y(n985) );
  AOI22X1TS U668 ( .A0(n985), .A1(n324), .B0(n1110), .B1(n323), .Y(n189) );
  OAI211XLTS U669 ( .A0(n212), .A1(n226), .B0(n190), .C0(n189), .Y(n2125) );
  INVX2TS U670 ( .A(n191), .Y(n1109) );
  AOI22X1TS U671 ( .A0(n192), .A1(\destinationAddressbuffer[2][8] ), .B0(n1109), .B1(n329), .Y(n194) );
  INVX2TS U672 ( .A(n201), .Y(n1788) );
  INVX2TS U673 ( .A(n195), .Y(n1351) );
  AOI22X1TS U674 ( .A0(n1788), .A1(n332), .B0(n1351), .B1(n331), .Y(n193) );
  OAI211XLTS U675 ( .A0(n205), .A1(n234), .B0(n194), .C0(n193), .Y(n2124) );
  CLKBUFX2TS U676 ( .A(n981), .Y(n1606) );
  INVX2TS U677 ( .A(n1606), .Y(n1805) );
  AOI22X1TS U678 ( .A0(n1805), .A1(writeOutbuffer[2]), .B0(n198), .B1(n343), 
        .Y(n197) );
  INVX2TS U679 ( .A(n195), .Y(n1362) );
  AOI22X1TS U680 ( .A0(n1111), .A1(n345), .B0(n1362), .B1(n344), .Y(n196) );
  OAI211XLTS U681 ( .A0(n212), .A1(n241), .B0(n197), .C0(n196), .Y(n2045) );
  INVX2TS U682 ( .A(n981), .Y(n209) );
  AOI22X1TS U683 ( .A0(n209), .A1(\destinationAddressbuffer[2][5] ), .B0(n198), 
        .B1(n367), .Y(n200) );
  AOI22X1TS U684 ( .A0(n1807), .A1(destinationAddressIn_NORTH[5]), .B0(n206), 
        .B1(n369), .Y(n199) );
  OAI211XLTS U685 ( .A0(n212), .A1(n258), .B0(n200), .C0(n199), .Y(n2121) );
  AOI22X1TS U686 ( .A0(n209), .A1(\destinationAddressbuffer[2][7] ), .B0(n1109), .B1(n354), .Y(n204) );
  INVX2TS U687 ( .A(n201), .Y(n202) );
  AOI22X1TS U688 ( .A0(n202), .A1(destinationAddressIn_NORTH[7]), .B0(n1362), 
        .B1(n356), .Y(n203) );
  OAI211XLTS U689 ( .A0(n205), .A1(n245), .B0(n204), .C0(n203), .Y(n2123) );
  AOI22X1TS U690 ( .A0(n209), .A1(\destinationAddressbuffer[2][4] ), .B0(n1787), .B1(n361), .Y(n208) );
  AOI22X1TS U691 ( .A0(n202), .A1(destinationAddressIn_NORTH[4]), .B0(n206), 
        .B1(n363), .Y(n207) );
  OAI211XLTS U692 ( .A0(n1344), .A1(n249), .B0(n208), .C0(n207), .Y(n2120) );
  AOI22X1TS U693 ( .A0(n209), .A1(\destinationAddressbuffer[2][6] ), .B0(n184), 
        .B1(n348), .Y(n211) );
  AOI22X1TS U694 ( .A0(n985), .A1(destinationAddressIn_NORTH[6]), .B0(n1351), 
        .B1(n349), .Y(n210) );
  OAI211XLTS U695 ( .A0(n212), .A1(n254), .B0(n211), .C0(n210), .Y(n2122) );
  INVX2TS U696 ( .A(n213), .Y(n304) );
  INVX2TS U697 ( .A(n1914), .Y(n381) );
  INVX2TS U698 ( .A(n1914), .Y(n308) );
  NAND2X1TS U699 ( .A(n219), .B(n1574), .Y(n221) );
  INVX2TS U700 ( .A(n216), .Y(n1435) );
  INVX2TS U701 ( .A(n1435), .Y(n917) );
  CLKBUFX2TS U702 ( .A(n917), .Y(n229) );
  INVX2TS U703 ( .A(n229), .Y(n253) );
  CLKBUFX2TS U704 ( .A(n217), .Y(n393) );
  INVX2TS U705 ( .A(n10), .Y(n1691) );
  CLKBUFX2TS U706 ( .A(n1423), .Y(n915) );
  INVX2TS U707 ( .A(n915), .Y(n237) );
  OR2X1TS U708 ( .A(n1571), .B(n221), .Y(n235) );
  INVX2TS U709 ( .A(n235), .Y(n1424) );
  AOI22X1TS U710 ( .A0(n237), .A1(\destinationAddressbuffer[5][10] ), .B0(
        n1424), .B1(n746), .Y(n225) );
  INVX2TS U711 ( .A(n1564), .Y(n1567) );
  NAND2BX1TS U712 ( .AN(n221), .B(n220), .Y(n223) );
  INVX2TS U713 ( .A(n246), .Y(n1696) );
  INVX2TS U714 ( .A(n1696), .Y(n260) );
  INVX2TS U715 ( .A(n260), .Y(n911) );
  OR2X1TS U716 ( .A(n1564), .B(n223), .Y(n242) );
  INVX2TS U717 ( .A(n242), .Y(n1447) );
  AOI22X1TS U718 ( .A0(n911), .A1(n390), .B0(n1447), .B1(n317), .Y(n224) );
  OAI211XLTS U719 ( .A0(n253), .A1(n393), .B0(n225), .C0(n224), .Y(n2090) );
  INVX2TS U720 ( .A(n229), .Y(n257) );
  CLKBUFX2TS U721 ( .A(n226), .Y(n398) );
  INVX2TS U722 ( .A(n235), .Y(n1720) );
  AOI22X1TS U723 ( .A0(n237), .A1(\destinationAddressbuffer[5][9] ), .B0(n1720), .B1(n729), .Y(n228) );
  INVX2TS U724 ( .A(n246), .Y(n1427) );
  INVX2TS U725 ( .A(n242), .Y(n1695) );
  AOI22X1TS U726 ( .A0(n1427), .A1(n395), .B0(n1695), .B1(n323), .Y(n227) );
  OAI211XLTS U727 ( .A0(n257), .A1(n398), .B0(n228), .C0(n227), .Y(n2089) );
  CLKBUFX2TS U728 ( .A(n230), .Y(n412) );
  INVX2TS U729 ( .A(n235), .Y(n1694) );
  AOI22X1TS U730 ( .A0(n237), .A1(\destinationAddressbuffer[5][11] ), .B0(
        n1694), .B1(n762), .Y(n233) );
  INVX2TS U731 ( .A(n246), .Y(n1449) );
  INVX2TS U732 ( .A(n242), .Y(n231) );
  INVX2TS U733 ( .A(n231), .Y(n904) );
  INVX2TS U734 ( .A(n904), .Y(n238) );
  AOI22X1TS U735 ( .A0(n1449), .A1(n408), .B0(n238), .B1(n339), .Y(n232) );
  OAI211XLTS U736 ( .A0(n253), .A1(n412), .B0(n233), .C0(n232), .Y(n2091) );
  CLKBUFX2TS U737 ( .A(n234), .Y(n405) );
  INVX2TS U738 ( .A(n235), .Y(n236) );
  INVX2TS U739 ( .A(n236), .Y(n916) );
  INVX2TS U740 ( .A(n916), .Y(n250) );
  AOI22X1TS U741 ( .A0(n237), .A1(\destinationAddressbuffer[5][8] ), .B0(n250), 
        .B1(n714), .Y(n240) );
  AOI22X1TS U742 ( .A0(n1437), .A1(n402), .B0(n238), .B1(n331), .Y(n239) );
  OAI211XLTS U743 ( .A0(n253), .A1(n405), .B0(n240), .C0(n239), .Y(n2088) );
  CLKBUFX2TS U744 ( .A(n241), .Y(n419) );
  INVX2TS U745 ( .A(n915), .Y(n1716) );
  AOI22X1TS U746 ( .A0(n1716), .A1(writeOutbuffer[5]), .B0(n250), .B1(n543), 
        .Y(n244) );
  INVX2TS U747 ( .A(n242), .Y(n1425) );
  AOI22X1TS U748 ( .A0(n1427), .A1(n416), .B0(n1425), .B1(n344), .Y(n243) );
  OAI211XLTS U749 ( .A0(n257), .A1(n419), .B0(n244), .C0(n243), .Y(n2042) );
  CLKBUFX2TS U750 ( .A(n245), .Y(n427) );
  INVX2TS U751 ( .A(n1423), .Y(n259) );
  AOI22X1TS U752 ( .A0(n259), .A1(\destinationAddressbuffer[5][7] ), .B0(n1694), .B1(n703), .Y(n248) );
  INVX2TS U753 ( .A(n246), .Y(n1437) );
  AOI22X1TS U754 ( .A0(n1437), .A1(n424), .B0(n1425), .B1(n356), .Y(n247) );
  OAI211XLTS U755 ( .A0(n257), .A1(n427), .B0(n248), .C0(n247), .Y(n2087) );
  CLKBUFX2TS U756 ( .A(n249), .Y(n423) );
  AOI22X1TS U757 ( .A0(n259), .A1(\destinationAddressbuffer[5][4] ), .B0(n250), 
        .B1(n657), .Y(n252) );
  AOI22X1TS U758 ( .A0(n1449), .A1(n420), .B0(n238), .B1(n363), .Y(n251) );
  OAI211XLTS U759 ( .A0(n253), .A1(n423), .B0(n252), .C0(n251), .Y(n2084) );
  CLKBUFX2TS U760 ( .A(n254), .Y(n439) );
  AOI22X1TS U761 ( .A0(n259), .A1(\destinationAddressbuffer[5][6] ), .B0(n236), 
        .B1(n689), .Y(n256) );
  AOI22X1TS U762 ( .A0(n1696), .A1(n435), .B0(n231), .B1(n349), .Y(n255) );
  OAI211XLTS U763 ( .A0(n257), .A1(n439), .B0(n256), .C0(n255), .Y(n2086) );
  CLKBUFX2TS U764 ( .A(n258), .Y(n433) );
  AOI22X1TS U765 ( .A0(n259), .A1(\destinationAddressbuffer[5][5] ), .B0(n1424), .B1(n669), .Y(n262) );
  INVX2TS U766 ( .A(n260), .Y(n1704) );
  AOI22X1TS U767 ( .A0(n1704), .A1(n430), .B0(n1447), .B1(n369), .Y(n261) );
  OAI211XLTS U768 ( .A0(n1435), .A1(n433), .B0(n262), .C0(n261), .Y(n2085) );
  INVX2TS U769 ( .A(n304), .Y(n375) );
  AOI31XLTS U770 ( .A0(n444), .A1(n378), .A2(n308), .B0(n1577), .Y(n265) );
  NAND2X1TS U771 ( .A(n269), .B(n1585), .Y(n271) );
  INVX2TS U772 ( .A(n267), .Y(n1401) );
  INVX2TS U773 ( .A(n1401), .Y(n940) );
  CLKBUFX2TS U774 ( .A(n940), .Y(n278) );
  INVX2TS U775 ( .A(n278), .Y(n294) );
  INVX2TS U776 ( .A(n268), .Y(n937) );
  INVX2TS U777 ( .A(n937), .Y(n1725) );
  CLKBUFX2TS U778 ( .A(n1390), .Y(n938) );
  INVX2TS U779 ( .A(n938), .Y(n284) );
  OR2X1TS U780 ( .A(n1581), .B(n271), .Y(n282) );
  INVX2TS U781 ( .A(n282), .Y(n1748) );
  AOI22X1TS U782 ( .A0(n284), .A1(\destinationAddressbuffer[4][9] ), .B0(n1748), .B1(n321), .Y(n274) );
  INVX2TS U783 ( .A(n3), .Y(n1750) );
  INVX2TS U784 ( .A(n8), .Y(n1749) );
  AOI22X1TS U785 ( .A0(n1750), .A1(n730), .B0(n275), .B1(n395), .Y(n273) );
  OAI211XLTS U786 ( .A0(n294), .A1(n398), .B0(n274), .C0(n273), .Y(n2101) );
  INVX2TS U787 ( .A(n278), .Y(n298) );
  INVX2TS U788 ( .A(n282), .Y(n1726) );
  AOI22X1TS U789 ( .A0(n284), .A1(\destinationAddressbuffer[4][11] ), .B0(
        n1726), .B1(n336), .Y(n277) );
  INVX2TS U790 ( .A(n3), .Y(n1741) );
  INVX2TS U791 ( .A(n8), .Y(n275) );
  INVX2TS U792 ( .A(n275), .Y(n279) );
  INVX2TS U793 ( .A(n279), .Y(n1413) );
  AOI22X1TS U794 ( .A0(n1741), .A1(n765), .B0(n1413), .B1(n408), .Y(n276) );
  OAI211XLTS U795 ( .A0(n298), .A1(n412), .B0(n277), .C0(n276), .Y(n2103) );
  INVX2TS U796 ( .A(n282), .Y(n1392) );
  AOI22X1TS U797 ( .A0(n284), .A1(\destinationAddressbuffer[4][10] ), .B0(
        n1392), .B1(n311), .Y(n281) );
  INVX2TS U798 ( .A(n279), .Y(n922) );
  AOI22X1TS U799 ( .A0(n300), .A1(n749), .B0(n922), .B1(n390), .Y(n280) );
  OAI211XLTS U800 ( .A0(n294), .A1(n393), .B0(n281), .C0(n280), .Y(n2102) );
  INVX2TS U801 ( .A(n282), .Y(n283) );
  INVX2TS U802 ( .A(n283), .Y(n939) );
  INVX2TS U803 ( .A(n939), .Y(n295) );
  AOI22X1TS U804 ( .A0(n284), .A1(\destinationAddressbuffer[4][8] ), .B0(n295), 
        .B1(n329), .Y(n287) );
  INVX2TS U805 ( .A(n3), .Y(n285) );
  INVX2TS U806 ( .A(n285), .Y(n942) );
  INVX2TS U807 ( .A(n942), .Y(n300) );
  INVX2TS U808 ( .A(n8), .Y(n1727) );
  AOI22X1TS U809 ( .A0(n300), .A1(n715), .B0(n1727), .B1(n402), .Y(n286) );
  OAI211XLTS U810 ( .A0(n294), .A1(n405), .B0(n287), .C0(n286), .Y(n2100) );
  INVX2TS U811 ( .A(n938), .Y(n1745) );
  AOI22X1TS U812 ( .A0(n1745), .A1(writeOutbuffer[4]), .B0(n295), .B1(n343), 
        .Y(n289) );
  INVX2TS U813 ( .A(n3), .Y(n1414) );
  INVX2TS U814 ( .A(n8), .Y(n1393) );
  AOI22X1TS U815 ( .A0(n1414), .A1(n545), .B0(n1393), .B1(n416), .Y(n288) );
  OAI211XLTS U816 ( .A0(n298), .A1(n419), .B0(n289), .C0(n288), .Y(n2043) );
  INVX2TS U817 ( .A(n1390), .Y(n299) );
  AOI22X1TS U818 ( .A0(n299), .A1(\destinationAddressbuffer[4][5] ), .B0(n1392), .B1(n367), .Y(n291) );
  AOI22X1TS U819 ( .A0(n1414), .A1(n671), .B0(n922), .B1(n430), .Y(n290) );
  OAI211XLTS U820 ( .A0(n298), .A1(n433), .B0(n291), .C0(n290), .Y(n2097) );
  AOI22X1TS U821 ( .A0(n299), .A1(\destinationAddressbuffer[4][7] ), .B0(n1726), .B1(n354), .Y(n293) );
  AOI22X1TS U822 ( .A0(n285), .A1(n704), .B0(n1393), .B1(n424), .Y(n292) );
  OAI211XLTS U823 ( .A0(n294), .A1(n427), .B0(n293), .C0(n292), .Y(n2099) );
  AOI22X1TS U824 ( .A0(n299), .A1(\destinationAddressbuffer[4][4] ), .B0(n295), 
        .B1(n361), .Y(n297) );
  AOI22X1TS U825 ( .A0(n285), .A1(n659), .B0(n1727), .B1(n420), .Y(n296) );
  OAI211XLTS U826 ( .A0(n298), .A1(n423), .B0(n297), .C0(n296), .Y(n2096) );
  AOI22X1TS U827 ( .A0(n299), .A1(\destinationAddressbuffer[4][6] ), .B0(n283), 
        .B1(n348), .Y(n302) );
  AOI22X1TS U828 ( .A0(n300), .A1(n691), .B0(n275), .B1(n435), .Y(n301) );
  OAI211XLTS U829 ( .A0(n1401), .A1(n439), .B0(n302), .C0(n301), .Y(n2098) );
  AOI31XLTS U830 ( .A0(n305), .A1(n381), .A2(n483), .B0(n1610), .Y(n307) );
  NAND2X1TS U831 ( .A(n310), .B(n1619), .Y(n313) );
  INVX2TS U832 ( .A(n309), .Y(n1089) );
  INVX2TS U833 ( .A(n1089), .Y(n1018) );
  CLKBUFX2TS U834 ( .A(n1018), .Y(n327) );
  INVX2TS U835 ( .A(n327), .Y(n360) );
  OR2X1TS U836 ( .A(n441), .B(n1619), .Y(n1084) );
  INVX2TS U837 ( .A(n1084), .Y(n1842) );
  OR2X1TS U838 ( .A(n310), .B(n1842), .Y(n1003) );
  INVX2TS U839 ( .A(n1003), .Y(n337) );
  OR2X1TS U840 ( .A(n1615), .B(n313), .Y(n335) );
  INVX2TS U841 ( .A(n335), .Y(n1078) );
  AOI22X1TS U842 ( .A0(n337), .A1(\destinationAddressbuffer[1][10] ), .B0(
        n1078), .B1(n311), .Y(n320) );
  INVX2TS U843 ( .A(n322), .Y(n355) );
  INVX2TS U844 ( .A(n355), .Y(n314) );
  INVX2TS U845 ( .A(n316), .Y(n338) );
  INVX2TS U846 ( .A(n338), .Y(n1094) );
  AOI22X1TS U847 ( .A0(n314), .A1(n318), .B0(n1094), .B1(n317), .Y(n319) );
  OAI211XLTS U848 ( .A0(n360), .A1(n393), .B0(n320), .C0(n319), .Y(n2138) );
  INVX2TS U849 ( .A(n335), .Y(n1845) );
  AOI22X1TS U850 ( .A0(n337), .A1(\destinationAddressbuffer[1][9] ), .B0(n1845), .B1(n321), .Y(n326) );
  INVX2TS U851 ( .A(n322), .Y(n1085) );
  INVX2TS U852 ( .A(n1085), .Y(n1011) );
  INVX2TS U853 ( .A(n338), .Y(n1079) );
  AOI22X1TS U854 ( .A0(n1011), .A1(n324), .B0(n350), .B1(n323), .Y(n325) );
  OAI211XLTS U855 ( .A0(n360), .A1(n398), .B0(n326), .C0(n325), .Y(n2137) );
  INVX2TS U856 ( .A(n327), .Y(n373) );
  INVX2TS U857 ( .A(n335), .Y(n328) );
  INVX2TS U858 ( .A(n328), .Y(n1017) );
  INVX2TS U859 ( .A(n1017), .Y(n362) );
  AOI22X1TS U860 ( .A0(n337), .A1(\destinationAddressbuffer[1][8] ), .B0(n362), 
        .B1(n329), .Y(n334) );
  INVX2TS U861 ( .A(n355), .Y(n1848) );
  INVX2TS U862 ( .A(n338), .Y(n330) );
  INVX2TS U863 ( .A(n330), .Y(n1020) );
  INVX2TS U864 ( .A(n1020), .Y(n350) );
  AOI22X1TS U865 ( .A0(n1848), .A1(n332), .B0(n350), .B1(n331), .Y(n333) );
  OAI211XLTS U866 ( .A0(n373), .A1(n405), .B0(n334), .C0(n333), .Y(n2136) );
  INVX2TS U867 ( .A(n335), .Y(n1813) );
  AOI22X1TS U868 ( .A0(n337), .A1(\destinationAddressbuffer[1][11] ), .B0(
        n1813), .B1(n336), .Y(n342) );
  INVX2TS U869 ( .A(n338), .Y(n1104) );
  AOI22X1TS U870 ( .A0(n314), .A1(n340), .B0(n1104), .B1(n339), .Y(n341) );
  OAI211XLTS U871 ( .A0(n360), .A1(n412), .B0(n342), .C0(n341), .Y(n2139) );
  CLKBUFX2TS U872 ( .A(n1003), .Y(n1620) );
  INVX2TS U873 ( .A(n1620), .Y(n1841) );
  AOI22X1TS U874 ( .A0(n1841), .A1(writeOutbuffer[1]), .B0(n362), .B1(n343), 
        .Y(n347) );
  INVX2TS U875 ( .A(n355), .Y(n1816) );
  AOI22X1TS U876 ( .A0(n1816), .A1(n345), .B0(n1094), .B1(n344), .Y(n346) );
  OAI211XLTS U877 ( .A0(n373), .A1(n419), .B0(n347), .C0(n346), .Y(n2046) );
  INVX2TS U878 ( .A(n1003), .Y(n368) );
  AOI22X1TS U879 ( .A0(n368), .A1(\destinationAddressbuffer[1][6] ), .B0(n328), 
        .B1(n348), .Y(n353) );
  AOI22X1TS U880 ( .A0(n1011), .A1(n351), .B0(n350), .B1(n349), .Y(n352) );
  OAI211XLTS U881 ( .A0(n373), .A1(n439), .B0(n353), .C0(n352), .Y(n2134) );
  AOI22X1TS U882 ( .A0(n368), .A1(\destinationAddressbuffer[1][7] ), .B0(n1813), .B1(n354), .Y(n359) );
  INVX2TS U883 ( .A(n355), .Y(n1080) );
  AOI22X1TS U884 ( .A0(n1080), .A1(n357), .B0(n1079), .B1(n356), .Y(n358) );
  OAI211XLTS U885 ( .A0(n360), .A1(n427), .B0(n359), .C0(n358), .Y(n2135) );
  AOI22X1TS U886 ( .A0(n368), .A1(\destinationAddressbuffer[1][4] ), .B0(n362), 
        .B1(n361), .Y(n366) );
  AOI22X1TS U887 ( .A0(n1848), .A1(n364), .B0(n1104), .B1(n363), .Y(n365) );
  OAI211XLTS U888 ( .A0(n1089), .A1(n423), .B0(n366), .C0(n365), .Y(n2132) );
  AOI22X1TS U889 ( .A0(n368), .A1(\destinationAddressbuffer[1][5] ), .B0(n1078), .B1(n367), .Y(n372) );
  AOI22X1TS U890 ( .A0(n1080), .A1(n370), .B0(n1079), .B1(n369), .Y(n371) );
  OAI211XLTS U891 ( .A0(n373), .A1(n433), .B0(n372), .C0(n371), .Y(n2133) );
  AOI31XLTS U892 ( .A0(n378), .A1(n381), .A2(n486), .B0(n1624), .Y(n380) );
  NAND2X1TS U893 ( .A(n384), .B(n1632), .Y(n387) );
  INVX2TS U894 ( .A(n383), .Y(n1060) );
  INVX2TS U895 ( .A(n1060), .Y(n1045) );
  CLKBUFX2TS U896 ( .A(n1045), .Y(n399) );
  INVX2TS U897 ( .A(n399), .Y(n428) );
  INVX2TS U898 ( .A(n11), .Y(n1852) );
  CLKBUFX2TS U899 ( .A(n1032), .Y(n1043) );
  INVX2TS U900 ( .A(n1043), .Y(n407) );
  OR2X1TS U901 ( .A(n1629), .B(n387), .Y(n413) );
  INVX2TS U902 ( .A(n413), .Y(n1854) );
  AOI22X1TS U903 ( .A0(n407), .A1(\destinationAddressbuffer[0][10] ), .B0(
        n1854), .B1(n385), .Y(n392) );
  INVX2TS U904 ( .A(n7), .Y(n389) );
  INVX2TS U905 ( .A(n389), .Y(n1027) );
  INVX2TS U906 ( .A(n1027), .Y(n409) );
  AOI22X1TS U907 ( .A0(n401), .A1(n749), .B0(n409), .B1(n390), .Y(n391) );
  OAI211XLTS U908 ( .A0(n428), .A1(n393), .B0(n392), .C0(n391), .Y(n2150) );
  INVX2TS U909 ( .A(n413), .Y(n1883) );
  AOI22X1TS U910 ( .A0(n407), .A1(\destinationAddressbuffer[0][9] ), .B0(n414), 
        .B1(n394), .Y(n397) );
  INVX2TS U911 ( .A(n4), .Y(n1887) );
  INVX2TS U912 ( .A(n7), .Y(n1885) );
  AOI22X1TS U913 ( .A0(n1887), .A1(n730), .B0(n389), .B1(n395), .Y(n396) );
  OAI211XLTS U914 ( .A0(n428), .A1(n398), .B0(n397), .C0(n396), .Y(n2149) );
  INVX2TS U915 ( .A(n399), .Y(n440) );
  INVX2TS U916 ( .A(n413), .Y(n1052) );
  AOI22X1TS U917 ( .A0(n407), .A1(\destinationAddressbuffer[0][8] ), .B0(n1052), .B1(n400), .Y(n404) );
  INVX2TS U918 ( .A(n4), .Y(n401) );
  INVX2TS U919 ( .A(n401), .Y(n1047) );
  INVX2TS U920 ( .A(n1047), .Y(n436) );
  INVX2TS U921 ( .A(n7), .Y(n1856) );
  AOI22X1TS U922 ( .A0(n436), .A1(n715), .B0(n1856), .B1(n402), .Y(n403) );
  OAI211XLTS U923 ( .A0(n440), .A1(n405), .B0(n404), .C0(n403), .Y(n2148) );
  AOI22X1TS U924 ( .A0(n407), .A1(\destinationAddressbuffer[0][11] ), .B0(n429), .B1(n406), .Y(n411) );
  INVX2TS U925 ( .A(n4), .Y(n1876) );
  AOI22X1TS U926 ( .A0(n1876), .A1(n765), .B0(n409), .B1(n408), .Y(n410) );
  OAI211XLTS U927 ( .A0(n428), .A1(n412), .B0(n411), .C0(n410), .Y(n2151) );
  INVX2TS U928 ( .A(n1032), .Y(n1880) );
  INVX2TS U929 ( .A(n413), .Y(n414) );
  INVX2TS U930 ( .A(n414), .Y(n1044) );
  INVX2TS U931 ( .A(n1044), .Y(n429) );
  AOI22X1TS U932 ( .A0(n1880), .A1(writeOutbuffer[0]), .B0(n429), .B1(n415), 
        .Y(n418) );
  INVX2TS U933 ( .A(n4), .Y(n1070) );
  INVX2TS U934 ( .A(n7), .Y(n1053) );
  AOI22X1TS U935 ( .A0(n1070), .A1(n545), .B0(n1053), .B1(n416), .Y(n417) );
  OAI211XLTS U936 ( .A0(n440), .A1(n419), .B0(n418), .C0(n417), .Y(n2047) );
  INVX2TS U937 ( .A(n1032), .Y(n434) );
  AOI22X1TS U938 ( .A0(n434), .A1(\destinationAddressbuffer[0][4] ), .B0(n1854), .B1(destinationAddressIn_WEST[4]), .Y(n422) );
  AOI22X1TS U939 ( .A0(n401), .A1(n659), .B0(n1856), .B1(n420), .Y(n421) );
  OAI211XLTS U940 ( .A0(n440), .A1(n423), .B0(n422), .C0(n421), .Y(n2144) );
  AOI22X1TS U941 ( .A0(n434), .A1(\destinationAddressbuffer[0][7] ), .B0(n1052), .B1(destinationAddressIn_WEST[7]), .Y(n426) );
  AOI22X1TS U942 ( .A0(n401), .A1(n704), .B0(n1053), .B1(n424), .Y(n425) );
  OAI211XLTS U943 ( .A0(n428), .A1(n427), .B0(n426), .C0(n425), .Y(n2147) );
  AOI22X1TS U944 ( .A0(n434), .A1(\destinationAddressbuffer[0][5] ), .B0(n429), 
        .B1(destinationAddressIn_WEST[5]), .Y(n432) );
  AOI22X1TS U945 ( .A0(n1070), .A1(n671), .B0(n409), .B1(n430), .Y(n431) );
  OAI211XLTS U946 ( .A0(n1060), .A1(n433), .B0(n432), .C0(n431), .Y(n2145) );
  AOI22X1TS U947 ( .A0(n434), .A1(\destinationAddressbuffer[0][6] ), .B0(n1883), .B1(destinationAddressIn_WEST[6]), .Y(n438) );
  AOI22X1TS U948 ( .A0(n436), .A1(n691), .B0(n389), .B1(n435), .Y(n437) );
  OAI211XLTS U949 ( .A0(n440), .A1(n439), .B0(n438), .C0(n437), .Y(n2146) );
  INVX2TS U950 ( .A(reset), .Y(n491) );
  NAND2X1TS U951 ( .A(n491), .B(n1908), .Y(n504) );
  INVX2TS U952 ( .A(n1912), .Y(n531) );
  INVX2TS U953 ( .A(n1914), .Y(n452) );
  INVX2TS U954 ( .A(n1915), .Y(n456) );
  INVX2TS U955 ( .A(n1906), .Y(n442) );
  NAND2X1TS U956 ( .A(n456), .B(n442), .Y(n455) );
  INVX2TS U957 ( .A(n1917), .Y(n444) );
  INVX2TS U958 ( .A(n1909), .Y(n527) );
  INVX2TS U959 ( .A(n1910), .Y(n530) );
  AOI22X1TS U960 ( .A0(n444), .A1(n527), .B0(n530), .B1(n443), .Y(n447) );
  INVX2TS U961 ( .A(n446), .Y(n451) );
  INVX2TS U962 ( .A(n466), .Y(n463) );
  INVX2TS U963 ( .A(n1918), .Y(n528) );
  AOI21X1TS U964 ( .A0(n528), .A1(n449), .B0(n448), .Y(n462) );
  ADDHX1TS U965 ( .A(n454), .B(n453), .CO(n466), .S(n468) );
  INVX2TS U966 ( .A(n468), .Y(n457) );
  OAI21XLTS U967 ( .A0(n456), .A1(n1918), .B0(n455), .Y(n488) );
  AOI21X1TS U968 ( .A0(n458), .A1(n457), .B0(n488), .Y(n460) );
  OAI22X1TS U969 ( .A0(n458), .A1(n457), .B0(n464), .B1(n463), .Y(n459) );
  AOI21X1TS U970 ( .A0(n467), .A1(n460), .B0(n459), .Y(n461) );
  AOI211X1TS U971 ( .A0(n464), .A1(n463), .B0(n462), .C0(n461), .Y(n465) );
  NAND2X1TS U972 ( .A(n469), .B(n466), .Y(n472) );
  XNOR2X1TS U973 ( .A(n1916), .B(n470), .Y(n471) );
  INVX2TS U974 ( .A(n496), .Y(n480) );
  INVX2TS U975 ( .A(n1910), .Y(n526) );
  INVX2TS U976 ( .A(n1918), .Y(n525) );
  ADDHXLTS U977 ( .A(n456), .B(n473), .CO(n476), .S(n492) );
  XNOR2X1TS U978 ( .A(n1913), .B(n494), .Y(n477) );
  NAND2X1TS U979 ( .A(n525), .B(n531), .Y(n529) );
  OAI21XLTS U980 ( .A0(n528), .A1(n1913), .B0(n529), .Y(n503) );
  INVX2TS U981 ( .A(n1909), .Y(n532) );
  NOR2XLTS U982 ( .A(n529), .B(n527), .Y(n835) );
  CLKBUFX2TS U983 ( .A(n835), .Y(n795) );
  CLKBUFX2TS U984 ( .A(n795), .Y(n815) );
  AOI21X1TS U985 ( .A0(n529), .A1(n532), .B0(n815), .Y(n500) );
  OAI22X1TS U986 ( .A0(n484), .A1(n503), .B0(n483), .B1(n500), .Y(n485) );
  AOI221XLTS U987 ( .A0(n503), .A1(n487), .B0(n486), .B1(n500), .C0(n485), .Y(
        n489) );
  AOI21X1TS U988 ( .A0(n489), .A1(n488), .B0(n1908), .Y(n490) );
  CLKBUFX2TS U989 ( .A(n1907), .Y(n641) );
  CLKBUFX2TS U990 ( .A(n641), .Y(n608) );
  NAND2X1TS U991 ( .A(n491), .B(n608), .Y(n502) );
  AOI22X1TS U992 ( .A0(n1906), .A1(n504), .B0(n502), .B1(n442), .Y(n1929) );
  INVX2TS U993 ( .A(n500), .Y(n501) );
  OAI22X1TS U994 ( .A0(n532), .A1(n504), .B0(n501), .B1(n502), .Y(n1934) );
  OAI22X1TS U995 ( .A0(n13), .A1(n504), .B0(n503), .B1(n502), .Y(n1935) );
  CLKBUFX2TS U996 ( .A(readIn_SOUTH), .Y(n1623) );
  CLKBUFX2TS U997 ( .A(n1623), .Y(n1566) );
  CLKBUFX2TS U998 ( .A(n1907), .Y(n841) );
  CLKBUFX2TS U999 ( .A(n544), .Y(n847) );
  CLKBUFX2TS U1000 ( .A(readIn_WEST), .Y(n1583) );
  CLKBUFX2TS U1001 ( .A(n1583), .Y(n1617) );
  INVX2TS U1002 ( .A(n1907), .Y(n521) );
  NOR4XLTS U1003 ( .A(readReady), .B(n515), .C(n446), .D(n509), .Y(n614) );
  CLKBUFX2TS U1004 ( .A(n614), .Y(n628) );
  CLKBUFX2TS U1005 ( .A(n628), .Y(n808) );
  CLKBUFX2TS U1006 ( .A(n808), .Y(n565) );
  AOI22X1TS U1007 ( .A0(n1566), .A1(n847), .B0(n1617), .B1(n565), .Y(n542) );
  CLKBUFX2TS U1008 ( .A(readIn_NORTH), .Y(n1597) );
  CLKBUFX2TS U1009 ( .A(n1597), .Y(n1565) );
  CLKBUFX2TS U1010 ( .A(n690), .Y(n564) );
  NOR4XLTS U1011 ( .A(n514), .B(n510), .C(n512), .D(n509), .Y(n590) );
  CLKBUFX2TS U1012 ( .A(n590), .Y(n601) );
  CLKBUFX2TS U1013 ( .A(n601), .Y(n776) );
  CLKBUFX2TS U1014 ( .A(n776), .Y(n825) );
  AOI22X1TS U1015 ( .A0(n1565), .A1(n564), .B0(readIn_EAST), .B1(n825), .Y(
        n541) );
  NOR3XLTS U1016 ( .A(n515), .B(n511), .C(n446), .Y(n517) );
  NOR3XLTS U1017 ( .A(n514), .B(n513), .C(n512), .Y(n516) );
  NAND4XLTS U1018 ( .A(n521), .B(n520), .C(n519), .D(n518), .Y(n733) );
  INVX2TS U1019 ( .A(n733), .Y(n522) );
  INVX2TS U1020 ( .A(n522), .Y(n581) );
  INVX2TS U1021 ( .A(n581), .Y(n523) );
  NOR3XLTS U1022 ( .A(n525), .B(n526), .C(n1912), .Y(n717) );
  CLKBUFX2TS U1023 ( .A(n717), .Y(n629) );
  CLKBUFX2TS U1024 ( .A(n629), .Y(n567) );
  NOR3XLTS U1025 ( .A(n528), .B(n1913), .C(n526), .Y(n692) );
  CLKBUFX2TS U1026 ( .A(n692), .Y(n630) );
  CLKBUFX2TS U1027 ( .A(n630), .Y(n566) );
  AOI22X1TS U1028 ( .A0(readOutbuffer[2]), .A1(n567), .B0(readOutbuffer[0]), 
        .B1(n566), .Y(n536) );
  NOR3XLTS U1029 ( .A(n525), .B(n13), .C(n527), .Y(n718) );
  CLKBUFX2TS U1030 ( .A(n718), .Y(n631) );
  CLKBUFX2TS U1031 ( .A(n631), .Y(n569) );
  NOR3XLTS U1032 ( .A(n528), .B(n531), .C(n532), .Y(n693) );
  CLKBUFX2TS U1033 ( .A(n693), .Y(n632) );
  CLKBUFX2TS U1034 ( .A(n632), .Y(n568) );
  AOI22X1TS U1035 ( .A0(readOutbuffer[6]), .A1(n569), .B0(readOutbuffer[4]), 
        .B1(n568), .Y(n535) );
  NOR2XLTS U1036 ( .A(n530), .B(n529), .Y(n719) );
  CLKBUFX2TS U1037 ( .A(n719), .Y(n633) );
  CLKBUFX2TS U1038 ( .A(n633), .Y(n571) );
  NOR3XLTS U1039 ( .A(n531), .B(n530), .C(n1918), .Y(n694) );
  CLKBUFX2TS U1040 ( .A(n694), .Y(n634) );
  CLKBUFX2TS U1041 ( .A(n634), .Y(n570) );
  AOI22X1TS U1042 ( .A0(readOutbuffer[3]), .A1(n571), .B0(readOutbuffer[1]), 
        .B1(n570), .Y(n534) );
  CLKBUFX2TS U1043 ( .A(n835), .Y(n856) );
  NOR3XLTS U1044 ( .A(n1913), .B(n442), .C(n532), .Y(n857) );
  CLKBUFX2TS U1045 ( .A(n857), .Y(n635) );
  CLKBUFX2TS U1046 ( .A(n635), .Y(n572) );
  AOI22X1TS U1047 ( .A0(readOutbuffer[7]), .A1(n856), .B0(readOutbuffer[5]), 
        .B1(n572), .Y(n533) );
  NAND4XLTS U1048 ( .A(n536), .B(n535), .C(n534), .D(n533), .Y(n537) );
  AOI22X1TS U1049 ( .A0(readOut), .A1(n552), .B0(n608), .B1(n537), .Y(n540) );
  INVX2TS U1050 ( .A(n12), .Y(n802) );
  CLKBUFX2TS U1051 ( .A(n776), .Y(n747) );
  AOI22X1TS U1052 ( .A0(writeIn_EAST), .A1(n747), .B0(n543), .B1(n565), .Y(
        n555) );
  CLKBUFX2TS U1053 ( .A(n544), .Y(n670) );
  CLKBUFX2TS U1054 ( .A(n670), .Y(n764) );
  AOI22X1TS U1055 ( .A0(n546), .A1(n564), .B0(n545), .B1(n764), .Y(n554) );
  AOI22X1TS U1056 ( .A0(writeOutbuffer[2]), .A1(n567), .B0(writeOutbuffer[0]), 
        .B1(n566), .Y(n550) );
  AOI22X1TS U1057 ( .A0(writeOutbuffer[6]), .A1(n569), .B0(writeOutbuffer[4]), 
        .B1(n568), .Y(n549) );
  AOI22X1TS U1058 ( .A0(writeOutbuffer[3]), .A1(n571), .B0(writeOutbuffer[1]), 
        .B1(n570), .Y(n548) );
  AOI22X1TS U1059 ( .A0(writeOutbuffer[7]), .A1(n856), .B0(writeOutbuffer[5]), 
        .B1(n572), .Y(n547) );
  NAND4XLTS U1060 ( .A(n550), .B(n549), .C(n548), .D(n547), .Y(n551) );
  AOI22X1TS U1061 ( .A0(writeOut), .A1(n552), .B0(n608), .B1(n551), .Y(n553)
         );
  CLKBUFX2TS U1062 ( .A(requesterAddressIn_NORTH[0]), .Y(n998) );
  CLKBUFX2TS U1063 ( .A(requesterAddressIn_EAST[0]), .Y(n1026) );
  CLKBUFX2TS U1064 ( .A(n1026), .Y(n997) );
  AOI22X1TS U1065 ( .A0(n998), .A1(n564), .B0(n997), .B1(n601), .Y(n563) );
  CLKBUFX2TS U1066 ( .A(requesterAddressIn_SOUTH[0]), .Y(n1028) );
  CLKBUFX2TS U1067 ( .A(n1028), .Y(n999) );
  CLKBUFX2TS U1068 ( .A(n670), .Y(n658) );
  CLKBUFX2TS U1069 ( .A(requesterAddressIn_WEST[0]), .Y(n921) );
  CLKBUFX2TS U1070 ( .A(n921), .Y(n948) );
  AOI22X1TS U1071 ( .A0(n999), .A1(n658), .B0(n948), .B1(n565), .Y(n562) );
  INVX2TS U1072 ( .A(n733), .Y(n685) );
  CLKBUFX2TS U1073 ( .A(n641), .Y(n596) );
  AOI22X1TS U1074 ( .A0(\requesterAddressbuffer[2][0] ), .A1(n567), .B0(
        \requesterAddressbuffer[0][0] ), .B1(n566), .Y(n559) );
  AOI22X1TS U1075 ( .A0(\requesterAddressbuffer[6][0] ), .A1(n569), .B0(
        \requesterAddressbuffer[4][0] ), .B1(n568), .Y(n558) );
  AOI22X1TS U1076 ( .A0(\requesterAddressbuffer[3][0] ), .A1(n571), .B0(
        \requesterAddressbuffer[1][0] ), .B1(n570), .Y(n557) );
  CLKBUFX2TS U1077 ( .A(n795), .Y(n751) );
  CLKBUFX2TS U1078 ( .A(n751), .Y(n602) );
  AOI22X1TS U1079 ( .A0(\requesterAddressbuffer[7][0] ), .A1(n602), .B0(
        \requesterAddressbuffer[5][0] ), .B1(n572), .Y(n556) );
  NAND4XLTS U1080 ( .A(n559), .B(n558), .C(n557), .D(n556), .Y(n560) );
  AOI22X1TS U1081 ( .A0(requesterAddressOut[0]), .A1(n685), .B0(n596), .B1(
        n560), .Y(n561) );
  INVX2TS U1082 ( .A(readRequesterAddress[0]), .Y(n947) );
  INVX2TS U1083 ( .A(n947), .Y(n996) );
  INVX2TS U1084 ( .A(n802), .Y(n597) );
  NAND2X1TS U1085 ( .A(n996), .B(n597), .Y(n609) );
  CLKBUFX2TS U1086 ( .A(requesterAddressIn_NORTH[1]), .Y(n1005) );
  CLKBUFX2TS U1087 ( .A(requesterAddressIn_EAST[1]), .Y(n1033) );
  CLKBUFX2TS U1088 ( .A(n1033), .Y(n1004) );
  AOI22X1TS U1089 ( .A0(n1005), .A1(n564), .B0(n1004), .B1(n590), .Y(n580) );
  CLKBUFX2TS U1090 ( .A(requesterAddressIn_SOUTH[1]), .Y(n1034) );
  CLKBUFX2TS U1091 ( .A(n1034), .Y(n1006) );
  CLKBUFX2TS U1092 ( .A(n544), .Y(n806) );
  CLKBUFX2TS U1093 ( .A(requesterAddressIn_WEST[1]), .Y(n927) );
  CLKBUFX2TS U1094 ( .A(n927), .Y(n956) );
  AOI22X1TS U1095 ( .A0(n1006), .A1(n806), .B0(n956), .B1(n565), .Y(n579) );
  INVX2TS U1096 ( .A(n733), .Y(n782) );
  AOI22X1TS U1097 ( .A0(\requesterAddressbuffer[2][1] ), .A1(n567), .B0(
        \requesterAddressbuffer[0][1] ), .B1(n566), .Y(n576) );
  AOI22X1TS U1098 ( .A0(\requesterAddressbuffer[6][1] ), .A1(n569), .B0(
        \requesterAddressbuffer[4][1] ), .B1(n568), .Y(n575) );
  AOI22X1TS U1099 ( .A0(\requesterAddressbuffer[3][1] ), .A1(n571), .B0(
        \requesterAddressbuffer[1][1] ), .B1(n570), .Y(n574) );
  AOI22X1TS U1100 ( .A0(\requesterAddressbuffer[7][1] ), .A1(n602), .B0(
        \requesterAddressbuffer[5][1] ), .B1(n572), .Y(n573) );
  NAND4XLTS U1101 ( .A(n576), .B(n575), .C(n574), .D(n573), .Y(n577) );
  AOI22X1TS U1102 ( .A0(requesterAddressOut[1]), .A1(n782), .B0(n596), .B1(
        n577), .Y(n578) );
  INVX2TS U1103 ( .A(readRequesterAddress[1]), .Y(n953) );
  INVX2TS U1104 ( .A(n953), .Y(n1639) );
  NAND2X1TS U1105 ( .A(n1639), .B(n597), .Y(n624) );
  CLKBUFX2TS U1106 ( .A(requesterAddressIn_NORTH[2]), .Y(n1012) );
  CLKBUFX2TS U1107 ( .A(n690), .Y(n613) );
  CLKBUFX2TS U1108 ( .A(requesterAddressIn_EAST[2]), .Y(n1038) );
  CLKBUFX2TS U1109 ( .A(n1038), .Y(n1010) );
  AOI22X1TS U1110 ( .A0(n1012), .A1(n613), .B0(n1010), .B1(n590), .Y(n589) );
  CLKBUFX2TS U1111 ( .A(requesterAddressIn_SOUTH[2]), .Y(n1039) );
  CLKBUFX2TS U1112 ( .A(n1039), .Y(n1013) );
  CLKBUFX2TS U1113 ( .A(requesterAddressIn_WEST[2]), .Y(n932) );
  CLKBUFX2TS U1114 ( .A(n932), .Y(n963) );
  AOI22X1TS U1115 ( .A0(n1013), .A1(n658), .B0(n963), .B1(n628), .Y(n588) );
  INVX2TS U1116 ( .A(n581), .Y(n758) );
  CLKBUFX2TS U1117 ( .A(n629), .Y(n615) );
  AOI22X1TS U1118 ( .A0(\requesterAddressbuffer[2][2] ), .A1(n615), .B0(
        \requesterAddressbuffer[0][2] ), .B1(n692), .Y(n585) );
  CLKBUFX2TS U1119 ( .A(n631), .Y(n616) );
  AOI22X1TS U1120 ( .A0(\requesterAddressbuffer[6][2] ), .A1(n616), .B0(
        \requesterAddressbuffer[4][2] ), .B1(n693), .Y(n584) );
  CLKBUFX2TS U1121 ( .A(n633), .Y(n617) );
  AOI22X1TS U1122 ( .A0(\requesterAddressbuffer[3][2] ), .A1(n617), .B0(
        \requesterAddressbuffer[1][2] ), .B1(n694), .Y(n583) );
  CLKBUFX2TS U1123 ( .A(n635), .Y(n618) );
  AOI22X1TS U1124 ( .A0(\requesterAddressbuffer[7][2] ), .A1(n602), .B0(
        \requesterAddressbuffer[5][2] ), .B1(n618), .Y(n582) );
  NAND4XLTS U1125 ( .A(n585), .B(n584), .C(n583), .D(n582), .Y(n586) );
  AOI22X1TS U1126 ( .A0(requesterAddressOut[2]), .A1(n758), .B0(n596), .B1(
        n586), .Y(n587) );
  INVX2TS U1127 ( .A(readRequesterAddress[2]), .Y(n962) );
  INVX2TS U1128 ( .A(n962), .Y(n1646) );
  NAND2X1TS U1129 ( .A(n1646), .B(n597), .Y(n642) );
  CLKBUFX2TS U1130 ( .A(requesterAddressIn_NORTH[3]), .Y(n1021) );
  CLKBUFX2TS U1131 ( .A(requesterAddressIn_EAST[3]), .Y(n1046) );
  CLKBUFX2TS U1132 ( .A(n1046), .Y(n1019) );
  AOI22X1TS U1133 ( .A0(n1021), .A1(n613), .B0(n1019), .B1(n590), .Y(n600) );
  CLKBUFX2TS U1134 ( .A(requesterAddressIn_SOUTH[3]), .Y(n1048) );
  CLKBUFX2TS U1135 ( .A(n1048), .Y(n1022) );
  CLKBUFX2TS U1136 ( .A(requesterAddressIn_WEST[3]), .Y(n941) );
  CLKBUFX2TS U1137 ( .A(n941), .Y(n973) );
  AOI22X1TS U1138 ( .A0(n1022), .A1(n806), .B0(n973), .B1(n614), .Y(n599) );
  AOI22X1TS U1139 ( .A0(\requesterAddressbuffer[2][3] ), .A1(n615), .B0(
        \requesterAddressbuffer[0][3] ), .B1(n692), .Y(n594) );
  AOI22X1TS U1140 ( .A0(\requesterAddressbuffer[6][3] ), .A1(n616), .B0(
        \requesterAddressbuffer[4][3] ), .B1(n693), .Y(n593) );
  AOI22X1TS U1141 ( .A0(\requesterAddressbuffer[3][3] ), .A1(n617), .B0(
        \requesterAddressbuffer[1][3] ), .B1(n694), .Y(n592) );
  CLKBUFX2TS U1142 ( .A(n751), .Y(n647) );
  AOI22X1TS U1143 ( .A0(\requesterAddressbuffer[7][3] ), .A1(n647), .B0(
        \requesterAddressbuffer[5][3] ), .B1(n618), .Y(n591) );
  NAND4XLTS U1144 ( .A(n594), .B(n593), .C(n592), .D(n591), .Y(n595) );
  AOI22X1TS U1145 ( .A0(requesterAddressOut[3]), .A1(n523), .B0(n596), .B1(
        n595), .Y(n598) );
  INVX2TS U1146 ( .A(readRequesterAddress[3]), .Y(n970) );
  INVX2TS U1147 ( .A(n970), .Y(n1653) );
  NAND2X1TS U1148 ( .A(n1653), .B(n597), .Y(n653) );
  CLKBUFX2TS U1149 ( .A(destinationAddressIn_NORTH[0]), .Y(n1664) );
  CLKBUFX2TS U1150 ( .A(destinationAddressIn_EAST[0]), .Y(n1812) );
  CLKBUFX2TS U1151 ( .A(n1812), .Y(n1692) );
  CLKBUFX2TS U1152 ( .A(n601), .Y(n646) );
  AOI22X1TS U1153 ( .A0(n1664), .A1(n613), .B0(n1692), .B1(n646), .Y(n612) );
  CLKBUFX2TS U1154 ( .A(destinationAddressIn_WEST[0]), .Y(n1693) );
  CLKBUFX2TS U1155 ( .A(n1693), .Y(n1756) );
  AOI22X1TS U1156 ( .A0(destinationAddressIn_SOUTH[0]), .A1(n658), .B0(n1756), 
        .B1(n614), .Y(n611) );
  AOI22X1TS U1157 ( .A0(\destinationAddressbuffer[2][0] ), .A1(n615), .B0(
        \destinationAddressbuffer[0][0] ), .B1(n630), .Y(n606) );
  AOI22X1TS U1158 ( .A0(\destinationAddressbuffer[6][0] ), .A1(n616), .B0(
        \destinationAddressbuffer[4][0] ), .B1(n632), .Y(n605) );
  AOI22X1TS U1159 ( .A0(\destinationAddressbuffer[3][0] ), .A1(n617), .B0(
        \destinationAddressbuffer[1][0] ), .B1(n634), .Y(n604) );
  AOI22X1TS U1160 ( .A0(\destinationAddressbuffer[7][0] ), .A1(n602), .B0(
        \destinationAddressbuffer[5][0] ), .B1(n618), .Y(n603) );
  NAND4XLTS U1161 ( .A(n606), .B(n605), .C(n604), .D(n603), .Y(n607) );
  AOI22X1TS U1162 ( .A0(destinationAddressOut[0]), .A1(n685), .B0(n608), .B1(
        n607), .Y(n610) );
  CLKBUFX2TS U1163 ( .A(destinationAddressIn_NORTH[1]), .Y(n1671) );
  CLKBUFX2TS U1164 ( .A(destinationAddressIn_EAST[1]), .Y(n1822) );
  CLKBUFX2TS U1165 ( .A(n1822), .Y(n1701) );
  AOI22X1TS U1166 ( .A0(n1671), .A1(n613), .B0(n1701), .B1(n646), .Y(n627) );
  CLKBUFX2TS U1167 ( .A(destinationAddressIn_WEST[1]), .Y(n1703) );
  CLKBUFX2TS U1168 ( .A(n1703), .Y(n1764) );
  AOI22X1TS U1169 ( .A0(destinationAddressIn_SOUTH[1]), .A1(n806), .B0(n1764), 
        .B1(n614), .Y(n626) );
  AOI22X1TS U1170 ( .A0(\destinationAddressbuffer[2][1] ), .A1(n615), .B0(
        \destinationAddressbuffer[0][1] ), .B1(n630), .Y(n622) );
  AOI22X1TS U1171 ( .A0(\destinationAddressbuffer[6][1] ), .A1(n616), .B0(
        \destinationAddressbuffer[4][1] ), .B1(n632), .Y(n621) );
  AOI22X1TS U1172 ( .A0(\destinationAddressbuffer[3][1] ), .A1(n617), .B0(
        \destinationAddressbuffer[1][1] ), .B1(n634), .Y(n620) );
  AOI22X1TS U1173 ( .A0(\destinationAddressbuffer[7][1] ), .A1(n647), .B0(
        \destinationAddressbuffer[5][1] ), .B1(n618), .Y(n619) );
  NAND4XLTS U1174 ( .A(n622), .B(n621), .C(n620), .D(n619), .Y(n623) );
  AOI22X1TS U1175 ( .A0(destinationAddressOut[1]), .A1(n685), .B0(n641), .B1(
        n623), .Y(n625) );
  CLKBUFX2TS U1176 ( .A(destinationAddressIn_NORTH[2]), .Y(n1677) );
  CLKBUFX2TS U1177 ( .A(n690), .Y(n672) );
  CLKBUFX2TS U1178 ( .A(destinationAddressIn_EAST[2]), .Y(n1833) );
  CLKBUFX2TS U1179 ( .A(n1833), .Y(n1710) );
  AOI22X1TS U1180 ( .A0(n1677), .A1(n672), .B0(n1710), .B1(n646), .Y(n645) );
  CLKBUFX2TS U1181 ( .A(n544), .Y(n786) );
  CLKBUFX2TS U1182 ( .A(destinationAddressIn_WEST[2]), .Y(n1712) );
  CLKBUFX2TS U1183 ( .A(n1712), .Y(n1771) );
  CLKBUFX2TS U1184 ( .A(n628), .Y(n668) );
  AOI22X1TS U1185 ( .A0(destinationAddressIn_SOUTH[2]), .A1(n786), .B0(n1771), 
        .B1(n668), .Y(n644) );
  CLKBUFX2TS U1186 ( .A(n629), .Y(n674) );
  CLKBUFX2TS U1187 ( .A(n630), .Y(n673) );
  AOI22X1TS U1188 ( .A0(\destinationAddressbuffer[2][2] ), .A1(n674), .B0(
        \destinationAddressbuffer[0][2] ), .B1(n673), .Y(n639) );
  CLKBUFX2TS U1189 ( .A(n631), .Y(n676) );
  CLKBUFX2TS U1190 ( .A(n632), .Y(n675) );
  AOI22X1TS U1191 ( .A0(\destinationAddressbuffer[6][2] ), .A1(n676), .B0(
        \destinationAddressbuffer[4][2] ), .B1(n675), .Y(n638) );
  CLKBUFX2TS U1192 ( .A(n633), .Y(n678) );
  CLKBUFX2TS U1193 ( .A(n634), .Y(n677) );
  AOI22X1TS U1194 ( .A0(\destinationAddressbuffer[3][2] ), .A1(n678), .B0(
        \destinationAddressbuffer[1][2] ), .B1(n677), .Y(n637) );
  CLKBUFX2TS U1195 ( .A(n635), .Y(n679) );
  AOI22X1TS U1196 ( .A0(\destinationAddressbuffer[7][2] ), .A1(n647), .B0(
        \destinationAddressbuffer[5][2] ), .B1(n679), .Y(n636) );
  NAND4XLTS U1197 ( .A(n639), .B(n638), .C(n637), .D(n636), .Y(n640) );
  AOI22X1TS U1198 ( .A0(destinationAddressOut[2]), .A1(n523), .B0(n641), .B1(
        n640), .Y(n643) );
  CLKBUFX2TS U1199 ( .A(destinationAddressIn_NORTH[3]), .Y(n1685) );
  CLKBUFX2TS U1200 ( .A(destinationAddressIn_EAST[3]), .Y(n1844) );
  CLKBUFX2TS U1201 ( .A(n1844), .Y(n1718) );
  AOI22X1TS U1202 ( .A0(n1685), .A1(n672), .B0(n1718), .B1(n646), .Y(n656) );
  CLKBUFX2TS U1203 ( .A(destinationAddressIn_WEST[3]), .Y(n1719) );
  CLKBUFX2TS U1204 ( .A(n1719), .Y(n1779) );
  AOI22X1TS U1205 ( .A0(destinationAddressIn_SOUTH[3]), .A1(n786), .B0(n1779), 
        .B1(n668), .Y(n655) );
  AOI22X1TS U1206 ( .A0(\destinationAddressbuffer[2][3] ), .A1(n674), .B0(
        \destinationAddressbuffer[0][3] ), .B1(n673), .Y(n651) );
  AOI22X1TS U1207 ( .A0(\destinationAddressbuffer[6][3] ), .A1(n676), .B0(
        \destinationAddressbuffer[4][3] ), .B1(n675), .Y(n650) );
  AOI22X1TS U1208 ( .A0(\destinationAddressbuffer[3][3] ), .A1(n678), .B0(
        \destinationAddressbuffer[1][3] ), .B1(n677), .Y(n649) );
  AOI22X1TS U1209 ( .A0(\destinationAddressbuffer[7][3] ), .A1(n647), .B0(
        \destinationAddressbuffer[5][3] ), .B1(n679), .Y(n648) );
  NAND4XLTS U1210 ( .A(n651), .B(n650), .C(n649), .D(n648), .Y(n652) );
  AOI22X1TS U1211 ( .A0(destinationAddressOut[3]), .A1(n758), .B0(n1907), .B1(
        n652), .Y(n654) );
  AOI22X1TS U1212 ( .A0(destinationAddressIn_EAST[4]), .A1(n747), .B0(n657), 
        .B1(n668), .Y(n667) );
  AOI22X1TS U1213 ( .A0(destinationAddressIn_NORTH[4]), .A1(n672), .B0(n659), 
        .B1(n658), .Y(n666) );
  INVX2TS U1214 ( .A(n1908), .Y(n767) );
  CLKBUFX2TS U1215 ( .A(n767), .Y(n863) );
  AOI22X1TS U1216 ( .A0(\destinationAddressbuffer[2][4] ), .A1(n674), .B0(
        \destinationAddressbuffer[0][4] ), .B1(n673), .Y(n663) );
  AOI22X1TS U1217 ( .A0(\destinationAddressbuffer[6][4] ), .A1(n676), .B0(
        \destinationAddressbuffer[4][4] ), .B1(n675), .Y(n662) );
  AOI22X1TS U1218 ( .A0(\destinationAddressbuffer[3][4] ), .A1(n678), .B0(
        \destinationAddressbuffer[1][4] ), .B1(n677), .Y(n661) );
  CLKBUFX2TS U1219 ( .A(n751), .Y(n705) );
  AOI22X1TS U1220 ( .A0(\destinationAddressbuffer[7][4] ), .A1(n705), .B0(
        \destinationAddressbuffer[5][4] ), .B1(n679), .Y(n660) );
  NAND4XLTS U1221 ( .A(n663), .B(n662), .C(n661), .D(n660), .Y(n664) );
  AOI22X1TS U1222 ( .A0(destinationAddressOut[4]), .A1(n782), .B0(n863), .B1(
        n664), .Y(n665) );
  CLKBUFX2TS U1223 ( .A(n776), .Y(n763) );
  AOI22X1TS U1224 ( .A0(destinationAddressIn_EAST[5]), .A1(n763), .B0(n669), 
        .B1(n668), .Y(n688) );
  CLKBUFX2TS U1225 ( .A(n670), .Y(n748) );
  AOI22X1TS U1226 ( .A0(destinationAddressIn_NORTH[5]), .A1(n672), .B0(n671), 
        .B1(n748), .Y(n687) );
  AOI22X1TS U1227 ( .A0(\destinationAddressbuffer[2][5] ), .A1(n674), .B0(
        \destinationAddressbuffer[0][5] ), .B1(n673), .Y(n683) );
  AOI22X1TS U1228 ( .A0(\destinationAddressbuffer[6][5] ), .A1(n676), .B0(
        \destinationAddressbuffer[4][5] ), .B1(n675), .Y(n682) );
  AOI22X1TS U1229 ( .A0(\destinationAddressbuffer[3][5] ), .A1(n678), .B0(
        \destinationAddressbuffer[1][5] ), .B1(n677), .Y(n681) );
  AOI22X1TS U1230 ( .A0(\destinationAddressbuffer[7][5] ), .A1(n705), .B0(
        \destinationAddressbuffer[5][5] ), .B1(n679), .Y(n680) );
  NAND4XLTS U1231 ( .A(n683), .B(n682), .C(n681), .D(n680), .Y(n684) );
  AOI22X1TS U1232 ( .A0(destinationAddressOut[5]), .A1(n685), .B0(n863), .B1(
        n684), .Y(n686) );
  CLKBUFX2TS U1233 ( .A(n808), .Y(n728) );
  AOI22X1TS U1234 ( .A0(destinationAddressIn_EAST[6]), .A1(n763), .B0(n689), 
        .B1(n728), .Y(n702) );
  CLKBUFX2TS U1235 ( .A(n690), .Y(n807) );
  CLKBUFX2TS U1236 ( .A(n807), .Y(n731) );
  AOI22X1TS U1237 ( .A0(destinationAddressIn_NORTH[6]), .A1(n731), .B0(n691), 
        .B1(n748), .Y(n701) );
  CLKBUFX2TS U1238 ( .A(n692), .Y(n809) );
  CLKBUFX2TS U1239 ( .A(n809), .Y(n734) );
  AOI22X1TS U1240 ( .A0(\destinationAddressbuffer[2][6] ), .A1(n717), .B0(
        \destinationAddressbuffer[0][6] ), .B1(n734), .Y(n698) );
  CLKBUFX2TS U1241 ( .A(n693), .Y(n811) );
  CLKBUFX2TS U1242 ( .A(n811), .Y(n735) );
  AOI22X1TS U1243 ( .A0(\destinationAddressbuffer[6][6] ), .A1(n718), .B0(
        \destinationAddressbuffer[4][6] ), .B1(n735), .Y(n697) );
  CLKBUFX2TS U1244 ( .A(n694), .Y(n813) );
  CLKBUFX2TS U1245 ( .A(n813), .Y(n736) );
  AOI22X1TS U1246 ( .A0(\destinationAddressbuffer[3][6] ), .A1(n719), .B0(
        \destinationAddressbuffer[1][6] ), .B1(n736), .Y(n696) );
  CLKBUFX2TS U1247 ( .A(n857), .Y(n826) );
  CLKBUFX2TS U1248 ( .A(n826), .Y(n737) );
  AOI22X1TS U1249 ( .A0(\destinationAddressbuffer[7][6] ), .A1(n705), .B0(
        \destinationAddressbuffer[5][6] ), .B1(n737), .Y(n695) );
  NAND4XLTS U1250 ( .A(n698), .B(n697), .C(n696), .D(n695), .Y(n699) );
  AOI22X1TS U1251 ( .A0(destinationAddressOut[6]), .A1(n782), .B0(n863), .B1(
        n699), .Y(n700) );
  AOI22X1TS U1252 ( .A0(destinationAddressIn_EAST[7]), .A1(n825), .B0(n703), 
        .B1(n728), .Y(n713) );
  AOI22X1TS U1253 ( .A0(destinationAddressIn_NORTH[7]), .A1(n731), .B0(n704), 
        .B1(n764), .Y(n712) );
  CLKBUFX2TS U1254 ( .A(n767), .Y(n757) );
  AOI22X1TS U1255 ( .A0(\destinationAddressbuffer[2][7] ), .A1(n717), .B0(
        \destinationAddressbuffer[0][7] ), .B1(n734), .Y(n709) );
  AOI22X1TS U1256 ( .A0(\destinationAddressbuffer[6][7] ), .A1(n718), .B0(
        \destinationAddressbuffer[4][7] ), .B1(n735), .Y(n708) );
  AOI22X1TS U1257 ( .A0(\destinationAddressbuffer[3][7] ), .A1(n719), .B0(
        \destinationAddressbuffer[1][7] ), .B1(n736), .Y(n707) );
  AOI22X1TS U1258 ( .A0(\destinationAddressbuffer[7][7] ), .A1(n705), .B0(
        \destinationAddressbuffer[5][7] ), .B1(n737), .Y(n706) );
  NAND4XLTS U1259 ( .A(n709), .B(n708), .C(n707), .D(n706), .Y(n710) );
  AOI22X1TS U1260 ( .A0(destinationAddressOut[7]), .A1(n522), .B0(n757), .B1(
        n710), .Y(n711) );
  AOI22X1TS U1261 ( .A0(destinationAddressIn_EAST[8]), .A1(n747), .B0(n714), 
        .B1(n728), .Y(n727) );
  AOI22X1TS U1262 ( .A0(n716), .A1(n731), .B0(n715), .B1(n748), .Y(n726) );
  CLKBUFX2TS U1263 ( .A(n717), .Y(n810) );
  AOI22X1TS U1264 ( .A0(\destinationAddressbuffer[2][8] ), .A1(n810), .B0(
        \destinationAddressbuffer[0][8] ), .B1(n734), .Y(n723) );
  CLKBUFX2TS U1265 ( .A(n718), .Y(n812) );
  AOI22X1TS U1266 ( .A0(\destinationAddressbuffer[6][8] ), .A1(n812), .B0(
        \destinationAddressbuffer[4][8] ), .B1(n735), .Y(n722) );
  CLKBUFX2TS U1267 ( .A(n719), .Y(n814) );
  AOI22X1TS U1268 ( .A0(\destinationAddressbuffer[3][8] ), .A1(n814), .B0(
        \destinationAddressbuffer[1][8] ), .B1(n736), .Y(n721) );
  AOI22X1TS U1269 ( .A0(\destinationAddressbuffer[7][8] ), .A1(n815), .B0(
        \destinationAddressbuffer[5][8] ), .B1(n737), .Y(n720) );
  NAND4XLTS U1270 ( .A(n723), .B(n722), .C(n721), .D(n720), .Y(n724) );
  AOI22X1TS U1271 ( .A0(destinationAddressOut[8]), .A1(n758), .B0(n757), .B1(
        n724), .Y(n725) );
  AOI22X1TS U1272 ( .A0(destinationAddressIn_EAST[9]), .A1(n763), .B0(n729), 
        .B1(n728), .Y(n745) );
  AOI22X1TS U1273 ( .A0(n732), .A1(n731), .B0(n730), .B1(n764), .Y(n744) );
  INVX2TS U1274 ( .A(n733), .Y(n842) );
  AOI22X1TS U1275 ( .A0(\destinationAddressbuffer[2][9] ), .A1(n810), .B0(
        \destinationAddressbuffer[0][9] ), .B1(n734), .Y(n741) );
  AOI22X1TS U1276 ( .A0(\destinationAddressbuffer[6][9] ), .A1(n812), .B0(
        \destinationAddressbuffer[4][9] ), .B1(n735), .Y(n740) );
  AOI22X1TS U1277 ( .A0(\destinationAddressbuffer[3][9] ), .A1(n814), .B0(
        \destinationAddressbuffer[1][9] ), .B1(n736), .Y(n739) );
  AOI22X1TS U1278 ( .A0(\destinationAddressbuffer[7][9] ), .A1(n815), .B0(
        \destinationAddressbuffer[5][9] ), .B1(n737), .Y(n738) );
  NAND4XLTS U1279 ( .A(n741), .B(n740), .C(n739), .D(n738), .Y(n742) );
  AOI22X1TS U1280 ( .A0(destinationAddressOut[9]), .A1(n842), .B0(n757), .B1(
        n742), .Y(n743) );
  CLKBUFX2TS U1281 ( .A(n808), .Y(n787) );
  AOI22X1TS U1282 ( .A0(destinationAddressIn_EAST[10]), .A1(n747), .B0(n746), 
        .B1(n787), .Y(n761) );
  CLKBUFX2TS U1283 ( .A(n807), .Y(n788) );
  AOI22X1TS U1284 ( .A0(n750), .A1(n788), .B0(n749), .B1(n748), .Y(n760) );
  CLKBUFX2TS U1285 ( .A(n810), .Y(n789) );
  CLKBUFX2TS U1286 ( .A(n809), .Y(n790) );
  AOI22X1TS U1287 ( .A0(\destinationAddressbuffer[2][10] ), .A1(n789), .B0(
        \destinationAddressbuffer[0][10] ), .B1(n790), .Y(n755) );
  CLKBUFX2TS U1288 ( .A(n812), .Y(n791) );
  CLKBUFX2TS U1289 ( .A(n811), .Y(n792) );
  AOI22X1TS U1290 ( .A0(\destinationAddressbuffer[6][10] ), .A1(n791), .B0(
        \destinationAddressbuffer[4][10] ), .B1(n792), .Y(n754) );
  CLKBUFX2TS U1291 ( .A(n814), .Y(n793) );
  CLKBUFX2TS U1292 ( .A(n813), .Y(n794) );
  AOI22X1TS U1293 ( .A0(\destinationAddressbuffer[3][10] ), .A1(n793), .B0(
        \destinationAddressbuffer[1][10] ), .B1(n794), .Y(n753) );
  CLKBUFX2TS U1294 ( .A(n826), .Y(n796) );
  AOI22X1TS U1295 ( .A0(\destinationAddressbuffer[7][10] ), .A1(n751), .B0(
        \destinationAddressbuffer[5][10] ), .B1(n796), .Y(n752) );
  NAND4XLTS U1296 ( .A(n755), .B(n754), .C(n753), .D(n752), .Y(n756) );
  AOI22X1TS U1297 ( .A0(destinationAddressOut[10]), .A1(n758), .B0(n757), .B1(
        n756), .Y(n759) );
  AOI22X1TS U1298 ( .A0(destinationAddressIn_EAST[11]), .A1(n763), .B0(n762), 
        .B1(n787), .Y(n775) );
  AOI22X1TS U1299 ( .A0(n766), .A1(n788), .B0(n765), .B1(n764), .Y(n774) );
  CLKBUFX2TS U1300 ( .A(n767), .Y(n821) );
  AOI22X1TS U1301 ( .A0(\destinationAddressbuffer[2][11] ), .A1(n789), .B0(
        \destinationAddressbuffer[0][11] ), .B1(n790), .Y(n771) );
  AOI22X1TS U1302 ( .A0(\destinationAddressbuffer[6][11] ), .A1(n791), .B0(
        \destinationAddressbuffer[4][11] ), .B1(n792), .Y(n770) );
  AOI22X1TS U1303 ( .A0(\destinationAddressbuffer[3][11] ), .A1(n793), .B0(
        \destinationAddressbuffer[1][11] ), .B1(n794), .Y(n769) );
  AOI22X1TS U1304 ( .A0(\destinationAddressbuffer[7][11] ), .A1(n795), .B0(
        \destinationAddressbuffer[5][11] ), .B1(n796), .Y(n768) );
  NAND4XLTS U1305 ( .A(n771), .B(n770), .C(n769), .D(n768), .Y(n772) );
  AOI22X1TS U1306 ( .A0(destinationAddressOut[11]), .A1(n522), .B0(n821), .B1(
        n772), .Y(n773) );
  CLKBUFX2TS U1307 ( .A(dataIn_EAST[0]), .Y(n1459) );
  CLKBUFX2TS U1308 ( .A(n1459), .Y(n1108) );
  CLKBUFX2TS U1309 ( .A(n776), .Y(n846) );
  AOI22X1TS U1310 ( .A0(dataIn_SOUTH[0]), .A1(n786), .B0(n1108), .B1(n846), 
        .Y(n785) );
  CLKBUFX2TS U1311 ( .A(dataIn_WEST[0]), .Y(n1499) );
  CLKBUFX2TS U1312 ( .A(n1499), .Y(n1391) );
  AOI22X1TS U1313 ( .A0(dataIn_NORTH[0]), .A1(n788), .B0(n1391), .B1(n787), 
        .Y(n784) );
  AOI22X1TS U1314 ( .A0(\dataoutbuffer[0][0] ), .A1(n790), .B0(
        \dataoutbuffer[2][0] ), .B1(n789), .Y(n780) );
  AOI22X1TS U1315 ( .A0(\dataoutbuffer[4][0] ), .A1(n792), .B0(
        \dataoutbuffer[6][0] ), .B1(n791), .Y(n779) );
  AOI22X1TS U1316 ( .A0(\dataoutbuffer[1][0] ), .A1(n794), .B0(
        \dataoutbuffer[3][0] ), .B1(n793), .Y(n778) );
  AOI22X1TS U1317 ( .A0(\dataoutbuffer[5][0] ), .A1(n796), .B0(
        \dataoutbuffer[7][0] ), .B1(n856), .Y(n777) );
  NAND4XLTS U1318 ( .A(n780), .B(n779), .C(n778), .D(n777), .Y(n781) );
  AOI22X1TS U1319 ( .A0(dataOut[0]), .A1(n782), .B0(n821), .B1(n781), .Y(n783)
         );
  CLKBUFX2TS U1320 ( .A(dataIn_EAST[1]), .Y(n1467) );
  CLKBUFX2TS U1321 ( .A(n1467), .Y(n1339) );
  AOI22X1TS U1322 ( .A0(dataIn_SOUTH[1]), .A1(n786), .B0(n1339), .B1(n825), 
        .Y(n805) );
  CLKBUFX2TS U1323 ( .A(dataIn_WEST[1]), .Y(n1506) );
  CLKBUFX2TS U1324 ( .A(n1506), .Y(n1397) );
  AOI22X1TS U1325 ( .A0(dataIn_NORTH[1]), .A1(n788), .B0(n1397), .B1(n787), 
        .Y(n804) );
  AOI22X1TS U1326 ( .A0(\dataoutbuffer[0][1] ), .A1(n790), .B0(
        \dataoutbuffer[2][1] ), .B1(n789), .Y(n800) );
  AOI22X1TS U1327 ( .A0(\dataoutbuffer[4][1] ), .A1(n792), .B0(
        \dataoutbuffer[6][1] ), .B1(n791), .Y(n799) );
  AOI22X1TS U1328 ( .A0(\dataoutbuffer[1][1] ), .A1(n794), .B0(
        \dataoutbuffer[3][1] ), .B1(n793), .Y(n798) );
  AOI22X1TS U1329 ( .A0(\dataoutbuffer[5][1] ), .A1(n796), .B0(
        \dataoutbuffer[7][1] ), .B1(n795), .Y(n797) );
  NAND4XLTS U1330 ( .A(n800), .B(n799), .C(n798), .D(n797), .Y(n801) );
  AOI22X1TS U1331 ( .A0(dataOut[1]), .A1(n523), .B0(n821), .B1(n801), .Y(n803)
         );
  CLKBUFX2TS U1332 ( .A(dataIn_EAST[2]), .Y(n1473) );
  CLKBUFX2TS U1333 ( .A(n1473), .Y(n1345) );
  AOI22X1TS U1334 ( .A0(dataIn_SOUTH[2]), .A1(n806), .B0(n1345), .B1(n846), 
        .Y(n824) );
  CLKBUFX2TS U1335 ( .A(n807), .Y(n849) );
  CLKBUFX2TS U1336 ( .A(dataIn_WEST[2]), .Y(n1513) );
  CLKBUFX2TS U1337 ( .A(n1513), .Y(n1402) );
  CLKBUFX2TS U1338 ( .A(n808), .Y(n848) );
  AOI22X1TS U1339 ( .A0(dataIn_NORTH[2]), .A1(n849), .B0(n1402), .B1(n848), 
        .Y(n823) );
  CLKBUFX2TS U1340 ( .A(n809), .Y(n851) );
  CLKBUFX2TS U1341 ( .A(n810), .Y(n850) );
  AOI22X1TS U1342 ( .A0(\dataoutbuffer[0][2] ), .A1(n851), .B0(
        \dataoutbuffer[2][2] ), .B1(n850), .Y(n819) );
  CLKBUFX2TS U1343 ( .A(n811), .Y(n853) );
  CLKBUFX2TS U1344 ( .A(n812), .Y(n852) );
  AOI22X1TS U1345 ( .A0(\dataoutbuffer[4][2] ), .A1(n853), .B0(
        \dataoutbuffer[6][2] ), .B1(n852), .Y(n818) );
  CLKBUFX2TS U1346 ( .A(n813), .Y(n855) );
  CLKBUFX2TS U1347 ( .A(n814), .Y(n854) );
  AOI22X1TS U1348 ( .A0(\dataoutbuffer[1][2] ), .A1(n855), .B0(
        \dataoutbuffer[3][2] ), .B1(n854), .Y(n817) );
  AOI22X1TS U1349 ( .A0(\dataoutbuffer[5][2] ), .A1(n826), .B0(
        \dataoutbuffer[7][2] ), .B1(n815), .Y(n816) );
  NAND4XLTS U1350 ( .A(n819), .B(n818), .C(n817), .D(n816), .Y(n820) );
  AOI22X1TS U1351 ( .A0(dataOut[2]), .A1(n842), .B0(n821), .B1(n820), .Y(n822)
         );
  INVX2TS U1352 ( .A(n12), .Y(n864) );
  CLKBUFX2TS U1353 ( .A(dataIn_EAST[3]), .Y(n1479) );
  CLKBUFX2TS U1354 ( .A(n1479), .Y(n1350) );
  AOI22X1TS U1355 ( .A0(dataIn_SOUTH[3]), .A1(n847), .B0(n1350), .B1(n825), 
        .Y(n834) );
  CLKBUFX2TS U1356 ( .A(dataIn_WEST[3]), .Y(n1522) );
  CLKBUFX2TS U1357 ( .A(n1522), .Y(n1407) );
  AOI22X1TS U1358 ( .A0(dataIn_NORTH[3]), .A1(n849), .B0(n1407), .B1(n848), 
        .Y(n833) );
  AOI22X1TS U1359 ( .A0(\dataoutbuffer[0][3] ), .A1(n851), .B0(
        \dataoutbuffer[2][3] ), .B1(n850), .Y(n830) );
  AOI22X1TS U1360 ( .A0(\dataoutbuffer[4][3] ), .A1(n853), .B0(
        \dataoutbuffer[6][3] ), .B1(n852), .Y(n829) );
  AOI22X1TS U1361 ( .A0(\dataoutbuffer[1][3] ), .A1(n855), .B0(
        \dataoutbuffer[3][3] ), .B1(n854), .Y(n828) );
  AOI22X1TS U1362 ( .A0(\dataoutbuffer[5][3] ), .A1(n826), .B0(
        \dataoutbuffer[7][3] ), .B1(n835), .Y(n827) );
  NAND4XLTS U1363 ( .A(n830), .B(n829), .C(n828), .D(n827), .Y(n831) );
  AOI22X1TS U1364 ( .A0(dataOut[3]), .A1(n842), .B0(n841), .B1(n831), .Y(n832)
         );
  CLKBUFX2TS U1365 ( .A(dataIn_EAST[4]), .Y(n1484) );
  CLKBUFX2TS U1366 ( .A(n1484), .Y(n1355) );
  AOI22X1TS U1367 ( .A0(dataIn_SOUTH[4]), .A1(n847), .B0(n1355), .B1(n846), 
        .Y(n845) );
  CLKBUFX2TS U1368 ( .A(dataIn_WEST[4]), .Y(n1529) );
  CLKBUFX2TS U1369 ( .A(n1529), .Y(n1411) );
  AOI22X1TS U1370 ( .A0(dataIn_NORTH[4]), .A1(n849), .B0(n1411), .B1(n848), 
        .Y(n844) );
  AOI22X1TS U1371 ( .A0(\dataoutbuffer[0][4] ), .A1(n851), .B0(
        \dataoutbuffer[2][4] ), .B1(n850), .Y(n839) );
  AOI22X1TS U1372 ( .A0(\dataoutbuffer[4][4] ), .A1(n853), .B0(
        \dataoutbuffer[6][4] ), .B1(n852), .Y(n838) );
  AOI22X1TS U1373 ( .A0(\dataoutbuffer[1][4] ), .A1(n855), .B0(
        \dataoutbuffer[3][4] ), .B1(n854), .Y(n837) );
  AOI22X1TS U1374 ( .A0(\dataoutbuffer[5][4] ), .A1(n857), .B0(
        \dataoutbuffer[7][4] ), .B1(n835), .Y(n836) );
  NAND4XLTS U1375 ( .A(n839), .B(n838), .C(n837), .D(n836), .Y(n840) );
  AOI22X1TS U1376 ( .A0(dataOut[4]), .A1(n842), .B0(n841), .B1(n840), .Y(n843)
         );
  CLKBUFX2TS U1377 ( .A(dataIn_EAST[5]), .Y(n1493) );
  CLKBUFX2TS U1378 ( .A(n1493), .Y(n1361) );
  AOI22X1TS U1379 ( .A0(dataIn_SOUTH[5]), .A1(n847), .B0(n1361), .B1(n846), 
        .Y(n867) );
  CLKBUFX2TS U1380 ( .A(dataIn_WEST[5]), .Y(n1537) );
  CLKBUFX2TS U1381 ( .A(n1537), .Y(n1419) );
  AOI22X1TS U1382 ( .A0(dataIn_NORTH[5]), .A1(n849), .B0(n1419), .B1(n848), 
        .Y(n866) );
  AOI22X1TS U1383 ( .A0(\dataoutbuffer[0][5] ), .A1(n851), .B0(
        \dataoutbuffer[2][5] ), .B1(n850), .Y(n861) );
  AOI22X1TS U1384 ( .A0(\dataoutbuffer[4][5] ), .A1(n853), .B0(
        \dataoutbuffer[6][5] ), .B1(n852), .Y(n860) );
  AOI22X1TS U1385 ( .A0(\dataoutbuffer[1][5] ), .A1(n855), .B0(
        \dataoutbuffer[3][5] ), .B1(n854), .Y(n859) );
  AOI22X1TS U1386 ( .A0(\dataoutbuffer[5][5] ), .A1(n857), .B0(
        \dataoutbuffer[7][5] ), .B1(n856), .Y(n858) );
  NAND4XLTS U1387 ( .A(n861), .B(n860), .C(n859), .D(n858), .Y(n862) );
  AOI22X1TS U1388 ( .A0(dataOut[5]), .A1(n523), .B0(n863), .B1(n862), .Y(n865)
         );
  INVX2TS U1389 ( .A(n947), .Y(n1755) );
  AOI22X1TS U1390 ( .A0(n1755), .A1(n1634), .B0(n1652), .B1(
        \requesterAddressbuffer[7][0] ), .Y(n870) );
  INVX2TS U1391 ( .A(n1512), .Y(n1641) );
  AOI22X1TS U1392 ( .A0(n52), .A1(n948), .B0(n1641), .B1(n1026), .Y(n869) );
  CLKBUFX2TS U1393 ( .A(n1028), .Y(n923) );
  CLKBUFX2TS U1394 ( .A(n998), .Y(n949) );
  AOI22X1TS U1395 ( .A0(n1517), .A1(n923), .B0(n871), .B1(n949), .Y(n868) );
  INVX2TS U1396 ( .A(n880), .Y(n1640) );
  INVX2TS U1397 ( .A(n1498), .Y(n1536) );
  AOI22X1TS U1398 ( .A0(n1640), .A1(n1639), .B0(n1536), .B1(
        \requesterAddressbuffer[7][1] ), .Y(n874) );
  AOI22X1TS U1399 ( .A0(n1656), .A1(n956), .B0(n875), .B1(n1033), .Y(n873) );
  CLKBUFX2TS U1400 ( .A(n1034), .Y(n928) );
  CLKBUFX2TS U1401 ( .A(n1005), .Y(n958) );
  AOI22X1TS U1402 ( .A0(n43), .A1(n928), .B0(n871), .B1(n958), .Y(n872) );
  AOI22X1TS U1403 ( .A0(n32), .A1(n1646), .B0(n1536), .B1(
        \requesterAddressbuffer[7][2] ), .Y(n879) );
  AOI22X1TS U1404 ( .A0(n1523), .A1(n963), .B0(n875), .B1(n1038), .Y(n878) );
  CLKBUFX2TS U1405 ( .A(n1039), .Y(n933) );
  INVX2TS U1406 ( .A(n876), .Y(n1515) );
  CLKBUFX2TS U1407 ( .A(n1012), .Y(n966) );
  AOI22X1TS U1408 ( .A0(n1517), .A1(n933), .B0(n1515), .B1(n966), .Y(n877) );
  INVX2TS U1409 ( .A(n880), .Y(n1654) );
  INVX2TS U1410 ( .A(n881), .Y(n1645) );
  AOI22X1TS U1411 ( .A0(n1654), .A1(n1653), .B0(n1645), .B1(
        \requesterAddressbuffer[7][3] ), .Y(n885) );
  INVX2TS U1412 ( .A(n1512), .Y(n1655) );
  AOI22X1TS U1413 ( .A0(n1647), .A1(n973), .B0(n1655), .B1(n1046), .Y(n884) );
  INVX2TS U1414 ( .A(n882), .Y(n1635) );
  CLKBUFX2TS U1415 ( .A(n1048), .Y(n943) );
  CLKBUFX2TS U1416 ( .A(n1021), .Y(n974) );
  AOI22X1TS U1417 ( .A0(n1635), .A1(n943), .B0(n1531), .B1(n974), .Y(n883) );
  INVX2TS U1418 ( .A(n947), .Y(n1811) );
  AOI22X1TS U1419 ( .A0(n1811), .A1(n1662), .B0(n1682), .B1(
        \requesterAddressbuffer[6][0] ), .Y(n888) );
  INVX2TS U1420 ( .A(n1472), .Y(n1670) );
  AOI22X1TS U1421 ( .A0(n921), .A1(n1684), .B0(requesterAddressIn_EAST[0]), 
        .B1(n1670), .Y(n887) );
  AOI22X1TS U1422 ( .A0(n923), .A1(n1462), .B0(n949), .B1(n1463), .Y(n886) );
  INVX2TS U1423 ( .A(n953), .Y(n1733) );
  INVX2TS U1424 ( .A(n896), .Y(n1669) );
  INVX2TS U1425 ( .A(n1458), .Y(n1492) );
  AOI22X1TS U1426 ( .A0(n1733), .A1(n1669), .B0(n1492), .B1(
        \requesterAddressbuffer[6][1] ), .Y(n892) );
  INVX2TS U1427 ( .A(n1472), .Y(n1676) );
  AOI22X1TS U1428 ( .A0(n927), .A1(n1485), .B0(requesterAddressIn_EAST[1]), 
        .B1(n1676), .Y(n891) );
  INVX2TS U1429 ( .A(n96), .Y(n1487) );
  INVX2TS U1430 ( .A(n889), .Y(n1488) );
  AOI22X1TS U1431 ( .A0(n928), .A1(n1487), .B0(n958), .B1(n1488), .Y(n890) );
  INVX2TS U1432 ( .A(n962), .Y(n1739) );
  AOI22X1TS U1433 ( .A0(n1739), .A1(n1662), .B0(n1492), .B1(
        \requesterAddressbuffer[6][2] ), .Y(n895) );
  AOI22X1TS U1434 ( .A0(n932), .A1(n1460), .B0(requesterAddressIn_EAST[2]), 
        .B1(n899), .Y(n894) );
  AOI22X1TS U1435 ( .A0(n933), .A1(n111), .B0(n966), .B1(n1488), .Y(n893) );
  INVX2TS U1436 ( .A(n970), .Y(n1747) );
  INVX2TS U1437 ( .A(n896), .Y(n1683) );
  INVX2TS U1438 ( .A(n897), .Y(n1675) );
  AOI22X1TS U1439 ( .A0(n1747), .A1(n1683), .B0(n1675), .B1(
        \requesterAddressbuffer[6][3] ), .Y(n903) );
  INVX2TS U1440 ( .A(n898), .Y(n1485) );
  AOI22X1TS U1441 ( .A0(n941), .A1(n1485), .B0(requesterAddressIn_EAST[3]), 
        .B1(n899), .Y(n902) );
  INVX2TS U1442 ( .A(n900), .Y(n1678) );
  AOI22X1TS U1443 ( .A0(n943), .A1(n1678), .B0(n974), .B1(n1665), .Y(n901) );
  AOI22X1TS U1444 ( .A0(n996), .A1(n1691), .B0(n1716), .B1(
        \requesterAddressbuffer[5][0] ), .Y(n907) );
  INVX2TS U1445 ( .A(n1435), .Y(n1702) );
  AOI22X1TS U1446 ( .A0(n921), .A1(n1720), .B0(requesterAddressIn_EAST[0]), 
        .B1(n1702), .Y(n906) );
  INVX2TS U1447 ( .A(n904), .Y(n1721) );
  AOI22X1TS U1448 ( .A0(n923), .A1(n1721), .B0(requesterAddressIn_NORTH[0]), 
        .B1(n1437), .Y(n905) );
  INVX2TS U1449 ( .A(n10), .Y(n1700) );
  INVX2TS U1450 ( .A(n1423), .Y(n1453) );
  AOI22X1TS U1451 ( .A0(n1639), .A1(n1700), .B0(n1453), .B1(
        \requesterAddressbuffer[5][1] ), .Y(n910) );
  INVX2TS U1452 ( .A(n1435), .Y(n1711) );
  AOI22X1TS U1453 ( .A0(n927), .A1(n1446), .B0(requesterAddressIn_EAST[1]), 
        .B1(n1711), .Y(n909) );
  AOI22X1TS U1454 ( .A0(n928), .A1(n1695), .B0(requesterAddressIn_NORTH[1]), 
        .B1(n1696), .Y(n908) );
  INVX2TS U1455 ( .A(n10), .Y(n1709) );
  AOI22X1TS U1456 ( .A0(n1646), .A1(n1709), .B0(n1453), .B1(
        \requesterAddressbuffer[5][2] ), .Y(n914) );
  AOI22X1TS U1457 ( .A0(n932), .A1(n1424), .B0(requesterAddressIn_EAST[2]), 
        .B1(n917), .Y(n913) );
  AOI22X1TS U1458 ( .A0(n933), .A1(n1425), .B0(requesterAddressIn_NORTH[2]), 
        .B1(n911), .Y(n912) );
  INVX2TS U1459 ( .A(n10), .Y(n1717) );
  INVX2TS U1460 ( .A(n915), .Y(n1708) );
  AOI22X1TS U1461 ( .A0(n1653), .A1(n1717), .B0(n1708), .B1(
        \requesterAddressbuffer[5][3] ), .Y(n920) );
  INVX2TS U1462 ( .A(n916), .Y(n1446) );
  AOI22X1TS U1463 ( .A0(n941), .A1(n1446), .B0(requesterAddressIn_EAST[3]), 
        .B1(n917), .Y(n919) );
  AOI22X1TS U1464 ( .A0(n943), .A1(n231), .B0(requesterAddressIn_NORTH[3]), 
        .B1(n1449), .Y(n918) );
  AOI22X1TS U1465 ( .A0(n996), .A1(n1725), .B0(n1745), .B1(
        \requesterAddressbuffer[4][0] ), .Y(n926) );
  INVX2TS U1466 ( .A(n1401), .Y(n1734) );
  AOI22X1TS U1467 ( .A0(n921), .A1(n1748), .B0(requesterAddressIn_EAST[0]), 
        .B1(n1734), .Y(n925) );
  AOI22X1TS U1468 ( .A0(n923), .A1(n1741), .B0(requesterAddressIn_NORTH[0]), 
        .B1(n922), .Y(n924) );
  INVX2TS U1469 ( .A(n953), .Y(n1863) );
  INVX2TS U1470 ( .A(n937), .Y(n1732) );
  INVX2TS U1471 ( .A(n1390), .Y(n1418) );
  AOI22X1TS U1472 ( .A0(n1863), .A1(n1732), .B0(n1418), .B1(
        \requesterAddressbuffer[4][1] ), .Y(n931) );
  INVX2TS U1473 ( .A(n1401), .Y(n1740) );
  AOI22X1TS U1474 ( .A0(n927), .A1(n1412), .B0(requesterAddressIn_EAST[1]), 
        .B1(n1740), .Y(n930) );
  AOI22X1TS U1475 ( .A0(n928), .A1(n1414), .B0(requesterAddressIn_NORTH[1]), 
        .B1(n1749), .Y(n929) );
  INVX2TS U1476 ( .A(n962), .Y(n1872) );
  AOI22X1TS U1477 ( .A0(n1872), .A1(n1725), .B0(n1418), .B1(
        \requesterAddressbuffer[4][2] ), .Y(n936) );
  AOI22X1TS U1478 ( .A0(n932), .A1(n1392), .B0(requesterAddressIn_EAST[2]), 
        .B1(n940), .Y(n935) );
  AOI22X1TS U1479 ( .A0(n933), .A1(n1750), .B0(requesterAddressIn_NORTH[2]), 
        .B1(n1749), .Y(n934) );
  INVX2TS U1480 ( .A(n970), .Y(n1882) );
  INVX2TS U1481 ( .A(n937), .Y(n1746) );
  INVX2TS U1482 ( .A(n938), .Y(n1738) );
  AOI22X1TS U1483 ( .A0(n1882), .A1(n1746), .B0(n1738), .B1(
        \requesterAddressbuffer[4][3] ), .Y(n946) );
  INVX2TS U1484 ( .A(n939), .Y(n1412) );
  AOI22X1TS U1485 ( .A0(n941), .A1(n1412), .B0(requesterAddressIn_EAST[3]), 
        .B1(n940), .Y(n945) );
  INVX2TS U1486 ( .A(n942), .Y(n1728) );
  AOI22X1TS U1487 ( .A0(n943), .A1(n1728), .B0(requesterAddressIn_NORTH[3]), 
        .B1(n1393), .Y(n944) );
  INVX2TS U1488 ( .A(n947), .Y(n1853) );
  AOI22X1TS U1489 ( .A0(n1853), .A1(n1754), .B0(n1776), .B1(
        \requesterAddressbuffer[3][0] ), .Y(n952) );
  AOI22X1TS U1490 ( .A0(n948), .A1(n141), .B0(n997), .B1(n128), .Y(n951) );
  INVX2TS U1491 ( .A(n964), .Y(n1772) );
  AOI22X1TS U1492 ( .A0(n999), .A1(n1772), .B0(n949), .B1(n1367), .Y(n950) );
  INVX2TS U1493 ( .A(n953), .Y(n1821) );
  INVX2TS U1494 ( .A(n971), .Y(n1762) );
  INVX2TS U1495 ( .A(n1366), .Y(n1385) );
  AOI22X1TS U1496 ( .A0(n1821), .A1(n1762), .B0(n1385), .B1(
        \requesterAddressbuffer[3][1] ), .Y(n961) );
  INVX2TS U1497 ( .A(n954), .Y(n1763) );
  AOI22X1TS U1498 ( .A0(n956), .A1(n955), .B0(n1004), .B1(n1763), .Y(n960) );
  INVX2TS U1499 ( .A(n964), .Y(n1781) );
  AOI22X1TS U1500 ( .A0(n1006), .A1(n1781), .B0(n958), .B1(n957), .Y(n959) );
  INVX2TS U1501 ( .A(n962), .Y(n1832) );
  AOI22X1TS U1502 ( .A0(n1832), .A1(n1754), .B0(n1385), .B1(
        \requesterAddressbuffer[3][2] ), .Y(n969) );
  AOI22X1TS U1503 ( .A0(n963), .A1(n1386), .B0(n1010), .B1(n1381), .Y(n968) );
  AOI22X1TS U1504 ( .A0(n1013), .A1(n125), .B0(n966), .B1(n965), .Y(n967) );
  INVX2TS U1505 ( .A(n970), .Y(n1843) );
  INVX2TS U1506 ( .A(n971), .Y(n1777) );
  INVX2TS U1507 ( .A(n1366), .Y(n1769) );
  AOI22X1TS U1508 ( .A0(n1843), .A1(n1777), .B0(n1769), .B1(
        \requesterAddressbuffer[3][3] ), .Y(n977) );
  AOI22X1TS U1509 ( .A0(n973), .A1(n141), .B0(n1019), .B1(n1778), .Y(n976) );
  AOI22X1TS U1510 ( .A0(n1022), .A1(n1772), .B0(n974), .B1(n1758), .Y(n975) );
  AOI22X1TS U1511 ( .A0(n1755), .A1(n1786), .B0(n1805), .B1(
        \requesterAddressbuffer[2][0] ), .Y(n980) );
  INVX2TS U1512 ( .A(n1344), .Y(n1793) );
  AOI22X1TS U1513 ( .A0(requesterAddressIn_WEST[0]), .A1(n1806), .B0(n997), 
        .B1(n1793), .Y(n979) );
  AOI22X1TS U1514 ( .A0(n999), .A1(n181), .B0(n998), .B1(n1111), .Y(n978) );
  INVX2TS U1515 ( .A(n989), .Y(n1792) );
  INVX2TS U1516 ( .A(n981), .Y(n1360) );
  AOI22X1TS U1517 ( .A0(n1863), .A1(n1792), .B0(n1360), .B1(
        \requesterAddressbuffer[2][1] ), .Y(n984) );
  INVX2TS U1518 ( .A(n1344), .Y(n1800) );
  AOI22X1TS U1519 ( .A0(requesterAddressIn_WEST[1]), .A1(n1356), .B0(n1004), 
        .B1(n1800), .Y(n983) );
  AOI22X1TS U1520 ( .A0(n1006), .A1(n1351), .B0(n1005), .B1(n1794), .Y(n982)
         );
  INVX2TS U1521 ( .A(n989), .Y(n1799) );
  AOI22X1TS U1522 ( .A0(n1872), .A1(n1799), .B0(n1360), .B1(
        \requesterAddressbuffer[2][2] ), .Y(n988) );
  AOI22X1TS U1523 ( .A0(requesterAddressIn_WEST[2]), .A1(n1109), .B0(n1010), 
        .B1(n991), .Y(n987) );
  AOI22X1TS U1524 ( .A0(n1013), .A1(n1110), .B0(n1012), .B1(n985), .Y(n986) );
  INVX2TS U1525 ( .A(n1606), .Y(n1798) );
  AOI22X1TS U1526 ( .A0(n1882), .A1(n1786), .B0(n1798), .B1(
        \requesterAddressbuffer[2][3] ), .Y(n995) );
  INVX2TS U1527 ( .A(n990), .Y(n1356) );
  AOI22X1TS U1528 ( .A0(requesterAddressIn_WEST[3]), .A1(n1356), .B0(n1019), 
        .B1(n991), .Y(n994) );
  INVX2TS U1529 ( .A(n992), .Y(n1801) );
  AOI22X1TS U1530 ( .A0(n1022), .A1(n1801), .B0(n1021), .B1(n1788), .Y(n993)
         );
  INVX2TS U1531 ( .A(n1084), .Y(n1098) );
  AOI22X1TS U1532 ( .A0(n996), .A1(n1098), .B0(n1841), .B1(
        \requesterAddressbuffer[1][0] ), .Y(n1002) );
  INVX2TS U1533 ( .A(n1089), .Y(n1823) );
  AOI22X1TS U1534 ( .A0(requesterAddressIn_WEST[0]), .A1(n1845), .B0(n997), 
        .B1(n1823), .Y(n1001) );
  AOI22X1TS U1535 ( .A0(n999), .A1(n1079), .B0(n998), .B1(n1080), .Y(n1000) );
  INVX2TS U1536 ( .A(n1084), .Y(n1831) );
  INVX2TS U1537 ( .A(n1003), .Y(n1103) );
  AOI22X1TS U1538 ( .A0(n1733), .A1(n1831), .B0(n1103), .B1(
        \requesterAddressbuffer[1][1] ), .Y(n1009) );
  INVX2TS U1539 ( .A(n1089), .Y(n1834) );
  AOI22X1TS U1540 ( .A0(requesterAddressIn_WEST[1]), .A1(n1099), .B0(n1004), 
        .B1(n1834), .Y(n1008) );
  AOI22X1TS U1541 ( .A0(n1006), .A1(n330), .B0(n1005), .B1(n1826), .Y(n1007)
         );
  AOI22X1TS U1542 ( .A0(n1739), .A1(n1842), .B0(n1103), .B1(
        \requesterAddressbuffer[1][2] ), .Y(n1016) );
  AOI22X1TS U1543 ( .A0(requesterAddressIn_WEST[2]), .A1(n1078), .B0(n1010), 
        .B1(n1018), .Y(n1015) );
  AOI22X1TS U1544 ( .A0(n1013), .A1(n1094), .B0(n1012), .B1(n1011), .Y(n1014)
         );
  INVX2TS U1545 ( .A(n1620), .Y(n1830) );
  AOI22X1TS U1546 ( .A0(n1747), .A1(n1098), .B0(n1830), .B1(
        \requesterAddressbuffer[1][3] ), .Y(n1025) );
  INVX2TS U1547 ( .A(n1017), .Y(n1099) );
  AOI22X1TS U1548 ( .A0(requesterAddressIn_WEST[3]), .A1(n1099), .B0(n1019), 
        .B1(n1018), .Y(n1024) );
  INVX2TS U1549 ( .A(n1020), .Y(n1836) );
  AOI22X1TS U1550 ( .A0(n1022), .A1(n1836), .B0(n1021), .B1(n1816), .Y(n1023)
         );
  AOI22X1TS U1551 ( .A0(readRequesterAddress[0]), .A1(n1852), .B0(n1880), .B1(
        \requesterAddressbuffer[0][0] ), .Y(n1031) );
  INVX2TS U1552 ( .A(n1060), .Y(n1864) );
  AOI22X1TS U1553 ( .A0(requesterAddressIn_WEST[0]), .A1(n1883), .B0(n1026), 
        .B1(n1864), .Y(n1030) );
  INVX2TS U1554 ( .A(n1027), .Y(n1069) );
  AOI22X1TS U1555 ( .A0(n1028), .A1(n1876), .B0(requesterAddressIn_NORTH[0]), 
        .B1(n1069), .Y(n1029) );
  INVX2TS U1556 ( .A(n11), .Y(n1862) );
  INVX2TS U1557 ( .A(n1032), .Y(n1074) );
  AOI22X1TS U1558 ( .A0(n1821), .A1(n1862), .B0(n1074), .B1(
        \requesterAddressbuffer[0][1] ), .Y(n1037) );
  INVX2TS U1559 ( .A(n1060), .Y(n1873) );
  AOI22X1TS U1560 ( .A0(requesterAddressIn_WEST[1]), .A1(n1068), .B0(n1033), 
        .B1(n1873), .Y(n1036) );
  AOI22X1TS U1561 ( .A0(n1034), .A1(n1070), .B0(requesterAddressIn_NORTH[1]), 
        .B1(n1885), .Y(n1035) );
  INVX2TS U1562 ( .A(n11), .Y(n1871) );
  AOI22X1TS U1563 ( .A0(n1832), .A1(n1871), .B0(n1074), .B1(
        \requesterAddressbuffer[0][2] ), .Y(n1042) );
  AOI22X1TS U1564 ( .A0(requesterAddressIn_WEST[2]), .A1(n1052), .B0(n1038), 
        .B1(n1045), .Y(n1041) );
  AOI22X1TS U1565 ( .A0(n1039), .A1(n1887), .B0(requesterAddressIn_NORTH[2]), 
        .B1(n1885), .Y(n1040) );
  INVX2TS U1566 ( .A(n11), .Y(n1881) );
  INVX2TS U1567 ( .A(n1043), .Y(n1870) );
  AOI22X1TS U1568 ( .A0(n1843), .A1(n1881), .B0(n1870), .B1(
        \requesterAddressbuffer[0][3] ), .Y(n1051) );
  INVX2TS U1569 ( .A(n1044), .Y(n1068) );
  AOI22X1TS U1570 ( .A0(requesterAddressIn_WEST[3]), .A1(n1068), .B0(n1046), 
        .B1(n1045), .Y(n1050) );
  INVX2TS U1571 ( .A(n1047), .Y(n1858) );
  AOI22X1TS U1572 ( .A0(n1048), .A1(n1858), .B0(requesterAddressIn_NORTH[3]), 
        .B1(n1053), .Y(n1049) );
  INVX2TS U1573 ( .A(n1043), .Y(n1064) );
  AOI21X1TS U1574 ( .A0(n1064), .A1(\dataoutbuffer[0][0] ), .B0(n1862), .Y(
        n1056) );
  AOI22X1TS U1575 ( .A0(n1052), .A1(n1391), .B0(n1864), .B1(n1108), .Y(n1055)
         );
  CLKBUFX2TS U1576 ( .A(dataIn_SOUTH[0]), .Y(n1501) );
  AOI22X1TS U1577 ( .A0(n1858), .A1(n1501), .B0(n1053), .B1(dataIn_NORTH[0]), 
        .Y(n1054) );
  AOI21X1TS U1578 ( .A0(n1064), .A1(\dataoutbuffer[0][1] ), .B0(n1871), .Y(
        n1059) );
  AOI22X1TS U1579 ( .A0(n414), .A1(n1397), .B0(n1873), .B1(n1339), .Y(n1058)
         );
  CLKBUFX2TS U1580 ( .A(dataIn_SOUTH[1]), .Y(n1508) );
  AOI22X1TS U1581 ( .A0(n1876), .A1(n1508), .B0(n409), .B1(dataIn_NORTH[1]), 
        .Y(n1057) );
  AOI21X1TS U1582 ( .A0(n1064), .A1(\dataoutbuffer[0][2] ), .B0(n1881), .Y(
        n1063) );
  AOI22X1TS U1583 ( .A0(n1068), .A1(n1402), .B0(n383), .B1(n1345), .Y(n1062)
         );
  CLKBUFX2TS U1584 ( .A(dataIn_SOUTH[2]), .Y(n1516) );
  AOI22X1TS U1585 ( .A0(n1887), .A1(n1516), .B0(n1069), .B1(dataIn_NORTH[2]), 
        .Y(n1061) );
  AOI21X1TS U1586 ( .A0(n1064), .A1(\dataoutbuffer[0][3] ), .B0(n1862), .Y(
        n1067) );
  AOI22X1TS U1587 ( .A0(n1854), .A1(n1407), .B0(n1864), .B1(n1350), .Y(n1066)
         );
  CLKBUFX2TS U1588 ( .A(dataIn_SOUTH[3]), .Y(n1525) );
  AOI22X1TS U1589 ( .A0(n436), .A1(n1525), .B0(n1856), .B1(dataIn_NORTH[3]), 
        .Y(n1065) );
  AOI21X1TS U1590 ( .A0(n1074), .A1(\dataoutbuffer[0][4] ), .B0(n1871), .Y(
        n1073) );
  AOI22X1TS U1591 ( .A0(n1068), .A1(n1411), .B0(n1873), .B1(n1355), .Y(n1072)
         );
  CLKBUFX2TS U1592 ( .A(dataIn_SOUTH[4]), .Y(n1532) );
  AOI22X1TS U1593 ( .A0(n1070), .A1(n1532), .B0(n1069), .B1(dataIn_NORTH[4]), 
        .Y(n1071) );
  AOI21X1TS U1594 ( .A0(n1074), .A1(\dataoutbuffer[0][5] ), .B0(n1881), .Y(
        n1077) );
  AOI22X1TS U1595 ( .A0(n414), .A1(n1419), .B0(n383), .B1(n1361), .Y(n1076) );
  CLKBUFX2TS U1596 ( .A(dataIn_SOUTH[5]), .Y(n1539) );
  AOI22X1TS U1597 ( .A0(n1858), .A1(n1539), .B0(n389), .B1(dataIn_NORTH[5]), 
        .Y(n1075) );
  INVX2TS U1598 ( .A(n1620), .Y(n1093) );
  AOI21X1TS U1599 ( .A0(n1093), .A1(\dataoutbuffer[1][0] ), .B0(n1098), .Y(
        n1083) );
  AOI22X1TS U1600 ( .A0(n1078), .A1(dataIn_WEST[0]), .B0(n1823), .B1(n1108), 
        .Y(n1082) );
  CLKBUFX2TS U1601 ( .A(dataIn_NORTH[0]), .Y(n1426) );
  CLKBUFX2TS U1602 ( .A(n1426), .Y(n1500) );
  CLKBUFX2TS U1603 ( .A(n1501), .Y(n1461) );
  AOI22X1TS U1604 ( .A0(n1080), .A1(n1500), .B0(n1079), .B1(n1461), .Y(n1081)
         );
  INVX2TS U1605 ( .A(n1084), .Y(n1820) );
  AOI21X1TS U1606 ( .A0(n1093), .A1(\dataoutbuffer[1][1] ), .B0(n1820), .Y(
        n1088) );
  AOI22X1TS U1607 ( .A0(n328), .A1(dataIn_WEST[1]), .B0(n1834), .B1(n1339), 
        .Y(n1087) );
  INVX2TS U1608 ( .A(n1085), .Y(n1826) );
  CLKBUFX2TS U1609 ( .A(dataIn_NORTH[1]), .Y(n1431) );
  CLKBUFX2TS U1610 ( .A(n1431), .Y(n1507) );
  CLKBUFX2TS U1611 ( .A(n1508), .Y(n1468) );
  AOI22X1TS U1612 ( .A0(n1826), .A1(n1507), .B0(n1104), .B1(n1468), .Y(n1086)
         );
  AOI21X1TS U1613 ( .A0(n1093), .A1(\dataoutbuffer[1][2] ), .B0(n1831), .Y(
        n1092) );
  AOI22X1TS U1614 ( .A0(n1099), .A1(dataIn_WEST[2]), .B0(n309), .B1(n1345), 
        .Y(n1091) );
  CLKBUFX2TS U1615 ( .A(dataIn_NORTH[2]), .Y(n1436) );
  CLKBUFX2TS U1616 ( .A(n1436), .Y(n1514) );
  CLKBUFX2TS U1617 ( .A(n1516), .Y(n1474) );
  AOI22X1TS U1618 ( .A0(n1011), .A1(n1514), .B0(n1836), .B1(n1474), .Y(n1090)
         );
  AOI21X1TS U1619 ( .A0(n1093), .A1(\dataoutbuffer[1][3] ), .B0(n1842), .Y(
        n1097) );
  AOI22X1TS U1620 ( .A0(n1813), .A1(dataIn_WEST[3]), .B0(n1823), .B1(n1350), 
        .Y(n1096) );
  CLKBUFX2TS U1621 ( .A(dataIn_NORTH[3]), .Y(n1442) );
  CLKBUFX2TS U1622 ( .A(n1442), .Y(n1524) );
  CLKBUFX2TS U1623 ( .A(n1525), .Y(n1480) );
  AOI22X1TS U1624 ( .A0(n1816), .A1(n1524), .B0(n1094), .B1(n1480), .Y(n1095)
         );
  AOI21X1TS U1625 ( .A0(n1103), .A1(\dataoutbuffer[1][4] ), .B0(n1098), .Y(
        n1102) );
  AOI22X1TS U1626 ( .A0(n1099), .A1(dataIn_WEST[4]), .B0(n1834), .B1(n1355), 
        .Y(n1101) );
  CLKBUFX2TS U1627 ( .A(dataIn_NORTH[4]), .Y(n1448) );
  CLKBUFX2TS U1628 ( .A(n1448), .Y(n1530) );
  CLKBUFX2TS U1629 ( .A(n1532), .Y(n1486) );
  AOI22X1TS U1630 ( .A0(n314), .A1(n1530), .B0(n350), .B1(n1486), .Y(n1100) );
  AOI21X1TS U1631 ( .A0(n1103), .A1(\dataoutbuffer[1][5] ), .B0(n1820), .Y(
        n1107) );
  AOI22X1TS U1632 ( .A0(n328), .A1(dataIn_WEST[5]), .B0(n309), .B1(n1361), .Y(
        n1106) );
  CLKBUFX2TS U1633 ( .A(dataIn_NORTH[5]), .Y(n1454) );
  CLKBUFX2TS U1634 ( .A(n1454), .Y(n1538) );
  CLKBUFX2TS U1635 ( .A(n1539), .Y(n1494) );
  AOI22X1TS U1636 ( .A0(n1826), .A1(n1538), .B0(n1104), .B1(n1494), .Y(n1105)
         );
  INVX2TS U1637 ( .A(n1606), .Y(n1349) );
  AOI21X1TS U1638 ( .A0(n1349), .A1(\dataoutbuffer[2][0] ), .B0(n1792), .Y(
        n1338) );
  AOI22X1TS U1639 ( .A0(n1109), .A1(dataIn_WEST[0]), .B0(n1793), .B1(n1108), 
        .Y(n1337) );
  AOI22X1TS U1640 ( .A0(n1111), .A1(n1500), .B0(n1110), .B1(dataIn_SOUTH[0]), 
        .Y(n1112) );
  AOI21X1TS U1641 ( .A0(n1349), .A1(\dataoutbuffer[2][1] ), .B0(n1799), .Y(
        n1343) );
  AOI22X1TS U1642 ( .A0(n184), .A1(dataIn_WEST[1]), .B0(n1800), .B1(n1339), 
        .Y(n1342) );
  INVX2TS U1643 ( .A(n1340), .Y(n1794) );
  AOI22X1TS U1644 ( .A0(n1794), .A1(n1507), .B0(n1362), .B1(dataIn_SOUTH[1]), 
        .Y(n1341) );
  AOI21X1TS U1645 ( .A0(n1349), .A1(\dataoutbuffer[2][2] ), .B0(n175), .Y(
        n1348) );
  AOI22X1TS U1646 ( .A0(n1356), .A1(dataIn_WEST[2]), .B0(n174), .B1(n1345), 
        .Y(n1347) );
  AOI22X1TS U1647 ( .A0(n985), .A1(n1514), .B0(n1801), .B1(dataIn_SOUTH[2]), 
        .Y(n1346) );
  AOI21X1TS U1648 ( .A0(n1349), .A1(\dataoutbuffer[2][3] ), .B0(n1792), .Y(
        n1354) );
  AOI22X1TS U1649 ( .A0(n1787), .A1(dataIn_WEST[3]), .B0(n1793), .B1(n1350), 
        .Y(n1353) );
  AOI22X1TS U1650 ( .A0(n1788), .A1(n1524), .B0(n1351), .B1(dataIn_SOUTH[3]), 
        .Y(n1352) );
  AOI21X1TS U1651 ( .A0(n1360), .A1(\dataoutbuffer[2][4] ), .B0(n1799), .Y(
        n1359) );
  AOI22X1TS U1652 ( .A0(n1356), .A1(dataIn_WEST[4]), .B0(n1800), .B1(n1355), 
        .Y(n1358) );
  AOI22X1TS U1653 ( .A0(n202), .A1(n1530), .B0(n206), .B1(dataIn_SOUTH[4]), 
        .Y(n1357) );
  AOI21X1TS U1654 ( .A0(n1360), .A1(\dataoutbuffer[2][5] ), .B0(n175), .Y(
        n1365) );
  AOI22X1TS U1655 ( .A0(n184), .A1(dataIn_WEST[5]), .B0(n174), .B1(n1361), .Y(
        n1364) );
  AOI22X1TS U1656 ( .A0(n1794), .A1(n1538), .B0(n1362), .B1(dataIn_SOUTH[5]), 
        .Y(n1363) );
  INVX2TS U1657 ( .A(n168), .Y(n1377) );
  AOI21X1TS U1658 ( .A0(n1377), .A1(\dataoutbuffer[3][0] ), .B0(n1762), .Y(
        n1370) );
  AOI22X1TS U1659 ( .A0(n134), .A1(dataIn_WEST[0]), .B0(n1770), .B1(
        dataIn_EAST[0]), .Y(n1369) );
  AOI22X1TS U1660 ( .A0(n1367), .A1(n1426), .B0(n1765), .B1(n1461), .Y(n1368)
         );
  AOI21X1TS U1661 ( .A0(n1377), .A1(\dataoutbuffer[3][1] ), .B0(n126), .Y(
        n1373) );
  AOI22X1TS U1662 ( .A0(n141), .A1(dataIn_WEST[1]), .B0(n1763), .B1(
        dataIn_EAST[1]), .Y(n1372) );
  AOI22X1TS U1663 ( .A0(n140), .A1(n1431), .B0(n1772), .B1(n1468), .Y(n1371)
         );
  AOI21X1TS U1664 ( .A0(n1377), .A1(\dataoutbuffer[3][2] ), .B0(n1777), .Y(
        n1376) );
  AOI22X1TS U1665 ( .A0(n134), .A1(dataIn_WEST[2]), .B0(n162), .B1(
        dataIn_EAST[2]), .Y(n1375) );
  AOI22X1TS U1666 ( .A0(n140), .A1(n1436), .B0(n1781), .B1(n1474), .Y(n1374)
         );
  AOI21X1TS U1667 ( .A0(n1377), .A1(\dataoutbuffer[3][3] ), .B0(n1762), .Y(
        n1380) );
  AOI22X1TS U1668 ( .A0(n1757), .A1(dataIn_WEST[3]), .B0(n128), .B1(
        dataIn_EAST[3]), .Y(n1379) );
  AOI22X1TS U1669 ( .A0(n1758), .A1(n1442), .B0(n125), .B1(n1480), .Y(n1378)
         );
  AOI21X1TS U1670 ( .A0(n1385), .A1(\dataoutbuffer[3][4] ), .B0(n126), .Y(
        n1384) );
  AOI22X1TS U1671 ( .A0(n955), .A1(dataIn_WEST[4]), .B0(n1381), .B1(
        dataIn_EAST[4]), .Y(n1383) );
  AOI22X1TS U1672 ( .A0(n140), .A1(n1448), .B0(n1781), .B1(n1486), .Y(n1382)
         );
  AOI21X1TS U1673 ( .A0(n1385), .A1(\dataoutbuffer[3][5] ), .B0(n1777), .Y(
        n1389) );
  AOI22X1TS U1674 ( .A0(n1386), .A1(dataIn_WEST[5]), .B0(n1763), .B1(
        dataIn_EAST[5]), .Y(n1388) );
  AOI22X1TS U1675 ( .A0(n957), .A1(n1454), .B0(n125), .B1(n1494), .Y(n1387) );
  INVX2TS U1676 ( .A(n938), .Y(n1406) );
  AOI21X1TS U1677 ( .A0(n1406), .A1(\dataoutbuffer[4][0] ), .B0(n1732), .Y(
        n1396) );
  AOI22X1TS U1678 ( .A0(n1392), .A1(n1391), .B0(n1734), .B1(dataIn_EAST[0]), 
        .Y(n1395) );
  AOI22X1TS U1679 ( .A0(n1728), .A1(dataIn_SOUTH[0]), .B0(n1393), .B1(n1500), 
        .Y(n1394) );
  AOI21X1TS U1680 ( .A0(n1406), .A1(\dataoutbuffer[4][1] ), .B0(n268), .Y(
        n1400) );
  AOI22X1TS U1681 ( .A0(n283), .A1(n1397), .B0(n1740), .B1(dataIn_EAST[1]), 
        .Y(n1399) );
  AOI22X1TS U1682 ( .A0(n1741), .A1(dataIn_SOUTH[1]), .B0(n1413), .B1(n1507), 
        .Y(n1398) );
  AOI21X1TS U1683 ( .A0(n1406), .A1(\dataoutbuffer[4][2] ), .B0(n1746), .Y(
        n1405) );
  AOI22X1TS U1684 ( .A0(n1412), .A1(n1402), .B0(n267), .B1(dataIn_EAST[2]), 
        .Y(n1404) );
  AOI22X1TS U1685 ( .A0(n1750), .A1(dataIn_SOUTH[2]), .B0(n1413), .B1(n1514), 
        .Y(n1403) );
  AOI21X1TS U1686 ( .A0(n1406), .A1(\dataoutbuffer[4][3] ), .B0(n1732), .Y(
        n1410) );
  AOI22X1TS U1687 ( .A0(n1726), .A1(n1407), .B0(n1734), .B1(dataIn_EAST[3]), 
        .Y(n1409) );
  AOI22X1TS U1688 ( .A0(n300), .A1(dataIn_SOUTH[3]), .B0(n1727), .B1(n1524), 
        .Y(n1408) );
  AOI21X1TS U1689 ( .A0(n1418), .A1(\dataoutbuffer[4][4] ), .B0(n268), .Y(
        n1417) );
  AOI22X1TS U1690 ( .A0(n1412), .A1(n1411), .B0(n1740), .B1(dataIn_EAST[4]), 
        .Y(n1416) );
  AOI22X1TS U1691 ( .A0(n1414), .A1(dataIn_SOUTH[4]), .B0(n1413), .B1(n1530), 
        .Y(n1415) );
  AOI21X1TS U1692 ( .A0(n1418), .A1(\dataoutbuffer[4][5] ), .B0(n1746), .Y(
        n1422) );
  AOI22X1TS U1693 ( .A0(n283), .A1(n1419), .B0(n267), .B1(dataIn_EAST[5]), .Y(
        n1421) );
  AOI22X1TS U1694 ( .A0(n1728), .A1(dataIn_SOUTH[5]), .B0(n275), .B1(n1538), 
        .Y(n1420) );
  INVX2TS U1695 ( .A(n915), .Y(n1441) );
  AOI21X1TS U1696 ( .A0(n1441), .A1(\dataoutbuffer[5][0] ), .B0(n1700), .Y(
        n1430) );
  AOI22X1TS U1697 ( .A0(n1424), .A1(n1499), .B0(n1702), .B1(n1459), .Y(n1429)
         );
  AOI22X1TS U1698 ( .A0(n1427), .A1(n1426), .B0(n1425), .B1(n1461), .Y(n1428)
         );
  AOI21X1TS U1699 ( .A0(n1441), .A1(\dataoutbuffer[5][1] ), .B0(n1709), .Y(
        n1434) );
  AOI22X1TS U1700 ( .A0(n236), .A1(n1506), .B0(n1711), .B1(n1467), .Y(n1433)
         );
  AOI22X1TS U1701 ( .A0(n1704), .A1(n1431), .B0(n1721), .B1(n1468), .Y(n1432)
         );
  AOI21X1TS U1702 ( .A0(n1441), .A1(\dataoutbuffer[5][2] ), .B0(n1717), .Y(
        n1440) );
  AOI22X1TS U1703 ( .A0(n1446), .A1(n1513), .B0(n216), .B1(n1473), .Y(n1439)
         );
  AOI22X1TS U1704 ( .A0(n1437), .A1(n1436), .B0(n1447), .B1(n1474), .Y(n1438)
         );
  AOI21X1TS U1705 ( .A0(n1441), .A1(\dataoutbuffer[5][3] ), .B0(n1700), .Y(
        n1445) );
  AOI22X1TS U1706 ( .A0(n1694), .A1(n1522), .B0(n1702), .B1(n1479), .Y(n1444)
         );
  AOI22X1TS U1707 ( .A0(n222), .A1(n1442), .B0(n1695), .B1(n1480), .Y(n1443)
         );
  AOI21X1TS U1708 ( .A0(n1453), .A1(\dataoutbuffer[5][4] ), .B0(n1709), .Y(
        n1452) );
  AOI22X1TS U1709 ( .A0(n1446), .A1(n1529), .B0(n1711), .B1(n1484), .Y(n1451)
         );
  AOI22X1TS U1710 ( .A0(n1449), .A1(n1448), .B0(n1447), .B1(n1486), .Y(n1450)
         );
  AOI21X1TS U1711 ( .A0(n1453), .A1(\dataoutbuffer[5][5] ), .B0(n1717), .Y(
        n1457) );
  AOI22X1TS U1712 ( .A0(n236), .A1(n1537), .B0(n216), .B1(n1493), .Y(n1456) );
  AOI22X1TS U1713 ( .A0(n1704), .A1(n1454), .B0(n238), .B1(n1494), .Y(n1455)
         );
  INVX2TS U1714 ( .A(n897), .Y(n1478) );
  AOI21X1TS U1715 ( .A0(n1478), .A1(\dataoutbuffer[6][0] ), .B0(n1669), .Y(
        n1466) );
  AOI22X1TS U1716 ( .A0(n1460), .A1(n1499), .B0(n1670), .B1(n1459), .Y(n1465)
         );
  AOI22X1TS U1717 ( .A0(n1463), .A1(dataIn_NORTH[0]), .B0(n1462), .B1(n1461), 
        .Y(n1464) );
  AOI21X1TS U1718 ( .A0(n1478), .A1(\dataoutbuffer[6][1] ), .B0(n78), .Y(n1471) );
  AOI22X1TS U1719 ( .A0(n80), .A1(n1506), .B0(n1676), .B1(n1467), .Y(n1470) );
  AOI22X1TS U1720 ( .A0(n99), .A1(dataIn_NORTH[1]), .B0(n1487), .B1(n1468), 
        .Y(n1469) );
  AOI21X1TS U1721 ( .A0(n1478), .A1(\dataoutbuffer[6][2] ), .B0(n1683), .Y(
        n1477) );
  AOI22X1TS U1722 ( .A0(n1485), .A1(n1513), .B0(n77), .B1(n1473), .Y(n1476) );
  AOI22X1TS U1723 ( .A0(n1488), .A1(dataIn_NORTH[2]), .B0(n1487), .B1(n1474), 
        .Y(n1475) );
  AOI21X1TS U1724 ( .A0(n1478), .A1(\dataoutbuffer[6][3] ), .B0(n1669), .Y(
        n1483) );
  AOI22X1TS U1725 ( .A0(n1663), .A1(n1522), .B0(n1670), .B1(n1479), .Y(n1482)
         );
  AOI22X1TS U1726 ( .A0(n1665), .A1(dataIn_NORTH[3]), .B0(n111), .B1(n1480), 
        .Y(n1481) );
  AOI21X1TS U1727 ( .A0(n1492), .A1(\dataoutbuffer[6][4] ), .B0(n78), .Y(n1491) );
  AOI22X1TS U1728 ( .A0(n1485), .A1(n1529), .B0(n1676), .B1(n1484), .Y(n1490)
         );
  AOI22X1TS U1729 ( .A0(n1488), .A1(dataIn_NORTH[4]), .B0(n1487), .B1(n1486), 
        .Y(n1489) );
  AOI21X1TS U1730 ( .A0(n1492), .A1(\dataoutbuffer[6][5] ), .B0(n1683), .Y(
        n1497) );
  AOI22X1TS U1731 ( .A0(n80), .A1(n1537), .B0(n77), .B1(n1493), .Y(n1496) );
  AOI22X1TS U1732 ( .A0(n99), .A1(dataIn_NORTH[5]), .B0(n105), .B1(n1494), .Y(
        n1495) );
  INVX2TS U1733 ( .A(n881), .Y(n1521) );
  AOI21X1TS U1734 ( .A0(n1521), .A1(\dataoutbuffer[7][0] ), .B0(n1640), .Y(
        n1504) );
  AOI22X1TS U1735 ( .A0(n47), .A1(n1499), .B0(n1655), .B1(dataIn_EAST[0]), .Y(
        n1503) );
  AOI22X1TS U1736 ( .A0(n68), .A1(n1501), .B0(n1515), .B1(n1500), .Y(n1502) );
  AOI21X1TS U1737 ( .A0(n1521), .A1(\dataoutbuffer[7][1] ), .B0(n32), .Y(n1511) );
  AOI22X1TS U1738 ( .A0(n52), .A1(n1506), .B0(n1641), .B1(dataIn_EAST[1]), .Y(
        n1510) );
  AOI22X1TS U1739 ( .A0(n1658), .A1(n1508), .B0(n49), .B1(n1507), .Y(n1509) );
  AOI21X1TS U1740 ( .A0(n1521), .A1(\dataoutbuffer[7][2] ), .B0(n1654), .Y(
        n1520) );
  AOI22X1TS U1741 ( .A0(n47), .A1(n1513), .B0(n31), .B1(dataIn_EAST[2]), .Y(
        n1519) );
  AOI22X1TS U1742 ( .A0(n1517), .A1(n1516), .B0(n1515), .B1(n1514), .Y(n1518)
         );
  AOI21X1TS U1743 ( .A0(n1521), .A1(\dataoutbuffer[7][3] ), .B0(n1640), .Y(
        n1528) );
  AOI22X1TS U1744 ( .A0(n1523), .A1(n1522), .B0(n1655), .B1(dataIn_EAST[3]), 
        .Y(n1527) );
  AOI22X1TS U1745 ( .A0(n1635), .A1(n1525), .B0(n1657), .B1(n1524), .Y(n1526)
         );
  AOI21X1TS U1746 ( .A0(n1536), .A1(\dataoutbuffer[7][4] ), .B0(n1634), .Y(
        n1535) );
  AOI22X1TS U1747 ( .A0(n1647), .A1(n1529), .B0(n1641), .B1(dataIn_EAST[4]), 
        .Y(n1534) );
  AOI22X1TS U1748 ( .A0(n1648), .A1(n1532), .B0(n1531), .B1(n1530), .Y(n1533)
         );
  AOI21X1TS U1749 ( .A0(n1536), .A1(\dataoutbuffer[7][5] ), .B0(n1654), .Y(
        n1542) );
  AOI22X1TS U1750 ( .A0(n61), .A1(n1537), .B0(n31), .B1(dataIn_EAST[5]), .Y(
        n1541) );
  AOI22X1TS U1751 ( .A0(n1635), .A1(n1539), .B0(n49), .B1(n1538), .Y(n1540) );
  INVX2TS U1752 ( .A(n1543), .Y(n1613) );
  AOI22X1TS U1753 ( .A0(n1545), .A1(n1566), .B0(n1565), .B1(n1544), .Y(n1547)
         );
  AOI22X1TS U1754 ( .A0(n1548), .A1(n1613), .B0(n1547), .B1(n1546), .Y(n1550)
         );
  AOI22X1TS U1755 ( .A0(n1551), .A1(n1617), .B0(n1550), .B1(n1549), .Y(n1553)
         );
  AOI32X1TS U1756 ( .A0(n1553), .A1(n1498), .A2(n1552), .B0(n1652), .B1(n1921), 
        .Y(n2048) );
  INVX2TS U1757 ( .A(n1543), .Y(n1627) );
  AOI22X1TS U1758 ( .A0(n1555), .A1(n1566), .B0(n1565), .B1(n1554), .Y(n1557)
         );
  AOI22X1TS U1759 ( .A0(n1558), .A1(n1627), .B0(n1557), .B1(n1556), .Y(n1560)
         );
  AOI22X1TS U1760 ( .A0(n1561), .A1(n1583), .B0(n1560), .B1(n1559), .Y(n1563)
         );
  AOI32X1TS U1761 ( .A0(n1563), .A1(n1458), .A2(n1562), .B0(n1682), .B1(n1922), 
        .Y(n2049) );
  AOI22X1TS U1762 ( .A0(n1567), .A1(n1566), .B0(n1565), .B1(n1564), .Y(n1569)
         );
  AOI22X1TS U1763 ( .A0(n1570), .A1(n1613), .B0(n1569), .B1(n1568), .Y(n1572)
         );
  AOI22X1TS U1764 ( .A0(n1573), .A1(n1583), .B0(n1572), .B1(n1571), .Y(n1575)
         );
  AOI32X1TS U1765 ( .A0(n1575), .A1(n1423), .A2(n1574), .B0(n1716), .B1(n1923), 
        .Y(n2050) );
  CLKBUFX2TS U1766 ( .A(n1623), .Y(n1609) );
  AOI22X1TS U1767 ( .A0(n1577), .A1(n1609), .B0(n1597), .B1(n1576), .Y(n1579)
         );
  AOI22X1TS U1768 ( .A0(n1580), .A1(n1627), .B0(n1579), .B1(n1578), .Y(n1582)
         );
  AOI22X1TS U1769 ( .A0(n1584), .A1(n1583), .B0(n1582), .B1(n1581), .Y(n1586)
         );
  AOI32X1TS U1770 ( .A0(n1586), .A1(n1390), .A2(n1585), .B0(n1745), .B1(n1924), 
        .Y(n2051) );
  AOI22X1TS U1771 ( .A0(n115), .A1(n1609), .B0(readIn_NORTH), .B1(n1587), .Y(
        n1589) );
  AOI22X1TS U1772 ( .A0(n1590), .A1(n1613), .B0(n1589), .B1(n1588), .Y(n1592)
         );
  AOI22X1TS U1773 ( .A0(n1593), .A1(readIn_WEST), .B0(n1592), .B1(n1591), .Y(
        n1595) );
  AOI32X1TS U1774 ( .A0(n1595), .A1(n1366), .A2(n1594), .B0(n1776), .B1(n1925), 
        .Y(n2052) );
  AOI22X1TS U1775 ( .A0(n1598), .A1(n1609), .B0(n1597), .B1(n1596), .Y(n1600)
         );
  AOI22X1TS U1776 ( .A0(n1601), .A1(n1627), .B0(n1600), .B1(n1599), .Y(n1603)
         );
  AOI22X1TS U1777 ( .A0(n1604), .A1(readIn_WEST), .B0(n1603), .B1(n1602), .Y(
        n1607) );
  AOI32X1TS U1778 ( .A0(n1607), .A1(n1606), .A2(n1605), .B0(n1805), .B1(n1926), 
        .Y(n2053) );
  AOI22X1TS U1779 ( .A0(n1610), .A1(n1609), .B0(readIn_NORTH), .B1(n1608), .Y(
        n1612) );
  AOI22X1TS U1780 ( .A0(n1614), .A1(n1613), .B0(n1612), .B1(n1611), .Y(n1616)
         );
  AOI22X1TS U1781 ( .A0(n1618), .A1(n1617), .B0(n1616), .B1(n1615), .Y(n1621)
         );
  AOI32X1TS U1782 ( .A0(n1621), .A1(n1620), .A2(n1619), .B0(n1841), .B1(n1927), 
        .Y(n2054) );
  AOI22X1TS U1783 ( .A0(n1624), .A1(n1623), .B0(readIn_NORTH), .B1(n1622), .Y(
        n1626) );
  AOI22X1TS U1784 ( .A0(n1628), .A1(n1627), .B0(n1626), .B1(n1625), .Y(n1630)
         );
  AOI22X1TS U1785 ( .A0(n1631), .A1(readIn_WEST), .B0(n1630), .B1(n1629), .Y(
        n1633) );
  AOI32X1TS U1786 ( .A0(n1633), .A1(n1043), .A2(n1632), .B0(n1880), .B1(n1928), 
        .Y(n2055) );
  AOI22X1TS U1787 ( .A0(n1811), .A1(n1634), .B0(n1645), .B1(
        \destinationAddressbuffer[7][0] ), .Y(n1638) );
  AOI22X1TS U1788 ( .A0(n52), .A1(n1693), .B0(n875), .B1(n1692), .Y(n1637) );
  CLKBUFX2TS U1789 ( .A(n1664), .Y(n1815) );
  AOI22X1TS U1790 ( .A0(n1635), .A1(destinationAddressIn_SOUTH[0]), .B0(n1531), 
        .B1(n1815), .Y(n1636) );
  AOI22X1TS U1791 ( .A0(n1640), .A1(n1639), .B0(n1645), .B1(
        \destinationAddressbuffer[7][1] ), .Y(n1644) );
  AOI22X1TS U1792 ( .A0(n61), .A1(n1703), .B0(n1641), .B1(n1701), .Y(n1643) );
  CLKBUFX2TS U1793 ( .A(n1671), .Y(n1825) );
  AOI22X1TS U1794 ( .A0(n39), .A1(destinationAddressIn_SOUTH[1]), .B0(n1515), 
        .B1(n1825), .Y(n1642) );
  AOI22X1TS U1795 ( .A0(n32), .A1(n1646), .B0(n1645), .B1(
        \destinationAddressbuffer[7][2] ), .Y(n1651) );
  AOI22X1TS U1796 ( .A0(n1647), .A1(n1712), .B0(n31), .B1(n1710), .Y(n1650) );
  CLKBUFX2TS U1797 ( .A(n1677), .Y(n1837) );
  AOI22X1TS U1798 ( .A0(n1648), .A1(destinationAddressIn_SOUTH[2]), .B0(n67), 
        .B1(n1837), .Y(n1649) );
  AOI22X1TS U1799 ( .A0(n1654), .A1(n1653), .B0(n1652), .B1(
        \destinationAddressbuffer[7][3] ), .Y(n1661) );
  AOI22X1TS U1800 ( .A0(n1656), .A1(n1719), .B0(n1655), .B1(n1718), .Y(n1660)
         );
  CLKBUFX2TS U1801 ( .A(n1685), .Y(n1847) );
  AOI22X1TS U1802 ( .A0(n1658), .A1(destinationAddressIn_SOUTH[3]), .B0(n1657), 
        .B1(n1847), .Y(n1659) );
  AOI22X1TS U1803 ( .A0(n1853), .A1(n1662), .B0(n1675), .B1(
        \destinationAddressbuffer[6][0] ), .Y(n1668) );
  AOI22X1TS U1804 ( .A0(n1663), .A1(n1693), .B0(n899), .B1(n1692), .Y(n1667)
         );
  CLKBUFX2TS U1805 ( .A(n1664), .Y(n1855) );
  CLKBUFX2TS U1806 ( .A(destinationAddressIn_SOUTH[0]), .Y(n1857) );
  CLKBUFX2TS U1807 ( .A(n1857), .Y(n1814) );
  AOI22X1TS U1808 ( .A0(n1665), .A1(n1855), .B0(n1686), .B1(n1814), .Y(n1666)
         );
  AOI22X1TS U1809 ( .A0(n1733), .A1(n1669), .B0(n1675), .B1(
        \destinationAddressbuffer[6][1] ), .Y(n1674) );
  AOI22X1TS U1810 ( .A0(n109), .A1(n1703), .B0(n1670), .B1(n1701), .Y(n1673)
         );
  CLKBUFX2TS U1811 ( .A(n1671), .Y(n1865) );
  CLKBUFX2TS U1812 ( .A(destinationAddressIn_SOUTH[1]), .Y(n1866) );
  CLKBUFX2TS U1813 ( .A(n1866), .Y(n1824) );
  AOI22X1TS U1814 ( .A0(n99), .A1(n1865), .B0(n1678), .B1(n1824), .Y(n1672) );
  AOI22X1TS U1815 ( .A0(n1739), .A1(n78), .B0(n1675), .B1(
        \destinationAddressbuffer[6][2] ), .Y(n1681) );
  AOI22X1TS U1816 ( .A0(n1684), .A1(n1712), .B0(n1676), .B1(n1710), .Y(n1680)
         );
  CLKBUFX2TS U1817 ( .A(n1677), .Y(n1874) );
  CLKBUFX2TS U1818 ( .A(destinationAddressIn_SOUTH[2]), .Y(n1875) );
  CLKBUFX2TS U1819 ( .A(n1875), .Y(n1835) );
  AOI22X1TS U1820 ( .A0(n1687), .A1(n1874), .B0(n1678), .B1(n1835), .Y(n1679)
         );
  AOI22X1TS U1821 ( .A0(n1747), .A1(n1683), .B0(n1682), .B1(
        \destinationAddressbuffer[6][3] ), .Y(n1690) );
  AOI22X1TS U1822 ( .A0(n1684), .A1(n1719), .B0(n77), .B1(n1718), .Y(n1689) );
  CLKBUFX2TS U1823 ( .A(n1685), .Y(n1884) );
  CLKBUFX2TS U1824 ( .A(destinationAddressIn_SOUTH[3]), .Y(n1886) );
  CLKBUFX2TS U1825 ( .A(n1886), .Y(n1846) );
  AOI22X1TS U1826 ( .A0(n1687), .A1(n1884), .B0(n1686), .B1(n1846), .Y(n1688)
         );
  AOI22X1TS U1827 ( .A0(n1853), .A1(n1691), .B0(n1708), .B1(
        \destinationAddressbuffer[5][0] ), .Y(n1699) );
  AOI22X1TS U1828 ( .A0(n1694), .A1(n1693), .B0(n917), .B1(n1692), .Y(n1698)
         );
  AOI22X1TS U1829 ( .A0(n1696), .A1(n1855), .B0(n1695), .B1(
        destinationAddressIn_SOUTH[0]), .Y(n1697) );
  AOI22X1TS U1830 ( .A0(readRequesterAddress[1]), .A1(n1700), .B0(n1708), .B1(
        \destinationAddressbuffer[5][1] ), .Y(n1707) );
  AOI22X1TS U1831 ( .A0(n250), .A1(n1703), .B0(n1702), .B1(n1701), .Y(n1706)
         );
  AOI22X1TS U1832 ( .A0(n1704), .A1(n1865), .B0(n231), .B1(
        destinationAddressIn_SOUTH[1]), .Y(n1705) );
  AOI22X1TS U1833 ( .A0(readRequesterAddress[2]), .A1(n1709), .B0(n1708), .B1(
        \destinationAddressbuffer[5][2] ), .Y(n1715) );
  AOI22X1TS U1834 ( .A0(n1720), .A1(n1712), .B0(n1711), .B1(n1710), .Y(n1714)
         );
  AOI22X1TS U1835 ( .A0(n1427), .A1(n1874), .B0(n1721), .B1(
        destinationAddressIn_SOUTH[2]), .Y(n1713) );
  AOI22X1TS U1836 ( .A0(readRequesterAddress[3]), .A1(n1717), .B0(n1716), .B1(
        \destinationAddressbuffer[5][3] ), .Y(n1724) );
  AOI22X1TS U1837 ( .A0(n1720), .A1(n1719), .B0(n216), .B1(n1718), .Y(n1723)
         );
  AOI22X1TS U1838 ( .A0(n222), .A1(n1884), .B0(n1721), .B1(
        destinationAddressIn_SOUTH[3]), .Y(n1722) );
  AOI22X1TS U1839 ( .A0(n1755), .A1(n1725), .B0(n1738), .B1(
        \destinationAddressbuffer[4][0] ), .Y(n1731) );
  AOI22X1TS U1840 ( .A0(n1726), .A1(n1756), .B0(n940), .B1(
        destinationAddressIn_EAST[0]), .Y(n1730) );
  AOI22X1TS U1841 ( .A0(n1728), .A1(n1857), .B0(n1727), .B1(n1855), .Y(n1729)
         );
  AOI22X1TS U1842 ( .A0(n1733), .A1(n1732), .B0(n1738), .B1(
        \destinationAddressbuffer[4][1] ), .Y(n1737) );
  AOI22X1TS U1843 ( .A0(n295), .A1(n1764), .B0(n1734), .B1(
        destinationAddressIn_EAST[1]), .Y(n1736) );
  AOI22X1TS U1844 ( .A0(n285), .A1(n1866), .B0(n922), .B1(n1865), .Y(n1735) );
  AOI22X1TS U1845 ( .A0(n1739), .A1(n268), .B0(n1738), .B1(
        \destinationAddressbuffer[4][2] ), .Y(n1744) );
  AOI22X1TS U1846 ( .A0(n1748), .A1(n1771), .B0(n1740), .B1(
        destinationAddressIn_EAST[2]), .Y(n1743) );
  AOI22X1TS U1847 ( .A0(n1741), .A1(n1875), .B0(n1749), .B1(n1874), .Y(n1742)
         );
  AOI22X1TS U1848 ( .A0(n1747), .A1(n1746), .B0(n1745), .B1(
        \destinationAddressbuffer[4][3] ), .Y(n1753) );
  AOI22X1TS U1849 ( .A0(n1748), .A1(n1779), .B0(n267), .B1(
        destinationAddressIn_EAST[3]), .Y(n1752) );
  AOI22X1TS U1850 ( .A0(n1750), .A1(n1886), .B0(n1749), .B1(n1884), .Y(n1751)
         );
  AOI22X1TS U1851 ( .A0(n1755), .A1(n1754), .B0(n1769), .B1(
        \destinationAddressbuffer[3][0] ), .Y(n1761) );
  AOI22X1TS U1852 ( .A0(n1757), .A1(n1756), .B0(n128), .B1(
        destinationAddressIn_EAST[0]), .Y(n1760) );
  AOI22X1TS U1853 ( .A0(n1758), .A1(n1815), .B0(n1765), .B1(n1814), .Y(n1759)
         );
  AOI22X1TS U1854 ( .A0(n1821), .A1(n1762), .B0(n1769), .B1(
        \destinationAddressbuffer[3][1] ), .Y(n1768) );
  AOI22X1TS U1855 ( .A0(n1780), .A1(n1764), .B0(n1763), .B1(
        destinationAddressIn_EAST[1]), .Y(n1767) );
  AOI22X1TS U1856 ( .A0(n1782), .A1(n1825), .B0(n1765), .B1(n1824), .Y(n1766)
         );
  AOI22X1TS U1857 ( .A0(n1832), .A1(n126), .B0(n1769), .B1(
        \destinationAddressbuffer[3][2] ), .Y(n1775) );
  AOI22X1TS U1858 ( .A0(n955), .A1(n1771), .B0(n1770), .B1(
        destinationAddressIn_EAST[2]), .Y(n1774) );
  AOI22X1TS U1859 ( .A0(n957), .A1(n1837), .B0(n1772), .B1(n1835), .Y(n1773)
         );
  AOI22X1TS U1860 ( .A0(n1843), .A1(n1777), .B0(n1776), .B1(
        \destinationAddressbuffer[3][3] ), .Y(n1785) );
  AOI22X1TS U1861 ( .A0(n1780), .A1(n1779), .B0(n1778), .B1(
        destinationAddressIn_EAST[3]), .Y(n1784) );
  AOI22X1TS U1862 ( .A0(n1782), .A1(n1847), .B0(n1781), .B1(n1846), .Y(n1783)
         );
  AOI22X1TS U1863 ( .A0(n1811), .A1(n1786), .B0(n1798), .B1(
        \destinationAddressbuffer[2][0] ), .Y(n1791) );
  AOI22X1TS U1864 ( .A0(n1787), .A1(destinationAddressIn_WEST[0]), .B0(n991), 
        .B1(n1812), .Y(n1790) );
  AOI22X1TS U1865 ( .A0(n1788), .A1(n1815), .B0(n180), .B1(n1814), .Y(n1789)
         );
  AOI22X1TS U1866 ( .A0(n1863), .A1(n1792), .B0(n1798), .B1(
        \destinationAddressbuffer[2][1] ), .Y(n1797) );
  AOI22X1TS U1867 ( .A0(n198), .A1(destinationAddressIn_WEST[1]), .B0(n1793), 
        .B1(n1822), .Y(n1796) );
  AOI22X1TS U1868 ( .A0(n1794), .A1(n1825), .B0(n1801), .B1(n1824), .Y(n1795)
         );
  AOI22X1TS U1869 ( .A0(n1872), .A1(n1799), .B0(n1798), .B1(
        \destinationAddressbuffer[2][2] ), .Y(n1804) );
  AOI22X1TS U1870 ( .A0(n1806), .A1(destinationAddressIn_WEST[2]), .B0(n1800), 
        .B1(n1833), .Y(n1803) );
  AOI22X1TS U1871 ( .A0(n1807), .A1(n1837), .B0(n1801), .B1(n1835), .Y(n1802)
         );
  AOI22X1TS U1872 ( .A0(n1882), .A1(n175), .B0(n1805), .B1(
        \destinationAddressbuffer[2][3] ), .Y(n1810) );
  AOI22X1TS U1873 ( .A0(n1806), .A1(destinationAddressIn_WEST[3]), .B0(n174), 
        .B1(n1844), .Y(n1809) );
  AOI22X1TS U1874 ( .A0(n1807), .A1(n1847), .B0(n180), .B1(n1846), .Y(n1808)
         );
  AOI22X1TS U1875 ( .A0(n1811), .A1(n1820), .B0(n1830), .B1(
        \destinationAddressbuffer[1][0] ), .Y(n1819) );
  AOI22X1TS U1876 ( .A0(n1813), .A1(destinationAddressIn_WEST[0]), .B0(n1018), 
        .B1(n1812), .Y(n1818) );
  AOI22X1TS U1877 ( .A0(n1816), .A1(n1815), .B0(n316), .B1(n1814), .Y(n1817)
         );
  AOI22X1TS U1878 ( .A0(n1821), .A1(n1820), .B0(n1830), .B1(
        \destinationAddressbuffer[1][1] ), .Y(n1829) );
  AOI22X1TS U1879 ( .A0(n362), .A1(destinationAddressIn_WEST[1]), .B0(n1823), 
        .B1(n1822), .Y(n1828) );
  AOI22X1TS U1880 ( .A0(n1826), .A1(n1825), .B0(n1836), .B1(n1824), .Y(n1827)
         );
  AOI22X1TS U1881 ( .A0(n1832), .A1(n1831), .B0(n1830), .B1(
        \destinationAddressbuffer[1][2] ), .Y(n1840) );
  AOI22X1TS U1882 ( .A0(n1845), .A1(destinationAddressIn_WEST[2]), .B0(n1834), 
        .B1(n1833), .Y(n1839) );
  AOI22X1TS U1883 ( .A0(n1848), .A1(n1837), .B0(n1836), .B1(n1835), .Y(n1838)
         );
  AOI22X1TS U1884 ( .A0(n1843), .A1(n1842), .B0(n1841), .B1(
        \destinationAddressbuffer[1][3] ), .Y(n1851) );
  AOI22X1TS U1885 ( .A0(n1845), .A1(destinationAddressIn_WEST[3]), .B0(n309), 
        .B1(n1844), .Y(n1850) );
  AOI22X1TS U1886 ( .A0(n1848), .A1(n1847), .B0(n316), .B1(n1846), .Y(n1849)
         );
  AOI22X1TS U1887 ( .A0(n1853), .A1(n1852), .B0(n1870), .B1(
        \destinationAddressbuffer[0][0] ), .Y(n1861) );
  AOI22X1TS U1888 ( .A0(n1854), .A1(destinationAddressIn_WEST[0]), .B0(n1045), 
        .B1(destinationAddressIn_EAST[0]), .Y(n1860) );
  AOI22X1TS U1889 ( .A0(n1858), .A1(n1857), .B0(n1856), .B1(n1855), .Y(n1859)
         );
  AOI22X1TS U1890 ( .A0(n1863), .A1(n1862), .B0(n1870), .B1(
        \destinationAddressbuffer[0][1] ), .Y(n1869) );
  AOI22X1TS U1891 ( .A0(n429), .A1(destinationAddressIn_WEST[1]), .B0(n1864), 
        .B1(destinationAddressIn_EAST[1]), .Y(n1868) );
  AOI22X1TS U1892 ( .A0(n436), .A1(n1866), .B0(n1069), .B1(n1865), .Y(n1867)
         );
  AOI22X1TS U1893 ( .A0(n1872), .A1(n1871), .B0(n1870), .B1(
        \destinationAddressbuffer[0][2] ), .Y(n1879) );
  AOI22X1TS U1894 ( .A0(n1883), .A1(destinationAddressIn_WEST[2]), .B0(n1873), 
        .B1(destinationAddressIn_EAST[2]), .Y(n1878) );
  AOI22X1TS U1895 ( .A0(n1876), .A1(n1875), .B0(n1885), .B1(n1874), .Y(n1877)
         );
  AOI22X1TS U1896 ( .A0(n1882), .A1(n1881), .B0(n1880), .B1(
        \destinationAddressbuffer[0][3] ), .Y(n1890) );
  AOI22X1TS U1897 ( .A0(n1883), .A1(destinationAddressIn_WEST[3]), .B0(n383), 
        .B1(destinationAddressIn_EAST[3]), .Y(n1889) );
  AOI22X1TS U1898 ( .A0(n1887), .A1(n1886), .B0(n1885), .B1(n1884), .Y(n1888)
         );
endmodule


module router ( clk, reset, localRouterAddress, destinationAddressIn_NORTH, 
        requesterAddressIn_NORTH, readIn_NORTH, writeIn_NORTH, dataIn_NORTH, 
        destinationAddressOut_NORTH, requesterAddressOut_NORTH, readOut_NORTH, 
        writeOut_NORTH, dataOut_NORTH, destinationAddressIn_SOUTH, 
        requesterAddressIn_SOUTH, readIn_SOUTH, writeIn_SOUTH, dataIn_SOUTH, 
        destinationAddressOut_SOUTH, requesterAddressOut_SOUTH, readOut_SOUTH, 
        writeOut_SOUTH, dataOut_SOUTH, destinationAddressIn_EAST, 
        requesterAddressIn_EAST, readIn_EAST, writeIn_EAST, dataIn_EAST, 
        destinationAddressOut_EAST, requesterAddressOut_EAST, readOut_EAST, 
        writeOut_EAST, dataOut_EAST, destinationAddressIn_WEST, 
        requesterAddressIn_WEST, readIn_WEST, writeIn_WEST, dataIn_WEST, 
        destinationAddressOut_WEST, requesterAddressOut_WEST, readOut_WEST, 
        writeOut_WEST, dataOut_WEST, cacheDataIn_A, cacheAddressIn_A, 
        cacheDataOut_A, memWrite_A, cacheDataIn_B, cacheAddressIn_B, 
        cacheDataOut_B, memWrite_B );
  input [3:0] localRouterAddress;
  input [11:0] destinationAddressIn_NORTH;
  input [3:0] requesterAddressIn_NORTH;
  input [5:0] dataIn_NORTH;
  output [11:0] destinationAddressOut_NORTH;
  output [3:0] requesterAddressOut_NORTH;
  output [5:0] dataOut_NORTH;
  input [11:0] destinationAddressIn_SOUTH;
  input [3:0] requesterAddressIn_SOUTH;
  input [5:0] dataIn_SOUTH;
  output [11:0] destinationAddressOut_SOUTH;
  output [3:0] requesterAddressOut_SOUTH;
  output [5:0] dataOut_SOUTH;
  input [11:0] destinationAddressIn_EAST;
  input [3:0] requesterAddressIn_EAST;
  input [5:0] dataIn_EAST;
  output [11:0] destinationAddressOut_EAST;
  output [3:0] requesterAddressOut_EAST;
  output [5:0] dataOut_EAST;
  input [11:0] destinationAddressIn_WEST;
  input [3:0] requesterAddressIn_WEST;
  input [5:0] dataIn_WEST;
  output [11:0] destinationAddressOut_WEST;
  output [3:0] requesterAddressOut_WEST;
  output [5:0] dataOut_WEST;
  output [5:0] cacheDataIn_A;
  output [7:0] cacheAddressIn_A;
  input [5:0] cacheDataOut_A;
  output [5:0] cacheDataIn_B;
  output [7:0] cacheAddressIn_B;
  input [5:0] cacheDataOut_B;
  input clk, reset, readIn_NORTH, writeIn_NORTH, readIn_SOUTH, writeIn_SOUTH,
         readIn_EAST, writeIn_EAST, readIn_WEST, writeIn_WEST;
  output readOut_NORTH, writeOut_NORTH, readOut_SOUTH, writeOut_SOUTH,
         readOut_EAST, writeOut_EAST, readOut_WEST, writeOut_WEST, memWrite_A,
         memWrite_B;
  wire   readInBuffer_NORTH, writeInBuffer_NORTH, memRead_NORTH,
         memWrite_NORTH, readInBuffer_SOUTH, writeInBuffer_SOUTH,
         memRead_SOUTH, memWrite_SOUTH, readInBuffer_EAST, writeInBuffer_EAST,
         memRead_EAST, memWrite_EAST, readInBuffer_WEST, writeInBuffer_WEST,
         memRead_WEST, memWrite_WEST, readReady_NORTH, readReady_SOUTH,
         readReady_EAST, readReady_WEST, N4, N5, N6, N7, N8, N9, N10, N11, N12,
         N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26,
         N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40,
         N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54,
         N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68,
         N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82,
         N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96,
         N97, N98, N99, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, net46966, net46967, net46968,
         net46969, net46970, net46971, net46972, net46973, net46974, net46975,
         net46976, net46977, net46978, net46979, net46980, net46981, net46982,
         net46983, net46984, net46985, net46986, net46987, net46988, net46989;
  wire   [3:0] outputPortSelect_NORTH;
  wire   [3:0] outputPortSelect_SOUTH;
  wire   [3:0] outputPortSelect_EAST;
  wire   [3:0] outputPortSelect_WEST;
  wire   [11:0] destinationAddressInBuffer_NORTH;
  wire   [3:0] requesterAddressInBuffer_NORTH;
  wire   [5:0] dataInBuffer_NORTH;
  wire   [3:0] cacheRequesterAddress_NORTH;
  wire   [11:0] destinationAddressInBuffer_SOUTH;
  wire   [3:0] requesterAddressInBuffer_SOUTH;
  wire   [5:0] dataInBuffer_SOUTH;
  wire   [3:0] cacheRequesterAddress_SOUTH;
  wire   [11:0] destinationAddressInBuffer_EAST;
  wire   [3:0] requesterAddressInBuffer_EAST;
  wire   [5:0] dataInBuffer_EAST;
  wire   [3:0] cacheRequesterAddress_EAST;
  wire   [11:0] destinationAddressInBuffer_WEST;
  wire   [3:0] requesterAddressInBuffer_WEST;
  wire   [5:0] dataInBuffer_WEST;
  wire   [3:0] cacheRequesterAddress_WEST;

  cacheAccessArbiter cacheController ( .clk(clk), .reset(n682), 
        .cacheAddressIn_NORTH({n419, n418, n417, n416, n415, n413, n411, n409}), .requesterAddressIn_NORTH({n653, n649, n645, n641}), .memRead_NORTH(
        memRead_NORTH), .memWrite_NORTH(memWrite_NORTH), .dataIn_NORTH(
        dataInBuffer_NORTH), .readReady_NORTH(readReady_NORTH), 
        .requesterAddressOut_NORTH(cacheRequesterAddress_NORTH), 
        .cacheAddressIn_SOUTH({n613, n611, n609, n607, n605, n600, n595, n590}), .requesterAddressIn_SOUTH({n407, n405, n403, n401}), .memRead_SOUTH(
        memRead_SOUTH), .memWrite_SOUTH(memWrite_SOUTH), .dataIn_SOUTH({n585, 
        n580, n575, n570, n565, n560}), .readReady_SOUTH(readReady_SOUTH), 
        .requesterAddressOut_SOUTH(cacheRequesterAddress_SOUTH), 
        .cacheAddressIn_EAST({n379, n377, n375, n373, n555, n550, n545, n540}), 
        .requesterAddressIn_EAST({n535, n534, n533, n532}), .memRead_EAST(
        memRead_EAST), .memWrite_EAST(n292), .dataIn_EAST({n531, n526, n521, 
        n516, n511, n506}), .readReady_EAST(readReady_EAST), 
        .requesterAddressOut_EAST(cacheRequesterAddress_EAST), 
        .cacheAddressIn_WEST({n501, n497, n493, n489, n485, n481, n477, n473}), 
        .requesterAddressIn_WEST({n469, n464, n459, n454}), .memRead_WEST(
        memRead_WEST), .memWrite_WEST(n328), .dataIn_WEST({n449, n445, n441, 
        n437, n433, n429}), .readReady_WEST(readReady_WEST), 
        .requesterAddressOut_WEST(cacheRequesterAddress_WEST), .cacheDataIn_A(
        cacheDataIn_A), .cacheAddressIn_A(cacheAddressIn_A), .cacheDataOut_A({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .memWrite_A(memWrite_A), 
        .cacheDataIn_B(cacheDataIn_B), .cacheAddressIn_B(cacheAddressIn_B), 
        .cacheDataOut_B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .memWrite_B(
        memWrite_B) );
  outputPortArbiter_0 outNorth ( .clk(clk), .reset(n680), .selectBit_NORTH(
        n351), .destinationAddressIn_NORTH({
        destinationAddressInBuffer_NORTH[11:8], n669, n665, n661, n657, 
        destinationAddressInBuffer_NORTH[3:0]}), .requesterAddressIn_NORTH({
        n653, n649, n645, n641}), .readIn_NORTH(n422), .writeIn_NORTH(n675), 
        .dataIn_NORTH({n637, n633, n629, n625, n621, n617}), .selectBit_SOUTH(
        n265), .destinationAddressIn_SOUTH({
        destinationAddressInBuffer_SOUTH[11:8], n612, n610, n608, n606, n604, 
        n599, n594, n589}), .requesterAddressIn_SOUTH(
        requesterAddressInBuffer_SOUTH), .readIn_SOUTH(n423), .writeIn_SOUTH(
        n674), .dataIn_SOUTH({n584, n579, n574, n569, n564, n559}), 
        .selectBit_EAST(n385), .destinationAddressIn_EAST({n372, n369, n366, 
        n363, n358, n356, n354, n352, n554, n549, n544, n539}), 
        .requesterAddressIn_EAST({n399, n397, n395, n393}), .readIn_EAST(n390), 
        .writeIn_EAST(n384), .dataIn_EAST({n530, n525, n520, n515, n510, n505}), .selectBit_WEST(outputPortSelect_WEST[0]), .destinationAddressIn_WEST({
        destinationAddressInBuffer_WEST[11:8], n501, n497, n493, n489, n485, 
        n481, n477, n473}), .requesterAddressIn_WEST({n468, n463, n458, n453}), 
        .readIn_WEST(n425), .writeIn_WEST(n670), .dataIn_WEST({n449, n445, 
        n441, n437, n433, n429}), .readReady(readReady_NORTH), 
        .readRequesterAddress(cacheRequesterAddress_NORTH), .cacheDataOut({
        net46984, net46985, net46986, net46987, net46988, net46989}), 
        .destinationAddressOut(destinationAddressOut_NORTH), 
        .requesterAddressOut(requesterAddressOut_NORTH), .readOut(
        readOut_NORTH), .writeOut(writeOut_NORTH), .dataOut(dataOut_NORTH) );
  outputPortArbiter_3 outSouth ( .clk(clk), .reset(n681), .selectBit_NORTH(
        n349), .destinationAddressIn_NORTH({
        destinationAddressInBuffer_NORTH[11:8], n666, n662, n658, n654, n414, 
        n412, n410, n408}), .requesterAddressIn_NORTH({n650, n646, n642, n638}), .readIn_NORTH(n677), .writeIn_NORTH(n421), .dataIn_NORTH({n634, n630, n626, 
        n622, n618, n614}), .selectBit_SOUTH(n270), 
        .destinationAddressIn_SOUTH({destinationAddressInBuffer_SOUTH[11:8], 
        n612, n610, n608, n606, n601, n596, n591, n586}), 
        .requesterAddressIn_SOUTH({n406, n404, n402, n400}), .readIn_SOUTH(
        n420), .writeIn_SOUTH(n674), .dataIn_SOUTH({n581, n576, n571, n566, 
        n561, n556}), .selectBit_EAST(n386), .destinationAddressIn_EAST({
        destinationAddressInBuffer_EAST[11:4], n551, n546, n541, n536}), 
        .requesterAddressIn_EAST({n398, n396, n394, n392}), .readIn_EAST(n389), 
        .writeIn_EAST(n382), .dataIn_EAST({n527, n522, n517, n512, n507, n502}), .selectBit_WEST(outputPortSelect_WEST[1]), .destinationAddressIn_WEST({
        destinationAddressInBuffer_WEST[11:8], n498, n494, n490, n486, n482, 
        n478, n474, n470}), .requesterAddressIn_WEST({n465, n460, n455, n450}), 
        .readIn_WEST(n672), .writeIn_WEST(n424), .dataIn_WEST({n446, n442, 
        n438, n434, n430, n426}), .readReady(readReady_SOUTH), 
        .readRequesterAddress(cacheRequesterAddress_SOUTH), .cacheDataOut({
        net46978, net46979, net46980, net46981, net46982, net46983}), 
        .destinationAddressOut(destinationAddressOut_SOUTH), 
        .requesterAddressOut(requesterAddressOut_SOUTH), .readOut(
        readOut_SOUTH), .writeOut(writeOut_SOUTH), .dataOut(dataOut_SOUTH) );
  outputPortArbiter_2 outEast ( .clk(clk), .reset(n682), .selectBit_NORTH(n348), .destinationAddressIn_NORTH({destinationAddressInBuffer_NORTH[11:8], n667, 
        n663, n659, n655, n414, n412, n410, n408}), .requesterAddressIn_NORTH(
        {n651, n647, n643, n639}), .readIn_NORTH(n678), .writeIn_NORTH(n421), 
        .dataIn_NORTH({n635, n631, n627, n623, n619, n615}), .selectBit_SOUTH(
        n360), .destinationAddressIn_SOUTH({
        destinationAddressInBuffer_SOUTH[11:8], n612, n610, n608, n606, n602, 
        n597, n592, n587}), .requesterAddressIn_SOUTH({n406, n404, n402, n400}), .readIn_SOUTH(n420), .writeIn_SOUTH(n674), .dataIn_SOUTH({n582, n577, n572, 
        n567, n562, n557}), .selectBit_EAST(n387), .destinationAddressIn_EAST(
        {n370, n367, n364, n361, n359, n357, n355, n353, n552, n547, n542, 
        n537}), .requesterAddressIn_EAST(requesterAddressInBuffer_EAST), 
        .readIn_EAST(n391), .writeIn_EAST(n381), .dataIn_EAST({n528, n523, 
        n518, n513, n508, n503}), .selectBit_WEST(outputPortSelect_WEST[2]), 
        .destinationAddressIn_WEST({destinationAddressInBuffer_WEST[11:8], 
        n499, n495, n491, n487, n483, n479, n475, n471}), 
        .requesterAddressIn_WEST({n466, n461, n456, n451}), .readIn_WEST(n673), 
        .writeIn_WEST(n424), .dataIn_WEST({n447, n443, n439, n435, n431, n427}), .readReady(readReady_EAST), .readRequesterAddress(cacheRequesterAddress_EAST), .cacheDataOut({net46972, net46973, net46974, net46975, net46976, net46977}), 
        .destinationAddressOut(destinationAddressOut_EAST), 
        .requesterAddressOut(requesterAddressOut_EAST), .readOut(readOut_EAST), 
        .writeOut(writeOut_EAST), .dataOut(dataOut_EAST) );
  outputPortArbiter_1 outWest ( .clk(clk), .reset(n679), .selectBit_NORTH(n350), .destinationAddressIn_NORTH({destinationAddressInBuffer_NORTH[11:8], n668, 
        n664, n660, n656, destinationAddressInBuffer_NORTH[3:0]}), 
        .requesterAddressIn_NORTH({n652, n648, n644, n640}), .readIn_NORTH(
        n422), .writeIn_NORTH(n676), .dataIn_NORTH({n636, n632, n628, n624, 
        n620, n616}), .selectBit_SOUTH(n281), .destinationAddressIn_SOUTH({
        destinationAddressInBuffer_SOUTH[11:8], n612, n610, n608, n606, n603, 
        n598, n593, n588}), .requesterAddressIn_SOUTH(
        requesterAddressInBuffer_SOUTH), .readIn_SOUTH(n423), .writeIn_SOUTH(
        n674), .dataIn_SOUTH({n583, n578, n573, n568, n563, n558}), 
        .selectBit_EAST(n388), .destinationAddressIn_EAST({n371, n368, n365, 
        n362, n380, n378, n376, n374, n553, n548, n543, n538}), 
        .requesterAddressIn_EAST(requesterAddressInBuffer_EAST), .readIn_EAST(
        n389), .writeIn_EAST(n383), .dataIn_EAST({n529, n524, n519, n514, n509, 
        n504}), .selectBit_WEST(outputPortSelect_WEST[3]), 
        .destinationAddressIn_WEST({destinationAddressInBuffer_WEST[11:8], 
        n500, n496, n492, n488, n484, n480, n476, n472}), 
        .requesterAddressIn_WEST({n467, n462, n457, n452}), .readIn_WEST(n425), 
        .writeIn_WEST(n671), .dataIn_WEST({n448, n444, n440, n436, n432, n428}), .readReady(readReady_WEST), .readRequesterAddress(cacheRequesterAddress_WEST), .cacheDataOut({net46966, net46967, net46968, net46969, net46970, net46971}), 
        .destinationAddressOut(destinationAddressOut_WEST), 
        .requesterAddressOut(requesterAddressOut_WEST), .readOut(readOut_WEST), 
        .writeOut(writeOut_WEST), .dataOut(dataOut_WEST) );
  DFFQX1TS writeInBuffer_SOUTH_reg ( .D(N45), .CK(clk), .Q(writeInBuffer_SOUTH) );
  DFFQX1TS \dataInBuffer_SOUTH_reg[5]  ( .D(N51), .CK(clk), .Q(
        dataInBuffer_SOUTH[5]) );
  DFFQX1TS \dataInBuffer_SOUTH_reg[4]  ( .D(N50), .CK(clk), .Q(
        dataInBuffer_SOUTH[4]) );
  DFFQX1TS \dataInBuffer_SOUTH_reg[3]  ( .D(N49), .CK(clk), .Q(
        dataInBuffer_SOUTH[3]) );
  DFFQX1TS \dataInBuffer_SOUTH_reg[2]  ( .D(N48), .CK(clk), .Q(
        dataInBuffer_SOUTH[2]) );
  DFFQX1TS \dataInBuffer_SOUTH_reg[1]  ( .D(N47), .CK(clk), .Q(
        dataInBuffer_SOUTH[1]) );
  DFFQX1TS \dataInBuffer_SOUTH_reg[0]  ( .D(N46), .CK(clk), .Q(
        dataInBuffer_SOUTH[0]) );
  DFFQX1TS \requesterAddressInBuffer_WEST_reg[3]  ( .D(N91), .CK(clk), .Q(
        requesterAddressInBuffer_WEST[3]) );
  DFFQX1TS \requesterAddressInBuffer_WEST_reg[2]  ( .D(N90), .CK(clk), .Q(
        requesterAddressInBuffer_WEST[2]) );
  DFFQX1TS \requesterAddressInBuffer_WEST_reg[1]  ( .D(N89), .CK(clk), .Q(
        requesterAddressInBuffer_WEST[1]) );
  DFFQX1TS \requesterAddressInBuffer_WEST_reg[0]  ( .D(N88), .CK(clk), .Q(
        requesterAddressInBuffer_WEST[0]) );
  DFFQX1TS \destinationAddressInBuffer_SOUTH_reg[3]  ( .D(N31), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[3]) );
  DFFQX1TS \destinationAddressInBuffer_EAST_reg[3]  ( .D(N55), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[3]) );
  DFFQX1TS \destinationAddressInBuffer_SOUTH_reg[2]  ( .D(N30), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[2]) );
  DFFQX1TS \destinationAddressInBuffer_EAST_reg[2]  ( .D(N54), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[2]) );
  DFFQX1TS \destinationAddressInBuffer_SOUTH_reg[1]  ( .D(N29), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[1]) );
  DFFQX1TS \destinationAddressInBuffer_EAST_reg[1]  ( .D(N53), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[1]) );
  DFFQX1TS \destinationAddressInBuffer_SOUTH_reg[0]  ( .D(N28), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[0]) );
  DFFQX1TS \destinationAddressInBuffer_EAST_reg[0]  ( .D(N52), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[0]) );
  DFFQX1TS \dataInBuffer_NORTH_reg[5]  ( .D(N27), .CK(clk), .Q(
        dataInBuffer_NORTH[5]) );
  DFFQX1TS \dataInBuffer_EAST_reg[5]  ( .D(N75), .CK(clk), .Q(
        dataInBuffer_EAST[5]) );
  DFFQX1TS \dataInBuffer_NORTH_reg[4]  ( .D(N26), .CK(clk), .Q(
        dataInBuffer_NORTH[4]) );
  DFFQX1TS \dataInBuffer_EAST_reg[4]  ( .D(N74), .CK(clk), .Q(
        dataInBuffer_EAST[4]) );
  DFFQX1TS \dataInBuffer_NORTH_reg[3]  ( .D(N25), .CK(clk), .Q(
        dataInBuffer_NORTH[3]) );
  DFFQX1TS \dataInBuffer_EAST_reg[3]  ( .D(N73), .CK(clk), .Q(
        dataInBuffer_EAST[3]) );
  DFFQX1TS \dataInBuffer_NORTH_reg[2]  ( .D(N24), .CK(clk), .Q(
        dataInBuffer_NORTH[2]) );
  DFFQX1TS \dataInBuffer_EAST_reg[2]  ( .D(N72), .CK(clk), .Q(
        dataInBuffer_EAST[2]) );
  DFFQX1TS \dataInBuffer_NORTH_reg[1]  ( .D(N23), .CK(clk), .Q(
        dataInBuffer_NORTH[1]) );
  DFFQX1TS \dataInBuffer_EAST_reg[1]  ( .D(N71), .CK(clk), .Q(
        dataInBuffer_EAST[1]) );
  DFFQX1TS \dataInBuffer_NORTH_reg[0]  ( .D(N22), .CK(clk), .Q(
        dataInBuffer_NORTH[0]) );
  DFFQX1TS \dataInBuffer_EAST_reg[0]  ( .D(N70), .CK(clk), .Q(
        dataInBuffer_EAST[0]) );
  DFFQX1TS \destinationAddressInBuffer_NORTH_reg[7]  ( .D(N11), .CK(clk), .Q(
        destinationAddressInBuffer_NORTH[7]) );
  DFFQX1TS \destinationAddressInBuffer_NORTH_reg[6]  ( .D(N10), .CK(clk), .Q(
        destinationAddressInBuffer_NORTH[6]) );
  DFFQX1TS \destinationAddressInBuffer_NORTH_reg[5]  ( .D(N9), .CK(clk), .Q(
        destinationAddressInBuffer_NORTH[5]) );
  DFFQX1TS \destinationAddressInBuffer_NORTH_reg[4]  ( .D(N8), .CK(clk), .Q(
        destinationAddressInBuffer_NORTH[4]) );
  DFFQX1TS writeInBuffer_NORTH_reg ( .D(N21), .CK(clk), .Q(writeInBuffer_NORTH) );
  DFFQX1TS writeInBuffer_WEST_reg ( .D(N93), .CK(clk), .Q(writeInBuffer_WEST)
         );
  DFFQX1TS readInBuffer_WEST_reg ( .D(N92), .CK(clk), .Q(readInBuffer_WEST) );
  DFFQX1TS readInBuffer_NORTH_reg ( .D(N20), .CK(clk), .Q(readInBuffer_NORTH)
         );
  DFFQX1TS \destinationAddressInBuffer_WEST_reg[11]  ( .D(N87), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[11]) );
  DFFQX1TS \destinationAddressInBuffer_WEST_reg[10]  ( .D(N86), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[10]) );
  DFFQX1TS \destinationAddressInBuffer_WEST_reg[9]  ( .D(N85), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[9]) );
  DFFQX1TS \destinationAddressInBuffer_WEST_reg[8]  ( .D(N84), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[8]) );
  DFFQX1TS readInBuffer_EAST_reg ( .D(N68), .CK(clk), .Q(readInBuffer_EAST) );
  DFFQX1TS \destinationAddressInBuffer_EAST_reg[11]  ( .D(N63), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[11]) );
  DFFQX1TS \destinationAddressInBuffer_EAST_reg[10]  ( .D(N62), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[10]) );
  DFFQX1TS \destinationAddressInBuffer_EAST_reg[9]  ( .D(N61), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[9]) );
  DFFQX1TS \destinationAddressInBuffer_EAST_reg[8]  ( .D(N60), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[8]) );
  DFFQX1TS \destinationAddressInBuffer_SOUTH_reg[7]  ( .D(N35), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[7]) );
  DFFQX1TS \destinationAddressInBuffer_SOUTH_reg[6]  ( .D(N34), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[6]) );
  DFFQX1TS \destinationAddressInBuffer_SOUTH_reg[5]  ( .D(N33), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[5]) );
  DFFQX1TS \destinationAddressInBuffer_SOUTH_reg[4]  ( .D(N32), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[4]) );
  DFFQX1TS writeInBuffer_EAST_reg ( .D(N69), .CK(clk), .Q(writeInBuffer_EAST)
         );
  DFFQX1TS \destinationAddressInBuffer_EAST_reg[7]  ( .D(N59), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[7]) );
  DFFQX1TS \destinationAddressInBuffer_EAST_reg[6]  ( .D(N58), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[6]) );
  DFFQX1TS \destinationAddressInBuffer_EAST_reg[5]  ( .D(N57), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[5]) );
  DFFQX1TS \destinationAddressInBuffer_EAST_reg[4]  ( .D(N56), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[4]) );
  DFFQX1TS \destinationAddressInBuffer_SOUTH_reg[11]  ( .D(N39), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[11]) );
  DFFQX1TS \destinationAddressInBuffer_SOUTH_reg[10]  ( .D(N38), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[10]) );
  DFFQX1TS \destinationAddressInBuffer_SOUTH_reg[9]  ( .D(N37), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[9]) );
  DFFQX1TS \destinationAddressInBuffer_SOUTH_reg[8]  ( .D(N36), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[8]) );
  DFFQX1TS \destinationAddressInBuffer_NORTH_reg[11]  ( .D(N15), .CK(clk), .Q(
        destinationAddressInBuffer_NORTH[11]) );
  DFFQX1TS \destinationAddressInBuffer_NORTH_reg[10]  ( .D(N14), .CK(clk), .Q(
        destinationAddressInBuffer_NORTH[10]) );
  DFFQX1TS \destinationAddressInBuffer_NORTH_reg[9]  ( .D(N13), .CK(clk), .Q(
        destinationAddressInBuffer_NORTH[9]) );
  DFFQX1TS \destinationAddressInBuffer_NORTH_reg[8]  ( .D(N12), .CK(clk), .Q(
        destinationAddressInBuffer_NORTH[8]) );
  DFFQX1TS \destinationAddressInBuffer_NORTH_reg[3]  ( .D(N7), .CK(clk), .Q(
        destinationAddressInBuffer_NORTH[3]) );
  DFFQX1TS \destinationAddressInBuffer_NORTH_reg[2]  ( .D(N6), .CK(clk), .Q(
        destinationAddressInBuffer_NORTH[2]) );
  DFFQX1TS \destinationAddressInBuffer_NORTH_reg[1]  ( .D(N5), .CK(clk), .Q(
        destinationAddressInBuffer_NORTH[1]) );
  DFFQX1TS \destinationAddressInBuffer_NORTH_reg[0]  ( .D(N4), .CK(clk), .Q(
        destinationAddressInBuffer_NORTH[0]) );
  DFFQX1TS \requesterAddressInBuffer_SOUTH_reg[3]  ( .D(N43), .CK(clk), .Q(
        requesterAddressInBuffer_SOUTH[3]) );
  DFFQX1TS \requesterAddressInBuffer_SOUTH_reg[2]  ( .D(N42), .CK(clk), .Q(
        requesterAddressInBuffer_SOUTH[2]) );
  DFFQX1TS \requesterAddressInBuffer_SOUTH_reg[1]  ( .D(N41), .CK(clk), .Q(
        requesterAddressInBuffer_SOUTH[1]) );
  DFFQX1TS \requesterAddressInBuffer_SOUTH_reg[0]  ( .D(N40), .CK(clk), .Q(
        requesterAddressInBuffer_SOUTH[0]) );
  DFFQX1TS \requesterAddressInBuffer_EAST_reg[3]  ( .D(N67), .CK(clk), .Q(
        requesterAddressInBuffer_EAST[3]) );
  DFFQX1TS \requesterAddressInBuffer_EAST_reg[2]  ( .D(N66), .CK(clk), .Q(
        requesterAddressInBuffer_EAST[2]) );
  DFFQX1TS \requesterAddressInBuffer_EAST_reg[1]  ( .D(N65), .CK(clk), .Q(
        requesterAddressInBuffer_EAST[1]) );
  DFFQX1TS \requesterAddressInBuffer_EAST_reg[0]  ( .D(N64), .CK(clk), .Q(
        requesterAddressInBuffer_EAST[0]) );
  DFFQX1TS readInBuffer_SOUTH_reg ( .D(N44), .CK(clk), .Q(readInBuffer_SOUTH)
         );
  DFFQX1TS \dataInBuffer_WEST_reg[5]  ( .D(N99), .CK(clk), .Q(
        dataInBuffer_WEST[5]) );
  DFFQX1TS \dataInBuffer_WEST_reg[4]  ( .D(N98), .CK(clk), .Q(
        dataInBuffer_WEST[4]) );
  DFFQX1TS \dataInBuffer_WEST_reg[3]  ( .D(N97), .CK(clk), .Q(
        dataInBuffer_WEST[3]) );
  DFFQX1TS \dataInBuffer_WEST_reg[2]  ( .D(N96), .CK(clk), .Q(
        dataInBuffer_WEST[2]) );
  DFFQX1TS \dataInBuffer_WEST_reg[1]  ( .D(N95), .CK(clk), .Q(
        dataInBuffer_WEST[1]) );
  DFFQX1TS \dataInBuffer_WEST_reg[0]  ( .D(N94), .CK(clk), .Q(
        dataInBuffer_WEST[0]) );
  DFFQX1TS \destinationAddressInBuffer_WEST_reg[3]  ( .D(N79), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[3]) );
  DFFQX1TS \destinationAddressInBuffer_WEST_reg[2]  ( .D(N78), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[2]) );
  DFFQX1TS \destinationAddressInBuffer_WEST_reg[1]  ( .D(N77), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[1]) );
  DFFQX1TS \destinationAddressInBuffer_WEST_reg[0]  ( .D(N76), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[0]) );
  DFFQX1TS \requesterAddressInBuffer_NORTH_reg[3]  ( .D(N19), .CK(clk), .Q(
        requesterAddressInBuffer_NORTH[3]) );
  DFFQX1TS \requesterAddressInBuffer_NORTH_reg[2]  ( .D(N18), .CK(clk), .Q(
        requesterAddressInBuffer_NORTH[2]) );
  DFFQX1TS \requesterAddressInBuffer_NORTH_reg[1]  ( .D(N17), .CK(clk), .Q(
        requesterAddressInBuffer_NORTH[1]) );
  DFFQX1TS \requesterAddressInBuffer_NORTH_reg[0]  ( .D(N16), .CK(clk), .Q(
        requesterAddressInBuffer_NORTH[0]) );
  DFFQX1TS \destinationAddressInBuffer_WEST_reg[7]  ( .D(N83), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[7]) );
  DFFQX1TS \destinationAddressInBuffer_WEST_reg[6]  ( .D(N82), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[6]) );
  DFFQX1TS \destinationAddressInBuffer_WEST_reg[5]  ( .D(N81), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[5]) );
  DFFQX1TS \destinationAddressInBuffer_WEST_reg[4]  ( .D(N80), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[4]) );
  DFFQX1TS \inWest/memRead_reg  ( .D(n73), .CK(clk), .Q(memRead_WEST) );
  DFFQX1TS \inEast/memRead_reg  ( .D(n79), .CK(clk), .Q(memRead_EAST) );
  DFFQX1TS \inNorth/memWrite_reg  ( .D(n96), .CK(clk), .Q(memWrite_NORTH) );
  DFFQX1TS \inWest/memWrite_reg  ( .D(n78), .CK(clk), .Q(memWrite_WEST) );
  DFFQX1TS \inNorth/memRead_reg  ( .D(n91), .CK(clk), .Q(memRead_NORTH) );
  DFFQX1TS \inEast/memWrite_reg  ( .D(n84), .CK(clk), .Q(memWrite_EAST) );
  DFFQX1TS \inSouth/memRead_reg  ( .D(n85), .CK(clk), .Q(memRead_SOUTH) );
  DFFQX1TS \inSouth/memWrite_reg  ( .D(n90), .CK(clk), .Q(memWrite_SOUTH) );
  DFFHQX1TS \inNorth/outputPortSelect_reg[0]  ( .D(n95), .CK(clk), .Q(
        outputPortSelect_NORTH[0]) );
  DFFHQX1TS \inNorth/outputPortSelect_reg[3]  ( .D(n92), .CK(clk), .Q(
        outputPortSelect_NORTH[3]) );
  DFFHQX1TS \inNorth/outputPortSelect_reg[1]  ( .D(n94), .CK(clk), .Q(
        outputPortSelect_NORTH[1]) );
  DFFHQX1TS \inNorth/outputPortSelect_reg[2]  ( .D(n93), .CK(clk), .Q(
        outputPortSelect_NORTH[2]) );
  DFFHQX1TS \inSouth/outputPortSelect_reg[0]  ( .D(n89), .CK(clk), .Q(
        outputPortSelect_SOUTH[0]) );
  DFFHQX1TS \inSouth/outputPortSelect_reg[3]  ( .D(n86), .CK(clk), .Q(
        outputPortSelect_SOUTH[3]) );
  DFFHQX1TS \inSouth/outputPortSelect_reg[1]  ( .D(n88), .CK(clk), .Q(
        outputPortSelect_SOUTH[1]) );
  DFFHQX1TS \inSouth/outputPortSelect_reg[2]  ( .D(n87), .CK(clk), .Q(
        outputPortSelect_SOUTH[2]) );
  DFFQX1TS \inEast/outputPortSelect_reg[1]  ( .D(n82), .CK(clk), .Q(
        outputPortSelect_EAST[1]) );
  DFFHQX1TS \inEast/outputPortSelect_reg[2]  ( .D(n81), .CK(clk), .Q(
        outputPortSelect_EAST[2]) );
  DFFQX1TS \inWest/outputPortSelect_reg[2]  ( .D(n75), .CK(clk), .Q(
        outputPortSelect_WEST[2]) );
  DFFQX1TS \inWest/outputPortSelect_reg[3]  ( .D(n74), .CK(clk), .Q(
        outputPortSelect_WEST[3]) );
  DFFQX1TS \inWest/outputPortSelect_reg[0]  ( .D(n77), .CK(clk), .Q(
        outputPortSelect_WEST[0]) );
  DFFQX1TS \inWest/outputPortSelect_reg[1]  ( .D(n76), .CK(clk), .Q(
        outputPortSelect_WEST[1]) );
  DFFQX1TS \inEast/outputPortSelect_reg[3]  ( .D(n80), .CK(clk), .Q(
        outputPortSelect_EAST[3]) );
  DFFQX1TS \inEast/outputPortSelect_reg[0]  ( .D(n83), .CK(clk), .Q(
        outputPortSelect_EAST[0]) );
  CLKBUFX2TS U258 ( .A(memWrite_WEST), .Y(n328) );
  CLKBUFX2TS U259 ( .A(memWrite_EAST), .Y(n292) );
  CLKBUFX2TS U260 ( .A(outputPortSelect_SOUTH[3]), .Y(n281) );
  CLKBUFX2TS U261 ( .A(outputPortSelect_SOUTH[0]), .Y(n265) );
  CLKBUFX2TS U262 ( .A(outputPortSelect_SOUTH[1]), .Y(n270) );
  INVX2TS U263 ( .A(n236), .Y(n326) );
  INVX2TS U264 ( .A(n236), .Y(n290) );
  INVX2TS U265 ( .A(n236), .Y(n680) );
  AO22XLTS U266 ( .A0(writeInBuffer_SOUTH), .A1(n285), .B0(n284), .B1(
        memWrite_SOUTH), .Y(n90) );
  CLKBUFX2TS U267 ( .A(n327), .Y(n330) );
  CLKBUFX2TS U268 ( .A(n291), .Y(n296) );
  CLKBUFX2TS U269 ( .A(n237), .Y(n241) );
  CLKBUFX2TS U270 ( .A(n212), .Y(n260) );
  CLKBUFX2TS U271 ( .A(n201), .Y(n286) );
  CLKBUFX2TS U272 ( .A(n190), .Y(n315) );
  CLKBUFX2TS U273 ( .A(n224), .Y(n230) );
  INVX2TS U274 ( .A(n310), .Y(n388) );
  INVX2TS U275 ( .A(n158), .Y(n194) );
  AO22XLTS U276 ( .A0(n345), .A1(n344), .B0(n327), .B1(
        outputPortSelect_WEST[2]), .Y(n75) );
  AO22XLTS U277 ( .A0(readInBuffer_SOUTH), .A1(n285), .B0(n284), .B1(
        memRead_SOUTH), .Y(n85) );
  AO22XLTS U278 ( .A0(n382), .A1(n313), .B0(n296), .B1(memWrite_EAST), .Y(n84)
         );
  AO22XLTS U279 ( .A0(readInBuffer_NORTH), .A1(n259), .B0(n237), .B1(
        memRead_NORTH), .Y(n91) );
  AO22XLTS U280 ( .A0(writeInBuffer_NORTH), .A1(n259), .B0(n241), .B1(
        memWrite_NORTH), .Y(n96) );
  AO22XLTS U281 ( .A0(n390), .A1(n313), .B0(n296), .B1(memRead_EAST), .Y(n79)
         );
  INVX2TS U282 ( .A(n231), .Y(n232) );
  INVX2TS U283 ( .A(outputPortSelect_EAST[3]), .Y(n310) );
  INVX2TS U284 ( .A(outputPortSelect_NORTH[2]), .Y(n254) );
  INVX2TS U285 ( .A(n187), .Y(n188) );
  INVX2TS U286 ( .A(n254), .Y(n348) );
  INVX2TS U287 ( .A(outputPortSelect_NORTH[1]), .Y(n246) );
  INVX2TS U288 ( .A(n246), .Y(n349) );
  INVX2TS U289 ( .A(outputPortSelect_NORTH[3]), .Y(n256) );
  INVX2TS U290 ( .A(n256), .Y(n350) );
  INVX2TS U291 ( .A(outputPortSelect_NORTH[0]), .Y(n240) );
  INVX2TS U292 ( .A(n240), .Y(n351) );
  INVX2TS U293 ( .A(destinationAddressInBuffer_EAST[4]), .Y(n152) );
  INVX2TS U294 ( .A(n152), .Y(n352) );
  INVX2TS U295 ( .A(n152), .Y(n353) );
  INVX2TS U296 ( .A(destinationAddressInBuffer_EAST[5]), .Y(n153) );
  INVX2TS U297 ( .A(n153), .Y(n354) );
  INVX2TS U298 ( .A(n153), .Y(n355) );
  INVX2TS U299 ( .A(destinationAddressInBuffer_EAST[6]), .Y(n154) );
  INVX2TS U300 ( .A(n154), .Y(n356) );
  INVX2TS U301 ( .A(n154), .Y(n357) );
  INVX2TS U302 ( .A(destinationAddressInBuffer_EAST[7]), .Y(n155) );
  INVX2TS U303 ( .A(n155), .Y(n358) );
  INVX2TS U304 ( .A(n155), .Y(n359) );
  INVX2TS U305 ( .A(outputPortSelect_SOUTH[2]), .Y(n278) );
  INVX2TS U306 ( .A(n278), .Y(n360) );
  INVX2TS U307 ( .A(destinationAddressInBuffer_EAST[8]), .Y(n148) );
  INVX2TS U308 ( .A(n148), .Y(n361) );
  INVX2TS U309 ( .A(n148), .Y(n362) );
  INVX2TS U310 ( .A(n148), .Y(n363) );
  INVX2TS U311 ( .A(destinationAddressInBuffer_EAST[9]), .Y(n149) );
  INVX2TS U312 ( .A(n149), .Y(n364) );
  INVX2TS U313 ( .A(n149), .Y(n365) );
  INVX2TS U314 ( .A(n149), .Y(n366) );
  INVX2TS U315 ( .A(destinationAddressInBuffer_EAST[10]), .Y(n150) );
  INVX2TS U316 ( .A(n150), .Y(n367) );
  INVX2TS U317 ( .A(n150), .Y(n368) );
  INVX2TS U318 ( .A(n150), .Y(n369) );
  INVX2TS U319 ( .A(destinationAddressInBuffer_EAST[11]), .Y(n151) );
  INVX2TS U320 ( .A(n151), .Y(n370) );
  INVX2TS U321 ( .A(n151), .Y(n371) );
  INVX2TS U322 ( .A(n151), .Y(n372) );
  INVX2TS U323 ( .A(n152), .Y(n373) );
  INVX2TS U324 ( .A(n152), .Y(n374) );
  INVX2TS U325 ( .A(n153), .Y(n375) );
  INVX2TS U326 ( .A(n153), .Y(n376) );
  INVX2TS U327 ( .A(n154), .Y(n377) );
  INVX2TS U328 ( .A(n154), .Y(n378) );
  INVX2TS U329 ( .A(n155), .Y(n379) );
  INVX2TS U330 ( .A(n155), .Y(n380) );
  INVX2TS U331 ( .A(writeInBuffer_EAST), .Y(n156) );
  INVX2TS U332 ( .A(n156), .Y(n381) );
  INVX2TS U333 ( .A(n156), .Y(n382) );
  INVX2TS U334 ( .A(n156), .Y(n383) );
  INVX2TS U335 ( .A(n156), .Y(n384) );
  INVX2TS U336 ( .A(outputPortSelect_EAST[0]), .Y(n295) );
  INVX2TS U337 ( .A(n295), .Y(n385) );
  INVX2TS U338 ( .A(outputPortSelect_EAST[1]), .Y(n300) );
  INVX2TS U339 ( .A(n300), .Y(n386) );
  CLKBUFX2TS U340 ( .A(outputPortSelect_EAST[2]), .Y(n387) );
  INVX2TS U341 ( .A(readInBuffer_EAST), .Y(n157) );
  INVX2TS U342 ( .A(n157), .Y(n389) );
  INVX2TS U343 ( .A(n157), .Y(n390) );
  INVX2TS U344 ( .A(n157), .Y(n391) );
  CLKBUFX2TS U345 ( .A(reset), .Y(n158) );
  CLKBUFX2TS U346 ( .A(n194), .Y(n220) );
  CLKBUFX2TS U347 ( .A(n220), .Y(n236) );
  INVX2TS U348 ( .A(n236), .Y(n682) );
  CLKBUFX2TS U349 ( .A(writeInBuffer_SOUTH), .Y(n674) );
  CLKBUFX2TS U350 ( .A(destinationAddressInBuffer_SOUTH[7]), .Y(n612) );
  CLKBUFX2TS U351 ( .A(destinationAddressInBuffer_SOUTH[6]), .Y(n610) );
  CLKBUFX2TS U352 ( .A(destinationAddressInBuffer_SOUTH[5]), .Y(n608) );
  CLKBUFX2TS U353 ( .A(destinationAddressInBuffer_SOUTH[4]), .Y(n606) );
  CLKBUFX2TS U354 ( .A(readInBuffer_SOUTH), .Y(n423) );
  CLKBUFX2TS U355 ( .A(dataInBuffer_SOUTH[5]), .Y(n584) );
  CLKBUFX2TS U356 ( .A(n584), .Y(n582) );
  CLKBUFX2TS U357 ( .A(dataInBuffer_SOUTH[4]), .Y(n579) );
  CLKBUFX2TS U358 ( .A(n579), .Y(n577) );
  CLKBUFX2TS U359 ( .A(requesterAddressInBuffer_WEST[2]), .Y(n176) );
  CLKBUFX2TS U360 ( .A(n176), .Y(n463) );
  CLKBUFX2TS U361 ( .A(requesterAddressInBuffer_WEST[1]), .Y(n175) );
  CLKBUFX2TS U362 ( .A(n175), .Y(n458) );
  CLKBUFX2TS U363 ( .A(dataInBuffer_SOUTH[2]), .Y(n569) );
  CLKBUFX2TS U364 ( .A(n569), .Y(n567) );
  CLKBUFX2TS U365 ( .A(dataInBuffer_SOUTH[3]), .Y(n574) );
  CLKBUFX2TS U366 ( .A(n574), .Y(n572) );
  CLKBUFX2TS U367 ( .A(dataInBuffer_SOUTH[1]), .Y(n564) );
  CLKBUFX2TS U368 ( .A(n564), .Y(n562) );
  CLKBUFX2TS U369 ( .A(dataInBuffer_SOUTH[0]), .Y(n559) );
  CLKBUFX2TS U370 ( .A(n559), .Y(n557) );
  CLKBUFX2TS U371 ( .A(dataInBuffer_SOUTH[4]), .Y(n578) );
  CLKBUFX2TS U372 ( .A(n578), .Y(n576) );
  CLKBUFX2TS U373 ( .A(dataInBuffer_SOUTH[5]), .Y(n583) );
  CLKBUFX2TS U374 ( .A(n583), .Y(n581) );
  CLKBUFX2TS U375 ( .A(n175), .Y(n457) );
  CLKBUFX2TS U376 ( .A(n176), .Y(n462) );
  CLKBUFX2TS U377 ( .A(n176), .Y(n460) );
  CLKBUFX2TS U378 ( .A(n175), .Y(n455) );
  CLKBUFX2TS U379 ( .A(destinationAddressInBuffer_SOUTH[1]), .Y(n180) );
  CLKBUFX2TS U380 ( .A(n180), .Y(n594) );
  CLKBUFX2TS U381 ( .A(destinationAddressInBuffer_SOUTH[2]), .Y(n181) );
  CLKBUFX2TS U382 ( .A(n181), .Y(n599) );
  CLKBUFX2TS U383 ( .A(requesterAddressInBuffer_WEST[3]), .Y(n177) );
  CLKBUFX2TS U384 ( .A(n177), .Y(n468) );
  CLKBUFX2TS U385 ( .A(destinationAddressInBuffer_SOUTH[0]), .Y(n182) );
  CLKBUFX2TS U386 ( .A(n182), .Y(n589) );
  CLKBUFX2TS U387 ( .A(destinationAddressInBuffer_SOUTH[3]), .Y(n179) );
  CLKBUFX2TS U388 ( .A(n179), .Y(n604) );
  CLKBUFX2TS U389 ( .A(requesterAddressInBuffer_WEST[0]), .Y(n178) );
  CLKBUFX2TS U390 ( .A(n178), .Y(n453) );
  CLKBUFX2TS U391 ( .A(dataInBuffer_SOUTH[0]), .Y(n558) );
  CLKBUFX2TS U392 ( .A(n558), .Y(n556) );
  CLKBUFX2TS U393 ( .A(dataInBuffer_SOUTH[2]), .Y(n568) );
  CLKBUFX2TS U394 ( .A(n568), .Y(n566) );
  CLKBUFX2TS U395 ( .A(dataInBuffer_SOUTH[3]), .Y(n573) );
  CLKBUFX2TS U396 ( .A(n573), .Y(n571) );
  CLKBUFX2TS U397 ( .A(dataInBuffer_SOUTH[1]), .Y(n563) );
  CLKBUFX2TS U398 ( .A(n563), .Y(n561) );
  CLKBUFX2TS U399 ( .A(n180), .Y(n593) );
  CLKBUFX2TS U400 ( .A(n181), .Y(n598) );
  CLKBUFX2TS U401 ( .A(n177), .Y(n467) );
  CLKBUFX2TS U402 ( .A(n182), .Y(n588) );
  CLKBUFX2TS U403 ( .A(n180), .Y(n591) );
  CLKBUFX2TS U404 ( .A(n177), .Y(n465) );
  CLKBUFX2TS U405 ( .A(n181), .Y(n596) );
  CLKBUFX2TS U406 ( .A(n182), .Y(n586) );
  CLKBUFX2TS U407 ( .A(n179), .Y(n603) );
  CLKBUFX2TS U408 ( .A(n178), .Y(n452) );
  CLKBUFX2TS U409 ( .A(n179), .Y(n601) );
  CLKBUFX2TS U410 ( .A(n178), .Y(n450) );
  CLKBUFX2TS U411 ( .A(readInBuffer_NORTH), .Y(n422) );
  CLKBUFX2TS U412 ( .A(writeInBuffer_NORTH), .Y(n421) );
  CLKBUFX2TS U413 ( .A(readInBuffer_WEST), .Y(n425) );
  CLKBUFX2TS U414 ( .A(writeInBuffer_WEST), .Y(n424) );
  CLKBUFX2TS U415 ( .A(dataInBuffer_NORTH[5]), .Y(n635) );
  CLKBUFX2TS U416 ( .A(dataInBuffer_EAST[5]), .Y(n528) );
  CLKBUFX2TS U417 ( .A(dataInBuffer_WEST[5]), .Y(n447) );
  CLKBUFX2TS U418 ( .A(dataInBuffer_NORTH[4]), .Y(n631) );
  CLKBUFX2TS U419 ( .A(dataInBuffer_EAST[4]), .Y(n523) );
  CLKBUFX2TS U420 ( .A(dataInBuffer_WEST[4]), .Y(n443) );
  CLKBUFX2TS U421 ( .A(requesterAddressInBuffer_NORTH[1]), .Y(n643) );
  CLKBUFX2TS U422 ( .A(requesterAddressInBuffer_WEST[1]), .Y(n456) );
  CLKBUFX2TS U423 ( .A(requesterAddressInBuffer_NORTH[2]), .Y(n647) );
  CLKBUFX2TS U424 ( .A(requesterAddressInBuffer_WEST[2]), .Y(n461) );
  CLKBUFX2TS U425 ( .A(dataInBuffer_WEST[5]), .Y(n448) );
  CLKBUFX2TS U426 ( .A(dataInBuffer_WEST[4]), .Y(n444) );
  CLKBUFX2TS U427 ( .A(dataInBuffer_NORTH[2]), .Y(n623) );
  CLKBUFX2TS U428 ( .A(dataInBuffer_EAST[2]), .Y(n513) );
  CLKBUFX2TS U429 ( .A(dataInBuffer_WEST[2]), .Y(n435) );
  CLKBUFX2TS U430 ( .A(dataInBuffer_NORTH[3]), .Y(n627) );
  CLKBUFX2TS U431 ( .A(dataInBuffer_EAST[3]), .Y(n518) );
  CLKBUFX2TS U432 ( .A(dataInBuffer_WEST[3]), .Y(n439) );
  CLKBUFX2TS U433 ( .A(dataInBuffer_NORTH[1]), .Y(n619) );
  CLKBUFX2TS U434 ( .A(dataInBuffer_EAST[1]), .Y(n508) );
  CLKBUFX2TS U435 ( .A(dataInBuffer_WEST[1]), .Y(n431) );
  CLKBUFX2TS U436 ( .A(dataInBuffer_NORTH[0]), .Y(n615) );
  CLKBUFX2TS U437 ( .A(dataInBuffer_EAST[0]), .Y(n503) );
  CLKBUFX2TS U438 ( .A(dataInBuffer_WEST[0]), .Y(n427) );
  CLKBUFX2TS U439 ( .A(dataInBuffer_WEST[4]), .Y(n442) );
  CLKBUFX2TS U440 ( .A(dataInBuffer_WEST[5]), .Y(n446) );
  CLKBUFX2TS U441 ( .A(requesterAddressInBuffer_NORTH[1]), .Y(n644) );
  CLKBUFX2TS U442 ( .A(requesterAddressInBuffer_NORTH[2]), .Y(n648) );
  CLKBUFX2TS U443 ( .A(requesterAddressInBuffer_NORTH[2]), .Y(n646) );
  CLKBUFX2TS U444 ( .A(requesterAddressInBuffer_SOUTH[2]), .Y(n404) );
  CLKBUFX2TS U445 ( .A(requesterAddressInBuffer_EAST[2]), .Y(n396) );
  CLKBUFX2TS U446 ( .A(requesterAddressInBuffer_NORTH[1]), .Y(n642) );
  CLKBUFX2TS U447 ( .A(requesterAddressInBuffer_SOUTH[1]), .Y(n402) );
  CLKBUFX2TS U448 ( .A(requesterAddressInBuffer_EAST[1]), .Y(n394) );
  CLKBUFX2TS U449 ( .A(readInBuffer_WEST), .Y(n672) );
  CLKBUFX2TS U450 ( .A(writeInBuffer_WEST), .Y(n670) );
  CLKBUFX2TS U451 ( .A(writeInBuffer_NORTH), .Y(n675) );
  CLKBUFX2TS U452 ( .A(destinationAddressInBuffer_WEST[4]), .Y(n487) );
  CLKBUFX2TS U453 ( .A(destinationAddressInBuffer_NORTH[4]), .Y(n655) );
  CLKBUFX2TS U454 ( .A(destinationAddressInBuffer_WEST[5]), .Y(n491) );
  CLKBUFX2TS U455 ( .A(destinationAddressInBuffer_NORTH[5]), .Y(n659) );
  CLKBUFX2TS U456 ( .A(destinationAddressInBuffer_WEST[7]), .Y(n499) );
  CLKBUFX2TS U457 ( .A(destinationAddressInBuffer_NORTH[7]), .Y(n667) );
  CLKBUFX2TS U458 ( .A(destinationAddressInBuffer_WEST[6]), .Y(n495) );
  CLKBUFX2TS U459 ( .A(destinationAddressInBuffer_NORTH[6]), .Y(n663) );
  CLKBUFX2TS U460 ( .A(requesterAddressInBuffer_NORTH[1]), .Y(n645) );
  CLKBUFX2TS U461 ( .A(requesterAddressInBuffer_EAST[1]), .Y(n395) );
  CLKBUFX2TS U462 ( .A(requesterAddressInBuffer_NORTH[2]), .Y(n649) );
  CLKBUFX2TS U463 ( .A(requesterAddressInBuffer_EAST[2]), .Y(n397) );
  CLKBUFX2TS U464 ( .A(requesterAddressInBuffer_NORTH[3]), .Y(n653) );
  CLKBUFX2TS U465 ( .A(requesterAddressInBuffer_EAST[3]), .Y(n399) );
  CLKBUFX2TS U466 ( .A(requesterAddressInBuffer_NORTH[0]), .Y(n641) );
  CLKBUFX2TS U467 ( .A(requesterAddressInBuffer_EAST[0]), .Y(n393) );
  CLKBUFX2TS U468 ( .A(destinationAddressInBuffer_SOUTH[1]), .Y(n592) );
  CLKBUFX2TS U469 ( .A(destinationAddressInBuffer_EAST[1]), .Y(n542) );
  CLKBUFX2TS U470 ( .A(destinationAddressInBuffer_WEST[1]), .Y(n475) );
  CLKBUFX2TS U471 ( .A(requesterAddressInBuffer_NORTH[3]), .Y(n651) );
  CLKBUFX2TS U472 ( .A(requesterAddressInBuffer_WEST[3]), .Y(n466) );
  CLKBUFX2TS U473 ( .A(destinationAddressInBuffer_SOUTH[2]), .Y(n597) );
  CLKBUFX2TS U474 ( .A(destinationAddressInBuffer_EAST[2]), .Y(n547) );
  CLKBUFX2TS U475 ( .A(destinationAddressInBuffer_WEST[2]), .Y(n479) );
  CLKBUFX2TS U476 ( .A(destinationAddressInBuffer_SOUTH[0]), .Y(n587) );
  CLKBUFX2TS U477 ( .A(destinationAddressInBuffer_EAST[0]), .Y(n537) );
  CLKBUFX2TS U478 ( .A(destinationAddressInBuffer_WEST[0]), .Y(n471) );
  CLKBUFX2TS U479 ( .A(destinationAddressInBuffer_SOUTH[3]), .Y(n602) );
  CLKBUFX2TS U480 ( .A(destinationAddressInBuffer_EAST[3]), .Y(n552) );
  CLKBUFX2TS U481 ( .A(destinationAddressInBuffer_WEST[3]), .Y(n483) );
  CLKBUFX2TS U482 ( .A(requesterAddressInBuffer_NORTH[0]), .Y(n639) );
  CLKBUFX2TS U483 ( .A(requesterAddressInBuffer_WEST[0]), .Y(n451) );
  CLKBUFX2TS U484 ( .A(destinationAddressInBuffer_WEST[5]), .Y(n493) );
  CLKBUFX2TS U485 ( .A(destinationAddressInBuffer_WEST[4]), .Y(n489) );
  CLKBUFX2TS U486 ( .A(destinationAddressInBuffer_WEST[6]), .Y(n497) );
  CLKBUFX2TS U487 ( .A(dataInBuffer_WEST[4]), .Y(n445) );
  CLKBUFX2TS U488 ( .A(destinationAddressInBuffer_WEST[7]), .Y(n501) );
  CLKBUFX2TS U489 ( .A(dataInBuffer_WEST[0]), .Y(n429) );
  CLKBUFX2TS U490 ( .A(dataInBuffer_WEST[1]), .Y(n433) );
  CLKBUFX2TS U491 ( .A(dataInBuffer_WEST[3]), .Y(n441) );
  CLKBUFX2TS U492 ( .A(dataInBuffer_WEST[5]), .Y(n449) );
  CLKBUFX2TS U493 ( .A(dataInBuffer_WEST[2]), .Y(n437) );
  CLKBUFX2TS U494 ( .A(destinationAddressInBuffer_WEST[3]), .Y(n485) );
  CLKBUFX2TS U495 ( .A(destinationAddressInBuffer_WEST[1]), .Y(n477) );
  CLKBUFX2TS U496 ( .A(destinationAddressInBuffer_WEST[2]), .Y(n481) );
  CLKBUFX2TS U497 ( .A(destinationAddressInBuffer_WEST[0]), .Y(n473) );
  CLKBUFX2TS U498 ( .A(dataInBuffer_WEST[0]), .Y(n428) );
  CLKBUFX2TS U499 ( .A(dataInBuffer_WEST[1]), .Y(n432) );
  CLKBUFX2TS U500 ( .A(dataInBuffer_WEST[3]), .Y(n440) );
  CLKBUFX2TS U501 ( .A(dataInBuffer_WEST[2]), .Y(n436) );
  CLKBUFX2TS U502 ( .A(dataInBuffer_WEST[0]), .Y(n426) );
  CLKBUFX2TS U503 ( .A(dataInBuffer_WEST[2]), .Y(n434) );
  CLKBUFX2TS U504 ( .A(dataInBuffer_WEST[3]), .Y(n438) );
  CLKBUFX2TS U505 ( .A(dataInBuffer_WEST[1]), .Y(n430) );
  CLKBUFX2TS U506 ( .A(destinationAddressInBuffer_WEST[1]), .Y(n476) );
  CLKBUFX2TS U507 ( .A(destinationAddressInBuffer_WEST[2]), .Y(n480) );
  CLKBUFX2TS U508 ( .A(requesterAddressInBuffer_NORTH[3]), .Y(n652) );
  CLKBUFX2TS U509 ( .A(destinationAddressInBuffer_WEST[0]), .Y(n472) );
  CLKBUFX2TS U510 ( .A(n220), .Y(n223) );
  INVX2TS U511 ( .A(n223), .Y(n679) );
  CLKBUFX2TS U512 ( .A(destinationAddressInBuffer_NORTH[1]), .Y(n410) );
  CLKBUFX2TS U513 ( .A(destinationAddressInBuffer_WEST[1]), .Y(n474) );
  CLKBUFX2TS U514 ( .A(requesterAddressInBuffer_NORTH[3]), .Y(n650) );
  CLKBUFX2TS U515 ( .A(requesterAddressInBuffer_SOUTH[3]), .Y(n406) );
  CLKBUFX2TS U516 ( .A(requesterAddressInBuffer_EAST[3]), .Y(n398) );
  CLKBUFX2TS U517 ( .A(destinationAddressInBuffer_NORTH[2]), .Y(n412) );
  CLKBUFX2TS U518 ( .A(destinationAddressInBuffer_WEST[2]), .Y(n478) );
  CLKBUFX2TS U519 ( .A(destinationAddressInBuffer_NORTH[0]), .Y(n408) );
  CLKBUFX2TS U520 ( .A(destinationAddressInBuffer_WEST[0]), .Y(n470) );
  INVX2TS U521 ( .A(n223), .Y(n681) );
  CLKBUFX2TS U522 ( .A(destinationAddressInBuffer_WEST[5]), .Y(n492) );
  CLKBUFX2TS U523 ( .A(destinationAddressInBuffer_NORTH[5]), .Y(n417) );
  CLKBUFX2TS U524 ( .A(destinationAddressInBuffer_WEST[7]), .Y(n500) );
  CLKBUFX2TS U525 ( .A(destinationAddressInBuffer_NORTH[7]), .Y(n419) );
  CLKBUFX2TS U526 ( .A(destinationAddressInBuffer_WEST[4]), .Y(n488) );
  CLKBUFX2TS U527 ( .A(destinationAddressInBuffer_NORTH[4]), .Y(n416) );
  CLKBUFX2TS U528 ( .A(destinationAddressInBuffer_WEST[6]), .Y(n496) );
  CLKBUFX2TS U529 ( .A(destinationAddressInBuffer_NORTH[6]), .Y(n418) );
  CLKBUFX2TS U530 ( .A(destinationAddressInBuffer_WEST[7]), .Y(n498) );
  CLKBUFX2TS U531 ( .A(destinationAddressInBuffer_NORTH[7]), .Y(n666) );
  CLKBUFX2TS U532 ( .A(destinationAddressInBuffer_WEST[6]), .Y(n494) );
  CLKBUFX2TS U533 ( .A(destinationAddressInBuffer_NORTH[6]), .Y(n662) );
  CLKBUFX2TS U534 ( .A(destinationAddressInBuffer_WEST[5]), .Y(n490) );
  CLKBUFX2TS U535 ( .A(destinationAddressInBuffer_NORTH[5]), .Y(n658) );
  CLKBUFX2TS U536 ( .A(destinationAddressInBuffer_WEST[4]), .Y(n486) );
  CLKBUFX2TS U537 ( .A(destinationAddressInBuffer_NORTH[4]), .Y(n654) );
  CLKBUFX2TS U538 ( .A(destinationAddressInBuffer_WEST[3]), .Y(n484) );
  CLKBUFX2TS U539 ( .A(requesterAddressInBuffer_NORTH[0]), .Y(n640) );
  CLKBUFX2TS U540 ( .A(destinationAddressInBuffer_NORTH[3]), .Y(n414) );
  CLKBUFX2TS U541 ( .A(destinationAddressInBuffer_WEST[3]), .Y(n482) );
  CLKBUFX2TS U542 ( .A(requesterAddressInBuffer_NORTH[0]), .Y(n638) );
  CLKBUFX2TS U543 ( .A(requesterAddressInBuffer_SOUTH[0]), .Y(n400) );
  CLKBUFX2TS U544 ( .A(requesterAddressInBuffer_EAST[0]), .Y(n392) );
  CLKBUFX2TS U545 ( .A(dataInBuffer_NORTH[4]), .Y(n159) );
  CLKBUFX2TS U546 ( .A(n159), .Y(n633) );
  CLKBUFX2TS U547 ( .A(dataInBuffer_EAST[4]), .Y(n161) );
  CLKBUFX2TS U548 ( .A(n161), .Y(n525) );
  CLKBUFX2TS U549 ( .A(dataInBuffer_NORTH[5]), .Y(n160) );
  CLKBUFX2TS U550 ( .A(n160), .Y(n637) );
  CLKBUFX2TS U551 ( .A(dataInBuffer_EAST[5]), .Y(n162) );
  CLKBUFX2TS U552 ( .A(n162), .Y(n530) );
  CLKBUFX2TS U553 ( .A(dataInBuffer_NORTH[3]), .Y(n167) );
  CLKBUFX2TS U554 ( .A(n167), .Y(n629) );
  CLKBUFX2TS U555 ( .A(dataInBuffer_EAST[3]), .Y(n168) );
  CLKBUFX2TS U556 ( .A(n168), .Y(n520) );
  CLKBUFX2TS U557 ( .A(dataInBuffer_NORTH[0]), .Y(n163) );
  CLKBUFX2TS U558 ( .A(n163), .Y(n617) );
  CLKBUFX2TS U559 ( .A(dataInBuffer_EAST[0]), .Y(n164) );
  CLKBUFX2TS U560 ( .A(n164), .Y(n505) );
  CLKBUFX2TS U561 ( .A(dataInBuffer_NORTH[1]), .Y(n169) );
  CLKBUFX2TS U562 ( .A(n169), .Y(n621) );
  CLKBUFX2TS U563 ( .A(dataInBuffer_EAST[1]), .Y(n170) );
  CLKBUFX2TS U564 ( .A(n170), .Y(n510) );
  CLKBUFX2TS U565 ( .A(dataInBuffer_NORTH[2]), .Y(n165) );
  CLKBUFX2TS U566 ( .A(n165), .Y(n625) );
  CLKBUFX2TS U567 ( .A(dataInBuffer_EAST[2]), .Y(n166) );
  CLKBUFX2TS U568 ( .A(n166), .Y(n515) );
  CLKBUFX2TS U569 ( .A(n160), .Y(n636) );
  CLKBUFX2TS U570 ( .A(n162), .Y(n529) );
  CLKBUFX2TS U571 ( .A(n159), .Y(n632) );
  CLKBUFX2TS U572 ( .A(n161), .Y(n524) );
  CLKBUFX2TS U573 ( .A(n159), .Y(n630) );
  CLKBUFX2TS U574 ( .A(n161), .Y(n522) );
  CLKBUFX2TS U575 ( .A(n160), .Y(n634) );
  CLKBUFX2TS U576 ( .A(n162), .Y(n527) );
  CLKBUFX2TS U577 ( .A(destinationAddressInBuffer_EAST[1]), .Y(n171) );
  CLKBUFX2TS U578 ( .A(n171), .Y(n544) );
  CLKBUFX2TS U579 ( .A(destinationAddressInBuffer_EAST[2]), .Y(n172) );
  CLKBUFX2TS U580 ( .A(n172), .Y(n549) );
  CLKBUFX2TS U581 ( .A(destinationAddressInBuffer_EAST[0]), .Y(n173) );
  CLKBUFX2TS U582 ( .A(n173), .Y(n539) );
  CLKBUFX2TS U583 ( .A(destinationAddressInBuffer_EAST[3]), .Y(n174) );
  CLKBUFX2TS U584 ( .A(n174), .Y(n554) );
  CLKBUFX2TS U585 ( .A(n161), .Y(n526) );
  CLKBUFX2TS U586 ( .A(n164), .Y(n506) );
  CLKBUFX2TS U587 ( .A(n170), .Y(n511) );
  CLKBUFX2TS U588 ( .A(n168), .Y(n521) );
  CLKBUFX2TS U589 ( .A(n162), .Y(n531) );
  CLKBUFX2TS U590 ( .A(n166), .Y(n516) );
  CLKBUFX2TS U591 ( .A(n174), .Y(n555) );
  CLKBUFX2TS U592 ( .A(n171), .Y(n545) );
  CLKBUFX2TS U593 ( .A(n172), .Y(n550) );
  CLKBUFX2TS U594 ( .A(n173), .Y(n540) );
  CLKBUFX2TS U595 ( .A(n163), .Y(n616) );
  CLKBUFX2TS U596 ( .A(n164), .Y(n504) );
  CLKBUFX2TS U597 ( .A(n169), .Y(n620) );
  CLKBUFX2TS U598 ( .A(n170), .Y(n509) );
  CLKBUFX2TS U599 ( .A(n167), .Y(n628) );
  CLKBUFX2TS U600 ( .A(n168), .Y(n519) );
  CLKBUFX2TS U601 ( .A(n165), .Y(n624) );
  CLKBUFX2TS U602 ( .A(n166), .Y(n514) );
  CLKBUFX2TS U603 ( .A(n163), .Y(n614) );
  CLKBUFX2TS U604 ( .A(n164), .Y(n502) );
  CLKBUFX2TS U605 ( .A(n165), .Y(n622) );
  CLKBUFX2TS U606 ( .A(n166), .Y(n512) );
  CLKBUFX2TS U607 ( .A(n167), .Y(n626) );
  CLKBUFX2TS U608 ( .A(n168), .Y(n517) );
  CLKBUFX2TS U609 ( .A(n169), .Y(n618) );
  CLKBUFX2TS U610 ( .A(n170), .Y(n507) );
  CLKBUFX2TS U611 ( .A(n171), .Y(n543) );
  CLKBUFX2TS U612 ( .A(n172), .Y(n548) );
  CLKBUFX2TS U613 ( .A(n173), .Y(n538) );
  CLKBUFX2TS U614 ( .A(n171), .Y(n541) );
  CLKBUFX2TS U615 ( .A(n172), .Y(n546) );
  CLKBUFX2TS U616 ( .A(n173), .Y(n536) );
  CLKBUFX2TS U617 ( .A(n174), .Y(n553) );
  CLKBUFX2TS U618 ( .A(n174), .Y(n551) );
  CLKBUFX2TS U619 ( .A(n422), .Y(n678) );
  CLKBUFX2TS U620 ( .A(n425), .Y(n673) );
  CLKBUFX2TS U621 ( .A(readInBuffer_NORTH), .Y(n677) );
  CLKBUFX2TS U622 ( .A(n416), .Y(n657) );
  CLKBUFX2TS U623 ( .A(n417), .Y(n661) );
  CLKBUFX2TS U624 ( .A(n419), .Y(n669) );
  CLKBUFX2TS U625 ( .A(n418), .Y(n665) );
  CLKBUFX2TS U626 ( .A(n395), .Y(n533) );
  CLKBUFX2TS U627 ( .A(n175), .Y(n459) );
  CLKBUFX2TS U628 ( .A(n397), .Y(n534) );
  CLKBUFX2TS U629 ( .A(n176), .Y(n464) );
  CLKBUFX2TS U630 ( .A(n399), .Y(n535) );
  CLKBUFX2TS U631 ( .A(n177), .Y(n469) );
  CLKBUFX2TS U632 ( .A(n393), .Y(n532) );
  CLKBUFX2TS U633 ( .A(n178), .Y(n454) );
  CLKBUFX2TS U634 ( .A(destinationAddressInBuffer_SOUTH[5]), .Y(n609) );
  CLKBUFX2TS U635 ( .A(destinationAddressInBuffer_SOUTH[4]), .Y(n607) );
  CLKBUFX2TS U636 ( .A(destinationAddressInBuffer_SOUTH[6]), .Y(n611) );
  CLKBUFX2TS U637 ( .A(dataInBuffer_SOUTH[4]), .Y(n580) );
  CLKBUFX2TS U638 ( .A(destinationAddressInBuffer_SOUTH[7]), .Y(n613) );
  CLKBUFX2TS U639 ( .A(dataInBuffer_SOUTH[0]), .Y(n560) );
  CLKBUFX2TS U640 ( .A(dataInBuffer_SOUTH[1]), .Y(n565) );
  CLKBUFX2TS U641 ( .A(dataInBuffer_SOUTH[3]), .Y(n575) );
  CLKBUFX2TS U642 ( .A(dataInBuffer_SOUTH[5]), .Y(n585) );
  CLKBUFX2TS U643 ( .A(dataInBuffer_SOUTH[2]), .Y(n570) );
  CLKBUFX2TS U644 ( .A(n179), .Y(n605) );
  CLKBUFX2TS U645 ( .A(n180), .Y(n595) );
  CLKBUFX2TS U646 ( .A(n181), .Y(n600) );
  CLKBUFX2TS U647 ( .A(n182), .Y(n590) );
  CLKBUFX2TS U648 ( .A(n424), .Y(n671) );
  CLKBUFX2TS U649 ( .A(n421), .Y(n676) );
  CLKBUFX2TS U650 ( .A(n417), .Y(n660) );
  CLKBUFX2TS U651 ( .A(n419), .Y(n668) );
  CLKBUFX2TS U652 ( .A(n416), .Y(n656) );
  CLKBUFX2TS U653 ( .A(n418), .Y(n664) );
  CLKBUFX2TS U654 ( .A(readInBuffer_SOUTH), .Y(n420) );
  CLKBUFX2TS U655 ( .A(requesterAddressInBuffer_SOUTH[0]), .Y(n401) );
  CLKBUFX2TS U656 ( .A(requesterAddressInBuffer_SOUTH[1]), .Y(n403) );
  CLKBUFX2TS U657 ( .A(requesterAddressInBuffer_SOUTH[2]), .Y(n405) );
  CLKBUFX2TS U658 ( .A(requesterAddressInBuffer_SOUTH[3]), .Y(n407) );
  CLKBUFX2TS U659 ( .A(destinationAddressInBuffer_NORTH[0]), .Y(n409) );
  CLKBUFX2TS U660 ( .A(destinationAddressInBuffer_NORTH[3]), .Y(n415) );
  CLKBUFX2TS U661 ( .A(destinationAddressInBuffer_NORTH[2]), .Y(n413) );
  CLKBUFX2TS U662 ( .A(destinationAddressInBuffer_NORTH[1]), .Y(n411) );
  NOR2BX1TS U664 ( .AN(dataIn_WEST[0]), .B(n290), .Y(N94) );
  CLKBUFX2TS U665 ( .A(n194), .Y(n206) );
  CLKBUFX2TS U666 ( .A(n206), .Y(n238) );
  INVX2TS U667 ( .A(n238), .Y(n183) );
  NOR2BX1TS U668 ( .AN(dataIn_WEST[1]), .B(n183), .Y(N95) );
  NOR2BX1TS U669 ( .AN(dataIn_WEST[2]), .B(n183), .Y(N96) );
  NOR2BX1TS U670 ( .AN(dataIn_WEST[3]), .B(n183), .Y(N97) );
  NOR2BX1TS U671 ( .AN(dataIn_WEST[4]), .B(n183), .Y(N98) );
  INVX2TS U672 ( .A(n238), .Y(n184) );
  NOR2BX1TS U673 ( .AN(dataIn_WEST[5]), .B(n184), .Y(N99) );
  NOR2BX1TS U674 ( .AN(writeIn_WEST), .B(n184), .Y(N93) );
  NOR2BX1TS U675 ( .AN(readIn_WEST), .B(n184), .Y(N92) );
  NOR2BX1TS U676 ( .AN(requesterAddressIn_WEST[0]), .B(n184), .Y(N88) );
  INVX2TS U677 ( .A(n238), .Y(n185) );
  NOR2BX1TS U678 ( .AN(requesterAddressIn_WEST[1]), .B(n185), .Y(N89) );
  NOR2BX1TS U679 ( .AN(requesterAddressIn_WEST[2]), .B(n185), .Y(N90) );
  NOR2BX1TS U680 ( .AN(requesterAddressIn_WEST[3]), .B(n185), .Y(N91) );
  NOR2BX1TS U681 ( .AN(destinationAddressIn_WEST[0]), .B(n185), .Y(N76) );
  CLKBUFX2TS U682 ( .A(n194), .Y(n218) );
  CLKBUFX2TS U683 ( .A(n218), .Y(n263) );
  INVX2TS U684 ( .A(n263), .Y(n186) );
  NOR2BX1TS U685 ( .AN(destinationAddressIn_WEST[1]), .B(n186), .Y(N77) );
  NOR2BX1TS U686 ( .AN(destinationAddressIn_WEST[2]), .B(n186), .Y(N78) );
  NOR2BX1TS U687 ( .AN(destinationAddressIn_WEST[3]), .B(n186), .Y(N79) );
  NOR2BX1TS U688 ( .AN(destinationAddressIn_WEST[4]), .B(n186), .Y(N80) );
  INVX2TS U689 ( .A(n263), .Y(n189) );
  NOR2BX1TS U690 ( .AN(destinationAddressIn_WEST[5]), .B(n189), .Y(N81) );
  NOR2BX1TS U691 ( .AN(destinationAddressIn_WEST[6]), .B(n189), .Y(N82) );
  NOR2BX1TS U692 ( .AN(destinationAddressIn_WEST[7]), .B(n189), .Y(N83) );
  CLKBUFX2TS U693 ( .A(destinationAddressIn_WEST[8]), .Y(n187) );
  NOR2BX1TS U694 ( .AN(n187), .B(n189), .Y(N84) );
  CLKBUFX2TS U695 ( .A(destinationAddressIn_WEST[9]), .Y(n190) );
  INVX2TS U696 ( .A(n263), .Y(n193) );
  NOR2BX1TS U697 ( .AN(n190), .B(n193), .Y(N85) );
  CLKBUFX2TS U698 ( .A(destinationAddressIn_WEST[10]), .Y(n191) );
  NOR2BX1TS U699 ( .AN(n191), .B(n193), .Y(N86) );
  CLKBUFX2TS U700 ( .A(destinationAddressIn_WEST[11]), .Y(n192) );
  NOR2BX1TS U701 ( .AN(n192), .B(n193), .Y(N87) );
  NOR2BX1TS U702 ( .AN(dataIn_EAST[0]), .B(n193), .Y(N70) );
  CLKBUFX2TS U703 ( .A(n194), .Y(n211) );
  CLKBUFX2TS U704 ( .A(n211), .Y(n293) );
  INVX2TS U705 ( .A(n293), .Y(n195) );
  NOR2BX1TS U706 ( .AN(dataIn_EAST[1]), .B(n195), .Y(N71) );
  NOR2BX1TS U707 ( .AN(dataIn_EAST[2]), .B(n195), .Y(N72) );
  NOR2BX1TS U708 ( .AN(dataIn_EAST[3]), .B(n195), .Y(N73) );
  NOR2BX1TS U709 ( .AN(dataIn_EAST[4]), .B(n195), .Y(N74) );
  INVX2TS U710 ( .A(n293), .Y(n196) );
  NOR2BX1TS U711 ( .AN(dataIn_EAST[5]), .B(n196), .Y(N75) );
  NOR2BX1TS U712 ( .AN(writeIn_EAST), .B(n196), .Y(N69) );
  NOR2BX1TS U713 ( .AN(readIn_EAST), .B(n196), .Y(N68) );
  NOR2BX1TS U714 ( .AN(requesterAddressIn_EAST[0]), .B(n196), .Y(N64) );
  INVX2TS U715 ( .A(n293), .Y(n197) );
  NOR2BX1TS U716 ( .AN(requesterAddressIn_EAST[1]), .B(n197), .Y(N65) );
  NOR2BX1TS U717 ( .AN(requesterAddressIn_EAST[2]), .B(n197), .Y(N66) );
  NOR2BX1TS U718 ( .AN(requesterAddressIn_EAST[3]), .B(n197), .Y(N67) );
  NOR2BX1TS U719 ( .AN(destinationAddressIn_EAST[0]), .B(n197), .Y(N52) );
  CLKBUFX2TS U720 ( .A(n220), .Y(n329) );
  INVX2TS U721 ( .A(n329), .Y(n198) );
  NOR2BX1TS U722 ( .AN(destinationAddressIn_EAST[1]), .B(n198), .Y(N53) );
  NOR2BX1TS U723 ( .AN(destinationAddressIn_EAST[2]), .B(n198), .Y(N54) );
  NOR2BX1TS U724 ( .AN(destinationAddressIn_EAST[3]), .B(n198), .Y(N55) );
  NOR2BX1TS U725 ( .AN(destinationAddressIn_EAST[4]), .B(n198), .Y(N56) );
  INVX2TS U726 ( .A(n329), .Y(n200) );
  NOR2BX1TS U727 ( .AN(destinationAddressIn_EAST[5]), .B(n200), .Y(N57) );
  NOR2BX1TS U728 ( .AN(destinationAddressIn_EAST[6]), .B(n200), .Y(N58) );
  NOR2BX1TS U729 ( .AN(destinationAddressIn_EAST[7]), .B(n200), .Y(N59) );
  CLKBUFX2TS U730 ( .A(destinationAddressIn_EAST[8]), .Y(n199) );
  NOR2BX1TS U731 ( .AN(n199), .B(n200), .Y(N60) );
  CLKBUFX2TS U732 ( .A(destinationAddressIn_EAST[9]), .Y(n201) );
  INVX2TS U733 ( .A(n329), .Y(n204) );
  NOR2BX1TS U734 ( .AN(n201), .B(n204), .Y(N61) );
  CLKBUFX2TS U735 ( .A(destinationAddressIn_EAST[10]), .Y(n202) );
  NOR2BX1TS U736 ( .AN(n202), .B(n204), .Y(N62) );
  CLKBUFX2TS U737 ( .A(destinationAddressIn_EAST[11]), .Y(n203) );
  NOR2BX1TS U738 ( .AN(n203), .B(n204), .Y(N63) );
  NOR2BX1TS U739 ( .AN(dataIn_SOUTH[0]), .B(n204), .Y(N46) );
  INVX2TS U740 ( .A(n206), .Y(n217) );
  NOR2BX1TS U741 ( .AN(dataIn_SOUTH[1]), .B(n217), .Y(N47) );
  NOR2BX1TS U742 ( .AN(dataIn_SOUTH[2]), .B(n217), .Y(N48) );
  NOR2BX1TS U743 ( .AN(dataIn_SOUTH[3]), .B(n217), .Y(N49) );
  INVX2TS U744 ( .A(n206), .Y(n205) );
  NOR2BX1TS U745 ( .AN(dataIn_SOUTH[4]), .B(n205), .Y(N50) );
  NOR2BX1TS U746 ( .AN(dataIn_SOUTH[5]), .B(n205), .Y(N51) );
  NOR2BX1TS U747 ( .AN(writeIn_SOUTH), .B(n205), .Y(N45) );
  NOR2BX1TS U748 ( .AN(readIn_SOUTH), .B(n205), .Y(N44) );
  INVX2TS U749 ( .A(n206), .Y(n207) );
  NOR2BX1TS U750 ( .AN(requesterAddressIn_SOUTH[0]), .B(n207), .Y(N40) );
  NOR2BX1TS U751 ( .AN(requesterAddressIn_SOUTH[1]), .B(n207), .Y(N41) );
  NOR2BX1TS U752 ( .AN(requesterAddressIn_SOUTH[2]), .B(n207), .Y(N42) );
  NOR2BX1TS U753 ( .AN(requesterAddressIn_SOUTH[3]), .B(n207), .Y(N43) );
  INVX2TS U754 ( .A(n211), .Y(n208) );
  NOR2BX1TS U755 ( .AN(destinationAddressIn_SOUTH[0]), .B(n208), .Y(N28) );
  NOR2BX1TS U756 ( .AN(destinationAddressIn_SOUTH[1]), .B(n208), .Y(N29) );
  NOR2BX1TS U757 ( .AN(destinationAddressIn_SOUTH[2]), .B(n208), .Y(N30) );
  NOR2BX1TS U758 ( .AN(destinationAddressIn_SOUTH[3]), .B(n208), .Y(N31) );
  INVX2TS U759 ( .A(n211), .Y(n209) );
  NOR2BX1TS U760 ( .AN(destinationAddressIn_SOUTH[4]), .B(n209), .Y(N32) );
  NOR2BX1TS U761 ( .AN(destinationAddressIn_SOUTH[5]), .B(n209), .Y(N33) );
  NOR2BX1TS U762 ( .AN(destinationAddressIn_SOUTH[6]), .B(n209), .Y(N34) );
  NOR2BX1TS U763 ( .AN(destinationAddressIn_SOUTH[7]), .B(n209), .Y(N35) );
  CLKBUFX2TS U764 ( .A(destinationAddressIn_SOUTH[8]), .Y(n210) );
  INVX2TS U765 ( .A(n211), .Y(n215) );
  NOR2BX1TS U766 ( .AN(n210), .B(n215), .Y(N36) );
  CLKBUFX2TS U767 ( .A(destinationAddressIn_SOUTH[9]), .Y(n212) );
  NOR2BX1TS U768 ( .AN(n212), .B(n215), .Y(N37) );
  CLKBUFX2TS U769 ( .A(destinationAddressIn_SOUTH[10]), .Y(n213) );
  NOR2BX1TS U770 ( .AN(n213), .B(n215), .Y(N38) );
  CLKBUFX2TS U771 ( .A(destinationAddressIn_SOUTH[11]), .Y(n214) );
  NOR2BX1TS U772 ( .AN(n214), .B(n215), .Y(N39) );
  INVX2TS U773 ( .A(n218), .Y(n216) );
  NOR2BX1TS U774 ( .AN(dataIn_NORTH[0]), .B(n216), .Y(N22) );
  NOR2BX1TS U775 ( .AN(dataIn_NORTH[1]), .B(n216), .Y(N23) );
  NOR2BX1TS U776 ( .AN(dataIn_NORTH[2]), .B(n216), .Y(N24) );
  NOR2BX1TS U777 ( .AN(dataIn_NORTH[3]), .B(n216), .Y(N25) );
  INVX2TS U778 ( .A(n218), .Y(n325) );
  NOR2BX1TS U779 ( .AN(dataIn_NORTH[4]), .B(n325), .Y(N26) );
  NOR2BX1TS U780 ( .AN(dataIn_NORTH[5]), .B(n217), .Y(N27) );
  NOR2BX1TS U781 ( .AN(writeIn_NORTH), .B(n325), .Y(N21) );
  NOR2BX1TS U782 ( .AN(readIn_NORTH), .B(n325), .Y(N20) );
  INVX2TS U783 ( .A(n218), .Y(n219) );
  NOR2BX1TS U784 ( .AN(requesterAddressIn_NORTH[0]), .B(n219), .Y(N16) );
  NOR2BX1TS U785 ( .AN(requesterAddressIn_NORTH[1]), .B(n219), .Y(N17) );
  NOR2BX1TS U786 ( .AN(requesterAddressIn_NORTH[2]), .B(n219), .Y(N18) );
  NOR2BX1TS U787 ( .AN(requesterAddressIn_NORTH[3]), .B(n219), .Y(N19) );
  NOR2BX1TS U788 ( .AN(destinationAddressIn_NORTH[0]), .B(n679), .Y(N4) );
  NOR2BX1TS U789 ( .AN(destinationAddressIn_NORTH[1]), .B(n680), .Y(N5) );
  NOR2BX1TS U790 ( .AN(destinationAddressIn_NORTH[2]), .B(n681), .Y(N6) );
  NOR2BX1TS U791 ( .AN(destinationAddressIn_NORTH[3]), .B(n158), .Y(N7) );
  INVX2TS U792 ( .A(n223), .Y(n221) );
  NOR2BX1TS U793 ( .AN(destinationAddressIn_NORTH[4]), .B(n221), .Y(N8) );
  NOR2BX1TS U794 ( .AN(destinationAddressIn_NORTH[5]), .B(n221), .Y(N9) );
  NOR2BX1TS U795 ( .AN(destinationAddressIn_NORTH[6]), .B(n221), .Y(N10) );
  NOR2BX1TS U796 ( .AN(destinationAddressIn_NORTH[7]), .B(n221), .Y(N11) );
  CLKBUFX2TS U797 ( .A(destinationAddressIn_NORTH[8]), .Y(n222) );
  INVX2TS U798 ( .A(n223), .Y(n227) );
  NOR2BX1TS U799 ( .AN(n222), .B(n227), .Y(N12) );
  CLKBUFX2TS U800 ( .A(destinationAddressIn_NORTH[9]), .Y(n224) );
  NOR2BX1TS U801 ( .AN(n224), .B(n227), .Y(N13) );
  CLKBUFX2TS U802 ( .A(destinationAddressIn_NORTH[10]), .Y(n225) );
  NOR2BX1TS U803 ( .AN(n225), .B(n227), .Y(N14) );
  CLKBUFX2TS U804 ( .A(destinationAddressIn_NORTH[11]), .Y(n226) );
  NOR2BX1TS U805 ( .AN(n226), .B(n227), .Y(N15) );
  CLKBUFX2TS U806 ( .A(localRouterAddress[2]), .Y(n243) );
  INVX2TS U807 ( .A(n243), .Y(n269) );
  CLKBUFX2TS U808 ( .A(localRouterAddress[3]), .Y(n228) );
  INVX2TS U809 ( .A(n228), .Y(n229) );
  INVX2TS U810 ( .A(n229), .Y(n317) );
  INVX2TS U811 ( .A(n317), .Y(n332) );
  CLKAND2X2TS U812 ( .A(n226), .B(n332), .Y(n244) );
  INVX2TS U813 ( .A(n243), .Y(n314) );
  OAI22X1TS U814 ( .A0(n225), .A1(n314), .B0(n226), .B1(n229), .Y(n239) );
  AOI211XLTS U815 ( .A0(n225), .A1(n269), .B0(n244), .C0(n239), .Y(n253) );
  CLKBUFX2TS U816 ( .A(localRouterAddress[1]), .Y(n231) );
  INVX2TS U817 ( .A(n232), .Y(n303) );
  INVX2TS U818 ( .A(n303), .Y(n316) );
  OR2X1TS U819 ( .A(n230), .B(n316), .Y(n235) );
  CLKBUFX2TS U820 ( .A(localRouterAddress[0]), .Y(n233) );
  INVX2TS U821 ( .A(n233), .Y(n324) );
  INVX2TS U822 ( .A(n303), .Y(n336) );
  AOI22X1TS U823 ( .A0(n222), .A1(n324), .B0(n230), .B1(n336), .Y(n234) );
  INVX2TS U824 ( .A(n233), .Y(n322) );
  OR2X1TS U825 ( .A(n222), .B(n322), .Y(n249) );
  NAND4XLTS U826 ( .A(n253), .B(n235), .C(n234), .D(n249), .Y(n251) );
  NOR2XLTS U827 ( .A(n290), .B(n251), .Y(n259) );
  NOR3XLTS U828 ( .A(n326), .B(n422), .C(n421), .Y(n237) );
  OAI21XLTS U829 ( .A0(readInBuffer_NORTH), .A1(writeInBuffer_NORTH), .B0(n238), .Y(n247) );
  INVX2TS U830 ( .A(n247), .Y(n252) );
  NAND2X1TS U831 ( .A(n252), .B(n239), .Y(n242) );
  OAI2BB2XLTS U832 ( .B0(n244), .B1(n242), .A0N(outputPortSelect_NORTH[0]), 
        .A1N(n241), .Y(n95) );
  INVX2TS U833 ( .A(n243), .Y(n318) );
  OR2X1TS U834 ( .A(n226), .B(n229), .Y(n245) );
  AOI31XLTS U835 ( .A0(n225), .A1(n318), .A2(n245), .B0(n244), .Y(n248) );
  OAI2BB2XLTS U836 ( .B0(n248), .B1(n247), .A0N(n237), .A1N(
        outputPortSelect_NORTH[1]), .Y(n94) );
  INVX2TS U837 ( .A(n231), .Y(n287) );
  CLKAND2X2TS U838 ( .A(n224), .B(n316), .Y(n250) );
  OAI22X1TS U839 ( .A0(n224), .A1(n287), .B0(n250), .B1(n249), .Y(n255) );
  NAND3XLTS U840 ( .A(n253), .B(n252), .C(n251), .Y(n258) );
  OAI2BB2XLTS U841 ( .B0(n255), .B1(n258), .A0N(n241), .A1N(
        outputPortSelect_NORTH[2]), .Y(n93) );
  INVX2TS U842 ( .A(n255), .Y(n257) );
  OAI2BB2XLTS U843 ( .B0(n258), .B1(n257), .A0N(outputPortSelect_NORTH[3]), 
        .A1N(n241), .Y(n92) );
  NOR2BX1TS U844 ( .AN(n214), .B(n228), .Y(n267) );
  OAI22X1TS U845 ( .A0(n213), .A1(n269), .B0(n214), .B1(n229), .Y(n264) );
  AOI211XLTS U846 ( .A0(n213), .A1(n318), .B0(n267), .C0(n264), .Y(n277) );
  AOI22X1TS U847 ( .A0(n210), .A1(n324), .B0(n260), .B1(n232), .Y(n262) );
  OR2X1TS U848 ( .A(n260), .B(n287), .Y(n261) );
  OR2X1TS U849 ( .A(n210), .B(n322), .Y(n273) );
  NAND4XLTS U850 ( .A(n277), .B(n262), .C(n261), .D(n273), .Y(n275) );
  NOR2XLTS U851 ( .A(n290), .B(n275), .Y(n285) );
  NOR3XLTS U852 ( .A(n326), .B(n423), .C(writeInBuffer_SOUTH), .Y(n279) );
  CLKBUFX2TS U853 ( .A(n279), .Y(n284) );
  OAI21XLTS U854 ( .A0(readInBuffer_SOUTH), .A1(writeInBuffer_SOUTH), .B0(n263), .Y(n271) );
  INVX2TS U855 ( .A(n271), .Y(n276) );
  NAND2X1TS U856 ( .A(n276), .B(n264), .Y(n266) );
  OAI2BB2XLTS U857 ( .B0(n267), .B1(n266), .A0N(outputPortSelect_SOUTH[0]), 
        .A1N(n279), .Y(n89) );
  OR2X1TS U858 ( .A(n214), .B(n332), .Y(n268) );
  AOI31XLTS U859 ( .A0(n213), .A1(n269), .A2(n268), .B0(n267), .Y(n272) );
  OAI2BB2XLTS U860 ( .B0(n272), .B1(n271), .A0N(n279), .A1N(
        outputPortSelect_SOUTH[1]), .Y(n88) );
  NOR2BX1TS U861 ( .AN(n212), .B(n303), .Y(n274) );
  OAI22X1TS U862 ( .A0(n212), .A1(n316), .B0(n274), .B1(n273), .Y(n280) );
  NAND3XLTS U863 ( .A(n277), .B(n276), .C(n275), .Y(n283) );
  OAI2BB2XLTS U864 ( .B0(n280), .B1(n283), .A0N(n279), .A1N(
        outputPortSelect_SOUTH[2]), .Y(n87) );
  INVX2TS U865 ( .A(n280), .Y(n282) );
  OAI2BB2XLTS U866 ( .B0(n283), .B1(n282), .A0N(outputPortSelect_SOUTH[3]), 
        .A1N(n284), .Y(n86) );
  NOR2BX1TS U867 ( .AN(n203), .B(n228), .Y(n298) );
  OAI22X1TS U868 ( .A0(n202), .A1(n318), .B0(n203), .B1(n332), .Y(n294) );
  AOI211XLTS U869 ( .A0(n202), .A1(n314), .B0(n298), .C0(n294), .Y(n308) );
  AOI22X1TS U870 ( .A0(n199), .A1(n324), .B0(n286), .B1(n287), .Y(n289) );
  OR2X1TS U871 ( .A(n286), .B(n287), .Y(n288) );
  OR2X1TS U872 ( .A(n199), .B(n322), .Y(n304) );
  NAND4XLTS U873 ( .A(n308), .B(n289), .C(n288), .D(n304), .Y(n306) );
  NOR2XLTS U874 ( .A(n290), .B(n306), .Y(n313) );
  NOR3XLTS U875 ( .A(n326), .B(n391), .C(n384), .Y(n291) );
  OAI21XLTS U876 ( .A0(n390), .A1(n383), .B0(n293), .Y(n301) );
  INVX2TS U877 ( .A(n301), .Y(n307) );
  NAND2X1TS U878 ( .A(n307), .B(n294), .Y(n297) );
  OAI2BB2XLTS U879 ( .B0(n298), .B1(n297), .A0N(outputPortSelect_EAST[0]), 
        .A1N(n291), .Y(n83) );
  OR2X1TS U880 ( .A(n203), .B(n320), .Y(n299) );
  AOI31XLTS U881 ( .A0(n202), .A1(n314), .A2(n299), .B0(n298), .Y(n302) );
  OAI2BB2XLTS U882 ( .B0(n302), .B1(n301), .A0N(n296), .A1N(
        outputPortSelect_EAST[1]), .Y(n82) );
  NOR2BX1TS U883 ( .AN(n201), .B(n303), .Y(n305) );
  OAI22X1TS U884 ( .A0(n201), .A1(n336), .B0(n305), .B1(n304), .Y(n309) );
  NAND3XLTS U885 ( .A(n308), .B(n307), .C(n306), .Y(n312) );
  OAI2BB2XLTS U886 ( .B0(n309), .B1(n312), .A0N(n296), .A1N(
        outputPortSelect_EAST[2]), .Y(n81) );
  INVX2TS U887 ( .A(n309), .Y(n311) );
  OAI2BB2XLTS U888 ( .B0(n312), .B1(n311), .A0N(outputPortSelect_EAST[3]), 
        .A1N(n291), .Y(n80) );
  NAND2X1TS U889 ( .A(n191), .B(n314), .Y(n338) );
  INVX2TS U890 ( .A(n338), .Y(n334) );
  NOR2XLTS U891 ( .A(n315), .B(n316), .Y(n319) );
  INVX2TS U892 ( .A(n317), .Y(n320) );
  OAI22X1TS U893 ( .A0(n191), .A1(n318), .B0(n192), .B1(n320), .Y(n342) );
  AOI211XLTS U894 ( .A0(n315), .A1(n336), .B0(n319), .C0(n342), .Y(n321) );
  NAND2X1TS U895 ( .A(n192), .B(n320), .Y(n339) );
  OAI211XLTS U896 ( .A0(n187), .A1(n322), .B0(n321), .C0(n339), .Y(n323) );
  AOI211XLTS U897 ( .A0(n187), .A1(n324), .B0(n334), .C0(n323), .Y(n343) );
  NOR2BX1TS U898 ( .AN(n343), .B(n325), .Y(n347) );
  NOR3XLTS U899 ( .A(n326), .B(n425), .C(n424), .Y(n327) );
  AO22XLTS U900 ( .A0(writeInBuffer_WEST), .A1(n347), .B0(n330), .B1(
        memWrite_WEST), .Y(n78) );
  OAI21XLTS U901 ( .A0(readInBuffer_WEST), .A1(writeInBuffer_WEST), .B0(n329), 
        .Y(n341) );
  NAND2X1TS U902 ( .A(n342), .B(n339), .Y(n331) );
  OAI2BB2XLTS U903 ( .B0(n341), .B1(n331), .A0N(n330), .A1N(
        outputPortSelect_WEST[0]), .Y(n77) );
  INVX2TS U904 ( .A(n339), .Y(n333) );
  OAI22X1TS U905 ( .A0(n334), .A1(n333), .B0(n192), .B1(n332), .Y(n335) );
  OAI2BB2XLTS U906 ( .B0(n335), .B1(n341), .A0N(n330), .A1N(
        outputPortSelect_WEST[1]), .Y(n76) );
  NAND2X1TS U907 ( .A(n315), .B(n232), .Y(n337) );
  AOI2BB2XLTS U908 ( .B0(n188), .B1(n337), .A0N(n315), .A1N(n336), .Y(n345) );
  NAND2X1TS U909 ( .A(n339), .B(n338), .Y(n340) );
  NOR4XLTS U910 ( .A(n343), .B(n342), .C(n341), .D(n340), .Y(n344) );
  INVX2TS U911 ( .A(n344), .Y(n346) );
  OAI2BB2XLTS U912 ( .B0(n346), .B1(n345), .A0N(outputPortSelect_WEST[3]), 
        .A1N(n330), .Y(n74) );
  AO22XLTS U913 ( .A0(readInBuffer_WEST), .A1(n347), .B0(n327), .B1(
        memRead_WEST), .Y(n73) );
endmodule

