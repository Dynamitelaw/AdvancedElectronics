

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO cacheBank 
  PIN clk 
    ANTENNAPARTIALMETALAREA 12.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 45.584 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.7016 LAYER M3 ; 
    ANTENNAMAXAREACAR 9.73625 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 36.3655 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0470146 LAYER VL ;
  END clk
  PIN reset 
    ANTENNADIFFAREA 0.32 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.14 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.178 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.078 LAYER M3 ; 
    ANTENNAMAXAREACAR 159.385 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 559.415 LAYER M3 ;
    ANTENNAMAXCUTCAR 2.05128 LAYER VL ;
    ANTENNADIFFAREA 0.32 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.72 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 3.168 LAYER MQ ;
    ANTENNAGATEAREA 0.078 LAYER MQ ; 
    ANTENNAMAXAREACAR 168.615 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 600.031 LAYER MQ ;
    ANTENNAMAXCUTCAR 2.05128 LAYER VQ ;
  END reset
  PIN cacheDataIn_A[31] 
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.368 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 40.6667 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 118.262 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 49.8974 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 158.877 LAYER MQ ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ ;
  END cacheDataIn_A[31]
  PIN cacheDataIn_A[30] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.706 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.8202 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 129.897 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 452.21 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 139.128 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 474.979 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 148.359 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 515.595 LAYER MQ ;
  END cacheDataIn_A[30]
  PIN cacheDataIn_A[29] 
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 38.6154 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 110.672 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 47.8462 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 151.287 LAYER MQ ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ ;
  END cacheDataIn_A[29]
  PIN cacheDataIn_A[28] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.566 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.3022 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 126.308 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 438.928 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 135.538 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 461.697 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 144.769 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 502.313 LAYER MQ ;
  END cacheDataIn_A[28]
  PIN cacheDataIn_A[27] 
    ANTENNAPARTIALMETALAREA 3.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.322 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.516 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 68.359 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 220.723 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 77.5897 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 261.338 LAYER MQ ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ ;
  END cacheDataIn_A[27]
  PIN cacheDataIn_A[26] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.746 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.9682 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 130.923 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 456.005 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 140.154 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 478.774 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 149.385 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 519.39 LAYER MQ ;
  END cacheDataIn_A[26]
  PIN cacheDataIn_A[25] 
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.22 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 39.641 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 114.467 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 48.8718 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 155.082 LAYER MQ ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ ;
  END cacheDataIn_A[25]
  PIN cacheDataIn_A[24] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.626 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5242 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 127.846 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 444.621 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 137.077 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 467.39 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 146.308 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 508.005 LAYER MQ ;
  END cacheDataIn_A[24]
  PIN cacheDataIn_A[23] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.806 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.1902 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 132.462 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 461.697 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 141.692 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 484.467 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 150.923 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 525.082 LAYER MQ ;
  END cacheDataIn_A[23]
  PIN cacheDataIn_A[22] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.786 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.1162 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 131.949 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 459.8 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 141.179 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 482.569 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 150.41 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 523.185 LAYER MQ ;
  END cacheDataIn_A[22]
  PIN cacheDataIn_A[21] 
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.368 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 40.6667 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 118.262 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 49.8974 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 158.877 LAYER MQ ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ ;
  END cacheDataIn_A[21]
  PIN cacheDataIn_A[20] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.706 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.8202 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 129.897 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 452.21 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 139.128 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 474.979 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 148.359 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 515.595 LAYER MQ ;
  END cacheDataIn_A[20]
  PIN cacheDataIn_A[19] 
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 38.6154 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 110.672 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 47.8462 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 151.287 LAYER MQ ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ ;
  END cacheDataIn_A[19]
  PIN cacheDataIn_A[18] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 139.128 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 482.569 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 148.359 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 523.185 LAYER MQ ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ ;
  END cacheDataIn_A[18]
  PIN cacheDataIn_A[17] 
    ANTENNAPARTIALMETALAREA 3.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.322 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.516 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 68.359 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 220.723 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 77.5897 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 261.338 LAYER MQ ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ ;
  END cacheDataIn_A[17]
  PIN cacheDataIn_A[16] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.746 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.9682 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 130.923 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 456.005 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 140.154 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 478.774 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 149.385 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 519.39 LAYER MQ ;
  END cacheDataIn_A[16]
  PIN cacheDataIn_A[15] 
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.22 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 39.641 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 114.467 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 48.8718 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 155.082 LAYER MQ ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ ;
  END cacheDataIn_A[15]
  PIN cacheDataIn_A[14] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.61 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.465 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 127.436 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 443.103 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 136.667 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 465.872 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 145.897 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 506.487 LAYER MQ ;
  END cacheDataIn_A[14]
  PIN cacheDataIn_A[13] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.806 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.1902 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 132.462 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 461.697 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 141.692 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 484.467 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 150.923 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 525.082 LAYER MQ ;
  END cacheDataIn_A[13]
  PIN cacheDataIn_A[12] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.77 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.057 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 131.538 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 458.282 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 140.769 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 481.051 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 150 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 521.667 LAYER MQ ;
  END cacheDataIn_A[12]
  PIN cacheDataIn_A[11] 
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.368 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 40.6667 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 118.262 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 49.8974 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 158.877 LAYER MQ ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ ;
  END cacheDataIn_A[11]
  PIN cacheDataIn_A[10] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.69 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.761 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 129.487 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 450.692 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 138.718 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 473.462 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 147.949 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 514.077 LAYER MQ ;
  END cacheDataIn_A[10]
  PIN cacheDataIn_A[9] 
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 38.6154 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 110.672 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 47.8462 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 151.287 LAYER MQ ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ ;
  END cacheDataIn_A[9]
  PIN cacheDataIn_A[8] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.566 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.3022 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 126.308 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 438.928 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 135.538 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 461.697 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 144.769 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 502.313 LAYER MQ ;
  END cacheDataIn_A[8]
  PIN cacheDataIn_A[7] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 127.333 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 446.518 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 136.564 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 469.287 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 145.795 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 509.903 LAYER MQ ;
  END cacheDataIn_A[7]
  PIN cacheDataIn_A[6] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.73 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.909 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 130.513 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 454.487 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 139.744 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 477.256 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 148.974 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 517.872 LAYER MQ ;
  END cacheDataIn_A[6]
  PIN cacheDataIn_A[5] 
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.22 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 39.641 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 114.467 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 48.8718 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 155.082 LAYER MQ ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ ;
  END cacheDataIn_A[5]
  PIN cacheDataIn_A[4] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 127.333 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 446.518 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 136.564 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 469.287 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 145.795 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 509.903 LAYER MQ ;
  END cacheDataIn_A[4]
  PIN cacheDataIn_A[3] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 127.333 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 446.518 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 136.564 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 469.287 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 145.795 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 509.903 LAYER MQ ;
  END cacheDataIn_A[3]
  PIN cacheDataIn_A[2] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.77 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.057 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 131.538 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 458.282 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 140.769 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 481.051 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 150 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 521.667 LAYER MQ ;
  END cacheDataIn_A[2]
  PIN cacheDataIn_A[1] 
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.368 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 40.6667 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 118.262 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 49.8974 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 158.877 LAYER MQ ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ ;
  END cacheDataIn_A[1]
  PIN cacheDataIn_A[0] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.69 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.761 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 129.487 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 450.692 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 138.718 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 473.462 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 147.949 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 514.077 LAYER MQ ;
  END cacheDataIn_A[0]
  PIN cacheAddressIn_A[7] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 127.333 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 446.518 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 136.564 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 469.287 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 145.795 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 509.903 LAYER MQ ;
  END cacheAddressIn_A[7]
  PIN cacheAddressIn_A[6] 
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.368 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 40.6667 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 118.262 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 49.8974 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 158.877 LAYER MQ ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ ;
  END cacheAddressIn_A[6]
  PIN cacheAddressIn_A[5] 
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.884 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 58.1026 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 182.774 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 67.3333 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 223.39 LAYER MQ ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ ;
  END cacheAddressIn_A[5]
  PIN cacheAddressIn_A[4] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 127.333 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 446.518 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 136.564 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 469.287 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 145.795 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 509.903 LAYER MQ ;
  END cacheAddressIn_A[4]
  PIN cacheAddressIn_A[3] 
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.18 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 60.1538 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 190.364 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 69.3846 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 230.979 LAYER MQ ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ ;
  END cacheAddressIn_A[3]
  PIN cacheAddressIn_A[2] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 127.333 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 446.518 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 136.564 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 469.287 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 145.795 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 509.903 LAYER MQ ;
  END cacheAddressIn_A[2]
  PIN cacheAddressIn_A[1] 
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.548 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 76.5641 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 251.082 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 85.7949 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 291.697 LAYER MQ ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ ;
  END cacheAddressIn_A[1]
  PIN cacheAddressIn_A[0] 
    ANTENNAPARTIALMETALAREA 3.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.322 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.064 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 120.667 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 414.262 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 129.897 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 454.877 LAYER MQ ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ ;
  END cacheAddressIn_A[0]
  PIN memWrite_A 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 127.333 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 446.518 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 136.564 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 469.287 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 145.795 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 509.903 LAYER MQ ;
  END memWrite_A
  PIN cacheDataOut_A[31] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_A[31]
  PIN cacheDataOut_A[30] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.726 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.8942 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_A[30]
  PIN cacheDataOut_A[29] 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.37 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_A[29]
  PIN cacheDataOut_A[28] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.4502 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_A[28]
  PIN cacheDataOut_A[27] 
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.85 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.701 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_A[27]
  PIN cacheDataOut_A[26] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.766 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.0422 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_A[26]
  PIN cacheDataOut_A[25] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_A[25]
  PIN cacheDataOut_A[24] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.646 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_A[24]
  PIN cacheDataOut_A[23] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.79 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.131 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_A[23]
  PIN cacheDataOut_A[22] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.806 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.1902 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_A[22]
  PIN cacheDataOut_A[21] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_A[21]
  PIN cacheDataOut_A[20] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.726 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.8942 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_A[20]
  PIN cacheDataOut_A[19] 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.37 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_A[19]
  PIN cacheDataOut_A[18] 
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_A[18]
  PIN cacheDataOut_A[17] 
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.85 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.701 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_A[17]
  PIN cacheDataOut_A[16] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.766 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.0422 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_A[16]
  PIN cacheDataOut_A[15] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_A[15]
  PIN cacheDataOut_A[14] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.646 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_A[14]
  PIN cacheDataOut_A[13] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.774 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.0718 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_A[13]
  PIN cacheDataOut_A[12] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.806 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.1902 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_A[12]
  PIN cacheDataOut_A[11] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_A[11]
  PIN cacheDataOut_A[10] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.726 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.8942 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_A[10]
  PIN cacheDataOut_A[9] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_A[9]
  PIN cacheDataOut_A[8] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.4502 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_A[8]
  PIN cacheDataOut_A[7] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_A[7]
  PIN cacheDataOut_A[6] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.766 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.0422 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_A[6]
  PIN cacheDataOut_A[5] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_A[5]
  PIN cacheDataOut_A[4] 
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.22 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_A[4]
  PIN cacheDataOut_A[3] 
    ANTENNAPARTIALMETALAREA 1.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.178 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.664 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_A[3]
  PIN cacheDataOut_A[2] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.806 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.1902 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_A[2]
  PIN cacheDataOut_A[1] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_A[1]
  PIN cacheDataOut_A[0] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.726 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.8942 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_A[0]
  PIN portA_writtenTo 
  END portA_writtenTo
  PIN cacheDataIn_B[31] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.746 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.9682 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 130.923 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 456.005 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 140.154 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 478.774 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 149.385 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 519.39 LAYER MQ ;
  END cacheDataIn_B[31]
  PIN cacheDataIn_B[30] 
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.22 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 39.641 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 114.467 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 48.8718 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 155.082 LAYER MQ ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ ;
  END cacheDataIn_B[30]
  PIN cacheDataIn_B[29] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.626 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5242 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 127.846 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 444.621 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 137.077 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 467.39 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 146.308 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 508.005 LAYER MQ ;
  END cacheDataIn_B[29]
  PIN cacheDataIn_B[28] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.806 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.1902 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 132.462 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 461.697 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 141.692 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 484.467 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 150.923 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 525.082 LAYER MQ ;
  END cacheDataIn_B[28]
  PIN cacheDataIn_B[27] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.786 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.1162 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 131.949 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 459.8 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 141.179 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 482.569 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 150.41 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 523.185 LAYER MQ ;
  END cacheDataIn_B[27]
  PIN cacheDataIn_B[26] 
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.368 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 40.6667 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 118.262 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 49.8974 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 158.877 LAYER MQ ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ ;
  END cacheDataIn_B[26]
  PIN cacheDataIn_B[25] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.706 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.8202 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 129.897 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 452.21 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 139.128 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 474.979 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 148.359 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 515.595 LAYER MQ ;
  END cacheDataIn_B[25]
  PIN cacheDataIn_B[24] 
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 38.6154 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 110.672 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 47.8462 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 151.287 LAYER MQ ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ ;
  END cacheDataIn_B[24]
  PIN cacheDataIn_B[23] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.566 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.3022 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 126.308 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 438.928 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 135.538 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 461.697 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 144.769 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 502.313 LAYER MQ ;
  END cacheDataIn_B[23]
  PIN cacheDataIn_B[22] 
    ANTENNAPARTIALMETALAREA 3.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.322 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.516 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 68.359 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 220.723 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 77.5897 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 261.338 LAYER MQ ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ ;
  END cacheDataIn_B[22]
  PIN cacheDataIn_B[21] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.746 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.9682 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 130.923 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 456.005 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 140.154 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 478.774 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 149.385 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 519.39 LAYER MQ ;
  END cacheDataIn_B[21]
  PIN cacheDataIn_B[20] 
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.22 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 39.641 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 114.467 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 48.8718 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 155.082 LAYER MQ ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ ;
  END cacheDataIn_B[20]
  PIN cacheDataIn_B[19] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.626 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5242 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 127.846 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 444.621 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 137.077 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 467.39 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 146.308 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 508.005 LAYER MQ ;
  END cacheDataIn_B[19]
  PIN cacheDataIn_B[18] 
    ANTENNAPARTIALMETALAREA 0.98 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.626 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.664 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 122.718 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 421.851 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 131.949 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 462.467 LAYER MQ ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ ;
  END cacheDataIn_B[18]
  PIN cacheDataIn_B[17] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.786 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.1162 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 131.949 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 459.8 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 141.179 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 482.569 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 150.41 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 523.185 LAYER MQ ;
  END cacheDataIn_B[17]
  PIN cacheDataIn_B[16] 
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.368 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 40.6667 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 118.262 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 49.8974 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 158.877 LAYER MQ ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ ;
  END cacheDataIn_B[16]
  PIN cacheDataIn_B[15] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.69 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.761 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 129.487 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 450.692 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 138.718 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 473.462 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 147.949 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 514.077 LAYER MQ ;
  END cacheDataIn_B[15]
  PIN cacheDataIn_B[14] 
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 38.6154 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 110.672 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 47.8462 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 151.287 LAYER MQ ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ ;
  END cacheDataIn_B[14]
  PIN cacheDataIn_B[13] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.566 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.3022 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 126.308 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 438.928 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 135.538 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 461.697 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 144.769 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 502.313 LAYER MQ ;
  END cacheDataIn_B[13]
  PIN cacheDataIn_B[12] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 127.333 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 446.518 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 136.564 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 469.287 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 145.795 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 509.903 LAYER MQ ;
  END cacheDataIn_B[12]
  PIN cacheDataIn_B[11] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.73 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.909 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 130.513 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 454.487 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 139.744 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 477.256 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 148.974 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 517.872 LAYER MQ ;
  END cacheDataIn_B[11]
  PIN cacheDataIn_B[10] 
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.22 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 39.641 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 114.467 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 48.8718 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 155.082 LAYER MQ ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ ;
  END cacheDataIn_B[10]
  PIN cacheDataIn_B[9] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.61 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.465 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 127.436 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 443.103 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 136.667 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 465.872 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 145.897 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 506.487 LAYER MQ ;
  END cacheDataIn_B[9]
  PIN cacheDataIn_B[8] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.806 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.1902 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 132.462 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 461.697 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 141.692 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 484.467 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 150.923 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 525.082 LAYER MQ ;
  END cacheDataIn_B[8]
  PIN cacheDataIn_B[7] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.77 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.057 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 131.538 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 458.282 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 140.769 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 481.051 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 150 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 521.667 LAYER MQ ;
  END cacheDataIn_B[7]
  PIN cacheDataIn_B[6] 
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.368 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 40.6667 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 118.262 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 49.8974 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 158.877 LAYER MQ ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ ;
  END cacheDataIn_B[6]
  PIN cacheDataIn_B[5] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.69 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.761 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 129.487 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 450.692 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 138.718 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 473.462 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 147.949 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 514.077 LAYER MQ ;
  END cacheDataIn_B[5]
  PIN cacheDataIn_B[4] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 127.333 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 446.518 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 136.564 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 469.287 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 145.795 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 509.903 LAYER MQ ;
  END cacheDataIn_B[4]
  PIN cacheDataIn_B[3] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 127.333 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 446.518 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 136.564 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 469.287 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 145.795 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 509.903 LAYER MQ ;
  END cacheDataIn_B[3]
  PIN cacheDataIn_B[2] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 127.333 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 446.518 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 136.564 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 469.287 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 145.795 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 509.903 LAYER MQ ;
  END cacheDataIn_B[2]
  PIN cacheDataIn_B[1] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.73 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.909 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 130.513 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 454.487 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 139.744 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 477.256 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 148.974 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 517.872 LAYER MQ ;
  END cacheDataIn_B[1]
  PIN cacheDataIn_B[0] 
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.22 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 39.641 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 114.467 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 48.8718 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 155.082 LAYER MQ ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ ;
  END cacheDataIn_B[0]
  PIN cacheAddressIn_B[7] 
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.916 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 92.9744 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 311.8 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 102.205 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 352.415 LAYER MQ ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ ;
  END cacheAddressIn_B[7]
  PIN cacheAddressIn_B[6] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 127.333 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 446.518 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 136.564 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 469.287 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 145.795 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 509.903 LAYER MQ ;
  END cacheAddressIn_B[6]
  PIN cacheAddressIn_B[5] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 127.333 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 446.518 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 136.564 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 469.287 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 145.795 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 509.903 LAYER MQ ;
  END cacheAddressIn_B[5]
  PIN cacheAddressIn_B[4] 
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.104 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 73.4872 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 239.697 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 82.7179 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 280.313 LAYER MQ ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ ;
  END cacheAddressIn_B[4]
  PIN cacheAddressIn_B[3] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 127.333 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 446.518 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 136.564 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 469.287 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 145.795 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 509.903 LAYER MQ ;
  END cacheAddressIn_B[3]
  PIN cacheAddressIn_B[2] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 127.333 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 446.518 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 136.564 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 469.287 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 145.795 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 509.903 LAYER MQ ;
  END cacheAddressIn_B[2]
  PIN cacheAddressIn_B[1] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 127.333 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 446.518 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 136.564 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 469.287 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 145.795 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 509.903 LAYER MQ ;
  END cacheAddressIn_B[1]
  PIN cacheAddressIn_B[0] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 127.333 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 446.518 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 136.564 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 469.287 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 145.795 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 509.903 LAYER MQ ;
  END cacheAddressIn_B[0]
  PIN memWrite_B 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.754 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.9978 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2 ; 
    ANTENNAMAXAREACAR 131.128 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 456.764 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAGATEAREA 0.039 LAYER M3 ; 
    ANTENNAMAXAREACAR 140.359 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 479.533 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
    ANTENNAGATEAREA 0.039 LAYER MQ ; 
    ANTENNAMAXAREACAR 149.59 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 520.149 LAYER MQ ;
  END memWrite_B
  PIN cacheDataOut_B[31] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.766 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.0422 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_B[31]
  PIN cacheDataOut_B[30] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_B[30]
  PIN cacheDataOut_B[29] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.646 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_B[29]
  PIN cacheDataOut_B[28] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.79 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.131 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_B[28]
  PIN cacheDataOut_B[27] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.806 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.1902 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_B[27]
  PIN cacheDataOut_B[26] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_B[26]
  PIN cacheDataOut_B[25] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.726 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.8942 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_B[25]
  PIN cacheDataOut_B[24] 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.37 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_B[24]
  PIN cacheDataOut_B[23] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.4502 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_B[23]
  PIN cacheDataOut_B[22] 
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.85 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.701 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_B[22]
  PIN cacheDataOut_B[21] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.766 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.0422 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_B[21]
  PIN cacheDataOut_B[20] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_B[20]
  PIN cacheDataOut_B[19] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.646 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_B[19]
  PIN cacheDataOut_B[18] 
    ANTENNAPARTIALMETALAREA 1.86 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.882 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.664 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_B[18]
  PIN cacheDataOut_B[17] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.806 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.1902 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_B[17]
  PIN cacheDataOut_B[16] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_B[16]
  PIN cacheDataOut_B[15] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.726 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.8942 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_B[15]
  PIN cacheDataOut_B[14] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_B[14]
  PIN cacheDataOut_B[13] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.4502 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_B[13]
  PIN cacheDataOut_B[12] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_B[12]
  PIN cacheDataOut_B[11] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.766 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.0422 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_B[11]
  PIN cacheDataOut_B[10] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_B[10]
  PIN cacheDataOut_B[9] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.646 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_B[9]
  PIN cacheDataOut_B[8] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.774 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.0718 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_B[8]
  PIN cacheDataOut_B[7] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.806 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.1902 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_B[7]
  PIN cacheDataOut_B[6] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_B[6]
  PIN cacheDataOut_B[5] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.726 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.8942 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_B[5]
  PIN cacheDataOut_B[4] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_B[4]
  PIN cacheDataOut_B[3] 
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_B[3]
  PIN cacheDataOut_B[2] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_B[2]
  PIN cacheDataOut_B[1] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.766 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.0422 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_B[1]
  PIN cacheDataOut_B[0] 
    ANTENNADIFFAREA 0.16 LAYER M2 ; 
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2 ;
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNADIFFAREA 0.16 LAYER MQ ; 
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ ;
  END cacheDataOut_B[0]
  PIN portB_writtenTo 
  END portB_writtenTo
END cacheBank

END LIBRARY
