
module outputPortArbiter ( clk, reset, selectBit_NORTH, 
        destinationAddressIn_NORTH, requesterAddressIn_NORTH, readIn_NORTH, 
        writeIn_NORTH, dataIn_NORTH, selectBit_SOUTH, 
        destinationAddressIn_SOUTH, requesterAddressIn_SOUTH, readIn_SOUTH, 
        writeIn_SOUTH, dataIn_SOUTH, selectBit_EAST, destinationAddressIn_EAST, 
        requesterAddressIn_EAST, readIn_EAST, writeIn_EAST, dataIn_EAST, 
        selectBit_WEST, destinationAddressIn_WEST, requesterAddressIn_WEST, 
        readIn_WEST, writeIn_WEST, dataIn_WEST, readReady, 
        readRequesterAddress, cacheDataOut, destinationAddressOut, 
        requesterAddressOut, readOut, writeOut, dataOut );
  input [13:0] destinationAddressIn_NORTH;
  input [5:0] requesterAddressIn_NORTH;
  input [31:0] dataIn_NORTH;
  input [13:0] destinationAddressIn_SOUTH;
  input [5:0] requesterAddressIn_SOUTH;
  input [31:0] dataIn_SOUTH;
  input [13:0] destinationAddressIn_EAST;
  input [5:0] requesterAddressIn_EAST;
  input [31:0] dataIn_EAST;
  input [13:0] destinationAddressIn_WEST;
  input [5:0] requesterAddressIn_WEST;
  input [31:0] dataIn_WEST;
  input [5:0] readRequesterAddress;
  input [31:0] cacheDataOut;
  output [13:0] destinationAddressOut;
  output [5:0] requesterAddressOut;
  output [31:0] dataOut;
  input clk, reset, selectBit_NORTH, readIn_NORTH, writeIn_NORTH,
         selectBit_SOUTH, readIn_SOUTH, writeIn_SOUTH, selectBit_EAST,
         readIn_EAST, writeIn_EAST, selectBit_WEST, readIn_WEST, writeIn_WEST,
         readReady;
  output readOut, writeOut;
  wire   N373, N374, N375, \requesterAddressbuffer[0][5] ,
         \requesterAddressbuffer[0][4] , \requesterAddressbuffer[0][3] ,
         \requesterAddressbuffer[0][2] , \requesterAddressbuffer[0][1] ,
         \requesterAddressbuffer[0][0] , \requesterAddressbuffer[1][5] ,
         \requesterAddressbuffer[1][4] , \requesterAddressbuffer[1][3] ,
         \requesterAddressbuffer[1][2] , \requesterAddressbuffer[1][1] ,
         \requesterAddressbuffer[1][0] , \requesterAddressbuffer[2][5] ,
         \requesterAddressbuffer[2][4] , \requesterAddressbuffer[2][3] ,
         \requesterAddressbuffer[2][2] , \requesterAddressbuffer[2][1] ,
         \requesterAddressbuffer[2][0] , \requesterAddressbuffer[3][5] ,
         \requesterAddressbuffer[3][4] , \requesterAddressbuffer[3][3] ,
         \requesterAddressbuffer[3][2] , \requesterAddressbuffer[3][1] ,
         \requesterAddressbuffer[3][0] , \requesterAddressbuffer[4][5] ,
         \requesterAddressbuffer[4][4] , \requesterAddressbuffer[4][3] ,
         \requesterAddressbuffer[4][2] , \requesterAddressbuffer[4][1] ,
         \requesterAddressbuffer[4][0] , \requesterAddressbuffer[5][5] ,
         \requesterAddressbuffer[5][4] , \requesterAddressbuffer[5][3] ,
         \requesterAddressbuffer[5][2] , \requesterAddressbuffer[5][1] ,
         \requesterAddressbuffer[5][0] , \requesterAddressbuffer[6][5] ,
         \requesterAddressbuffer[6][4] , \requesterAddressbuffer[6][3] ,
         \requesterAddressbuffer[6][2] , \requesterAddressbuffer[6][1] ,
         \requesterAddressbuffer[6][0] , \requesterAddressbuffer[7][5] ,
         \requesterAddressbuffer[7][4] , \requesterAddressbuffer[7][3] ,
         \requesterAddressbuffer[7][2] , \requesterAddressbuffer[7][1] ,
         \requesterAddressbuffer[7][0] , \destinationAddressbuffer[0][13] ,
         \destinationAddressbuffer[0][12] , \destinationAddressbuffer[0][11] ,
         \destinationAddressbuffer[0][10] , \destinationAddressbuffer[0][9] ,
         \destinationAddressbuffer[0][8] , \destinationAddressbuffer[0][7] ,
         \destinationAddressbuffer[0][6] , \destinationAddressbuffer[0][5] ,
         \destinationAddressbuffer[0][4] , \destinationAddressbuffer[0][3] ,
         \destinationAddressbuffer[0][2] , \destinationAddressbuffer[0][1] ,
         \destinationAddressbuffer[0][0] , \destinationAddressbuffer[1][13] ,
         \destinationAddressbuffer[1][12] , \destinationAddressbuffer[1][11] ,
         \destinationAddressbuffer[1][10] , \destinationAddressbuffer[1][9] ,
         \destinationAddressbuffer[1][8] , \destinationAddressbuffer[1][7] ,
         \destinationAddressbuffer[1][6] , \destinationAddressbuffer[1][5] ,
         \destinationAddressbuffer[1][4] , \destinationAddressbuffer[1][3] ,
         \destinationAddressbuffer[1][2] , \destinationAddressbuffer[1][1] ,
         \destinationAddressbuffer[1][0] , \destinationAddressbuffer[2][13] ,
         \destinationAddressbuffer[2][12] , \destinationAddressbuffer[2][11] ,
         \destinationAddressbuffer[2][10] , \destinationAddressbuffer[2][9] ,
         \destinationAddressbuffer[2][8] , \destinationAddressbuffer[2][7] ,
         \destinationAddressbuffer[2][6] , \destinationAddressbuffer[2][5] ,
         \destinationAddressbuffer[2][4] , \destinationAddressbuffer[2][3] ,
         \destinationAddressbuffer[2][2] , \destinationAddressbuffer[2][1] ,
         \destinationAddressbuffer[2][0] , \destinationAddressbuffer[3][13] ,
         \destinationAddressbuffer[3][12] , \destinationAddressbuffer[3][11] ,
         \destinationAddressbuffer[3][10] , \destinationAddressbuffer[3][9] ,
         \destinationAddressbuffer[3][8] , \destinationAddressbuffer[3][7] ,
         \destinationAddressbuffer[3][6] , \destinationAddressbuffer[3][5] ,
         \destinationAddressbuffer[3][4] , \destinationAddressbuffer[3][3] ,
         \destinationAddressbuffer[3][2] , \destinationAddressbuffer[3][1] ,
         \destinationAddressbuffer[3][0] , \destinationAddressbuffer[4][13] ,
         \destinationAddressbuffer[4][12] , \destinationAddressbuffer[4][11] ,
         \destinationAddressbuffer[4][10] , \destinationAddressbuffer[4][9] ,
         \destinationAddressbuffer[4][8] , \destinationAddressbuffer[4][7] ,
         \destinationAddressbuffer[4][6] , \destinationAddressbuffer[4][5] ,
         \destinationAddressbuffer[4][4] , \destinationAddressbuffer[4][3] ,
         \destinationAddressbuffer[4][2] , \destinationAddressbuffer[4][1] ,
         \destinationAddressbuffer[4][0] , \destinationAddressbuffer[5][13] ,
         \destinationAddressbuffer[5][12] , \destinationAddressbuffer[5][11] ,
         \destinationAddressbuffer[5][10] , \destinationAddressbuffer[5][9] ,
         \destinationAddressbuffer[5][8] , \destinationAddressbuffer[5][7] ,
         \destinationAddressbuffer[5][6] , \destinationAddressbuffer[5][5] ,
         \destinationAddressbuffer[5][4] , \destinationAddressbuffer[5][3] ,
         \destinationAddressbuffer[5][2] , \destinationAddressbuffer[5][1] ,
         \destinationAddressbuffer[5][0] , \destinationAddressbuffer[6][13] ,
         \destinationAddressbuffer[6][12] , \destinationAddressbuffer[6][11] ,
         \destinationAddressbuffer[6][10] , \destinationAddressbuffer[6][9] ,
         \destinationAddressbuffer[6][8] , \destinationAddressbuffer[6][7] ,
         \destinationAddressbuffer[6][6] , \destinationAddressbuffer[6][5] ,
         \destinationAddressbuffer[6][4] , \destinationAddressbuffer[6][3] ,
         \destinationAddressbuffer[6][2] , \destinationAddressbuffer[6][1] ,
         \destinationAddressbuffer[6][0] , \destinationAddressbuffer[7][13] ,
         \destinationAddressbuffer[7][12] , \destinationAddressbuffer[7][11] ,
         \destinationAddressbuffer[7][10] , \destinationAddressbuffer[7][9] ,
         \destinationAddressbuffer[7][8] , \destinationAddressbuffer[7][7] ,
         \destinationAddressbuffer[7][6] , \destinationAddressbuffer[7][5] ,
         \destinationAddressbuffer[7][4] , \destinationAddressbuffer[7][3] ,
         \destinationAddressbuffer[7][2] , \destinationAddressbuffer[7][1] ,
         \destinationAddressbuffer[7][0] , \dataoutbuffer[7][31] ,
         \dataoutbuffer[7][30] , \dataoutbuffer[7][29] ,
         \dataoutbuffer[7][28] , \dataoutbuffer[7][27] ,
         \dataoutbuffer[7][26] , \dataoutbuffer[7][25] ,
         \dataoutbuffer[7][24] , \dataoutbuffer[7][23] ,
         \dataoutbuffer[7][22] , \dataoutbuffer[7][21] ,
         \dataoutbuffer[7][20] , \dataoutbuffer[7][19] ,
         \dataoutbuffer[7][18] , \dataoutbuffer[7][17] ,
         \dataoutbuffer[7][16] , \dataoutbuffer[7][15] ,
         \dataoutbuffer[7][14] , \dataoutbuffer[7][13] ,
         \dataoutbuffer[7][12] , \dataoutbuffer[7][11] ,
         \dataoutbuffer[7][10] , \dataoutbuffer[7][9] , \dataoutbuffer[7][8] ,
         \dataoutbuffer[7][7] , \dataoutbuffer[7][6] , \dataoutbuffer[7][5] ,
         \dataoutbuffer[7][4] , \dataoutbuffer[7][3] , \dataoutbuffer[7][2] ,
         \dataoutbuffer[7][1] , \dataoutbuffer[7][0] , \dataoutbuffer[6][31] ,
         \dataoutbuffer[6][30] , \dataoutbuffer[6][29] ,
         \dataoutbuffer[6][28] , \dataoutbuffer[6][27] ,
         \dataoutbuffer[6][26] , \dataoutbuffer[6][25] ,
         \dataoutbuffer[6][24] , \dataoutbuffer[6][23] ,
         \dataoutbuffer[6][22] , \dataoutbuffer[6][21] ,
         \dataoutbuffer[6][20] , \dataoutbuffer[6][19] ,
         \dataoutbuffer[6][18] , \dataoutbuffer[6][17] ,
         \dataoutbuffer[6][16] , \dataoutbuffer[6][15] ,
         \dataoutbuffer[6][14] , \dataoutbuffer[6][13] ,
         \dataoutbuffer[6][12] , \dataoutbuffer[6][11] ,
         \dataoutbuffer[6][10] , \dataoutbuffer[6][9] , \dataoutbuffer[6][8] ,
         \dataoutbuffer[6][7] , \dataoutbuffer[6][6] , \dataoutbuffer[6][5] ,
         \dataoutbuffer[6][4] , \dataoutbuffer[6][3] , \dataoutbuffer[6][2] ,
         \dataoutbuffer[6][1] , \dataoutbuffer[6][0] , \dataoutbuffer[5][31] ,
         \dataoutbuffer[5][30] , \dataoutbuffer[5][29] ,
         \dataoutbuffer[5][28] , \dataoutbuffer[5][27] ,
         \dataoutbuffer[5][26] , \dataoutbuffer[5][25] ,
         \dataoutbuffer[5][24] , \dataoutbuffer[5][23] ,
         \dataoutbuffer[5][22] , \dataoutbuffer[5][21] ,
         \dataoutbuffer[5][20] , \dataoutbuffer[5][19] ,
         \dataoutbuffer[5][18] , \dataoutbuffer[5][17] ,
         \dataoutbuffer[5][16] , \dataoutbuffer[5][15] ,
         \dataoutbuffer[5][14] , \dataoutbuffer[5][13] ,
         \dataoutbuffer[5][12] , \dataoutbuffer[5][11] ,
         \dataoutbuffer[5][10] , \dataoutbuffer[5][9] , \dataoutbuffer[5][8] ,
         \dataoutbuffer[5][7] , \dataoutbuffer[5][6] , \dataoutbuffer[5][5] ,
         \dataoutbuffer[5][4] , \dataoutbuffer[5][3] , \dataoutbuffer[5][2] ,
         \dataoutbuffer[5][1] , \dataoutbuffer[5][0] , \dataoutbuffer[4][31] ,
         \dataoutbuffer[4][30] , \dataoutbuffer[4][29] ,
         \dataoutbuffer[4][28] , \dataoutbuffer[4][27] ,
         \dataoutbuffer[4][26] , \dataoutbuffer[4][25] ,
         \dataoutbuffer[4][24] , \dataoutbuffer[4][23] ,
         \dataoutbuffer[4][22] , \dataoutbuffer[4][21] ,
         \dataoutbuffer[4][20] , \dataoutbuffer[4][19] ,
         \dataoutbuffer[4][18] , \dataoutbuffer[4][17] ,
         \dataoutbuffer[4][16] , \dataoutbuffer[4][15] ,
         \dataoutbuffer[4][14] , \dataoutbuffer[4][13] ,
         \dataoutbuffer[4][12] , \dataoutbuffer[4][11] ,
         \dataoutbuffer[4][10] , \dataoutbuffer[4][9] , \dataoutbuffer[4][8] ,
         \dataoutbuffer[4][7] , \dataoutbuffer[4][6] , \dataoutbuffer[4][5] ,
         \dataoutbuffer[4][4] , \dataoutbuffer[4][3] , \dataoutbuffer[4][2] ,
         \dataoutbuffer[4][1] , \dataoutbuffer[4][0] , \dataoutbuffer[3][31] ,
         \dataoutbuffer[3][30] , \dataoutbuffer[3][29] ,
         \dataoutbuffer[3][28] , \dataoutbuffer[3][27] ,
         \dataoutbuffer[3][26] , \dataoutbuffer[3][25] ,
         \dataoutbuffer[3][24] , \dataoutbuffer[3][23] ,
         \dataoutbuffer[3][22] , \dataoutbuffer[3][21] ,
         \dataoutbuffer[3][20] , \dataoutbuffer[3][19] ,
         \dataoutbuffer[3][18] , \dataoutbuffer[3][17] ,
         \dataoutbuffer[3][16] , \dataoutbuffer[3][15] ,
         \dataoutbuffer[3][14] , \dataoutbuffer[3][13] ,
         \dataoutbuffer[3][12] , \dataoutbuffer[3][11] ,
         \dataoutbuffer[3][10] , \dataoutbuffer[3][9] , \dataoutbuffer[3][8] ,
         \dataoutbuffer[3][7] , \dataoutbuffer[3][6] , \dataoutbuffer[3][5] ,
         \dataoutbuffer[3][4] , \dataoutbuffer[3][3] , \dataoutbuffer[3][2] ,
         \dataoutbuffer[3][1] , \dataoutbuffer[3][0] , \dataoutbuffer[2][31] ,
         \dataoutbuffer[2][30] , \dataoutbuffer[2][29] ,
         \dataoutbuffer[2][28] , \dataoutbuffer[2][27] ,
         \dataoutbuffer[2][26] , \dataoutbuffer[2][25] ,
         \dataoutbuffer[2][24] , \dataoutbuffer[2][23] ,
         \dataoutbuffer[2][22] , \dataoutbuffer[2][21] ,
         \dataoutbuffer[2][20] , \dataoutbuffer[2][19] ,
         \dataoutbuffer[2][18] , \dataoutbuffer[2][17] ,
         \dataoutbuffer[2][16] , \dataoutbuffer[2][15] ,
         \dataoutbuffer[2][14] , \dataoutbuffer[2][13] ,
         \dataoutbuffer[2][12] , \dataoutbuffer[2][11] ,
         \dataoutbuffer[2][10] , \dataoutbuffer[2][9] , \dataoutbuffer[2][8] ,
         \dataoutbuffer[2][7] , \dataoutbuffer[2][6] , \dataoutbuffer[2][5] ,
         \dataoutbuffer[2][4] , \dataoutbuffer[2][3] , \dataoutbuffer[2][2] ,
         \dataoutbuffer[2][1] , \dataoutbuffer[2][0] , \dataoutbuffer[1][31] ,
         \dataoutbuffer[1][30] , \dataoutbuffer[1][29] ,
         \dataoutbuffer[1][28] , \dataoutbuffer[1][27] ,
         \dataoutbuffer[1][26] , \dataoutbuffer[1][25] ,
         \dataoutbuffer[1][24] , \dataoutbuffer[1][23] ,
         \dataoutbuffer[1][22] , \dataoutbuffer[1][21] ,
         \dataoutbuffer[1][20] , \dataoutbuffer[1][19] ,
         \dataoutbuffer[1][18] , \dataoutbuffer[1][17] ,
         \dataoutbuffer[1][16] , \dataoutbuffer[1][15] ,
         \dataoutbuffer[1][14] , \dataoutbuffer[1][13] ,
         \dataoutbuffer[1][12] , \dataoutbuffer[1][11] ,
         \dataoutbuffer[1][10] , \dataoutbuffer[1][9] , \dataoutbuffer[1][8] ,
         \dataoutbuffer[1][7] , \dataoutbuffer[1][6] , \dataoutbuffer[1][5] ,
         \dataoutbuffer[1][4] , \dataoutbuffer[1][3] , \dataoutbuffer[1][2] ,
         \dataoutbuffer[1][1] , \dataoutbuffer[1][0] , \dataoutbuffer[0][31] ,
         \dataoutbuffer[0][30] , \dataoutbuffer[0][29] ,
         \dataoutbuffer[0][28] , \dataoutbuffer[0][27] ,
         \dataoutbuffer[0][26] , \dataoutbuffer[0][25] ,
         \dataoutbuffer[0][24] , \dataoutbuffer[0][23] ,
         \dataoutbuffer[0][22] , \dataoutbuffer[0][21] ,
         \dataoutbuffer[0][20] , \dataoutbuffer[0][19] ,
         \dataoutbuffer[0][18] , \dataoutbuffer[0][17] ,
         \dataoutbuffer[0][16] , \dataoutbuffer[0][15] ,
         \dataoutbuffer[0][14] , \dataoutbuffer[0][13] ,
         \dataoutbuffer[0][12] , \dataoutbuffer[0][11] ,
         \dataoutbuffer[0][10] , \dataoutbuffer[0][9] , \dataoutbuffer[0][8] ,
         \dataoutbuffer[0][7] , \dataoutbuffer[0][6] , \dataoutbuffer[0][5] ,
         \dataoutbuffer[0][4] , \dataoutbuffer[0][3] , \dataoutbuffer[0][2] ,
         \dataoutbuffer[0][1] , \dataoutbuffer[0][0] , empty_reg, N4718, n2397,
         n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
         n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
         n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
         n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
         n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
         n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
         n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
         n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
         n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
         n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
         n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
         n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
         n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
         n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
         n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
         n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997,
         n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007,
         n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
         n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
         n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
         n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
         n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057,
         n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067,
         n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077,
         n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087,
         n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
         n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107,
         n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
         n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329;
  wire   [0:7] writeOutbuffer;
  wire   [0:7] readOutbuffer;
  wire   [2:0] read_reg;

  DFFNSRX1TS full_reg_reg ( .D(N4718), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(
        n5328) );
  DFFNSRX1TS \write_reg_reg[0]  ( .D(n2888), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(N373), .QN(n5327) );
  DFFNSRX1TS \write_reg_reg[2]  ( .D(n2886), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(N375), .QN(n5326) );
  DFFNSRX1TS \read_reg_reg[0]  ( .D(n2889), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(read_reg[0]), .QN(n5325) );
  DFFNSRX1TS \read_reg_reg[1]  ( .D(n2883), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(read_reg[1]), .QN(n5324) );
  DFFNSRX1TS \write_reg_reg[1]  ( .D(n2887), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(N374), .QN(n5323) );
  DFFNSRX1TS \readOutbuffer_reg[6]  ( .D(n2569), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[6]) );
  DFFNSRX1TS \readOutbuffer_reg[4]  ( .D(n2567), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[4]) );
  DFFNSRX1TS \readOutbuffer_reg[3]  ( .D(n2566), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[3]) );
  DFFNSRX1TS \writeOutbuffer_reg[7]  ( .D(n2578), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[7]) );
  DFFNSRX1TS \dataoutbuffer_reg[6][4]  ( .D(n2638), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][18]  ( .D(n2624), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[6][18] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][25]  ( .D(n2617), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[6][25] ) );
  DFFNSRX1TS \writeOutbuffer_reg[6]  ( .D(n2577), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[6]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][4]  ( .D(n2544), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][7]  ( .D(n2541), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][8]  ( .D(n2540), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][11]  ( .D(n2537), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][11] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][13]  ( .D(n2535), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][13] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][3]  ( .D(n2703), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][14]  ( .D(n2692), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[4][14] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][15]  ( .D(n2691), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[4][15] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][17]  ( .D(n2689), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[4][17] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][9]  ( .D(n2511), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][13]  ( .D(n2507), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][13] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][7]  ( .D(n2731), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][7] ) );
  DFFNSRX1TS \writeOutbuffer_reg[3]  ( .D(n2574), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[3]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][7]  ( .D(n2499), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][10]  ( .D(n2496), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][13]  ( .D(n2493), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][13] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][0]  ( .D(n2770), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][2]  ( .D(n2768), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][6]  ( .D(n2764), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][6] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][16]  ( .D(n2754), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[2][16] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][22]  ( .D(n2748), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[2][22] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][24]  ( .D(n2746), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[2][24] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][31]  ( .D(n2739), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[2][31] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][6]  ( .D(n2486), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][8]  ( .D(n2484), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][10]  ( .D(n2482), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][12]  ( .D(n2480), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][12] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][0]  ( .D(n2802), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][0]  ( .D(n2834), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][1]  ( .D(n2833), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][2]  ( .D(n2832), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][5]  ( .D(n2829), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][9]  ( .D(n2825), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][9] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][20]  ( .D(n2814), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[0][20] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][23]  ( .D(n2811), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[0][23] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][27]  ( .D(n2807), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[0][27] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][28]  ( .D(n2806), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[0][28] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][7]  ( .D(n2457), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][9]  ( .D(n2455), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][11]  ( .D(n2453), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][11] ) );
  DFFNSRX1TS \readOutbuffer_reg[7]  ( .D(n2570), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[7]) );
  DFFNSRX1TS \readOutbuffer_reg[2]  ( .D(n2565), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[2]) );
  DFFNSRX1TS \writeOutbuffer_reg[2]  ( .D(n2573), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[2]) );
  DFFNSRX1TS \readOutbuffer_reg[5]  ( .D(n2568), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[5]) );
  DFFNSRX1TS \readOutbuffer_reg[1]  ( .D(n2564), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[1]) );
  DFFNSRX1TS \readOutbuffer_reg[0]  ( .D(n2563), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[0]) );
  DFFNSRX1TS \writeOutbuffer_reg[4]  ( .D(n2575), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[4]) );
  DFFNSRX1TS \requesterAddressbuffer_reg[7][0]  ( .D(n2882), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[7][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[7][1]  ( .D(n2881), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[7][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[7][3]  ( .D(n2879), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[7][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][0]  ( .D(n2610), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][1]  ( .D(n2609), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][2]  ( .D(n2608), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][3]  ( .D(n2607), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][4]  ( .D(n2606), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][5]  ( .D(n2605), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][6]  ( .D(n2604), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][6] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][7]  ( .D(n2603), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][7] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][8]  ( .D(n2602), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][8] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][9]  ( .D(n2601), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][9] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][10]  ( .D(n2600), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[7][10] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][11]  ( .D(n2599), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[7][11] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][12]  ( .D(n2598), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[7][12] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][13]  ( .D(n2597), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[7][13] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][14]  ( .D(n2596), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[7][14] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][15]  ( .D(n2595), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[7][15] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][16]  ( .D(n2594), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[7][16] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][17]  ( .D(n2593), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[7][17] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][18]  ( .D(n2592), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[7][18] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][19]  ( .D(n2591), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[7][19] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][20]  ( .D(n2590), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[7][20] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][21]  ( .D(n2589), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[7][21] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][22]  ( .D(n2588), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[7][22] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][23]  ( .D(n2587), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[7][23] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][24]  ( .D(n2586), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[7][24] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][25]  ( .D(n2585), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[7][25] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][26]  ( .D(n2584), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[7][26] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][27]  ( .D(n2583), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[7][27] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][28]  ( .D(n2582), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[7][28] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][29]  ( .D(n2581), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[7][29] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][30]  ( .D(n2580), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[7][30] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][31]  ( .D(n2579), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[7][31] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][1]  ( .D(n2561), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][2]  ( .D(n2560), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][3]  ( .D(n2559), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][5]  ( .D(n2557), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][6]  ( .D(n2556), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][7]  ( .D(n2555), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][8]  ( .D(n2554), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][10]  ( .D(n2552), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][11]  ( .D(n2551), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][11] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][12]  ( .D(n2550), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][12] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][13]  ( .D(n2549), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][13] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][0]  ( .D(n2642), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][2]  ( .D(n2640), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][3]  ( .D(n2639), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][5]  ( .D(n2637), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][7]  ( .D(n2635), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][7] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][8]  ( .D(n2634), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][8] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][9]  ( .D(n2633), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][9] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][11]  ( .D(n2631), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[6][11] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][14]  ( .D(n2628), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[6][14] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][15]  ( .D(n2627), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[6][15] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][16]  ( .D(n2626), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[6][16] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][17]  ( .D(n2625), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[6][17] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][19]  ( .D(n2623), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[6][19] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][22]  ( .D(n2620), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[6][22] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][24]  ( .D(n2618), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[6][24] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][26]  ( .D(n2616), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[6][26] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][27]  ( .D(n2615), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[6][27] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][28]  ( .D(n2614), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[6][28] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][30]  ( .D(n2612), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[6][30] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][31]  ( .D(n2611), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[6][31] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[5][0]  ( .D(n2870), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[5][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[5][1]  ( .D(n2869), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[5][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[5][2]  ( .D(n2868), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[5][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[5][3]  ( .D(n2867), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[5][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[5][4]  ( .D(n2866), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[5][4] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[5][5]  ( .D(n2865), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[5][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][0]  ( .D(n2674), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][2]  ( .D(n2672), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][3]  ( .D(n2671), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][4]  ( .D(n2670), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][5]  ( .D(n2669), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][6]  ( .D(n2668), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][6] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][7]  ( .D(n2667), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][7] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][8]  ( .D(n2666), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][8] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][9]  ( .D(n2665), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][9] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][10]  ( .D(n2664), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[5][10] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][12]  ( .D(n2662), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[5][12] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][13]  ( .D(n2661), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[5][13] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][14]  ( .D(n2660), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[5][14] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][17]  ( .D(n2657), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[5][17] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][18]  ( .D(n2656), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[5][18] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][19]  ( .D(n2655), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[5][19] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][20]  ( .D(n2654), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[5][20] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][21]  ( .D(n2653), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[5][21] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][22]  ( .D(n2652), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[5][22] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][23]  ( .D(n2651), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[5][23] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][24]  ( .D(n2650), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[5][24] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][25]  ( .D(n2649), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[5][25] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][26]  ( .D(n2648), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[5][26] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][27]  ( .D(n2647), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[5][27] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][28]  ( .D(n2646), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[5][28] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][29]  ( .D(n2645), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[5][29] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][30]  ( .D(n2644), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[5][30] ) );
  DFFNSRX1TS \writeOutbuffer_reg[5]  ( .D(n2576), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[5]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][0]  ( .D(n2534), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][1]  ( .D(n2533), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][2]  ( .D(n2532), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][3]  ( .D(n2531), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][4]  ( .D(n2530), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][5]  ( .D(n2529), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][6]  ( .D(n2528), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][7]  ( .D(n2527), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][8]  ( .D(n2526), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][9]  ( .D(n2525), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][10]  ( .D(n2524), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][11]  ( .D(n2523), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][11] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][12]  ( .D(n2522), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][12] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][13]  ( .D(n2521), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][13] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[4][4]  ( .D(n2860), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[4][4] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[4][5]  ( .D(n2859), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[4][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][0]  ( .D(n2706), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][1]  ( .D(n2705), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][6]  ( .D(n2700), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][6] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][8]  ( .D(n2698), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][8] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][10]  ( .D(n2696), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[4][10] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][11]  ( .D(n2695), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[4][11] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][12]  ( .D(n2694), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[4][12] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][16]  ( .D(n2690), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[4][16] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][19]  ( .D(n2687), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[4][19] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][20]  ( .D(n2686), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[4][20] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][21]  ( .D(n2685), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[4][21] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][22]  ( .D(n2684), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[4][22] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][29]  ( .D(n2677), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[4][29] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][31]  ( .D(n2675), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[4][31] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][2]  ( .D(n2736), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][4]  ( .D(n2734), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][5]  ( .D(n2733), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][13]  ( .D(n2725), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[3][13] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][15]  ( .D(n2723), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[3][15] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][18]  ( .D(n2720), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[3][18] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][20]  ( .D(n2718), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[3][20] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][23]  ( .D(n2715), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[3][23] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][25]  ( .D(n2713), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[3][25] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][2]  ( .D(n2504), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][8]  ( .D(n2498), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][9]  ( .D(n2497), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][12]  ( .D(n2494), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][12] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[2][2]  ( .D(n2850), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[2][3]  ( .D(n2849), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[2][5]  ( .D(n2847), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][1]  ( .D(n2769), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][10]  ( .D(n2760), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[2][10] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][27]  ( .D(n2743), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[2][27] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][0]  ( .D(n2492), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][1]  ( .D(n2491), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][3]  ( .D(n2489), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][4]  ( .D(n2488), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][5]  ( .D(n2487), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][7]  ( .D(n2485), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][9]  ( .D(n2483), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][11]  ( .D(n2481), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][11] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[1][0]  ( .D(n2846), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[1][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[1][1]  ( .D(n2845), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[1][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[1][2]  ( .D(n2844), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[1][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[1][3]  ( .D(n2843), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[1][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[1][4]  ( .D(n2842), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[1][4] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[1][5]  ( .D(n2841), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[1][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][1]  ( .D(n2801), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][3]  ( .D(n2799), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][4]  ( .D(n2798), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][6]  ( .D(n2796), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][6] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][7]  ( .D(n2795), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][7] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][9]  ( .D(n2793), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][9] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][11]  ( .D(n2791), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[1][11] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][12]  ( .D(n2790), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[1][12] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][13]  ( .D(n2789), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[1][13] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][14]  ( .D(n2788), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[1][14] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][15]  ( .D(n2787), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[1][15] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][16]  ( .D(n2786), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[1][16] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][17]  ( .D(n2785), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[1][17] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][18]  ( .D(n2784), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[1][18] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][21]  ( .D(n2781), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[1][21] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][23]  ( .D(n2779), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[1][23] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][24]  ( .D(n2778), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[1][24] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][25]  ( .D(n2777), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[1][25] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][26]  ( .D(n2776), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[1][26] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][28]  ( .D(n2774), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[1][28] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][29]  ( .D(n2773), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[1][29] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][30]  ( .D(n2772), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[1][30] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][31]  ( .D(n2771), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[1][31] ) );
  DFFNSRX1TS \writeOutbuffer_reg[1]  ( .D(n2572), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[1]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][0]  ( .D(n2478), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][1]  ( .D(n2477), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][2]  ( .D(n2476), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][3]  ( .D(n2475), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][4]  ( .D(n2474), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][5]  ( .D(n2473), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][6]  ( .D(n2472), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][7]  ( .D(n2471), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][8]  ( .D(n2470), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][9]  ( .D(n2469), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][10]  ( .D(n2468), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][11]  ( .D(n2467), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][11] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][12]  ( .D(n2466), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][12] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][13]  ( .D(n2465), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][13] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[0][0]  ( .D(n2840), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[0][1]  ( .D(n2839), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[0][2]  ( .D(n2838), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[0][4]  ( .D(n2836), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][4] ) );
  DFFNSRX1TS \writeOutbuffer_reg[0]  ( .D(n2571), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[0]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][0]  ( .D(n2464), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][4]  ( .D(n2460), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][6]  ( .D(n2458), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][10]  ( .D(n2454), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][13]  ( .D(n2451), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][13] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[7][2]  ( .D(n2880), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[7][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[7][4]  ( .D(n2878), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[7][4] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[7][5]  ( .D(n2877), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[7][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][0]  ( .D(n2562), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][4]  ( .D(n2558), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][9]  ( .D(n2553), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][9] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[6][0]  ( .D(n2876), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[6][1]  ( .D(n2875), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[6][2]  ( .D(n2874), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[6][3]  ( .D(n2873), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[6][4]  ( .D(n2872), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][4] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[6][5]  ( .D(n2871), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][1]  ( .D(n2641), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][6]  ( .D(n2636), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][6] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][10]  ( .D(n2632), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[6][10] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][12]  ( .D(n2630), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[6][12] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][13]  ( .D(n2629), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[6][13] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][20]  ( .D(n2622), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[6][20] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][21]  ( .D(n2621), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[6][21] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][23]  ( .D(n2619), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[6][23] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][29]  ( .D(n2613), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[6][29] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][0]  ( .D(n2548), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][1]  ( .D(n2547), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][2]  ( .D(n2546), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][3]  ( .D(n2545), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][5]  ( .D(n2543), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][6]  ( .D(n2542), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][9]  ( .D(n2539), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][10]  ( .D(n2538), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][12]  ( .D(n2536), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][12] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][1]  ( .D(n2673), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][11]  ( .D(n2663), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[5][11] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][15]  ( .D(n2659), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[5][15] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][16]  ( .D(n2658), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[5][16] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][31]  ( .D(n2643), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[5][31] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[4][0]  ( .D(n2864), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[4][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[4][1]  ( .D(n2863), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[4][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[4][2]  ( .D(n2862), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[4][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[4][3]  ( .D(n2861), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[4][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][2]  ( .D(n2704), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][4]  ( .D(n2702), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][5]  ( .D(n2701), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][7]  ( .D(n2699), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][7] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][9]  ( .D(n2697), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][9] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][13]  ( .D(n2693), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[4][13] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][18]  ( .D(n2688), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[4][18] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][23]  ( .D(n2683), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[4][23] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][24]  ( .D(n2682), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[4][24] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][25]  ( .D(n2681), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[4][25] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][26]  ( .D(n2680), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[4][26] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][27]  ( .D(n2679), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[4][27] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][28]  ( .D(n2678), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[4][28] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][30]  ( .D(n2676), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[4][30] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][0]  ( .D(n2520), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][1]  ( .D(n2519), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][2]  ( .D(n2518), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][3]  ( .D(n2517), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][4]  ( .D(n2516), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][5]  ( .D(n2515), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][6]  ( .D(n2514), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][7]  ( .D(n2513), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][8]  ( .D(n2512), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][10]  ( .D(n2510), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][11]  ( .D(n2509), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][11] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][12]  ( .D(n2508), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][12] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[3][0]  ( .D(n2858), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[3][1]  ( .D(n2857), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[3][2]  ( .D(n2856), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[3][3]  ( .D(n2855), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[3][4]  ( .D(n2854), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][4] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[3][5]  ( .D(n2853), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][0]  ( .D(n2738), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][1]  ( .D(n2737), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][3]  ( .D(n2735), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][6]  ( .D(n2732), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][6] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][8]  ( .D(n2730), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][8] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][9]  ( .D(n2729), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][9] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][10]  ( .D(n2728), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[3][10] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][11]  ( .D(n2727), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[3][11] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][12]  ( .D(n2726), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[3][12] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][14]  ( .D(n2724), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[3][14] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][16]  ( .D(n2722), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[3][16] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][17]  ( .D(n2721), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[3][17] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][19]  ( .D(n2719), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[3][19] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][21]  ( .D(n2717), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[3][21] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][22]  ( .D(n2716), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[3][22] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][24]  ( .D(n2714), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[3][24] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][26]  ( .D(n2712), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[3][26] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][27]  ( .D(n2711), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[3][27] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][28]  ( .D(n2710), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[3][28] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][29]  ( .D(n2709), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[3][29] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][30]  ( .D(n2708), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[3][30] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][31]  ( .D(n2707), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[3][31] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][0]  ( .D(n2506), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][1]  ( .D(n2505), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][3]  ( .D(n2503), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][4]  ( .D(n2502), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][5]  ( .D(n2501), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][6]  ( .D(n2500), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][11]  ( .D(n2495), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][11] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[2][0]  ( .D(n2852), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[2][1]  ( .D(n2851), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[2][4]  ( .D(n2848), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][3]  ( .D(n2767), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][4]  ( .D(n2766), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][5]  ( .D(n2765), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][7]  ( .D(n2763), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][7] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][8]  ( .D(n2762), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][8] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][9]  ( .D(n2761), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][9] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][11]  ( .D(n2759), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[2][11] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][12]  ( .D(n2758), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[2][12] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][13]  ( .D(n2757), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[2][13] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][14]  ( .D(n2756), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[2][14] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][15]  ( .D(n2755), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[2][15] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][17]  ( .D(n2753), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[2][17] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][18]  ( .D(n2752), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[2][18] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][19]  ( .D(n2751), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[2][19] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][20]  ( .D(n2750), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[2][20] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][21]  ( .D(n2749), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[2][21] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][23]  ( .D(n2747), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[2][23] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][25]  ( .D(n2745), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[2][25] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][26]  ( .D(n2744), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[2][26] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][28]  ( .D(n2742), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[2][28] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][29]  ( .D(n2741), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[2][29] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][30]  ( .D(n2740), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[2][30] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][2]  ( .D(n2490), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][13]  ( .D(n2479), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][13] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][2]  ( .D(n2800), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][5]  ( .D(n2797), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][8]  ( .D(n2794), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][8] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][10]  ( .D(n2792), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[1][10] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][19]  ( .D(n2783), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[1][19] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][20]  ( .D(n2782), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[1][20] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][22]  ( .D(n2780), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[1][22] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][27]  ( .D(n2775), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[1][27] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[0][3]  ( .D(n2837), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[0][5]  ( .D(n2835), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][3]  ( .D(n2831), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][4]  ( .D(n2830), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][6]  ( .D(n2828), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][6] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][7]  ( .D(n2827), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][7] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][8]  ( .D(n2826), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][8] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][10]  ( .D(n2824), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[0][10] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][11]  ( .D(n2823), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[0][11] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][12]  ( .D(n2822), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[0][12] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][13]  ( .D(n2821), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[0][13] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][14]  ( .D(n2820), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[0][14] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][15]  ( .D(n2819), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[0][15] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][16]  ( .D(n2818), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[0][16] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][17]  ( .D(n2817), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[0][17] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][18]  ( .D(n2816), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[0][18] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][19]  ( .D(n2815), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[0][19] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][21]  ( .D(n2813), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[0][21] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][22]  ( .D(n2812), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[0][22] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][24]  ( .D(n2810), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[0][24] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][25]  ( .D(n2809), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[0][25] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][26]  ( .D(n2808), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[0][26] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][29]  ( .D(n2805), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[0][29] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][30]  ( .D(n2804), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[0][30] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][31]  ( .D(n2803), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataoutbuffer[0][31] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][1]  ( .D(n2463), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][2]  ( .D(n2462), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][3]  ( .D(n2461), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][5]  ( .D(n2459), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][8]  ( .D(n2456), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][12]  ( .D(n2452), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][12] ) );
  DFFNSRX1TS empty_reg_reg ( .D(n2885), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        empty_reg) );
  DFFNSRX1TS writeOut_reg ( .D(n2449), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        writeOut) );
  DFFNSRX1TS \requesterAddressOut_reg[0]  ( .D(n2434), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[0]) );
  DFFNSRX1TS \requesterAddressOut_reg[3]  ( .D(n2431), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[3]) );
  DFFNSRX1TS readOut_reg ( .D(n2450), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        readOut) );
  DFFNSRX1TS \destinationAddressOut_reg[6]  ( .D(n2448), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[6]) );
  DFFNSRX1TS \destinationAddressOut_reg[7]  ( .D(n2447), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[7]) );
  DFFNSRX1TS \destinationAddressOut_reg[8]  ( .D(n2446), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[8]) );
  DFFNSRX1TS \destinationAddressOut_reg[9]  ( .D(n2445), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[9]) );
  DFFNSRX1TS \destinationAddressOut_reg[10]  ( .D(n2444), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[10]) );
  DFFNSRX1TS \destinationAddressOut_reg[11]  ( .D(n2443), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[11]) );
  DFFNSRX1TS \destinationAddressOut_reg[12]  ( .D(n2442), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[12]) );
  DFFNSRX1TS \destinationAddressOut_reg[13]  ( .D(n2441), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[13]) );
  DFFNSRX1TS \destinationAddressOut_reg[0]  ( .D(n2440), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[0]) );
  DFFNSRX1TS \destinationAddressOut_reg[1]  ( .D(n2439), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[1]) );
  DFFNSRX1TS \destinationAddressOut_reg[2]  ( .D(n2438), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[2]) );
  DFFNSRX1TS \destinationAddressOut_reg[3]  ( .D(n2437), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[3]) );
  DFFNSRX1TS \destinationAddressOut_reg[4]  ( .D(n2436), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[4]) );
  DFFNSRX1TS \destinationAddressOut_reg[5]  ( .D(n2435), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[5]) );
  DFFNSRX1TS \requesterAddressOut_reg[1]  ( .D(n2433), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[1]) );
  DFFNSRX1TS \requesterAddressOut_reg[2]  ( .D(n2432), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[2]) );
  DFFNSRX1TS \requesterAddressOut_reg[4]  ( .D(n2430), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[4]) );
  DFFNSRX1TS \requesterAddressOut_reg[5]  ( .D(n2429), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[5]) );
  DFFNSRX1TS \dataOut_reg[0]  ( .D(n2428), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[0]) );
  DFFNSRX1TS \dataOut_reg[1]  ( .D(n2427), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[1]) );
  DFFNSRX1TS \dataOut_reg[2]  ( .D(n2426), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[2]) );
  DFFNSRX1TS \dataOut_reg[3]  ( .D(n2425), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[3]) );
  DFFNSRX1TS \dataOut_reg[4]  ( .D(n2424), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[4]) );
  DFFNSRX1TS \dataOut_reg[5]  ( .D(n2423), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[5]) );
  DFFNSRX1TS \dataOut_reg[6]  ( .D(n2422), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[6]) );
  DFFNSRX1TS \dataOut_reg[7]  ( .D(n2421), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[7]) );
  DFFNSRX1TS \dataOut_reg[8]  ( .D(n2420), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[8]) );
  DFFNSRX1TS \dataOut_reg[9]  ( .D(n2419), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[9]) );
  DFFNSRX1TS \dataOut_reg[10]  ( .D(n2418), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[10]) );
  DFFNSRX1TS \dataOut_reg[11]  ( .D(n2417), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[11]) );
  DFFNSRX1TS \dataOut_reg[12]  ( .D(n2416), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[12]) );
  DFFNSRX1TS \dataOut_reg[13]  ( .D(n2415), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[13]) );
  DFFNSRX1TS \dataOut_reg[14]  ( .D(n2414), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[14]) );
  DFFNSRX1TS \dataOut_reg[15]  ( .D(n2413), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[15]) );
  DFFNSRX1TS \dataOut_reg[16]  ( .D(n2412), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[16]) );
  DFFNSRX1TS \dataOut_reg[17]  ( .D(n2411), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[17]) );
  DFFNSRX1TS \dataOut_reg[18]  ( .D(n2410), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[18]) );
  DFFNSRX1TS \dataOut_reg[19]  ( .D(n2409), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[19]) );
  DFFNSRX1TS \dataOut_reg[20]  ( .D(n2408), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[20]) );
  DFFNSRX1TS \dataOut_reg[21]  ( .D(n2407), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[21]) );
  DFFNSRX1TS \dataOut_reg[22]  ( .D(n2406), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[22]) );
  DFFNSRX1TS \dataOut_reg[23]  ( .D(n2405), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[23]) );
  DFFNSRX1TS \dataOut_reg[24]  ( .D(n2404), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[24]) );
  DFFNSRX1TS \dataOut_reg[25]  ( .D(n2403), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[25]) );
  DFFNSRX1TS \dataOut_reg[26]  ( .D(n2402), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[26]) );
  DFFNSRX1TS \dataOut_reg[27]  ( .D(n2401), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[27]) );
  DFFNSRX1TS \dataOut_reg[28]  ( .D(n2400), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[28]) );
  DFFNSRX1TS \dataOut_reg[29]  ( .D(n2399), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[29]) );
  DFFNSRX1TS \dataOut_reg[30]  ( .D(n2398), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[30]) );
  DFFNSRX1TS \dataOut_reg[31]  ( .D(n2397), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[31]) );
  DFFNSRX1TS \read_reg_reg[2]  ( .D(n2884), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(read_reg[2]), .QN(n5329) );
  NOR2BX2TS U2896 ( .AN(n4496), .B(n4495), .Y(n4674) );
  CMPR32X2TS U2897 ( .A(n4267), .B(N374), .C(n4266), .CO(n4262), .S(n4275) );
  XOR2X1TS U2898 ( .A(N375), .B(n2939), .Y(n3089) );
  CMPR32X2TS U2899 ( .A(read_reg[1]), .B(n5323), .C(n4246), .CO(n4245), .S(
        n4280) );
  CMPR32X2TS U2900 ( .A(n4249), .B(N374), .C(n2938), .CO(n2939), .S(n3317) );
  NAND2X1TS U2901 ( .A(N374), .B(n2946), .Y(n2944) );
  NOR2XLTS U2902 ( .A(n2900), .B(n2945), .Y(n2946) );
  INVX2TS U2903 ( .A(n2946), .Y(n3315) );
  INVX2TS U2904 ( .A(n3085), .Y(n4532) );
  NOR2XLTS U2905 ( .A(n3089), .B(n2902), .Y(n3380) );
  AND2X2TS U2906 ( .A(n3089), .B(n2901), .Y(n3608) );
  BUFX3TS U2907 ( .A(n4932), .Y(n5318) );
  NOR2XLTS U2908 ( .A(n3315), .B(N374), .Y(n4484) );
  OAI21XLTS U2909 ( .A0(n3708), .A1(n3614), .B0(n4491), .Y(n4488) );
  NOR2X1TS U2910 ( .A(n4480), .B(n4477), .Y(n4607) );
  NOR2X2TS U2911 ( .A(n4477), .B(n4474), .Y(n4613) );
  OAI21XLTS U2912 ( .A0(n2904), .A1(n2898), .B0(n5327), .Y(n3109) );
  CLKINVX3TS U2913 ( .A(n4278), .Y(n2890) );
  OR2X1TS U2914 ( .A(n4484), .B(n3386), .Y(n3875) );
  OR2X1TS U2915 ( .A(n4484), .B(n3617), .Y(n4077) );
  OR2X1TS U2916 ( .A(n4463), .B(n3320), .Y(n3968) );
  OR2X1TS U2917 ( .A(n4462), .B(n3320), .Y(n3969) );
  NAND2X1TS U2918 ( .A(n3615), .B(n2897), .Y(n4277) );
  AND2X2TS U2919 ( .A(n4513), .B(n4519), .Y(n2952) );
  NOR2X2TS U2920 ( .A(n4508), .B(n4504), .Y(n4696) );
  NOR2X2TS U2921 ( .A(n4501), .B(n4508), .Y(n4687) );
  INVX3TS U2922 ( .A(n4482), .Y(n4612) );
  NAND2BX1TS U2923 ( .AN(n4524), .B(n4526), .Y(n3386) );
  NOR2X2TS U2924 ( .A(n4502), .B(n2998), .Y(n4703) );
  INVX3TS U2925 ( .A(n4537), .Y(n4787) );
  OAI21X1TS U2926 ( .A0(n3877), .A1(n2993), .B0(n4518), .Y(n2956) );
  NAND2BX1TS U2927 ( .AN(n4469), .B(n4471), .Y(n3320) );
  INVX3TS U2928 ( .A(n4518), .Y(n4728) );
  INVX3TS U2929 ( .A(n4511), .Y(n4701) );
  NOR2X4TS U2930 ( .A(n4495), .B(n4492), .Y(n4672) );
  NAND2BX1TS U2931 ( .AN(n4488), .B(n4489), .Y(n3617) );
  INVX3TS U2932 ( .A(n4500), .Y(n4671) );
  OAI21X1TS U2933 ( .A0(n3877), .A1(n3708), .B0(n4500), .Y(n4495) );
  OAI21X1TS U2934 ( .A0(n3876), .A1(n3614), .B0(n4473), .Y(n4469) );
  NAND2BX1TS U2935 ( .AN(n3084), .B(n3091), .Y(n4531) );
  NOR2X1TS U2936 ( .A(n2996), .B(n4506), .Y(n2995) );
  AOI31X1TS U2937 ( .A0(n3383), .A1(n3619), .A2(n3618), .B0(n3382), .Y(n4526)
         );
  AOI31X1TS U2938 ( .A0(n3091), .A1(n3619), .A2(n4502), .B0(n3084), .Y(n3085)
         );
  OAI21X1TS U2939 ( .A0(n3381), .A1(n4512), .B0(n2947), .Y(n2948) );
  AOI31X1TS U2940 ( .A0(n3091), .A1(n4503), .A2(n3619), .B0(n3092), .Y(n4496)
         );
  AOI31X1TS U2941 ( .A0(n3612), .A1(n3619), .A2(n3618), .B0(n3611), .Y(n4489)
         );
  NOR2X1TS U2942 ( .A(n4512), .B(n3610), .Y(n3110) );
  INVX1TS U2943 ( .A(n3610), .Y(n3612) );
  NOR3X1TS U2944 ( .A(n3318), .B(n3619), .C(n3610), .Y(n3319) );
  INVX1TS U2945 ( .A(n3088), .Y(n2994) );
  INVX1TS U2946 ( .A(n4522), .Y(n3382) );
  INVX1TS U2947 ( .A(n4486), .Y(n3611) );
  INVX1TS U2948 ( .A(n4501), .Y(n4509) );
  NAND3X1TS U2949 ( .A(n3106), .B(n3317), .C(n3608), .Y(n4475) );
  NAND3X1TS U2950 ( .A(n3317), .B(n3380), .C(n3106), .Y(n2947) );
  NAND3X1TS U2951 ( .A(n3380), .B(n3607), .C(n3106), .Y(n4530) );
  NAND3X1TS U2952 ( .A(n3607), .B(n3106), .C(n3608), .Y(n4493) );
  NAND3X1TS U2953 ( .A(n3317), .B(n3609), .C(n3380), .Y(n4501) );
  NAND3X1TS U2954 ( .A(n3607), .B(n3609), .C(n3380), .Y(n4522) );
  NAND3X1TS U2955 ( .A(n3317), .B(n3609), .C(n3608), .Y(n4467) );
  NAND3X1TS U2956 ( .A(N374), .B(n2946), .C(n4503), .Y(n4462) );
  INVX1TS U2957 ( .A(n3107), .Y(n4514) );
  NOR2X4TS U2958 ( .A(n3615), .B(n3231), .Y(n3232) );
  NOR2X1TS U2959 ( .A(n3619), .B(n3083), .Y(n3107) );
  INVX1TS U2960 ( .A(n3083), .Y(n3091) );
  INVX1TS U2961 ( .A(n2996), .Y(n3231) );
  INVX1TS U2962 ( .A(n3609), .Y(n3106) );
  NOR2X4TS U2963 ( .A(n4273), .B(n4821), .Y(n2908) );
  NOR2X4TS U2964 ( .A(n4273), .B(n4798), .Y(n2922) );
  NAND2X2TS U2965 ( .A(n5328), .B(n4809), .Y(n3615) );
  NOR3X1TS U2966 ( .A(N375), .B(n5323), .C(n3614), .Y(n2996) );
  NOR2X1TS U2967 ( .A(n5323), .B(n3316), .Y(n2943) );
  CLKBUFX3TS U2968 ( .A(n5249), .Y(n5295) );
  CLKBUFX3TS U2969 ( .A(n4875), .Y(n2891) );
  CLKBUFX3TS U2970 ( .A(n4802), .Y(n2892) );
  CLKBUFX3TS U2971 ( .A(n5311), .Y(n2893) );
  CLKBUFX3TS U2972 ( .A(n4803), .Y(n2894) );
  CLKBUFX3TS U2973 ( .A(n4884), .Y(n2895) );
  NOR3X1TS U2974 ( .A(n2899), .B(n2904), .C(n2898), .Y(n2941) );
  NOR2X1TS U2975 ( .A(n2901), .B(n2903), .Y(n2940) );
  INVX1TS U2976 ( .A(n2904), .Y(n2942) );
  INVX1TS U2977 ( .A(n2899), .Y(n2900) );
  OAI21X1TS U2978 ( .A0(n3614), .A1(n3384), .B0(n4528), .Y(n4524) );
  NAND4BXLTS U2979 ( .AN(n2898), .B(n2940), .C(n2900), .D(n2904), .Y(n4795) );
  NAND4XLTS U2980 ( .A(n2898), .B(n2940), .C(n2900), .D(n2942), .Y(n4798) );
  NAND4BXLTS U2981 ( .AN(n2898), .B(n2899), .C(n2940), .D(n2942), .Y(n4815) );
  NAND3XLTS U2982 ( .A(n2903), .B(n2941), .C(n2902), .Y(n4816) );
  NAND3BXLTS U2983 ( .AN(n2903), .B(n2901), .C(n2941), .Y(n4821) );
  NAND2X1TS U2984 ( .A(n2994), .B(n2903), .Y(n3381) );
  AND3X1TS U2985 ( .A(n3316), .B(n3315), .C(n3614), .Y(n3613) );
  NOR3XLTS U2986 ( .A(n2956), .B(n4517), .C(n4512), .Y(n3029) );
  NAND2X1TS U2987 ( .A(n3108), .B(n4480), .Y(n3111) );
  NOR2BX1TS U2988 ( .AN(n4475), .B(n3110), .Y(n3108) );
  AO22XLTS U2989 ( .A0(n2927), .A1(n5304), .B0(n2928), .B1(n5280), .Y(n2935)
         );
  NAND4XLTS U2990 ( .A(n4815), .B(n4795), .C(n4798), .D(n4821), .Y(n2911) );
  AO22XLTS U2991 ( .A0(n2909), .A1(n5280), .B0(n2910), .B1(n5290), .Y(n2920)
         );
  OR2X2TS U2992 ( .A(n4483), .B(n3386), .Y(n4228) );
  OR2X2TS U2993 ( .A(n4483), .B(n3617), .Y(n4243) );
  INVX2TS U2994 ( .A(n4243), .Y(n4644) );
  INVX2TS U2995 ( .A(n3158), .Y(n5085) );
  OAI21X1TS U2996 ( .A0(n3877), .A1(n3384), .B0(n4537), .Y(n4535) );
  INVX2TS U2997 ( .A(n3381), .Y(n3383) );
  NAND3XLTS U2998 ( .A(n3619), .B(n4522), .C(n3618), .Y(n4521) );
  NAND3X1TS U2999 ( .A(n3609), .B(n3608), .C(n3607), .Y(n4486) );
  NAND3XLTS U3000 ( .A(n3619), .B(n4486), .C(n3618), .Y(n4485) );
  INVX2TS U3001 ( .A(n2947), .Y(n4517) );
  NOR2BX1TS U3002 ( .AN(n4467), .B(n3319), .Y(n4471) );
  INVX2TS U3003 ( .A(n2955), .Y(n5217) );
  INVX2TS U3004 ( .A(n3700), .Y(n4788) );
  INVX2TS U3005 ( .A(n3243), .Y(n5188) );
  INVX2TS U3006 ( .A(n3060), .Y(n5074) );
  INVX2TS U3007 ( .A(n3065), .Y(n5075) );
  INVX2TS U3008 ( .A(n3526), .Y(n5033) );
  INVX2TS U3009 ( .A(n4782), .Y(n3704) );
  INVX2TS U3010 ( .A(n4790), .Y(n3699) );
  INVX2TS U3011 ( .A(n3141), .Y(n5308) );
  INVX2TS U3012 ( .A(n3136), .Y(n5306) );
  INVX2TS U3013 ( .A(n3042), .Y(n5145) );
  INVX2TS U3014 ( .A(n3272), .Y(n5044) );
  INVX2TS U3015 ( .A(n3495), .Y(n5001) );
  INVX2TS U3016 ( .A(n3537), .Y(n4730) );
  INVX2TS U3017 ( .A(n2952), .Y(n3538) );
  INVX2TS U3018 ( .A(n3202), .Y(n5055) );
  OR2X2TS U3019 ( .A(n4503), .B(n2998), .Y(n3567) );
  INVX2TS U3020 ( .A(n3197), .Y(n5054) );
  OR2X2TS U3021 ( .A(n4495), .B(n4498), .Y(n3807) );
  INVX2TS U3022 ( .A(n3358), .Y(n5123) );
  INVX2TS U3023 ( .A(n3353), .Y(n5124) );
  INVX2TS U3024 ( .A(n3445), .Y(n5012) );
  INVX2TS U3025 ( .A(n3446), .Y(n5011) );
  INVX2TS U3026 ( .A(n3807), .Y(n4673) );
  CLKBUFX2TS U3027 ( .A(n4607), .Y(n4615) );
  INVX2TS U3028 ( .A(n3168), .Y(n5023) );
  INVX2TS U3029 ( .A(n4076), .Y(n4616) );
  INVX2TS U3030 ( .A(n4614), .Y(n4071) );
  INVX2TS U3031 ( .A(n4613), .Y(n4072) );
  NAND2BXLTS U3032 ( .AN(n3092), .B(n3091), .Y(n4498) );
  INVX2TS U3033 ( .A(n3110), .Y(n4474) );
  INVX2TS U3034 ( .A(n4465), .Y(n4796) );
  OAI21X1TS U3035 ( .A0(n3877), .A1(n3876), .B0(n4482), .Y(n4477) );
  XOR2XLTS U3036 ( .A(n4264), .B(n4263), .Y(n4276) );
  CLKAND2X2TS U3037 ( .A(n4261), .B(n4259), .Y(n4265) );
  NOR2XLTS U3038 ( .A(n2896), .B(n3615), .Y(n4284) );
  AOI21X1TS U3039 ( .A0(n4502), .A1(n2944), .B0(n4463), .Y(n3088) );
  ADDFX1TS U3040 ( .A(n2899), .B(n2904), .CI(n2903), .CO(n4249), .S(n4247) );
  NAND2X1TS U3041 ( .A(n2903), .B(n3088), .Y(n3610) );
  ADDFX1TS U3042 ( .A(n2901), .B(n2898), .CI(n4247), .CO(n4248), .S(n4259) );
  AOI211XLTS U3043 ( .A0(n4256), .A1(n4255), .B0(n4254), .C0(n4253), .Y(n4257)
         );
  NOR3XLTS U3044 ( .A(n4280), .B(n4282), .C(n4279), .Y(n4254) );
  INVX2TS U3045 ( .A(n3875), .Y(n4761) );
  INVX2TS U3046 ( .A(n4077), .Y(n4645) );
  CLKBUFX2TS U3047 ( .A(n4128), .Y(n4641) );
  INVX2TS U3048 ( .A(n3698), .Y(n4789) );
  INVX2TS U3049 ( .A(n4228), .Y(n4759) );
  CLKBUFX2TS U3050 ( .A(n4744), .Y(n4757) );
  INVX2TS U3051 ( .A(n3533), .Y(n4731) );
  INVX2TS U3052 ( .A(n3567), .Y(n4702) );
  INVX2TS U3053 ( .A(n3969), .Y(n4586) );
  INVX2TS U3054 ( .A(n3968), .Y(n4584) );
  CLKBUFX2TS U3055 ( .A(n4579), .Y(n4318) );
  CLKAND2X2TS U3056 ( .A(n4261), .B(n4260), .Y(n4266) );
  NAND3XLTS U3057 ( .A(n5321), .B(n5320), .C(n5319), .Y(n2397) );
  NAND3XLTS U3058 ( .A(n5303), .B(n5302), .C(n5301), .Y(n2398) );
  NAND4XLTS U3059 ( .A(n5289), .B(n5288), .C(n5287), .D(n5286), .Y(n2399) );
  NAND3XLTS U3060 ( .A(n5279), .B(n5278), .C(n5277), .Y(n2400) );
  NAND3XLTS U3061 ( .A(n5269), .B(n5268), .C(n5267), .Y(n2401) );
  NAND4XLTS U3062 ( .A(n5258), .B(n5257), .C(n5256), .D(n5255), .Y(n2402) );
  NAND3XLTS U3063 ( .A(n5248), .B(n5247), .C(n5246), .Y(n2403) );
  NAND3XLTS U3064 ( .A(n5237), .B(n5236), .C(n5235), .Y(n2404) );
  NAND3XLTS U3065 ( .A(n5226), .B(n5225), .C(n5224), .Y(n2405) );
  NAND3XLTS U3066 ( .A(n5216), .B(n5215), .C(n5214), .Y(n2406) );
  NAND4XLTS U3067 ( .A(n5206), .B(n5205), .C(n5204), .D(n5203), .Y(n2407) );
  NAND3XLTS U3068 ( .A(n5197), .B(n5196), .C(n5195), .Y(n2408) );
  NAND3XLTS U3069 ( .A(n5186), .B(n5185), .C(n5184), .Y(n2409) );
  NAND3XLTS U3070 ( .A(n5175), .B(n5174), .C(n5173), .Y(n2410) );
  NAND3XLTS U3071 ( .A(n5165), .B(n5164), .C(n5163), .Y(n2411) );
  NAND3XLTS U3072 ( .A(n5155), .B(n5154), .C(n5153), .Y(n2412) );
  NAND3XLTS U3073 ( .A(n5144), .B(n5143), .C(n5142), .Y(n2413) );
  NAND3XLTS U3074 ( .A(n5133), .B(n5132), .C(n5131), .Y(n2414) );
  NAND4XLTS U3075 ( .A(n5122), .B(n5121), .C(n5120), .D(n5119), .Y(n2415) );
  NAND4XLTS U3076 ( .A(n5113), .B(n5112), .C(n5111), .D(n5110), .Y(n2416) );
  NAND4XLTS U3077 ( .A(n5104), .B(n5103), .C(n5102), .D(n5101), .Y(n2417) );
  NAND3XLTS U3078 ( .A(n5095), .B(n5094), .C(n5093), .Y(n2418) );
  NAND3XLTS U3079 ( .A(n5084), .B(n5083), .C(n5082), .Y(n2419) );
  NAND4XLTS U3080 ( .A(n5073), .B(n5072), .C(n5071), .D(n5070), .Y(n2420) );
  NAND3XLTS U3081 ( .A(n5064), .B(n5063), .C(n5062), .Y(n2421) );
  NAND3XLTS U3082 ( .A(n5053), .B(n5052), .C(n5051), .Y(n2422) );
  NAND3XLTS U3083 ( .A(n5042), .B(n5041), .C(n5040), .Y(n2423) );
  NAND3XLTS U3084 ( .A(n5032), .B(n5031), .C(n5030), .Y(n2424) );
  NAND3XLTS U3085 ( .A(n5021), .B(n5020), .C(n5019), .Y(n2425) );
  NAND3XLTS U3086 ( .A(n5010), .B(n5009), .C(n5008), .Y(n2426) );
  NAND3XLTS U3087 ( .A(n5000), .B(n4999), .C(n4998), .Y(n2427) );
  NAND3XLTS U3088 ( .A(n4989), .B(n4988), .C(n4987), .Y(n2428) );
  NAND4XLTS U3089 ( .A(n4979), .B(n4978), .C(n4977), .D(n4976), .Y(n2429) );
  NAND4XLTS U3090 ( .A(n4970), .B(n4969), .C(n4968), .D(n4967), .Y(n2430) );
  NAND4XLTS U3091 ( .A(n4961), .B(n4960), .C(n4959), .D(n4958), .Y(n2432) );
  NAND4XLTS U3092 ( .A(n4952), .B(n4951), .C(n4950), .D(n4949), .Y(n2433) );
  NAND4XLTS U3093 ( .A(n4943), .B(n4942), .C(n4941), .D(n4976), .Y(n2435) );
  NAND4XLTS U3094 ( .A(n4935), .B(n4934), .C(n4933), .D(n4967), .Y(n2436) );
  NAND4XLTS U3095 ( .A(n4926), .B(n4925), .C(n4924), .D(n4923), .Y(n2437) );
  NAND4XLTS U3096 ( .A(n4917), .B(n4916), .C(n4915), .D(n4958), .Y(n2438) );
  NAND4XLTS U3097 ( .A(n4909), .B(n4908), .C(n4907), .D(n4949), .Y(n2439) );
  NAND4XLTS U3098 ( .A(n4901), .B(n4900), .C(n4899), .D(n4898), .Y(n2440) );
  NAND3XLTS U3099 ( .A(n4892), .B(n4891), .C(n4890), .Y(n2441) );
  NAND3XLTS U3100 ( .A(n4883), .B(n4882), .C(n4881), .Y(n2442) );
  NAND3XLTS U3101 ( .A(n4874), .B(n4873), .C(n4872), .Y(n2443) );
  NAND3XLTS U3102 ( .A(n4866), .B(n4865), .C(n4864), .Y(n2444) );
  NAND3XLTS U3103 ( .A(n4858), .B(n4857), .C(n4856), .Y(n2445) );
  NAND3XLTS U3104 ( .A(n4850), .B(n4849), .C(n4848), .Y(n2446) );
  NAND3XLTS U3105 ( .A(n4842), .B(n4841), .C(n4840), .Y(n2447) );
  NAND3XLTS U3106 ( .A(n4834), .B(n4833), .C(n4832), .Y(n2448) );
  OAI31X1TS U3107 ( .A0(empty_reg), .A1(n4808), .A2(n4807), .B0(n2897), .Y(
        n4810) );
  OAI211XLTS U3108 ( .A0(n5305), .A1(n2925), .B0(n2937), .C0(n4923), .Y(n2431)
         );
  AOI211XLTS U3109 ( .A0(n2926), .A1(n2908), .B0(n2935), .C0(n2934), .Y(n2937)
         );
  AO22XLTS U3110 ( .A0(n5318), .A1(requesterAddressOut[3]), .B0(n2890), .B1(
        n2933), .Y(n2934) );
  OAI211XLTS U3111 ( .A0(n5291), .A1(n2906), .B0(n2923), .C0(n4898), .Y(n2434)
         );
  AOI211XLTS U3112 ( .A0(n2907), .A1(n2908), .B0(n2920), .C0(n2919), .Y(n2923)
         );
  OAI31X1TS U3113 ( .A0(empty_reg), .A1(n4824), .A2(n4823), .B0(n4822), .Y(
        n4826) );
  OAI211XLTS U3114 ( .A0(n3704), .A1(n3036), .B0(n3177), .C0(n3176), .Y(n2452)
         );
  OAI211XLTS U3115 ( .A0(n3704), .A1(n4235), .B0(n3183), .C0(n3182), .Y(n2456)
         );
  NAND4XLTS U3116 ( .A(n4794), .B(n4793), .C(n4792), .D(n4791), .Y(n2459) );
  NAND4XLTS U3117 ( .A(n4781), .B(n4780), .C(n4779), .D(n4778), .Y(n2461) );
  NAND4XLTS U3118 ( .A(n4777), .B(n4776), .C(n4775), .D(n4774), .Y(n2462) );
  NAND4XLTS U3119 ( .A(n4773), .B(n4772), .C(n4771), .D(n4770), .Y(n2463) );
  OAI211XLTS U3120 ( .A0(n3699), .A1(n5306), .B0(n3655), .C0(n3654), .Y(n2803)
         );
  OAI211XLTS U3121 ( .A0(n3698), .A1(n5292), .B0(n3694), .C0(n3693), .Y(n2804)
         );
  OAI211XLTS U3122 ( .A0(n3704), .A1(n4171), .B0(n3703), .C0(n3702), .Y(n2805)
         );
  OAI211XLTS U3123 ( .A0(n3699), .A1(n4060), .B0(n3652), .C0(n3651), .Y(n2808)
         );
  OAI211XLTS U3124 ( .A0(n3700), .A1(n4183), .B0(n3600), .C0(n3599), .Y(n2809)
         );
  OAI211XLTS U3125 ( .A0(n3698), .A1(n3150), .B0(n3646), .C0(n3645), .Y(n2810)
         );
  OAI211XLTS U3126 ( .A0(n3700), .A1(n4223), .B0(n3667), .C0(n3666), .Y(n2812)
         );
  OAI211XLTS U3127 ( .A0(n3699), .A1(n4039), .B0(n3594), .C0(n3593), .Y(n2813)
         );
  OAI211XLTS U3128 ( .A0(n3698), .A1(n5176), .B0(n3673), .C0(n3672), .Y(n2815)
         );
  OAI211XLTS U3129 ( .A0(n3704), .A1(n4205), .B0(n3603), .C0(n3602), .Y(n2816)
         );
  OAI211XLTS U3130 ( .A0(n3699), .A1(n5156), .B0(n3214), .C0(n3213), .Y(n2817)
         );
  OAI211XLTS U3131 ( .A0(n3704), .A1(n5145), .B0(n3188), .C0(n3187), .Y(n2818)
         );
  OAI211XLTS U3132 ( .A0(n3699), .A1(n3346), .B0(n3591), .C0(n3590), .Y(n2819)
         );
  OAI211XLTS U3133 ( .A0(n3699), .A1(n5123), .B0(n3658), .C0(n3657), .Y(n2820)
         );
  OAI211XLTS U3134 ( .A0(n3699), .A1(n2966), .B0(n3649), .C0(n3648), .Y(n2821)
         );
  OAI211XLTS U3135 ( .A0(n3699), .A1(n4044), .B0(n3588), .C0(n3587), .Y(n2822)
         );
  OAI211XLTS U3136 ( .A0(n3699), .A1(n4029), .B0(n3597), .C0(n3596), .Y(n2823)
         );
  OAI211XLTS U3137 ( .A0(n3699), .A1(n4022), .B0(n3585), .C0(n3584), .Y(n2824)
         );
  OAI211XLTS U3138 ( .A0(n3704), .A1(n4166), .B0(n3181), .C0(n3180), .Y(n2826)
         );
  OAI211XLTS U3139 ( .A0(n3699), .A1(n5054), .B0(n3205), .C0(n3204), .Y(n2827)
         );
  OAI211XLTS U3140 ( .A0(n3698), .A1(n5043), .B0(n3697), .C0(n3696), .Y(n2828)
         );
  OAI211XLTS U3141 ( .A0(n3700), .A1(n4136), .B0(n3685), .C0(n3684), .Y(n2830)
         );
  OAI211XLTS U3142 ( .A0(n3700), .A1(n3985), .B0(n3688), .C0(n3687), .Y(n2831)
         );
  NAND4XLTS U3143 ( .A(n4458), .B(n4457), .C(n4456), .D(n4792), .Y(n2835) );
  NAND4XLTS U3144 ( .A(n4451), .B(n4450), .C(n4449), .D(n4779), .Y(n2837) );
  OAI211XLTS U3145 ( .A0(n3299), .A1(n4229), .B0(n3843), .C0(n3842), .Y(n2775)
         );
  OAI211XLTS U3146 ( .A0(n4227), .A1(n4240), .B0(n4226), .C0(n4225), .Y(n2780)
         );
  OAI211XLTS U3147 ( .A0(n5188), .A1(n4240), .B0(n4232), .C0(n4231), .Y(n2782)
         );
  OAI211XLTS U3148 ( .A0(n5177), .A1(n4240), .B0(n3867), .C0(n3866), .Y(n2783)
         );
  OAI211XLTS U3149 ( .A0(n3157), .A1(n4229), .B0(n4160), .C0(n4159), .Y(n2792)
         );
  OAI211XLTS U3150 ( .A0(n4170), .A1(n4229), .B0(n4169), .C0(n4168), .Y(n2794)
         );
  OAI211XLTS U3151 ( .A0(n4141), .A1(n4229), .B0(n3837), .C0(n3836), .Y(n2797)
         );
  OAI211XLTS U3152 ( .A0(n5001), .A1(n4240), .B0(n3858), .C0(n3857), .Y(n2800)
         );
  OAI211XLTS U3153 ( .A0(n3538), .A1(n3893), .B0(n3175), .C0(n3174), .Y(n2479)
         );
  NAND4XLTS U3154 ( .A(n4719), .B(n4718), .C(n4717), .D(n4716), .Y(n2490) );
  OAI211XLTS U3155 ( .A0(n3537), .A1(n5292), .B0(n3464), .C0(n3463), .Y(n2740)
         );
  OAI211XLTS U3156 ( .A0(n3538), .A1(n3127), .B0(n3135), .C0(n3134), .Y(n2741)
         );
  OAI211XLTS U3157 ( .A0(n3542), .A1(n5270), .B0(n3522), .C0(n3521), .Y(n2742)
         );
  OAI211XLTS U3158 ( .A0(n3533), .A1(n4089), .B0(n3504), .C0(n3503), .Y(n2744)
         );
  OAI211XLTS U3159 ( .A0(n3542), .A1(n5239), .B0(n3541), .C0(n3540), .Y(n2745)
         );
  OAI211XLTS U3160 ( .A0(n3533), .A1(n4215), .B0(n2961), .C0(n2960), .Y(n2747)
         );
  OAI211XLTS U3161 ( .A0(n3542), .A1(n4043), .B0(n3516), .C0(n3515), .Y(n2749)
         );
  OAI211XLTS U3162 ( .A0(n3537), .A1(n5187), .B0(n3473), .C0(n3472), .Y(n2750)
         );
  OAI211XLTS U3163 ( .A0(n3537), .A1(n5176), .B0(n3470), .C0(n3469), .Y(n2751)
         );
  OAI211XLTS U3164 ( .A0(n3537), .A1(n5166), .B0(n3476), .C0(n3475), .Y(n2752)
         );
  OAI211XLTS U3165 ( .A0(n3537), .A1(n4207), .B0(n3467), .C0(n3466), .Y(n2753)
         );
  OAI211XLTS U3166 ( .A0(n3537), .A1(n5134), .B0(n3501), .C0(n3500), .Y(n2755)
         );
  OAI211XLTS U3167 ( .A0(n3542), .A1(n5124), .B0(n3525), .C0(n3524), .Y(n2756)
         );
  OAI211XLTS U3168 ( .A0(n3537), .A1(n2963), .B0(n2971), .C0(n2970), .Y(n2757)
         );
  OAI211XLTS U3169 ( .A0(n3542), .A1(n4162), .B0(n3510), .C0(n3509), .Y(n2758)
         );
  OAI211XLTS U3170 ( .A0(n3533), .A1(n4102), .B0(n3479), .C0(n3478), .Y(n2759)
         );
  OAI211XLTS U3171 ( .A0(n3542), .A1(n5074), .B0(n3068), .C0(n3067), .Y(n2761)
         );
  OAI211XLTS U3172 ( .A0(n3542), .A1(n4166), .B0(n3059), .C0(n3058), .Y(n2762)
         );
  OAI211XLTS U3173 ( .A0(n3537), .A1(n5055), .B0(n3455), .C0(n3454), .Y(n2763)
         );
  OAI211XLTS U3174 ( .A0(n3542), .A1(n5033), .B0(n3536), .C0(n3535), .Y(n2765)
         );
  OAI211XLTS U3175 ( .A0(n3538), .A1(n5022), .B0(n3171), .C0(n3170), .Y(n2766)
         );
  OAI211XLTS U3176 ( .A0(n3542), .A1(n5011), .B0(n3513), .C0(n3512), .Y(n2767)
         );
  NAND4XLTS U3177 ( .A(n4416), .B(n4415), .C(n4414), .D(n4725), .Y(n2848) );
  NAND4XLTS U3178 ( .A(n4407), .B(n4406), .C(n4405), .D(n4713), .Y(n2851) );
  NAND4XLTS U3179 ( .A(n4404), .B(n4403), .C(n4402), .D(n4709), .Y(n2852) );
  OAI211XLTS U3180 ( .A0(n3574), .A1(n3074), .B0(n3196), .C0(n3195), .Y(n2495)
         );
  OAI211XLTS U3181 ( .A0(n3567), .A1(n4244), .B0(n3007), .C0(n3006), .Y(n2500)
         );
  NAND4XLTS U3182 ( .A(n4707), .B(n4706), .C(n4705), .D(n4704), .Y(n2501) );
  NAND4XLTS U3183 ( .A(n4700), .B(n4699), .C(n4698), .D(n4697), .Y(n2502) );
  NAND4XLTS U3184 ( .A(n4695), .B(n4694), .C(n4693), .D(n4692), .Y(n2503) );
  NAND4XLTS U3185 ( .A(n4686), .B(n4685), .C(n4684), .D(n4683), .Y(n2505) );
  NAND4XLTS U3186 ( .A(n4682), .B(n4681), .C(n4680), .D(n4679), .Y(n2506) );
  OAI211XLTS U3187 ( .A0(n3579), .A1(n5306), .B0(n3573), .C0(n3572), .Y(n2707)
         );
  OAI211XLTS U3188 ( .A0(n3575), .A1(n5293), .B0(n3557), .C0(n3556), .Y(n2708)
         );
  OAI211XLTS U3189 ( .A0(n3574), .A1(n4175), .B0(n3452), .C0(n3451), .Y(n2709)
         );
  OAI211XLTS U3190 ( .A0(n3574), .A1(n3951), .B0(n3404), .C0(n3403), .Y(n2710)
         );
  OAI211XLTS U3191 ( .A0(n3575), .A1(n5259), .B0(n3304), .C0(n3303), .Y(n2711)
         );
  OAI211XLTS U3192 ( .A0(n3574), .A1(n4089), .B0(n3435), .C0(n3434), .Y(n2712)
         );
  OAI211XLTS U3193 ( .A0(n3574), .A1(n4179), .B0(n3242), .C0(n3241), .Y(n2714)
         );
  OAI211XLTS U3194 ( .A0(n3567), .A1(n5207), .B0(n3566), .C0(n3565), .Y(n2716)
         );
  OAI211XLTS U3195 ( .A0(n3575), .A1(n4043), .B0(n3295), .C0(n3294), .Y(n2717)
         );
  OAI211XLTS U3196 ( .A0(n3575), .A1(n5177), .B0(n3267), .C0(n3266), .Y(n2719)
         );
  OAI211XLTS U3197 ( .A0(n3574), .A1(n4206), .B0(n3258), .C0(n3257), .Y(n2721)
         );
  OAI211XLTS U3198 ( .A0(n3575), .A1(n5145), .B0(n3548), .C0(n3547), .Y(n2722)
         );
  OAI211XLTS U3199 ( .A0(n3574), .A1(n3357), .B0(n3441), .C0(n3440), .Y(n2724)
         );
  OAI211XLTS U3200 ( .A0(n3575), .A1(n4162), .B0(n3285), .C0(n3284), .Y(n2726)
         );
  OAI211XLTS U3201 ( .A0(n3567), .A1(n3365), .B0(n3554), .C0(n3553), .Y(n2727)
         );
  OAI211XLTS U3202 ( .A0(n3575), .A1(n5085), .B0(n3255), .C0(n3254), .Y(n2728)
         );
  OAI211XLTS U3203 ( .A0(n3574), .A1(n3064), .B0(n3417), .C0(n3416), .Y(n2729)
         );
  OAI211XLTS U3204 ( .A0(n3575), .A1(n4166), .B0(n3551), .C0(n3550), .Y(n2730)
         );
  OAI211XLTS U3205 ( .A0(n3574), .A1(n4018), .B0(n3276), .C0(n3275), .Y(n2732)
         );
  OAI211XLTS U3206 ( .A0(n3574), .A1(n3985), .B0(n3449), .C0(n3448), .Y(n2735)
         );
  OAI211XLTS U3207 ( .A0(n3574), .A1(n4084), .B0(n3426), .C0(n3425), .Y(n2737)
         );
  OAI211XLTS U3208 ( .A0(n3574), .A1(n4118), .B0(n3423), .C0(n3422), .Y(n2738)
         );
  NAND4XLTS U3209 ( .A(n4401), .B(n4400), .C(n4399), .D(n4705), .Y(n2853) );
  NAND4XLTS U3210 ( .A(n4398), .B(n4397), .C(n4396), .D(n4698), .Y(n2854) );
  NAND4XLTS U3211 ( .A(n4395), .B(n4394), .C(n4393), .D(n4693), .Y(n2855) );
  NAND4XLTS U3212 ( .A(n4392), .B(n4391), .C(n4390), .D(n4689), .Y(n2856) );
  NAND4XLTS U3213 ( .A(n4389), .B(n4388), .C(n4387), .D(n4684), .Y(n2857) );
  NAND4XLTS U3214 ( .A(n4386), .B(n4385), .C(n4384), .D(n4680), .Y(n2858) );
  OAI211XLTS U3215 ( .A0(n3807), .A1(n4189), .B0(n3099), .C0(n3098), .Y(n2508)
         );
  OAI211XLTS U3216 ( .A0(n3831), .A1(n3074), .B0(n3224), .C0(n3223), .Y(n2509)
         );
  OAI211XLTS U3217 ( .A0(n3807), .A1(n4195), .B0(n3101), .C0(n3100), .Y(n2510)
         );
  OAI211XLTS U3218 ( .A0(n3827), .A1(n4235), .B0(n3222), .C0(n3221), .Y(n2512)
         );
  OAI211XLTS U3219 ( .A0(n3807), .A1(n4192), .B0(n3095), .C0(n3094), .Y(n2513)
         );
  OAI211XLTS U3220 ( .A0(n3807), .A1(n4244), .B0(n3097), .C0(n3096), .Y(n2514)
         );
  NAND4XLTS U3221 ( .A(n4678), .B(n4677), .C(n4676), .D(n4675), .Y(n2515) );
  NAND4XLTS U3222 ( .A(n4670), .B(n4669), .C(n4668), .D(n4667), .Y(n2516) );
  NAND4XLTS U3223 ( .A(n4665), .B(n4664), .C(n4663), .D(n4662), .Y(n2517) );
  NAND4XLTS U3224 ( .A(n4661), .B(n4660), .C(n4659), .D(n4658), .Y(n2518) );
  NAND4XLTS U3225 ( .A(n4657), .B(n4656), .C(n4655), .D(n4654), .Y(n2519) );
  NAND4XLTS U3226 ( .A(n4653), .B(n4652), .C(n4651), .D(n4650), .Y(n2520) );
  OAI211XLTS U3227 ( .A0(n3831), .A1(n4198), .B0(n3813), .C0(n3812), .Y(n2676)
         );
  OAI211XLTS U3228 ( .A0(n3826), .A1(n3947), .B0(n3764), .C0(n3763), .Y(n2678)
         );
  OAI211XLTS U3229 ( .A0(n3831), .A1(n3299), .B0(n3819), .C0(n3818), .Y(n2679)
         );
  OAI211XLTS U3230 ( .A0(n3831), .A1(n4089), .B0(n3830), .C0(n3829), .Y(n2680)
         );
  OAI211XLTS U3231 ( .A0(n3807), .A1(n3236), .B0(n3788), .C0(n3787), .Y(n2681)
         );
  OAI211XLTS U3232 ( .A0(n3831), .A1(n4179), .B0(n3810), .C0(n3809), .Y(n2682)
         );
  OAI211XLTS U3233 ( .A0(n3807), .A1(n2958), .B0(n3797), .C0(n3796), .Y(n2683)
         );
  OAI211XLTS U3234 ( .A0(n3826), .A1(n3409), .B0(n3773), .C0(n3772), .Y(n2688)
         );
  OAI211XLTS U3235 ( .A0(n3831), .A1(n4113), .B0(n3718), .C0(n3717), .Y(n2693)
         );
  OAI211XLTS U3236 ( .A0(n3831), .A1(n3064), .B0(n3721), .C0(n3720), .Y(n2697)
         );
  OAI211XLTS U3237 ( .A0(n3826), .A1(n5054), .B0(n3724), .C0(n3723), .Y(n2699)
         );
  OAI211XLTS U3238 ( .A0(n3807), .A1(n3529), .B0(n3758), .C0(n3757), .Y(n2701)
         );
  OAI211XLTS U3239 ( .A0(n3831), .A1(n4136), .B0(n3816), .C0(n3815), .Y(n2702)
         );
  OAI211XLTS U3240 ( .A0(n3831), .A1(n4132), .B0(n3825), .C0(n3824), .Y(n2704)
         );
  NAND4XLTS U3241 ( .A(n4376), .B(n4375), .C(n4374), .D(n4663), .Y(n2861) );
  NAND4XLTS U3242 ( .A(n4373), .B(n4372), .C(n4371), .D(n4659), .Y(n2862) );
  NAND4XLTS U3243 ( .A(n4370), .B(n4369), .C(n4368), .D(n4655), .Y(n2863) );
  NAND4XLTS U3244 ( .A(n4367), .B(n4366), .C(n4365), .D(n4651), .Y(n2864) );
  OAI211XLTS U3245 ( .A0(n5308), .A1(n4157), .B0(n3745), .C0(n3744), .Y(n2643)
         );
  OAI211XLTS U3246 ( .A0(n5145), .A1(n4157), .B0(n3643), .C0(n3642), .Y(n2658)
         );
  OAI211XLTS U3247 ( .A0(n5135), .A1(n4157), .B0(n4109), .C0(n4108), .Y(n2659)
         );
  OAI211XLTS U3248 ( .A0(n4106), .A1(n4157), .B0(n4105), .C0(n4104), .Y(n2663)
         );
  OAI211XLTS U3249 ( .A0(n4084), .A1(n4140), .B0(n4083), .C0(n4082), .Y(n2673)
         );
  OAI211XLTS U3250 ( .A0(n4064), .A1(n4189), .B0(n3377), .C0(n3376), .Y(n2536)
         );
  OAI211XLTS U3251 ( .A0(n4064), .A1(n4195), .B0(n3379), .C0(n3378), .Y(n2538)
         );
  OAI211XLTS U3252 ( .A0(n4071), .A1(n3890), .B0(n3314), .C0(n3313), .Y(n2539)
         );
  OAI211XLTS U3253 ( .A0(n4072), .A1(n3003), .B0(n3306), .C0(n3305), .Y(n2542)
         );
  NAND4XLTS U3254 ( .A(n4620), .B(n4619), .C(n4618), .D(n4617), .Y(n2543) );
  NAND4XLTS U3255 ( .A(n4606), .B(n4605), .C(n4604), .D(n4603), .Y(n2545) );
  NAND4XLTS U3256 ( .A(n4602), .B(n4601), .C(n4600), .D(n4599), .Y(n2546) );
  NAND4XLTS U3257 ( .A(n4598), .B(n4597), .C(n4596), .D(n4595), .Y(n2547) );
  NAND4XLTS U3258 ( .A(n4594), .B(n4593), .C(n4592), .D(n4591), .Y(n2548) );
  OAI211XLTS U3259 ( .A0(n4064), .A1(n3130), .B0(n4003), .C0(n4002), .Y(n2613)
         );
  OAI211XLTS U3260 ( .A0(n4076), .A1(n4215), .B0(n4067), .C0(n4066), .Y(n2619)
         );
  OAI211XLTS U3261 ( .A0(n4072), .A1(n4043), .B0(n4042), .C0(n4041), .Y(n2621)
         );
  OAI211XLTS U3262 ( .A0(n4076), .A1(n3246), .B0(n4050), .C0(n4049), .Y(n2622)
         );
  OAI211XLTS U3263 ( .A0(n4076), .A1(n4113), .B0(n4075), .C0(n4074), .Y(n2629)
         );
  OAI211XLTS U3264 ( .A0(n4076), .A1(n3280), .B0(n4047), .C0(n4046), .Y(n2630)
         );
  OAI211XLTS U3265 ( .A0(n4072), .A1(n5085), .B0(n4025), .C0(n4024), .Y(n2632)
         );
  OAI211XLTS U3266 ( .A0(n4064), .A1(n5043), .B0(n4021), .C0(n4020), .Y(n2636)
         );
  OAI211XLTS U3267 ( .A0(n4064), .A1(n3009), .B0(n4059), .C0(n4058), .Y(n2641)
         );
  NAND4XLTS U3268 ( .A(n4345), .B(n4344), .C(n4343), .D(n4618), .Y(n2871) );
  NAND4XLTS U3269 ( .A(n4341), .B(n4340), .C(n4339), .D(n4609), .Y(n2872) );
  NAND4XLTS U3270 ( .A(n4338), .B(n4337), .C(n4336), .D(n4604), .Y(n2873) );
  NAND4XLTS U3271 ( .A(n4335), .B(n4334), .C(n4333), .D(n4600), .Y(n2874) );
  NAND4XLTS U3272 ( .A(n4332), .B(n4331), .C(n4330), .D(n4596), .Y(n2875) );
  NAND4XLTS U3273 ( .A(n4329), .B(n4328), .C(n4327), .D(n4592), .Y(n2876) );
  OAI211XLTS U3274 ( .A0(n3890), .A1(n3968), .B0(n3889), .C0(n3888), .Y(n2553)
         );
  NAND4XLTS U3275 ( .A(n4577), .B(n4576), .C(n4575), .D(n4574), .Y(n2558) );
  NAND4XLTS U3276 ( .A(n4545), .B(n4544), .C(n4543), .D(n4542), .Y(n2562) );
  NAND4XLTS U3277 ( .A(n4326), .B(n4325), .C(n4324), .D(n4588), .Y(n2877) );
  NAND4XLTS U3278 ( .A(n4316), .B(n4315), .C(n4314), .D(n4575), .Y(n2878) );
  NAND4XLTS U3279 ( .A(n4305), .B(n4304), .C(n4303), .D(n4559), .Y(n2880) );
  OAI211XLTS U3280 ( .A0(n3699), .A1(n3893), .B0(n3216), .C0(n3215), .Y(n2451)
         );
  OAI211XLTS U3281 ( .A0(n3700), .A1(n3032), .B0(n3087), .C0(n3086), .Y(n2454)
         );
  OAI211XLTS U3282 ( .A0(n3698), .A1(n4244), .B0(n3103), .C0(n3102), .Y(n2458)
         );
  NAND4XLTS U3283 ( .A(n4786), .B(n4785), .C(n4784), .D(n4783), .Y(n2460) );
  NAND4XLTS U3284 ( .A(n4769), .B(n4768), .C(n4767), .D(n4766), .Y(n2464) );
  OAI211XLTS U3285 ( .A0(n3704), .A1(n4817), .B0(n3190), .C0(n3189), .Y(n2571)
         );
  NAND4XLTS U3286 ( .A(n4454), .B(n4453), .C(n4452), .D(n4784), .Y(n2836) );
  NAND4XLTS U3287 ( .A(n4448), .B(n4447), .C(n4446), .D(n4775), .Y(n2838) );
  NAND4XLTS U3288 ( .A(n4445), .B(n4444), .C(n4443), .D(n4771), .Y(n2839) );
  NAND4XLTS U3289 ( .A(n4442), .B(n4441), .C(n4440), .D(n4767), .Y(n2840) );
  OAI211XLTS U3290 ( .A0(n3893), .A1(n3875), .B0(n3872), .C0(n3871), .Y(n2465)
         );
  OAI211XLTS U3291 ( .A0(n4189), .A1(n4228), .B0(n4188), .C0(n4187), .Y(n2466)
         );
  OAI211XLTS U3292 ( .A0(n3076), .A1(n4240), .B0(n4237), .C0(n4236), .Y(n2467)
         );
  OAI211XLTS U3293 ( .A0(n4195), .A1(n4228), .B0(n4194), .C0(n4193), .Y(n2468)
         );
  OAI211XLTS U3294 ( .A0(n3890), .A1(n3875), .B0(n3874), .C0(n3873), .Y(n2469)
         );
  OAI211XLTS U3295 ( .A0(n4235), .A1(n4240), .B0(n4234), .C0(n4233), .Y(n2470)
         );
  OAI211XLTS U3296 ( .A0(n4192), .A1(n4228), .B0(n4191), .C0(n4190), .Y(n2471)
         );
  OAI211XLTS U3297 ( .A0(n4244), .A1(n4228), .B0(n4197), .C0(n4196), .Y(n2472)
         );
  NAND4XLTS U3298 ( .A(n4765), .B(n4764), .C(n4763), .D(n4762), .Y(n2473) );
  NAND4XLTS U3299 ( .A(n4756), .B(n4755), .C(n4754), .D(n4753), .Y(n2474) );
  NAND4XLTS U3300 ( .A(n4752), .B(n4751), .C(n4750), .D(n4749), .Y(n2475) );
  NAND4XLTS U3301 ( .A(n4748), .B(n4747), .C(n4746), .D(n4745), .Y(n2476) );
  NAND4XLTS U3302 ( .A(n4743), .B(n4742), .C(n4741), .D(n4740), .Y(n2477) );
  NAND4XLTS U3303 ( .A(n4739), .B(n4738), .C(n4737), .D(n4736), .Y(n2478) );
  OAI211XLTS U3304 ( .A0(n4817), .A1(n4240), .B0(n4239), .C0(n4238), .Y(n2572)
         );
  OAI211XLTS U3305 ( .A0(n5308), .A1(n4240), .B0(n3395), .C0(n3394), .Y(n2771)
         );
  OAI211XLTS U3306 ( .A0(n5293), .A1(n4240), .B0(n4201), .C0(n4200), .Y(n2772)
         );
  OAI211XLTS U3307 ( .A0(n4175), .A1(n4229), .B0(n4174), .C0(n4173), .Y(n2773)
         );
  OAI211XLTS U3308 ( .A0(n3951), .A1(n4229), .B0(n3834), .C0(n3833), .Y(n2774)
         );
  OAI211XLTS U3309 ( .A0(n4085), .A1(n4240), .B0(n3852), .C0(n3851), .Y(n2776)
         );
  OAI211XLTS U3310 ( .A0(n4183), .A1(n4229), .B0(n4182), .C0(n4181), .Y(n2777)
         );
  OAI211XLTS U3311 ( .A0(n4179), .A1(n4229), .B0(n4178), .C0(n4177), .Y(n2778)
         );
  OAI211XLTS U3312 ( .A0(n5217), .A1(n4240), .B0(n4218), .C0(n4217), .Y(n2779)
         );
  OAI211XLTS U3313 ( .A0(n4043), .A1(n4240), .B0(n3861), .C0(n3860), .Y(n2781)
         );
  OAI211XLTS U3314 ( .A0(n4205), .A1(n4240), .B0(n4204), .C0(n4203), .Y(n2784)
         );
  OAI211XLTS U3315 ( .A0(n3209), .A1(n4240), .B0(n4210), .C0(n4209), .Y(n2785)
         );
  OAI211XLTS U3316 ( .A0(n5145), .A1(n4240), .B0(n4222), .C0(n4221), .Y(n2786)
         );
  OAI211XLTS U3317 ( .A0(n5135), .A1(n4240), .B0(n4214), .C0(n4213), .Y(n2787)
         );
  OAI211XLTS U3318 ( .A0(n3357), .A1(n4229), .B0(n3389), .C0(n3388), .Y(n2788)
         );
  OAI211XLTS U3319 ( .A0(n4117), .A1(n4240), .B0(n3707), .C0(n3706), .Y(n2789)
         );
  OAI211XLTS U3320 ( .A0(n3280), .A1(n4229), .B0(n4165), .C0(n4164), .Y(n2790)
         );
  OAI211XLTS U3321 ( .A0(n4102), .A1(n4229), .B0(n3392), .C0(n3391), .Y(n2791)
         );
  OAI211XLTS U3322 ( .A0(n3064), .A1(n4229), .B0(n4186), .C0(n4185), .Y(n2793)
         );
  OAI211XLTS U3323 ( .A0(n3201), .A1(n4229), .B0(n3840), .C0(n3839), .Y(n2795)
         );
  OAI211XLTS U3324 ( .A0(n4018), .A1(n4229), .B0(n3846), .C0(n3845), .Y(n2796)
         );
  OAI211XLTS U3325 ( .A0(n5023), .A1(n4240), .B0(n3855), .C0(n3854), .Y(n2798)
         );
  OAI211XLTS U3326 ( .A0(n3985), .A1(n4229), .B0(n3849), .C0(n3848), .Y(n2799)
         );
  OAI211XLTS U3327 ( .A0(n4990), .A1(n4240), .B0(n3864), .C0(n3863), .Y(n2801)
         );
  NAND4XLTS U3328 ( .A(n4439), .B(n4438), .C(n4437), .D(n4763), .Y(n2841) );
  NAND4XLTS U3329 ( .A(n4435), .B(n4434), .C(n4433), .D(n4754), .Y(n2842) );
  NAND4XLTS U3330 ( .A(n4432), .B(n4431), .C(n4430), .D(n4750), .Y(n2843) );
  NAND4XLTS U3331 ( .A(n4429), .B(n4428), .C(n4427), .D(n4746), .Y(n2844) );
  NAND4XLTS U3332 ( .A(n4426), .B(n4425), .C(n4424), .D(n4741), .Y(n2845) );
  NAND4XLTS U3333 ( .A(n4423), .B(n4422), .C(n4421), .D(n4737), .Y(n2846) );
  OAI211XLTS U3334 ( .A0(n3533), .A1(n3074), .B0(n3080), .C0(n3079), .Y(n2481)
         );
  OAI211XLTS U3335 ( .A0(n3538), .A1(n3890), .B0(n3173), .C0(n3172), .Y(n2483)
         );
  OAI211XLTS U3336 ( .A0(n3542), .A1(n2973), .B0(n2978), .C0(n2977), .Y(n2485)
         );
  NAND4XLTS U3337 ( .A(n4735), .B(n4734), .C(n4733), .D(n4732), .Y(n2487) );
  NAND4XLTS U3338 ( .A(n4727), .B(n4726), .C(n4725), .D(n4724), .Y(n2488) );
  NAND4XLTS U3339 ( .A(n4723), .B(n4722), .C(n4721), .D(n4720), .Y(n2489) );
  NAND4XLTS U3340 ( .A(n4715), .B(n4714), .C(n4713), .D(n4712), .Y(n2491) );
  NAND4XLTS U3341 ( .A(n4711), .B(n4710), .C(n4709), .D(n4708), .Y(n2492) );
  OAI211XLTS U3342 ( .A0(n3542), .A1(n5259), .B0(n3519), .C0(n3518), .Y(n2743)
         );
  OAI211XLTS U3343 ( .A0(n3538), .A1(n4022), .B0(n3162), .C0(n3161), .Y(n2760)
         );
  OAI211XLTS U3344 ( .A0(n3537), .A1(n3009), .B0(n3016), .C0(n3015), .Y(n2769)
         );
  NAND4XLTS U3345 ( .A(n4420), .B(n4419), .C(n4418), .D(n4733), .Y(n2847) );
  NAND4XLTS U3346 ( .A(n4413), .B(n4412), .C(n4411), .D(n4721), .Y(n2849) );
  NAND4XLTS U3347 ( .A(n4410), .B(n4409), .C(n4408), .D(n4717), .Y(n2850) );
  OAI211XLTS U3348 ( .A0(n3567), .A1(n4189), .B0(n3070), .C0(n3069), .Y(n2494)
         );
  OAI211XLTS U3349 ( .A0(n3579), .A1(n3890), .B0(n3125), .C0(n3124), .Y(n2497)
         );
  OAI211XLTS U3350 ( .A0(n3575), .A1(n4235), .B0(n3192), .C0(n3191), .Y(n2498)
         );
  NAND4XLTS U3351 ( .A(n4691), .B(n4690), .C(n4689), .D(n4688), .Y(n2504) );
  OAI211XLTS U3352 ( .A0(n3574), .A1(n4183), .B0(n3239), .C0(n3238), .Y(n2713)
         );
  OAI211XLTS U3353 ( .A0(n3579), .A1(n2954), .B0(n3578), .C0(n3577), .Y(n2715)
         );
  OAI211XLTS U3354 ( .A0(n3575), .A1(n5188), .B0(n3252), .C0(n3251), .Y(n2718)
         );
  OAI211XLTS U3355 ( .A0(n3574), .A1(n3406), .B0(n3414), .C0(n3413), .Y(n2720)
         );
  OAI211XLTS U3356 ( .A0(n3574), .A1(n4211), .B0(n3420), .C0(n3419), .Y(n2723)
         );
  OAI211XLTS U3357 ( .A0(n3575), .A1(n4117), .B0(n3563), .C0(n3562), .Y(n2725)
         );
  OAI211XLTS U3358 ( .A0(n3575), .A1(n5033), .B0(n3560), .C0(n3559), .Y(n2733)
         );
  OAI211XLTS U3359 ( .A0(n3574), .A1(n4136), .B0(n3438), .C0(n3437), .Y(n2734)
         );
  OAI211XLTS U3360 ( .A0(n3579), .A1(n3494), .B0(n3570), .C0(n3569), .Y(n2736)
         );
  OAI211XLTS U3361 ( .A0(n3826), .A1(n5306), .B0(n3767), .C0(n3766), .Y(n2675)
         );
  OAI211XLTS U3362 ( .A0(n3826), .A1(n3127), .B0(n3776), .C0(n3775), .Y(n2677)
         );
  OAI211XLTS U3363 ( .A0(n3807), .A1(n5207), .B0(n3761), .C0(n3760), .Y(n2684)
         );
  OAI211XLTS U3364 ( .A0(n3807), .A1(n3292), .B0(n3800), .C0(n3799), .Y(n2685)
         );
  OAI211XLTS U3365 ( .A0(n3831), .A1(n3246), .B0(n3715), .C0(n3714), .Y(n2686)
         );
  OAI211XLTS U3366 ( .A0(n3807), .A1(n5176), .B0(n3803), .C0(n3802), .Y(n2687)
         );
  OAI211XLTS U3367 ( .A0(n3831), .A1(n4219), .B0(n3712), .C0(n3711), .Y(n2690)
         );
  OAI211XLTS U3368 ( .A0(n3807), .A1(n4161), .B0(n3794), .C0(n3793), .Y(n2694)
         );
  OAI211XLTS U3369 ( .A0(n3831), .A1(n4102), .B0(n3822), .C0(n3821), .Y(n2695)
         );
  OAI211XLTS U3370 ( .A0(n3807), .A1(n5086), .B0(n3806), .C0(n3805), .Y(n2696)
         );
  OAI211XLTS U3371 ( .A0(n3827), .A1(n4166), .B0(n3733), .C0(n3732), .Y(n2698)
         );
  OAI211XLTS U3372 ( .A0(n3826), .A1(n5044), .B0(n3727), .C0(n3726), .Y(n2700)
         );
  OAI211XLTS U3373 ( .A0(n3807), .A1(n3009), .B0(n3779), .C0(n3778), .Y(n2705)
         );
  OAI211XLTS U3374 ( .A0(n3807), .A1(n3018), .B0(n3782), .C0(n3781), .Y(n2706)
         );
  NAND4XLTS U3375 ( .A(n4383), .B(n4382), .C(n4381), .D(n4676), .Y(n2859) );
  NAND4XLTS U3376 ( .A(n4379), .B(n4378), .C(n4377), .D(n4668), .Y(n2860) );
  OAI211XLTS U3377 ( .A0(n3893), .A1(n4077), .B0(n3753), .C0(n3752), .Y(n2521)
         );
  OAI211XLTS U3378 ( .A0(n4189), .A1(n4243), .B0(n4150), .C0(n4149), .Y(n2522)
         );
  OAI211XLTS U3379 ( .A0(n3076), .A1(n4157), .B0(n4154), .C0(n4153), .Y(n2523)
         );
  OAI211XLTS U3380 ( .A0(n4195), .A1(n4243), .B0(n4146), .C0(n4145), .Y(n2524)
         );
  OAI211XLTS U3381 ( .A0(n3890), .A1(n4077), .B0(n3755), .C0(n3754), .Y(n2525)
         );
  OAI211XLTS U3382 ( .A0(n4235), .A1(n4157), .B0(n4156), .C0(n4155), .Y(n2526)
         );
  OAI211XLTS U3383 ( .A0(n4192), .A1(n4243), .B0(n4148), .C0(n4147), .Y(n2527)
         );
  OAI211XLTS U3384 ( .A0(n4244), .A1(n4243), .B0(n4242), .C0(n4241), .Y(n2528)
         );
  NAND4XLTS U3385 ( .A(n4649), .B(n4648), .C(n4647), .D(n4646), .Y(n2529) );
  NAND4XLTS U3386 ( .A(n4640), .B(n4639), .C(n4638), .D(n4637), .Y(n2530) );
  NAND4XLTS U3387 ( .A(n4636), .B(n4635), .C(n4634), .D(n4633), .Y(n2531) );
  NAND4XLTS U3388 ( .A(n4632), .B(n4631), .C(n4630), .D(n4629), .Y(n2532) );
  NAND4XLTS U3389 ( .A(n4628), .B(n4627), .C(n4626), .D(n4625), .Y(n2533) );
  NAND4XLTS U3390 ( .A(n4624), .B(n4623), .C(n4622), .D(n4621), .Y(n2534) );
  OAI211XLTS U3391 ( .A0(n4817), .A1(n4157), .B0(n4152), .C0(n4151), .Y(n2576)
         );
  OAI211XLTS U3392 ( .A0(n4198), .A1(n4140), .B0(n4095), .C0(n4094), .Y(n2644)
         );
  OAI211XLTS U3393 ( .A0(n4175), .A1(n4140), .B0(n4080), .C0(n4079), .Y(n2645)
         );
  OAI211XLTS U3394 ( .A0(n3951), .A1(n4140), .B0(n3739), .C0(n3738), .Y(n2646)
         );
  OAI211XLTS U3395 ( .A0(n5259), .A1(n4157), .B0(n3640), .C0(n3639), .Y(n2647)
         );
  OAI211XLTS U3396 ( .A0(n4089), .A1(n4140), .B0(n4088), .C0(n4087), .Y(n2648)
         );
  OAI211XLTS U3397 ( .A0(n5239), .A1(n4157), .B0(n4131), .C0(n4130), .Y(n2649)
         );
  OAI211XLTS U3398 ( .A0(n5227), .A1(n4157), .B0(n4127), .C0(n4126), .Y(n2650)
         );
  OAI211XLTS U3399 ( .A0(n5217), .A1(n4157), .B0(n4124), .C0(n4123), .Y(n2651)
         );
  OAI211XLTS U3400 ( .A0(n4223), .A1(n4140), .B0(n4098), .C0(n4097), .Y(n2652)
         );
  OAI211XLTS U3401 ( .A0(n3289), .A1(n4140), .B0(n3628), .C0(n3627), .Y(n2653)
         );
  OAI211XLTS U3402 ( .A0(n3246), .A1(n4140), .B0(n3625), .C0(n3624), .Y(n2654)
         );
  OAI211XLTS U3403 ( .A0(n5177), .A1(n4157), .B0(n3748), .C0(n3747), .Y(n2655)
         );
  OAI211XLTS U3404 ( .A0(n3406), .A1(n4140), .B0(n3622), .C0(n3621), .Y(n2656)
         );
  OAI211XLTS U3405 ( .A0(n3209), .A1(n4157), .B0(n3637), .C0(n3636), .Y(n2657)
         );
  OAI211XLTS U3406 ( .A0(n5124), .A1(n4157), .B0(n3634), .C0(n3633), .Y(n2660)
         );
  OAI211XLTS U3407 ( .A0(n4117), .A1(n4157), .B0(n4116), .C0(n4115), .Y(n2661)
         );
  OAI211XLTS U3408 ( .A0(n4162), .A1(n4157), .B0(n4112), .C0(n4111), .Y(n2662)
         );
  OAI211XLTS U3409 ( .A0(n5085), .A1(n4157), .B0(n3631), .C0(n3630), .Y(n2664)
         );
  OAI211XLTS U3410 ( .A0(n3064), .A1(n4140), .B0(n4092), .C0(n4091), .Y(n2665)
         );
  OAI211XLTS U3411 ( .A0(n4170), .A1(n4140), .B0(n4101), .C0(n4100), .Y(n2666)
         );
  OAI211XLTS U3412 ( .A0(n3201), .A1(n4140), .B0(n3742), .C0(n3741), .Y(n2667)
         );
  OAI211XLTS U3413 ( .A0(n4018), .A1(n4140), .B0(n3736), .C0(n3735), .Y(n2668)
         );
  OAI211XLTS U3414 ( .A0(n5033), .A1(n4157), .B0(n4144), .C0(n4143), .Y(n2669)
         );
  OAI211XLTS U3415 ( .A0(n5023), .A1(n4157), .B0(n4139), .C0(n4138), .Y(n2670)
         );
  OAI211XLTS U3416 ( .A0(n5011), .A1(n4157), .B0(n3751), .C0(n3750), .Y(n2671)
         );
  OAI211XLTS U3417 ( .A0(n5001), .A1(n4157), .B0(n4135), .C0(n4134), .Y(n2672)
         );
  OAI211XLTS U3418 ( .A0(n3023), .A1(n4157), .B0(n4121), .C0(n4120), .Y(n2674)
         );
  NAND4XLTS U3419 ( .A(n4364), .B(n4363), .C(n4362), .D(n4647), .Y(n2865) );
  NAND4XLTS U3420 ( .A(n4360), .B(n4359), .C(n4358), .D(n4638), .Y(n2866) );
  NAND4XLTS U3421 ( .A(n4357), .B(n4356), .C(n4355), .D(n4634), .Y(n2867) );
  NAND4XLTS U3422 ( .A(n4354), .B(n4353), .C(n4352), .D(n4630), .Y(n2868) );
  NAND4XLTS U3423 ( .A(n4351), .B(n4350), .C(n4349), .D(n4626), .Y(n2869) );
  NAND4XLTS U3424 ( .A(n4348), .B(n4347), .C(n4346), .D(n4622), .Y(n2870) );
  OAI211XLTS U3425 ( .A0(n4071), .A1(n5306), .B0(n3981), .C0(n3980), .Y(n2611)
         );
  OAI211XLTS U3426 ( .A0(n4072), .A1(n5293), .B0(n4013), .C0(n4012), .Y(n2612)
         );
  OAI211XLTS U3427 ( .A0(n4072), .A1(n5270), .B0(n3881), .C0(n3880), .Y(n2614)
         );
  OAI211XLTS U3428 ( .A0(n4064), .A1(n5260), .B0(n4007), .C0(n4006), .Y(n2615)
         );
  OAI211XLTS U3429 ( .A0(n4064), .A1(n3430), .B0(n4063), .C0(n4062), .Y(n2616)
         );
  OAI211XLTS U3430 ( .A0(n4071), .A1(n5228), .B0(n3997), .C0(n3996), .Y(n2618)
         );
  OAI211XLTS U3431 ( .A0(n4072), .A1(n4227), .B0(n4038), .C0(n4037), .Y(n2620)
         );
  OAI211XLTS U3432 ( .A0(n4076), .A1(n3262), .B0(n4017), .C0(n4016), .Y(n2623)
         );
  OAI211XLTS U3433 ( .A0(n4076), .A1(n4206), .B0(n4035), .C0(n4034), .Y(n2625)
         );
  OAI211XLTS U3434 ( .A0(n4071), .A1(n3045), .B0(n4000), .C0(n3999), .Y(n2626)
         );
  OAI211XLTS U3435 ( .A0(n4064), .A1(n5134), .B0(n4010), .C0(n4009), .Y(n2627)
         );
  OAI211XLTS U3436 ( .A0(n4076), .A1(n3357), .B0(n4070), .C0(n4069), .Y(n2628)
         );
  OAI211XLTS U3437 ( .A0(n4076), .A1(n4102), .B0(n4032), .C0(n4031), .Y(n2631)
         );
  OAI211XLTS U3438 ( .A0(n4064), .A1(n5075), .B0(n3978), .C0(n3977), .Y(n2633)
         );
  OAI211XLTS U3439 ( .A0(n4076), .A1(n4170), .B0(n3994), .C0(n3993), .Y(n2634)
         );
  OAI211XLTS U3440 ( .A0(n4071), .A1(n5054), .B0(n3887), .C0(n3886), .Y(n2635)
         );
  OAI211XLTS U3441 ( .A0(n4076), .A1(n4141), .B0(n3991), .C0(n3990), .Y(n2637)
         );
  OAI211XLTS U3442 ( .A0(n4071), .A1(n5012), .B0(n3988), .C0(n3987), .Y(n2639)
         );
  OAI211XLTS U3443 ( .A0(n4064), .A1(n3492), .B0(n4056), .C0(n4055), .Y(n2640)
         );
  OAI211XLTS U3444 ( .A0(n4072), .A1(n3023), .B0(n4028), .C0(n4027), .Y(n2642)
         );
  OAI211XLTS U3445 ( .A0(n3893), .A1(n3968), .B0(n3892), .C0(n3891), .Y(n2549)
         );
  OAI211XLTS U3446 ( .A0(n4189), .A1(n3969), .B0(n3895), .C0(n3894), .Y(n2550)
         );
  OAI211XLTS U3447 ( .A0(n3076), .A1(n3964), .B0(n3914), .C0(n3913), .Y(n2551)
         );
  OAI211XLTS U3448 ( .A0(n4195), .A1(n3969), .B0(n3897), .C0(n3896), .Y(n2552)
         );
  OAI211XLTS U3449 ( .A0(n4235), .A1(n3964), .B0(n3922), .C0(n3921), .Y(n2554)
         );
  OAI211XLTS U3450 ( .A0(n4192), .A1(n3969), .B0(n3324), .C0(n3323), .Y(n2555)
         );
  OAI211XLTS U3451 ( .A0(n4244), .A1(n3969), .B0(n3322), .C0(n3321), .Y(n2556)
         );
  NAND4XLTS U3452 ( .A(n4590), .B(n4589), .C(n4588), .D(n4587), .Y(n2557) );
  NAND4XLTS U3453 ( .A(n4569), .B(n4568), .C(n4567), .D(n4566), .Y(n2559) );
  NAND4XLTS U3454 ( .A(n4561), .B(n4560), .C(n4559), .D(n4558), .Y(n2560) );
  NAND4XLTS U3455 ( .A(n4553), .B(n4552), .C(n4551), .D(n4550), .Y(n2561) );
  OAI211XLTS U3456 ( .A0(n5308), .A1(n3964), .B0(n3900), .C0(n3899), .Y(n2579)
         );
  OAI211XLTS U3457 ( .A0(n4198), .A1(n3975), .B0(n3943), .C0(n3942), .Y(n2580)
         );
  OAI211XLTS U3458 ( .A0(n4171), .A1(n3964), .B0(n3917), .C0(n3916), .Y(n2581)
         );
  OAI211XLTS U3459 ( .A0(n3951), .A1(n3975), .B0(n3950), .C0(n3949), .Y(n2582)
         );
  OAI211XLTS U3460 ( .A0(n3299), .A1(n3975), .B0(n3946), .C0(n3945), .Y(n2583)
         );
  OAI211XLTS U3461 ( .A0(n4085), .A1(n3964), .B0(n3925), .C0(n3924), .Y(n2584)
         );
  OAI211XLTS U3462 ( .A0(n5239), .A1(n3964), .B0(n3903), .C0(n3902), .Y(n2585)
         );
  OAI211XLTS U3463 ( .A0(n4179), .A1(n3975), .B0(n3928), .C0(n3927), .Y(n2586)
         );
  OAI211XLTS U3464 ( .A0(n4215), .A1(n3975), .B0(n3931), .C0(n3930), .Y(n2587)
         );
  OAI211XLTS U3465 ( .A0(n4227), .A1(n3964), .B0(n3906), .C0(n3905), .Y(n2588)
         );
  OAI211XLTS U3466 ( .A0(n3289), .A1(n3975), .B0(n3954), .C0(n3953), .Y(n2589)
         );
  OAI211XLTS U3467 ( .A0(n5188), .A1(n3964), .B0(n3912), .C0(n3911), .Y(n2590)
         );
  OAI211XLTS U3468 ( .A0(n5177), .A1(n3964), .B0(n3920), .C0(n3919), .Y(n2591)
         );
  OAI211XLTS U3469 ( .A0(n3406), .A1(n3975), .B0(n3934), .C0(n3933), .Y(n2592)
         );
  OAI211XLTS U3470 ( .A0(n4206), .A1(n3975), .B0(n3334), .C0(n3333), .Y(n2593)
         );
  OAI211XLTS U3471 ( .A0(n4219), .A1(n3975), .B0(n3373), .C0(n3372), .Y(n2594)
         );
  OAI211XLTS U3472 ( .A0(n5135), .A1(n3964), .B0(n3349), .C0(n3348), .Y(n2595)
         );
  OAI211XLTS U3473 ( .A0(n5124), .A1(n3964), .B0(n3361), .C0(n3360), .Y(n2596)
         );
  OAI211XLTS U3474 ( .A0(n4113), .A1(n3975), .B0(n3331), .C0(n3330), .Y(n2597)
         );
  OAI211XLTS U3475 ( .A0(n4162), .A1(n3964), .B0(n3352), .C0(n3351), .Y(n2598)
         );
  OAI211XLTS U3476 ( .A0(n4102), .A1(n3975), .B0(n3370), .C0(n3369), .Y(n2599)
         );
  OAI211XLTS U3477 ( .A0(n5085), .A1(n3964), .B0(n3328), .C0(n3327), .Y(n2600)
         );
  OAI211XLTS U3478 ( .A0(n3064), .A1(n3975), .B0(n3337), .C0(n3336), .Y(n2601)
         );
  OAI211XLTS U3479 ( .A0(n4170), .A1(n3975), .B0(n3340), .C0(n3339), .Y(n2602)
         );
  OAI211XLTS U3480 ( .A0(n3201), .A1(n3975), .B0(n3972), .C0(n3971), .Y(n2603)
         );
  OAI211XLTS U3481 ( .A0(n3271), .A1(n3964), .B0(n3909), .C0(n3908), .Y(n2604)
         );
  OAI211XLTS U3482 ( .A0(n4141), .A1(n3975), .B0(n3957), .C0(n3956), .Y(n2605)
         );
  OAI211XLTS U3483 ( .A0(n4136), .A1(n3975), .B0(n3967), .C0(n3966), .Y(n2606)
         );
  OAI211XLTS U3484 ( .A0(n3985), .A1(n3975), .B0(n3963), .C0(n3962), .Y(n2607)
         );
  OAI211XLTS U3485 ( .A0(n4132), .A1(n3975), .B0(n3940), .C0(n3939), .Y(n2608)
         );
  OAI211XLTS U3486 ( .A0(n4084), .A1(n3975), .B0(n3960), .C0(n3959), .Y(n2609)
         );
  OAI211XLTS U3487 ( .A0(n4118), .A1(n3975), .B0(n3937), .C0(n3936), .Y(n2610)
         );
  NAND4XLTS U3488 ( .A(n4308), .B(n4307), .C(n4306), .D(n4567), .Y(n2879) );
  NAND4XLTS U3489 ( .A(n4297), .B(n4296), .C(n4295), .D(n4551), .Y(n2881) );
  NAND4XLTS U3490 ( .A(n4289), .B(n4288), .C(n4287), .D(n4543), .Y(n2882) );
  OAI211XLTS U3491 ( .A0(n3827), .A1(n4817), .B0(n3220), .C0(n3219), .Y(n2575)
         );
  AOI2BB1XLTS U3492 ( .A0N(n4537), .A1N(readOutbuffer[0]), .B0(n4536), .Y(
        n2563) );
  AOI2BB1XLTS U3493 ( .A0N(n4528), .A1N(readOutbuffer[1]), .B0(n4527), .Y(
        n2564) );
  AOI2BB1XLTS U3494 ( .A0N(n4491), .A1N(readOutbuffer[5]), .B0(n4490), .Y(
        n2568) );
  OAI211XLTS U3495 ( .A0(n3542), .A1(n4817), .B0(n2986), .C0(n2985), .Y(n2573)
         );
  AOI2BB2XLTS U3496 ( .B0(n4520), .B1(n4519), .A0N(n4518), .A1N(
        readOutbuffer[2]), .Y(n2565) );
  AOI211XLTS U3497 ( .A0(n4464), .A1(n4517), .B0(n4516), .C0(n4515), .Y(n4520)
         );
  AOI2BB1XLTS U3498 ( .A0N(n4473), .A1N(readOutbuffer[7]), .B0(n4472), .Y(
        n2570) );
  OAI211XLTS U3499 ( .A0(n3700), .A1(n3074), .B0(n3105), .C0(n3104), .Y(n2453)
         );
  OAI211XLTS U3500 ( .A0(n3699), .A1(n3890), .B0(n3218), .C0(n3217), .Y(n2455)
         );
  OAI211XLTS U3501 ( .A0(n3704), .A1(n2973), .B0(n3185), .C0(n3184), .Y(n2457)
         );
  OAI211XLTS U3502 ( .A0(n3698), .A1(n3401), .B0(n3691), .C0(n3690), .Y(n2806)
         );
  OAI211XLTS U3503 ( .A0(n3704), .A1(n5259), .B0(n3606), .C0(n3605), .Y(n2807)
         );
  OAI211XLTS U3504 ( .A0(n3698), .A1(n2958), .B0(n3664), .C0(n3663), .Y(n2811)
         );
  OAI211XLTS U3505 ( .A0(n3698), .A1(n5187), .B0(n3670), .C0(n3669), .Y(n2814)
         );
  OAI211XLTS U3506 ( .A0(n3700), .A1(n3064), .B0(n3582), .C0(n3581), .Y(n2825)
         );
  OAI211XLTS U3507 ( .A0(n3699), .A1(n3531), .B0(n3661), .C0(n3660), .Y(n2829)
         );
  OAI211XLTS U3508 ( .A0(n3700), .A1(n4132), .B0(n3679), .C0(n3678), .Y(n2832)
         );
  OAI211XLTS U3509 ( .A0(n3700), .A1(n4084), .B0(n3682), .C0(n3681), .Y(n2833)
         );
  OAI211XLTS U3510 ( .A0(n3700), .A1(n4118), .B0(n3676), .C0(n3675), .Y(n2834)
         );
  OAI211XLTS U3511 ( .A0(n3023), .A1(n4240), .B0(n3870), .C0(n3869), .Y(n2802)
         );
  OAI211XLTS U3512 ( .A0(n3542), .A1(n3036), .B0(n3041), .C0(n3040), .Y(n2480)
         );
  OAI211XLTS U3513 ( .A0(n3537), .A1(n4195), .B0(n3034), .C0(n3033), .Y(n2482)
         );
  OAI211XLTS U3514 ( .A0(n3542), .A1(n4235), .B0(n2992), .C0(n2991), .Y(n2484)
         );
  OAI211XLTS U3515 ( .A0(n3542), .A1(n3003), .B0(n3082), .C0(n3081), .Y(n2486)
         );
  OAI211XLTS U3516 ( .A0(n3538), .A1(n5306), .B0(n3144), .C0(n3143), .Y(n2739)
         );
  OAI211XLTS U3517 ( .A0(n3538), .A1(n5228), .B0(n3153), .C0(n3152), .Y(n2746)
         );
  OAI211XLTS U3518 ( .A0(n3533), .A1(n4223), .B0(n3488), .C0(n3487), .Y(n2748)
         );
  OAI211XLTS U3519 ( .A0(n3542), .A1(n5145), .B0(n3050), .C0(n3049), .Y(n2754)
         );
  OAI211XLTS U3520 ( .A0(n3537), .A1(n5043), .B0(n3507), .C0(n3506), .Y(n2764)
         );
  OAI211XLTS U3521 ( .A0(n3533), .A1(n4132), .B0(n3498), .C0(n3497), .Y(n2768)
         );
  OAI211XLTS U3522 ( .A0(n3537), .A1(n3018), .B0(n3026), .C0(n3025), .Y(n2770)
         );
  OAI211XLTS U3523 ( .A0(n3579), .A1(n3893), .B0(n3119), .C0(n3118), .Y(n2493)
         );
  OAI211XLTS U3524 ( .A0(n3567), .A1(n4195), .B0(n3072), .C0(n3071), .Y(n2496)
         );
  OAI211XLTS U3525 ( .A0(n3567), .A1(n4192), .B0(n3000), .C0(n2999), .Y(n2499)
         );
  OAI211XLTS U3526 ( .A0(n3575), .A1(n4817), .B0(n3194), .C0(n3193), .Y(n2574)
         );
  OAI211XLTS U3527 ( .A0(n3579), .A1(n5054), .B0(n3545), .C0(n3544), .Y(n2731)
         );
  OAI211XLTS U3528 ( .A0(n3826), .A1(n3893), .B0(n3228), .C0(n3227), .Y(n2507)
         );
  OAI211XLTS U3529 ( .A0(n3826), .A1(n3890), .B0(n3226), .C0(n3225), .Y(n2511)
         );
  OAI211XLTS U3530 ( .A0(n3826), .A1(n5156), .B0(n3730), .C0(n3729), .Y(n2689)
         );
  OAI211XLTS U3531 ( .A0(n3807), .A1(n5134), .B0(n3791), .C0(n3790), .Y(n2691)
         );
  OAI211XLTS U3532 ( .A0(n3827), .A1(n5124), .B0(n3785), .C0(n3784), .Y(n2692)
         );
  OAI211XLTS U3533 ( .A0(n3826), .A1(n5012), .B0(n3770), .C0(n3769), .Y(n2703)
         );
  OAI211XLTS U3534 ( .A0(n4071), .A1(n3893), .B0(n3312), .C0(n3311), .Y(n2535)
         );
  OAI211XLTS U3535 ( .A0(n4076), .A1(n3074), .B0(n3113), .C0(n3112), .Y(n2537)
         );
  OAI211XLTS U3536 ( .A0(n4072), .A1(n4235), .B0(n3310), .C0(n3309), .Y(n2540)
         );
  OAI211XLTS U3537 ( .A0(n4064), .A1(n4192), .B0(n3375), .C0(n3374), .Y(n2541)
         );
  NAND4XLTS U3538 ( .A(n4611), .B(n4610), .C(n4609), .D(n4608), .Y(n2544) );
  OAI211XLTS U3539 ( .A0(n4072), .A1(n4817), .B0(n3308), .C0(n3307), .Y(n2577)
         );
  OAI211XLTS U3540 ( .A0(n4071), .A1(n5238), .B0(n3984), .C0(n3983), .Y(n2617)
         );
  OAI211XLTS U3541 ( .A0(n4072), .A1(n4205), .B0(n3884), .C0(n3883), .Y(n2624)
         );
  OAI211XLTS U3542 ( .A0(n4064), .A1(n3166), .B0(n4053), .C0(n4052), .Y(n2638)
         );
  OAI211XLTS U3543 ( .A0(n2984), .A1(n3975), .B0(n3974), .C0(n3973), .Y(n2578)
         );
  AOI2BB1XLTS U3544 ( .A0N(n4511), .A1N(readOutbuffer[3]), .B0(n4510), .Y(
        n2566) );
  OAI21XLTS U3545 ( .A0(n4498), .A1(n4797), .B0(n4497), .Y(n4499) );
  OAI21XLTS U3546 ( .A0(n4480), .A1(n4797), .B0(n4479), .Y(n4481) );
  OAI32X1TS U3547 ( .A0(n4286), .A1(n5325), .A2(n4278), .B0(n5324), .B1(n4286), 
        .Y(n2883) );
  AOI211XLTS U3548 ( .A0(n4271), .A1(read_reg[2]), .B0(n4270), .C0(n4269), .Y(
        n4272) );
  XOR2XLTS U3549 ( .A(read_reg[0]), .B(n4274), .Y(n4270) );
  OAI21XLTS U3550 ( .A0(n4271), .A1(read_reg[2]), .B0(n4268), .Y(n4269) );
  OR2X1TS U3551 ( .A(n4815), .B(n4273), .Y(n5291) );
  OR2X1TS U3552 ( .A(n4795), .B(n4273), .Y(n5305) );
  INVX2TS U3553 ( .A(n2896), .Y(n2897) );
  INVX2TS U3554 ( .A(n2901), .Y(n2902) );
  INVX2TS U3555 ( .A(n3063), .Y(n3064) );
  INVX2TS U3556 ( .A(n3200), .Y(n3201) );
  INVX2TS U3557 ( .A(n3139), .Y(n3140) );
  INVX2TS U3558 ( .A(n3356), .Y(n3357) );
  INVX2TS U3559 ( .A(n3055), .Y(n3056) );
  INVX2TS U3560 ( .A(n3493), .Y(n3494) );
  INVX2TS U3561 ( .A(n3022), .Y(n3023) );
  INVX2TS U3562 ( .A(n3235), .Y(n3236) );
  INVX2TS U3563 ( .A(n3291), .Y(n3292) );
  INVX2TS U3564 ( .A(n2957), .Y(n2958) );
  INVX2TS U3565 ( .A(n3345), .Y(n3346) );
  INVX2TS U3566 ( .A(n3405), .Y(n3406) );
  INVX2TS U3567 ( .A(n3149), .Y(n3150) );
  INVX2TS U3568 ( .A(n3298), .Y(n3299) );
  INVX2TS U3569 ( .A(n3530), .Y(n3531) );
  INVX2TS U3570 ( .A(n3483), .Y(n3484) );
  INVX2TS U3571 ( .A(n3247), .Y(n3248) );
  INVX2TS U3572 ( .A(n3364), .Y(n3365) );
  INVX2TS U3573 ( .A(n3400), .Y(n3401) );
  INVX2TS U3574 ( .A(n2953), .Y(n2954) );
  INVX2TS U3575 ( .A(n3126), .Y(n3127) );
  INVX2TS U3576 ( .A(n3459), .Y(n3460) );
  INVX2TS U3577 ( .A(n3528), .Y(n3529) );
  INVX2TS U3578 ( .A(n2965), .Y(n2966) );
  INVX2TS U3579 ( .A(n2962), .Y(n2963) );
  INVX2TS U3580 ( .A(n4460), .Y(n4461) );
  INVX2TS U3581 ( .A(n2983), .Y(n2984) );
  INVX2TS U3582 ( .A(n2980), .Y(n2981) );
  INVX2TS U3583 ( .A(n3245), .Y(n3246) );
  INVX2TS U3584 ( .A(n3408), .Y(n3409) );
  INVX2TS U3585 ( .A(n3017), .Y(n3018) );
  INVX2TS U3586 ( .A(n3073), .Y(n3074) );
  INVX2TS U3587 ( .A(n3208), .Y(n3209) );
  INVX2TS U3588 ( .A(n3279), .Y(n3280) );
  INVX2TS U3589 ( .A(n3261), .Y(n3262) );
  INVX2TS U3590 ( .A(n3129), .Y(n3130) );
  INVX2TS U3591 ( .A(n3008), .Y(n3009) );
  INVX2TS U3592 ( .A(n3075), .Y(n3076) );
  INVX2TS U3593 ( .A(n3156), .Y(n3157) );
  INVX2TS U3594 ( .A(n3491), .Y(n3492) );
  INVX2TS U3595 ( .A(n3044), .Y(n3045) );
  INVX2TS U3596 ( .A(n3429), .Y(n3430) );
  INVX2TS U3597 ( .A(n3288), .Y(n3289) );
  INVX2TS U3598 ( .A(n3002), .Y(n3003) );
  INVX2TS U3599 ( .A(n2972), .Y(n2973) );
  INVX2TS U3600 ( .A(n3035), .Y(n3036) );
  INVX2TS U3601 ( .A(n3165), .Y(n3166) );
  INVX2TS U3602 ( .A(n2924), .Y(n2925) );
  INVX2TS U3603 ( .A(n2905), .Y(n2906) );
  INVX2TS U3604 ( .A(n3031), .Y(n3032) );
  INVX2TS U3605 ( .A(n3270), .Y(n3271) );
  NAND2X1TS U3607 ( .A(read_reg[1]), .B(read_reg[0]), .Y(n4283) );
  CLKBUFX2TS U3608 ( .A(reset), .Y(n2896) );
  OAI21XLTS U3609 ( .A0(empty_reg), .A1(n4283), .B0(n2897), .Y(n4286) );
  OR2X1TS U3610 ( .A(n2896), .B(empty_reg), .Y(n4278) );
  CLKBUFX2TS U3611 ( .A(readReady), .Y(n2898) );
  CLKBUFX2TS U3612 ( .A(selectBit_SOUTH), .Y(n2899) );
  CLKBUFX2TS U3613 ( .A(selectBit_WEST), .Y(n2901) );
  CLKBUFX2TS U3614 ( .A(selectBit_EAST), .Y(n2903) );
  CLKBUFX2TS U3615 ( .A(selectBit_NORTH), .Y(n2904) );
  NAND2X1TS U3616 ( .A(empty_reg), .B(n2897), .Y(n4273) );
  CLKBUFX2TS U3617 ( .A(requesterAddressIn_SOUTH[0]), .Y(n2905) );
  CLKBUFX2TS U3618 ( .A(requesterAddressIn_WEST[0]), .Y(n2907) );
  CLKBUFX2TS U3619 ( .A(requesterAddressIn_EAST[0]), .Y(n2909) );
  OR2X2TS U3620 ( .A(n4273), .B(n4816), .Y(n5307) );
  INVX2TS U3621 ( .A(n5307), .Y(n5280) );
  CLKBUFX2TS U3622 ( .A(requesterAddressIn_NORTH[0]), .Y(n2910) );
  INVX2TS U3623 ( .A(n5305), .Y(n5290) );
  NOR3BX1TS U3624 ( .AN(n4816), .B(n4273), .C(n2911), .Y(n4932) );
  NOR3XLTS U3625 ( .A(read_reg[2]), .B(n5324), .C(n5325), .Y(n4875) );
  NOR3XLTS U3626 ( .A(read_reg[1]), .B(read_reg[2]), .C(n5325), .Y(n4803) );
  AOI22X1TS U3627 ( .A0(\requesterAddressbuffer[3][0] ), .A1(n4875), .B0(
        \requesterAddressbuffer[1][0] ), .B1(n2894), .Y(n2917) );
  NOR3X1TS U3628 ( .A(read_reg[0]), .B(n5329), .C(n5324), .Y(n5311) );
  NOR3XLTS U3629 ( .A(read_reg[1]), .B(n5329), .C(n5325), .Y(n4802) );
  AOI22X1TS U3630 ( .A0(\requesterAddressbuffer[6][0] ), .A1(n2893), .B0(
        \requesterAddressbuffer[5][0] ), .B1(n2892), .Y(n2916) );
  NOR3X1TS U3631 ( .A(read_reg[1]), .B(read_reg[0]), .C(n5329), .Y(n5249) );
  NOR3XLTS U3632 ( .A(n5324), .B(n5329), .C(n5325), .Y(n4884) );
  AOI22X1TS U3633 ( .A0(\requesterAddressbuffer[4][0] ), .A1(n5249), .B0(
        \requesterAddressbuffer[7][0] ), .B1(n2895), .Y(n2915) );
  NOR3XLTS U3634 ( .A(read_reg[2]), .B(read_reg[0]), .C(n5324), .Y(n2912) );
  BUFX3TS U3635 ( .A(n2912), .Y(n5310) );
  NOR3XLTS U3636 ( .A(read_reg[1]), .B(read_reg[2]), .C(read_reg[0]), .Y(n2913) );
  BUFX3TS U3637 ( .A(n2913), .Y(n5312) );
  AOI22X1TS U3638 ( .A0(\requesterAddressbuffer[2][0] ), .A1(n5310), .B0(
        \requesterAddressbuffer[0][0] ), .B1(n5312), .Y(n2914) );
  NAND4XLTS U3639 ( .A(n2917), .B(n2916), .C(n2915), .D(n2914), .Y(n2918) );
  AO22XLTS U3640 ( .A0(n4932), .A1(requesterAddressOut[0]), .B0(n2890), .B1(
        n2918), .Y(n2919) );
  CLKBUFX2TS U3641 ( .A(readRequesterAddress[0]), .Y(n2921) );
  NAND2X1TS U3642 ( .A(n2921), .B(n2922), .Y(n4898) );
  CLKBUFX2TS U3643 ( .A(requesterAddressIn_NORTH[3]), .Y(n2924) );
  CLKBUFX2TS U3644 ( .A(requesterAddressIn_WEST[3]), .Y(n2926) );
  CLKBUFX2TS U3645 ( .A(requesterAddressIn_SOUTH[3]), .Y(n2927) );
  INVX2TS U3646 ( .A(n5291), .Y(n5304) );
  CLKBUFX2TS U3647 ( .A(requesterAddressIn_EAST[3]), .Y(n2928) );
  AOI22X1TS U3648 ( .A0(\requesterAddressbuffer[3][3] ), .A1(n4875), .B0(
        \requesterAddressbuffer[1][3] ), .B1(n2894), .Y(n2932) );
  AOI22X1TS U3649 ( .A0(\requesterAddressbuffer[6][3] ), .A1(n2893), .B0(
        \requesterAddressbuffer[7][3] ), .B1(n2895), .Y(n2931) );
  AOI22X1TS U3650 ( .A0(\requesterAddressbuffer[0][3] ), .A1(n5312), .B0(
        \requesterAddressbuffer[5][3] ), .B1(n2892), .Y(n2930) );
  AOI22X1TS U3651 ( .A0(\requesterAddressbuffer[4][3] ), .A1(n5295), .B0(
        \requesterAddressbuffer[2][3] ), .B1(n5310), .Y(n2929) );
  NAND4XLTS U3652 ( .A(n2932), .B(n2931), .C(n2930), .D(n2929), .Y(n2933) );
  CLKBUFX2TS U3653 ( .A(readRequesterAddress[3]), .Y(n2936) );
  NAND2X1TS U3654 ( .A(n2936), .B(n2922), .Y(n4923) );
  ADDHXLTS U3655 ( .A(N373), .B(n4247), .CO(n2938), .S(n3609) );
  NAND2X1TS U3656 ( .A(n2898), .B(n5327), .Y(n3877) );
  NAND2X1TS U3657 ( .A(N374), .B(n5326), .Y(n2993) );
  NAND2X1TS U3658 ( .A(n2941), .B(n2940), .Y(n4809) );
  NAND2X1TS U3659 ( .A(n2904), .B(N373), .Y(n3316) );
  AOI2BB2X1TS U3660 ( .B0(N374), .B1(n3316), .A0N(n3316), .A1N(N374), .Y(n3619) );
  OAI22X1TS U3661 ( .A0(n2942), .A1(n5327), .B0(N373), .B1(n2904), .Y(n2945)
         );
  NAND2X1TS U3662 ( .A(n2945), .B(n2899), .Y(n3083) );
  XOR2X1TS U3663 ( .A(n2943), .B(n5326), .Y(n4502) );
  INVX2TS U3664 ( .A(n4502), .Y(n4503) );
  INVX2TS U3665 ( .A(n4462), .Y(n4463) );
  OAI21X1TS U3666 ( .A0(n2945), .A1(n2899), .B0(n3083), .Y(n3618) );
  INVX2TS U3667 ( .A(n3618), .Y(n3318) );
  INVX2TS U3668 ( .A(n4484), .Y(n4483) );
  OAI21X1TS U3669 ( .A0(n2946), .A1(n3619), .B0(n4483), .Y(n3090) );
  NAND2X1TS U3670 ( .A(n3318), .B(n3090), .Y(n4512) );
  AOI21X1TS U3671 ( .A0(n3107), .A1(n5326), .B0(n2948), .Y(n4513) );
  OAI32X1TS U3672 ( .A0(n3615), .A1(n3109), .A2(n2993), .B0(n4513), .B1(n3615), 
        .Y(n4518) );
  INVX2TS U3673 ( .A(n2956), .Y(n4519) );
  NAND2X2TS U3674 ( .A(n4517), .B(n4519), .Y(n3533) );
  CLKBUFX2TS U3675 ( .A(dataIn_WEST[23]), .Y(n2949) );
  INVX2TS U3676 ( .A(n2949), .Y(n4215) );
  CLKBUFX2TS U3677 ( .A(cacheDataOut[23]), .Y(n2950) );
  NOR3XLTS U3678 ( .A(n3877), .B(n3615), .C(n2993), .Y(n2951) );
  BUFX3TS U3679 ( .A(n2951), .Y(n4417) );
  AOI22X1TS U3680 ( .A0(n2950), .A1(n4417), .B0(\dataoutbuffer[2][23] ), .B1(
        n4728), .Y(n2961) );
  CLKBUFX2TS U3681 ( .A(dataIn_NORTH[23]), .Y(n2953) );
  INVX2TS U3682 ( .A(n3029), .Y(n3542) );
  CLKBUFX2TS U3683 ( .A(dataIn_EAST[23]), .Y(n2955) );
  OR2X2TS U3684 ( .A(n2956), .B(n4514), .Y(n3537) );
  CLKBUFX2TS U3685 ( .A(dataIn_SOUTH[23]), .Y(n2957) );
  OAI22X1TS U3686 ( .A0(n3542), .A1(n5217), .B0(n3537), .B1(n2958), .Y(n2959)
         );
  AOI21X1TS U3687 ( .A0(n2952), .A1(n2953), .B0(n2959), .Y(n2960) );
  CLKBUFX2TS U3688 ( .A(dataIn_SOUTH[13]), .Y(n2962) );
  CLKBUFX2TS U3689 ( .A(cacheDataOut[13]), .Y(n2964) );
  AOI22X1TS U3690 ( .A0(n2964), .A1(n4417), .B0(\dataoutbuffer[2][13] ), .B1(
        n4728), .Y(n2971) );
  CLKBUFX2TS U3691 ( .A(dataIn_NORTH[13]), .Y(n2965) );
  CLKBUFX2TS U3692 ( .A(dataIn_WEST[13]), .Y(n2967) );
  INVX2TS U3693 ( .A(n2967), .Y(n4113) );
  CLKBUFX2TS U3694 ( .A(dataIn_EAST[13]), .Y(n2968) );
  INVX2TS U3695 ( .A(n2968), .Y(n4117) );
  OAI22X1TS U3696 ( .A0(n3533), .A1(n4113), .B0(n3542), .B1(n4117), .Y(n2969)
         );
  AOI21X1TS U3697 ( .A0(n2952), .A1(n2965), .B0(n2969), .Y(n2970) );
  CLKBUFX2TS U3698 ( .A(destinationAddressIn_EAST[7]), .Y(n2972) );
  CLKBUFX2TS U3699 ( .A(destinationAddressIn_SOUTH[7]), .Y(n2974) );
  AOI22X1TS U3700 ( .A0(n2974), .A1(n4730), .B0(
        \destinationAddressbuffer[2][7] ), .B1(n4728), .Y(n2978) );
  CLKBUFX2TS U3701 ( .A(destinationAddressIn_NORTH[7]), .Y(n2975) );
  CLKBUFX2TS U3702 ( .A(destinationAddressIn_WEST[7]), .Y(n2976) );
  AOI22X1TS U3703 ( .A0(n2952), .A1(n2975), .B0(n4731), .B1(n2976), .Y(n2977)
         );
  CLKBUFX2TS U3704 ( .A(writeIn_EAST), .Y(n2979) );
  INVX2TS U3705 ( .A(n2979), .Y(n4817) );
  CLKBUFX2TS U3706 ( .A(writeIn_SOUTH), .Y(n2980) );
  AOI22X1TS U3707 ( .A0(n2980), .A1(n4730), .B0(writeOutbuffer[2]), .B1(n4728), 
        .Y(n2986) );
  CLKBUFX2TS U3708 ( .A(writeIn_NORTH), .Y(n2982) );
  CLKBUFX2TS U3709 ( .A(writeIn_WEST), .Y(n2983) );
  AOI22X1TS U3710 ( .A0(n2952), .A1(n2982), .B0(n4731), .B1(n2983), .Y(n2985)
         );
  CLKBUFX2TS U3711 ( .A(destinationAddressIn_EAST[8]), .Y(n2987) );
  INVX2TS U3712 ( .A(n2987), .Y(n4235) );
  CLKBUFX2TS U3713 ( .A(destinationAddressIn_SOUTH[8]), .Y(n2988) );
  AOI22X1TS U3714 ( .A0(n2988), .A1(n4730), .B0(
        \destinationAddressbuffer[2][8] ), .B1(n4728), .Y(n2992) );
  CLKBUFX2TS U3715 ( .A(destinationAddressIn_NORTH[8]), .Y(n2989) );
  CLKBUFX2TS U3716 ( .A(destinationAddressIn_WEST[8]), .Y(n2990) );
  AOI22X1TS U3717 ( .A0(n2952), .A1(n2989), .B0(n4731), .B1(n2990), .Y(n2991)
         );
  NAND2X1TS U3718 ( .A(N373), .B(n2898), .Y(n3614) );
  OAI31X1TS U3719 ( .A0(n3318), .A1(n3619), .A2(n3381), .B0(n4501), .Y(n4506)
         );
  OAI32X1TS U3720 ( .A0(n3615), .A1(n2994), .A2(n2993), .B0(n2995), .B1(n3615), 
        .Y(n4511) );
  NAND2X1TS U3721 ( .A(n2995), .B(n4511), .Y(n2998) );
  INVX2TS U3722 ( .A(n2974), .Y(n4192) );
  NAND2X1TS U3723 ( .A(n4511), .B(n3231), .Y(n4508) );
  NOR2XLTS U3724 ( .A(n3318), .B(n3619), .Y(n2997) );
  NAND2X1TS U3725 ( .A(n2997), .B(n4501), .Y(n4504) );
  AOI22X1TS U3726 ( .A0(n2972), .A1(n4696), .B0(
        \destinationAddressbuffer[3][7] ), .B1(n4701), .Y(n3000) );
  AOI22X1TS U3727 ( .A0(n4703), .A1(n2975), .B0(n4687), .B1(n2976), .Y(n2999)
         );
  CLKBUFX2TS U3728 ( .A(destinationAddressIn_SOUTH[6]), .Y(n3001) );
  INVX2TS U3729 ( .A(n3001), .Y(n4244) );
  CLKBUFX2TS U3730 ( .A(destinationAddressIn_EAST[6]), .Y(n3002) );
  AOI22X1TS U3731 ( .A0(n3002), .A1(n4696), .B0(
        \destinationAddressbuffer[3][6] ), .B1(n4701), .Y(n3007) );
  CLKBUFX2TS U3732 ( .A(destinationAddressIn_NORTH[6]), .Y(n3004) );
  CLKBUFX2TS U3733 ( .A(destinationAddressIn_WEST[6]), .Y(n3005) );
  AOI22X1TS U3734 ( .A0(n4703), .A1(n3004), .B0(n4687), .B1(n3005), .Y(n3006)
         );
  CLKBUFX2TS U3735 ( .A(dataIn_SOUTH[1]), .Y(n3008) );
  CLKBUFX2TS U3736 ( .A(cacheDataOut[1]), .Y(n3010) );
  AOI22X1TS U3737 ( .A0(n3010), .A1(n4417), .B0(\dataoutbuffer[2][1] ), .B1(
        n4728), .Y(n3016) );
  CLKBUFX2TS U3738 ( .A(dataIn_NORTH[1]), .Y(n3011) );
  CLKBUFX2TS U3739 ( .A(dataIn_WEST[1]), .Y(n3012) );
  INVX2TS U3740 ( .A(n3012), .Y(n4084) );
  CLKBUFX2TS U3741 ( .A(dataIn_EAST[1]), .Y(n3013) );
  INVX2TS U3742 ( .A(n3013), .Y(n4990) );
  OAI22X1TS U3743 ( .A0(n3533), .A1(n4084), .B0(n3542), .B1(n4990), .Y(n3014)
         );
  AOI21X1TS U3744 ( .A0(n2952), .A1(n3011), .B0(n3014), .Y(n3015) );
  CLKBUFX2TS U3745 ( .A(dataIn_SOUTH[0]), .Y(n3017) );
  CLKBUFX2TS U3746 ( .A(cacheDataOut[0]), .Y(n3019) );
  AOI22X1TS U3747 ( .A0(n3019), .A1(n4417), .B0(\dataoutbuffer[2][0] ), .B1(
        n4728), .Y(n3026) );
  CLKBUFX2TS U3748 ( .A(dataIn_NORTH[0]), .Y(n3020) );
  CLKBUFX2TS U3749 ( .A(dataIn_WEST[0]), .Y(n3021) );
  INVX2TS U3750 ( .A(n3021), .Y(n4118) );
  CLKBUFX2TS U3751 ( .A(dataIn_EAST[0]), .Y(n3022) );
  OAI22X1TS U3752 ( .A0(n3533), .A1(n4118), .B0(n3542), .B1(n3023), .Y(n3024)
         );
  AOI21X1TS U3753 ( .A0(n2952), .A1(n3020), .B0(n3024), .Y(n3025) );
  CLKBUFX2TS U3754 ( .A(destinationAddressIn_SOUTH[10]), .Y(n3027) );
  INVX2TS U3755 ( .A(n3027), .Y(n4195) );
  CLKBUFX2TS U3756 ( .A(destinationAddressIn_EAST[10]), .Y(n3028) );
  CLKBUFX2TS U3757 ( .A(n3029), .Y(n4729) );
  AOI22X1TS U3758 ( .A0(n3028), .A1(n4729), .B0(
        \destinationAddressbuffer[2][10] ), .B1(n4728), .Y(n3034) );
  CLKBUFX2TS U3759 ( .A(destinationAddressIn_NORTH[10]), .Y(n3030) );
  CLKBUFX2TS U3760 ( .A(destinationAddressIn_WEST[10]), .Y(n3031) );
  AOI22X1TS U3761 ( .A0(n2952), .A1(n3030), .B0(n4731), .B1(n3031), .Y(n3033)
         );
  CLKBUFX2TS U3762 ( .A(destinationAddressIn_EAST[12]), .Y(n3035) );
  CLKBUFX2TS U3763 ( .A(destinationAddressIn_SOUTH[12]), .Y(n3037) );
  AOI22X1TS U3764 ( .A0(n3037), .A1(n4730), .B0(
        \destinationAddressbuffer[2][12] ), .B1(n4728), .Y(n3041) );
  CLKBUFX2TS U3765 ( .A(destinationAddressIn_NORTH[12]), .Y(n3038) );
  CLKBUFX2TS U3766 ( .A(destinationAddressIn_WEST[12]), .Y(n3039) );
  AOI22X1TS U3767 ( .A0(n2952), .A1(n3038), .B0(n4731), .B1(n3039), .Y(n3040)
         );
  CLKBUFX2TS U3768 ( .A(dataIn_EAST[16]), .Y(n3042) );
  CLKBUFX2TS U3769 ( .A(cacheDataOut[16]), .Y(n3043) );
  AOI22X1TS U3770 ( .A0(n3043), .A1(n4417), .B0(\dataoutbuffer[2][16] ), .B1(
        n4728), .Y(n3050) );
  CLKBUFX2TS U3771 ( .A(dataIn_NORTH[16]), .Y(n3044) );
  CLKBUFX2TS U3772 ( .A(dataIn_WEST[16]), .Y(n3046) );
  INVX2TS U3773 ( .A(n3046), .Y(n4219) );
  CLKBUFX2TS U3774 ( .A(dataIn_SOUTH[16]), .Y(n3047) );
  INVX2TS U3775 ( .A(n3047), .Y(n5146) );
  OAI22X1TS U3776 ( .A0(n3533), .A1(n4219), .B0(n3537), .B1(n5146), .Y(n3048)
         );
  AOI21X1TS U3777 ( .A0(n2952), .A1(n3044), .B0(n3048), .Y(n3049) );
  CLKBUFX2TS U3778 ( .A(dataIn_EAST[8]), .Y(n3051) );
  INVX2TS U3779 ( .A(n3051), .Y(n4166) );
  CLKBUFX2TS U3780 ( .A(cacheDataOut[8]), .Y(n3052) );
  AOI22X1TS U3781 ( .A0(n3052), .A1(n4417), .B0(\dataoutbuffer[2][8] ), .B1(
        n4728), .Y(n3059) );
  CLKBUFX2TS U3782 ( .A(dataIn_NORTH[8]), .Y(n3053) );
  CLKBUFX2TS U3783 ( .A(dataIn_WEST[8]), .Y(n3054) );
  INVX2TS U3784 ( .A(n3054), .Y(n4170) );
  CLKBUFX2TS U3785 ( .A(dataIn_SOUTH[8]), .Y(n3055) );
  OAI22X1TS U3786 ( .A0(n3533), .A1(n4170), .B0(n3537), .B1(n3056), .Y(n3057)
         );
  AOI21X1TS U3787 ( .A0(n2952), .A1(n3053), .B0(n3057), .Y(n3058) );
  CLKBUFX2TS U3788 ( .A(dataIn_EAST[9]), .Y(n3060) );
  CLKBUFX2TS U3789 ( .A(cacheDataOut[9]), .Y(n3061) );
  AOI22X1TS U3790 ( .A0(n3061), .A1(n4417), .B0(\dataoutbuffer[2][9] ), .B1(
        n4728), .Y(n3068) );
  CLKBUFX2TS U3791 ( .A(dataIn_NORTH[9]), .Y(n3062) );
  CLKBUFX2TS U3792 ( .A(dataIn_WEST[9]), .Y(n3063) );
  CLKBUFX2TS U3793 ( .A(dataIn_SOUTH[9]), .Y(n3065) );
  OAI22X1TS U3794 ( .A0(n3533), .A1(n3064), .B0(n3537), .B1(n5075), .Y(n3066)
         );
  AOI21X1TS U3795 ( .A0(n2952), .A1(n3062), .B0(n3066), .Y(n3067) );
  INVX2TS U3796 ( .A(n3037), .Y(n4189) );
  AOI22X1TS U3797 ( .A0(n3039), .A1(n4687), .B0(
        \destinationAddressbuffer[3][12] ), .B1(n4701), .Y(n3070) );
  AOI22X1TS U3798 ( .A0(n4703), .A1(n3038), .B0(n4696), .B1(n3035), .Y(n3069)
         );
  AOI22X1TS U3799 ( .A0(n3030), .A1(n4703), .B0(
        \destinationAddressbuffer[3][10] ), .B1(n4701), .Y(n3072) );
  AOI22X1TS U3800 ( .A0(n4696), .A1(n3028), .B0(n4687), .B1(n3031), .Y(n3071)
         );
  CLKBUFX2TS U3801 ( .A(destinationAddressIn_WEST[11]), .Y(n3073) );
  CLKBUFX2TS U3802 ( .A(destinationAddressIn_EAST[11]), .Y(n3075) );
  AOI22X1TS U3803 ( .A0(n3075), .A1(n4729), .B0(
        \destinationAddressbuffer[2][11] ), .B1(n4728), .Y(n3080) );
  CLKBUFX2TS U3804 ( .A(destinationAddressIn_NORTH[11]), .Y(n3077) );
  CLKBUFX2TS U3805 ( .A(destinationAddressIn_SOUTH[11]), .Y(n3078) );
  AOI22X1TS U3806 ( .A0(n2952), .A1(n3077), .B0(n4730), .B1(n3078), .Y(n3079)
         );
  AOI22X1TS U3807 ( .A0(n3004), .A1(n2952), .B0(
        \destinationAddressbuffer[2][6] ), .B1(n4728), .Y(n3082) );
  AOI22X1TS U3808 ( .A0(n4731), .A1(n3005), .B0(n4730), .B1(n3001), .Y(n3081)
         );
  INVX2TS U3809 ( .A(n3317), .Y(n3607) );
  NAND2X1TS U3810 ( .A(n5323), .B(n5326), .Y(n3384) );
  OAI31X1TS U3811 ( .A0(n3618), .A1(n3090), .A2(n3381), .B0(n4530), .Y(n3084)
         );
  OAI32X1TS U3812 ( .A0(n3615), .A1(n3109), .A2(n3384), .B0(n3085), .B1(n3615), 
        .Y(n4537) );
  OR2X2TS U3813 ( .A(n4530), .B(n4535), .Y(n3700) );
  OR2X2TS U3814 ( .A(n4535), .B(n4531), .Y(n3698) );
  AOI22X1TS U3815 ( .A0(n3027), .A1(n4789), .B0(
        \destinationAddressbuffer[0][10] ), .B1(n4787), .Y(n3087) );
  NOR2X2TS U3816 ( .A(n4532), .B(n4535), .Y(n4790) );
  NOR2XLTS U3817 ( .A(n3090), .B(n3618), .Y(n3093) );
  NAND2X1TS U3818 ( .A(n3093), .B(n4530), .Y(n4529) );
  NOR2X2TS U3819 ( .A(n4535), .B(n4529), .Y(n4782) );
  AOI22X1TS U3820 ( .A0(n4790), .A1(n3030), .B0(n4782), .B1(n3028), .Y(n3086)
         );
  NAND2X1TS U3821 ( .A(N375), .B(n5323), .Y(n3708) );
  OAI31X1TS U3822 ( .A0(n3618), .A1(n3090), .A2(n3610), .B0(n4493), .Y(n3092)
         );
  OAI32X1TS U3823 ( .A0(n3615), .A1(n3109), .A2(n3708), .B0(n4496), .B1(n3615), 
        .Y(n4500) );
  NOR2X2TS U3824 ( .A(n4493), .B(n4495), .Y(n4666) );
  AOI22X1TS U3825 ( .A0(n2976), .A1(n4666), .B0(
        \destinationAddressbuffer[4][7] ), .B1(n4671), .Y(n3095) );
  NAND2X1TS U3826 ( .A(n3093), .B(n4493), .Y(n4492) );
  AOI22X1TS U3827 ( .A0(n4672), .A1(n2972), .B0(n4674), .B1(n2975), .Y(n3094)
         );
  AOI22X1TS U3828 ( .A0(n3002), .A1(n4672), .B0(
        \destinationAddressbuffer[4][6] ), .B1(n4671), .Y(n3097) );
  AOI22X1TS U3829 ( .A0(n4674), .A1(n3004), .B0(n4666), .B1(n3005), .Y(n3096)
         );
  AOI22X1TS U3830 ( .A0(n3035), .A1(n4672), .B0(
        \destinationAddressbuffer[4][12] ), .B1(n4671), .Y(n3099) );
  AOI22X1TS U3831 ( .A0(n4674), .A1(n3038), .B0(n4666), .B1(n3039), .Y(n3098)
         );
  AOI22X1TS U3832 ( .A0(n3028), .A1(n4672), .B0(
        \destinationAddressbuffer[4][10] ), .B1(n4671), .Y(n3101) );
  AOI22X1TS U3833 ( .A0(n4674), .A1(n3030), .B0(n4666), .B1(n3031), .Y(n3100)
         );
  AOI22X1TS U3834 ( .A0(n3005), .A1(n4788), .B0(
        \destinationAddressbuffer[0][6] ), .B1(n4787), .Y(n3103) );
  AOI22X1TS U3835 ( .A0(n4790), .A1(n3004), .B0(n4782), .B1(n3002), .Y(n3102)
         );
  AOI22X1TS U3836 ( .A0(n3075), .A1(n4782), .B0(
        \destinationAddressbuffer[0][11] ), .B1(n4787), .Y(n3105) );
  AOI22X1TS U3837 ( .A0(n4790), .A1(n3077), .B0(n4789), .B1(n3078), .Y(n3104)
         );
  NAND2X1TS U3838 ( .A(N374), .B(N375), .Y(n3876) );
  NAND2X1TS U3839 ( .A(N375), .B(n3107), .Y(n4480) );
  INVX2TS U3840 ( .A(n3111), .Y(n4478) );
  OAI32X1TS U3841 ( .A0(n3615), .A1(n3109), .A2(n3876), .B0(n4478), .B1(n3615), 
        .Y(n4482) );
  OR2X2TS U3842 ( .A(n4475), .B(n4477), .Y(n4076) );
  AOI22X1TS U3843 ( .A0(n3078), .A1(n4615), .B0(
        \destinationAddressbuffer[6][11] ), .B1(n4612), .Y(n3113) );
  NOR2X2TS U3844 ( .A(n3111), .B(n4477), .Y(n4614) );
  AOI22X1TS U3845 ( .A0(n4613), .A1(n3075), .B0(n4614), .B1(n3077), .Y(n3112)
         );
  INVX2TS U3846 ( .A(n4703), .Y(n3579) );
  CLKBUFX2TS U3847 ( .A(destinationAddressIn_NORTH[13]), .Y(n3114) );
  INVX2TS U3848 ( .A(n3114), .Y(n3893) );
  CLKBUFX2TS U3849 ( .A(destinationAddressIn_WEST[13]), .Y(n3115) );
  AOI22X1TS U3850 ( .A0(n3115), .A1(n4687), .B0(
        \destinationAddressbuffer[3][13] ), .B1(n4701), .Y(n3119) );
  CLKBUFX2TS U3851 ( .A(destinationAddressIn_EAST[13]), .Y(n3116) );
  CLKBUFX2TS U3852 ( .A(destinationAddressIn_SOUTH[13]), .Y(n3117) );
  AOI22X1TS U3853 ( .A0(n4696), .A1(n3116), .B0(n4702), .B1(n3117), .Y(n3118)
         );
  CLKBUFX2TS U3854 ( .A(destinationAddressIn_NORTH[9]), .Y(n3120) );
  INVX2TS U3855 ( .A(n3120), .Y(n3890) );
  CLKBUFX2TS U3856 ( .A(destinationAddressIn_SOUTH[9]), .Y(n3121) );
  AOI22X1TS U3857 ( .A0(n3121), .A1(n4702), .B0(
        \destinationAddressbuffer[3][9] ), .B1(n4701), .Y(n3125) );
  CLKBUFX2TS U3858 ( .A(destinationAddressIn_EAST[9]), .Y(n3122) );
  CLKBUFX2TS U3859 ( .A(destinationAddressIn_WEST[9]), .Y(n3123) );
  AOI22X1TS U3860 ( .A0(n4696), .A1(n3122), .B0(n4687), .B1(n3123), .Y(n3124)
         );
  CLKBUFX2TS U3861 ( .A(dataIn_NORTH[29]), .Y(n3126) );
  CLKBUFX2TS U3862 ( .A(cacheDataOut[29]), .Y(n3128) );
  AOI22X1TS U3863 ( .A0(n3128), .A1(n4417), .B0(\dataoutbuffer[2][29] ), .B1(
        n4728), .Y(n3135) );
  CLKBUFX2TS U3864 ( .A(dataIn_SOUTH[29]), .Y(n3129) );
  CLKBUFX2TS U3865 ( .A(dataIn_WEST[29]), .Y(n3131) );
  INVX2TS U3866 ( .A(n3131), .Y(n4175) );
  CLKBUFX2TS U3867 ( .A(dataIn_EAST[29]), .Y(n3132) );
  INVX2TS U3868 ( .A(n3132), .Y(n4171) );
  OAI22X1TS U3869 ( .A0(n3533), .A1(n4175), .B0(n3542), .B1(n4171), .Y(n3133)
         );
  AOI21X1TS U3870 ( .A0(n4730), .A1(n3129), .B0(n3133), .Y(n3134) );
  CLKBUFX2TS U3871 ( .A(dataIn_NORTH[31]), .Y(n3136) );
  CLKBUFX2TS U3872 ( .A(cacheDataOut[31]), .Y(n3137) );
  AOI22X1TS U3873 ( .A0(n3137), .A1(n4417), .B0(\dataoutbuffer[2][31] ), .B1(
        n4728), .Y(n3144) );
  CLKBUFX2TS U3874 ( .A(dataIn_SOUTH[31]), .Y(n3138) );
  CLKBUFX2TS U3875 ( .A(dataIn_WEST[31]), .Y(n3139) );
  CLKBUFX2TS U3876 ( .A(dataIn_EAST[31]), .Y(n3141) );
  OAI22X1TS U3877 ( .A0(n3533), .A1(n3140), .B0(n3542), .B1(n5308), .Y(n3142)
         );
  AOI21X1TS U3878 ( .A0(n4730), .A1(n3138), .B0(n3142), .Y(n3143) );
  CLKBUFX2TS U3879 ( .A(dataIn_NORTH[24]), .Y(n3145) );
  INVX2TS U3880 ( .A(n3145), .Y(n5228) );
  CLKBUFX2TS U3881 ( .A(cacheDataOut[24]), .Y(n3146) );
  AOI22X1TS U3882 ( .A0(n3146), .A1(n4417), .B0(\dataoutbuffer[2][24] ), .B1(
        n4728), .Y(n3153) );
  CLKBUFX2TS U3883 ( .A(dataIn_WEST[24]), .Y(n3147) );
  CLKBUFX2TS U3884 ( .A(dataIn_EAST[24]), .Y(n3148) );
  INVX2TS U3885 ( .A(n3148), .Y(n5227) );
  CLKBUFX2TS U3886 ( .A(dataIn_SOUTH[24]), .Y(n3149) );
  OAI22X1TS U3887 ( .A0(n3542), .A1(n5227), .B0(n3537), .B1(n3150), .Y(n3151)
         );
  AOI21X1TS U3888 ( .A0(n4731), .A1(n3147), .B0(n3151), .Y(n3152) );
  CLKBUFX2TS U3889 ( .A(dataIn_NORTH[10]), .Y(n3154) );
  INVX2TS U3890 ( .A(n3154), .Y(n4022) );
  CLKBUFX2TS U3891 ( .A(cacheDataOut[10]), .Y(n3155) );
  AOI22X1TS U3892 ( .A0(n3155), .A1(n4417), .B0(\dataoutbuffer[2][10] ), .B1(
        n4728), .Y(n3162) );
  CLKBUFX2TS U3893 ( .A(dataIn_WEST[10]), .Y(n3156) );
  CLKBUFX2TS U3894 ( .A(dataIn_EAST[10]), .Y(n3158) );
  CLKBUFX2TS U3895 ( .A(dataIn_SOUTH[10]), .Y(n3159) );
  INVX2TS U3896 ( .A(n3159), .Y(n5086) );
  OAI22X1TS U3897 ( .A0(n3542), .A1(n5085), .B0(n3537), .B1(n5086), .Y(n3160)
         );
  AOI21X1TS U3898 ( .A0(n4731), .A1(n3156), .B0(n3160), .Y(n3161) );
  CLKBUFX2TS U3899 ( .A(dataIn_NORTH[4]), .Y(n3163) );
  INVX2TS U3900 ( .A(n3163), .Y(n5022) );
  CLKBUFX2TS U3901 ( .A(cacheDataOut[4]), .Y(n3164) );
  AOI22X1TS U3902 ( .A0(n3164), .A1(n4417), .B0(\dataoutbuffer[2][4] ), .B1(
        n4728), .Y(n3171) );
  CLKBUFX2TS U3903 ( .A(dataIn_SOUTH[4]), .Y(n3165) );
  CLKBUFX2TS U3904 ( .A(dataIn_WEST[4]), .Y(n3167) );
  INVX2TS U3905 ( .A(n3167), .Y(n4136) );
  CLKBUFX2TS U3906 ( .A(dataIn_EAST[4]), .Y(n3168) );
  OAI22X1TS U3907 ( .A0(n3533), .A1(n4136), .B0(n3542), .B1(n5023), .Y(n3169)
         );
  AOI21X1TS U3908 ( .A0(n4730), .A1(n3165), .B0(n3169), .Y(n3170) );
  AOI22X1TS U3909 ( .A0(n3122), .A1(n4729), .B0(
        \destinationAddressbuffer[2][9] ), .B1(n4728), .Y(n3173) );
  AOI22X1TS U3910 ( .A0(n4731), .A1(n3123), .B0(n4730), .B1(n3121), .Y(n3172)
         );
  AOI22X1TS U3911 ( .A0(n3117), .A1(n4730), .B0(
        \destinationAddressbuffer[2][13] ), .B1(n4728), .Y(n3175) );
  AOI22X1TS U3912 ( .A0(n4731), .A1(n3115), .B0(n4729), .B1(n3116), .Y(n3174)
         );
  AOI22X1TS U3913 ( .A0(n3038), .A1(n4790), .B0(
        \destinationAddressbuffer[0][12] ), .B1(n4787), .Y(n3177) );
  AOI22X1TS U3914 ( .A0(n4788), .A1(n3039), .B0(n4789), .B1(n3037), .Y(n3176)
         );
  NOR3XLTS U3915 ( .A(n3877), .B(n3615), .C(n3384), .Y(n3178) );
  BUFX3TS U3916 ( .A(n3178), .Y(n4455) );
  AOI22X1TS U3917 ( .A0(n3052), .A1(n4455), .B0(\dataoutbuffer[0][8] ), .B1(
        n4787), .Y(n3181) );
  OAI22X1TS U3918 ( .A0(n3700), .A1(n4170), .B0(n3698), .B1(n3056), .Y(n3179)
         );
  AOI21X1TS U3919 ( .A0(n4790), .A1(n3053), .B0(n3179), .Y(n3180) );
  AOI22X1TS U3920 ( .A0(n2988), .A1(n4789), .B0(
        \destinationAddressbuffer[0][8] ), .B1(n4787), .Y(n3183) );
  AOI22X1TS U3921 ( .A0(n4788), .A1(n2990), .B0(n4790), .B1(n2989), .Y(n3182)
         );
  AOI22X1TS U3922 ( .A0(n2975), .A1(n4790), .B0(
        \destinationAddressbuffer[0][7] ), .B1(n4787), .Y(n3185) );
  AOI22X1TS U3923 ( .A0(n4788), .A1(n2976), .B0(n4789), .B1(n2974), .Y(n3184)
         );
  AOI22X1TS U3924 ( .A0(n3043), .A1(n4455), .B0(\dataoutbuffer[0][16] ), .B1(
        n4787), .Y(n3188) );
  OAI22X1TS U3925 ( .A0(n3700), .A1(n4219), .B0(n3698), .B1(n5146), .Y(n3186)
         );
  AOI21X1TS U3926 ( .A0(n4790), .A1(n3044), .B0(n3186), .Y(n3187) );
  AOI22X1TS U3927 ( .A0(n2982), .A1(n4790), .B0(writeOutbuffer[0]), .B1(n4787), 
        .Y(n3190) );
  AOI22X1TS U3928 ( .A0(n4788), .A1(n2983), .B0(n4789), .B1(n2980), .Y(n3189)
         );
  INVX2TS U3929 ( .A(n4696), .Y(n3575) );
  AOI22X1TS U3930 ( .A0(n2990), .A1(n4687), .B0(
        \destinationAddressbuffer[3][8] ), .B1(n4701), .Y(n3192) );
  AOI22X1TS U3931 ( .A0(n4703), .A1(n2989), .B0(n4702), .B1(n2988), .Y(n3191)
         );
  AOI22X1TS U3932 ( .A0(n2983), .A1(n4687), .B0(writeOutbuffer[3]), .B1(n4701), 
        .Y(n3194) );
  AOI22X1TS U3933 ( .A0(n4703), .A1(n2982), .B0(n4702), .B1(n2980), .Y(n3193)
         );
  INVX2TS U3934 ( .A(n4687), .Y(n3574) );
  AOI22X1TS U3935 ( .A0(n3078), .A1(n4702), .B0(
        \destinationAddressbuffer[3][11] ), .B1(n4701), .Y(n3196) );
  AOI22X1TS U3936 ( .A0(n4703), .A1(n3077), .B0(n4696), .B1(n3075), .Y(n3195)
         );
  CLKBUFX2TS U3937 ( .A(dataIn_NORTH[7]), .Y(n3197) );
  CLKBUFX2TS U3938 ( .A(cacheDataOut[7]), .Y(n3198) );
  AOI22X1TS U3939 ( .A0(n3198), .A1(n4455), .B0(\dataoutbuffer[0][7] ), .B1(
        n4787), .Y(n3205) );
  CLKBUFX2TS U3940 ( .A(dataIn_EAST[7]), .Y(n3199) );
  CLKBUFX2TS U3941 ( .A(dataIn_WEST[7]), .Y(n3200) );
  CLKBUFX2TS U3942 ( .A(dataIn_SOUTH[7]), .Y(n3202) );
  OAI22X1TS U3943 ( .A0(n3700), .A1(n3201), .B0(n3698), .B1(n5055), .Y(n3203)
         );
  AOI21X1TS U3944 ( .A0(n4782), .A1(n3199), .B0(n3203), .Y(n3204) );
  CLKBUFX2TS U3945 ( .A(dataIn_NORTH[17]), .Y(n3206) );
  INVX2TS U3946 ( .A(n3206), .Y(n5156) );
  CLKBUFX2TS U3947 ( .A(cacheDataOut[17]), .Y(n3207) );
  AOI22X1TS U3948 ( .A0(n3207), .A1(n4455), .B0(\dataoutbuffer[0][17] ), .B1(
        n4787), .Y(n3214) );
  CLKBUFX2TS U3949 ( .A(dataIn_EAST[17]), .Y(n3208) );
  CLKBUFX2TS U3950 ( .A(dataIn_WEST[17]), .Y(n3210) );
  INVX2TS U3951 ( .A(n3210), .Y(n4206) );
  CLKBUFX2TS U3952 ( .A(dataIn_SOUTH[17]), .Y(n3211) );
  INVX2TS U3953 ( .A(n3211), .Y(n4207) );
  OAI22X1TS U3954 ( .A0(n3700), .A1(n4206), .B0(n3698), .B1(n4207), .Y(n3212)
         );
  AOI21X1TS U3955 ( .A0(n4782), .A1(n3208), .B0(n3212), .Y(n3213) );
  AOI22X1TS U3956 ( .A0(n3115), .A1(n4788), .B0(
        \destinationAddressbuffer[0][13] ), .B1(n4787), .Y(n3216) );
  AOI22X1TS U3957 ( .A0(n4782), .A1(n3116), .B0(n4789), .B1(n3117), .Y(n3215)
         );
  AOI22X1TS U3958 ( .A0(n3123), .A1(n4788), .B0(
        \destinationAddressbuffer[0][9] ), .B1(n4787), .Y(n3218) );
  AOI22X1TS U3959 ( .A0(n4782), .A1(n3122), .B0(n4789), .B1(n3121), .Y(n3217)
         );
  INVX2TS U3960 ( .A(n4672), .Y(n3827) );
  AOI22X1TS U3961 ( .A0(n2982), .A1(n4674), .B0(writeOutbuffer[4]), .B1(n4671), 
        .Y(n3220) );
  AOI22X1TS U3962 ( .A0(n4666), .A1(n2983), .B0(n4673), .B1(n2980), .Y(n3219)
         );
  AOI22X1TS U3963 ( .A0(n2990), .A1(n4666), .B0(
        \destinationAddressbuffer[4][8] ), .B1(n4671), .Y(n3222) );
  AOI22X1TS U3964 ( .A0(n4674), .A1(n2989), .B0(n4673), .B1(n2988), .Y(n3221)
         );
  INVX2TS U3965 ( .A(n4666), .Y(n3831) );
  AOI22X1TS U3966 ( .A0(n3075), .A1(n4672), .B0(
        \destinationAddressbuffer[4][11] ), .B1(n4671), .Y(n3224) );
  AOI22X1TS U3967 ( .A0(n4674), .A1(n3077), .B0(n4673), .B1(n3078), .Y(n3223)
         );
  INVX2TS U3968 ( .A(n4674), .Y(n3826) );
  AOI22X1TS U3969 ( .A0(n3123), .A1(n4666), .B0(
        \destinationAddressbuffer[4][9] ), .B1(n4671), .Y(n3226) );
  AOI22X1TS U3970 ( .A0(n4672), .A1(n3122), .B0(n4673), .B1(n3121), .Y(n3225)
         );
  AOI22X1TS U3971 ( .A0(n3117), .A1(n4673), .B0(
        \destinationAddressbuffer[4][13] ), .B1(n4671), .Y(n3228) );
  AOI22X1TS U3972 ( .A0(n4672), .A1(n3116), .B0(n4666), .B1(n3115), .Y(n3227)
         );
  CLKBUFX2TS U3973 ( .A(dataIn_WEST[25]), .Y(n3229) );
  INVX2TS U3974 ( .A(n3229), .Y(n4183) );
  CLKBUFX2TS U3975 ( .A(cacheDataOut[25]), .Y(n3230) );
  AOI22X1TS U3976 ( .A0(n3230), .A1(n3232), .B0(\dataoutbuffer[3][25] ), .B1(
        n4701), .Y(n3239) );
  CLKBUFX2TS U3977 ( .A(dataIn_EAST[25]), .Y(n3233) );
  CLKBUFX2TS U3978 ( .A(dataIn_NORTH[25]), .Y(n3234) );
  INVX2TS U3979 ( .A(n3234), .Y(n5238) );
  CLKBUFX2TS U3980 ( .A(dataIn_SOUTH[25]), .Y(n3235) );
  OAI22X1TS U3981 ( .A0(n3579), .A1(n5238), .B0(n3567), .B1(n3236), .Y(n3237)
         );
  AOI21X1TS U3982 ( .A0(n4696), .A1(n3233), .B0(n3237), .Y(n3238) );
  INVX2TS U3983 ( .A(n3147), .Y(n4179) );
  AOI22X1TS U3984 ( .A0(n3146), .A1(n3232), .B0(\dataoutbuffer[3][24] ), .B1(
        n4701), .Y(n3242) );
  OAI22X1TS U3985 ( .A0(n3579), .A1(n5228), .B0(n3567), .B1(n3150), .Y(n3240)
         );
  AOI21X1TS U3986 ( .A0(n4696), .A1(n3148), .B0(n3240), .Y(n3241) );
  CLKBUFX2TS U3987 ( .A(dataIn_EAST[20]), .Y(n3243) );
  CLKBUFX2TS U3988 ( .A(cacheDataOut[20]), .Y(n3244) );
  AOI22X1TS U3989 ( .A0(n3244), .A1(n3232), .B0(\dataoutbuffer[3][20] ), .B1(
        n4701), .Y(n3252) );
  CLKBUFX2TS U3990 ( .A(dataIn_WEST[20]), .Y(n3245) );
  CLKBUFX2TS U3991 ( .A(dataIn_NORTH[20]), .Y(n3247) );
  CLKBUFX2TS U3992 ( .A(dataIn_SOUTH[20]), .Y(n3249) );
  INVX2TS U3993 ( .A(n3249), .Y(n5187) );
  OAI22X1TS U3994 ( .A0(n3579), .A1(n3248), .B0(n3567), .B1(n5187), .Y(n3250)
         );
  AOI21X1TS U3995 ( .A0(n4687), .A1(n3245), .B0(n3250), .Y(n3251) );
  AOI22X1TS U3996 ( .A0(n3155), .A1(n3232), .B0(\dataoutbuffer[3][10] ), .B1(
        n4701), .Y(n3255) );
  OAI22X1TS U3997 ( .A0(n3579), .A1(n4022), .B0(n3567), .B1(n5086), .Y(n3253)
         );
  AOI21X1TS U3998 ( .A0(n4687), .A1(n3156), .B0(n3253), .Y(n3254) );
  AOI22X1TS U3999 ( .A0(n3207), .A1(n3232), .B0(\dataoutbuffer[3][17] ), .B1(
        n4701), .Y(n3258) );
  OAI22X1TS U4000 ( .A0(n3579), .A1(n5156), .B0(n3567), .B1(n4207), .Y(n3256)
         );
  AOI21X1TS U4001 ( .A0(n4696), .A1(n3208), .B0(n3256), .Y(n3257) );
  CLKBUFX2TS U4002 ( .A(dataIn_EAST[19]), .Y(n3259) );
  INVX2TS U4003 ( .A(n3259), .Y(n5177) );
  CLKBUFX2TS U4004 ( .A(cacheDataOut[19]), .Y(n3260) );
  AOI22X1TS U4005 ( .A0(n3260), .A1(n3232), .B0(\dataoutbuffer[3][19] ), .B1(
        n4701), .Y(n3267) );
  CLKBUFX2TS U4006 ( .A(dataIn_WEST[19]), .Y(n3261) );
  CLKBUFX2TS U4007 ( .A(dataIn_NORTH[19]), .Y(n3263) );
  INVX2TS U4008 ( .A(n3263), .Y(n4014) );
  CLKBUFX2TS U4009 ( .A(dataIn_SOUTH[19]), .Y(n3264) );
  INVX2TS U4010 ( .A(n3264), .Y(n5176) );
  OAI22X1TS U4011 ( .A0(n3579), .A1(n4014), .B0(n3567), .B1(n5176), .Y(n3265)
         );
  AOI21X1TS U4012 ( .A0(n4687), .A1(n3261), .B0(n3265), .Y(n3266) );
  CLKBUFX2TS U4013 ( .A(dataIn_WEST[6]), .Y(n3268) );
  INVX2TS U4014 ( .A(n3268), .Y(n4018) );
  CLKBUFX2TS U4015 ( .A(cacheDataOut[6]), .Y(n3269) );
  AOI22X1TS U4016 ( .A0(n3269), .A1(n3232), .B0(\dataoutbuffer[3][6] ), .B1(
        n4701), .Y(n3276) );
  CLKBUFX2TS U4017 ( .A(dataIn_EAST[6]), .Y(n3270) );
  CLKBUFX2TS U4018 ( .A(dataIn_NORTH[6]), .Y(n3272) );
  CLKBUFX2TS U4019 ( .A(dataIn_SOUTH[6]), .Y(n3273) );
  INVX2TS U4020 ( .A(n3273), .Y(n5043) );
  OAI22X1TS U4021 ( .A0(n3579), .A1(n5044), .B0(n3567), .B1(n5043), .Y(n3274)
         );
  AOI21X1TS U4022 ( .A0(n4696), .A1(n3270), .B0(n3274), .Y(n3275) );
  CLKBUFX2TS U4023 ( .A(dataIn_EAST[12]), .Y(n3277) );
  INVX2TS U4024 ( .A(n3277), .Y(n4162) );
  CLKBUFX2TS U4025 ( .A(cacheDataOut[12]), .Y(n3278) );
  AOI22X1TS U4026 ( .A0(n3278), .A1(n3232), .B0(\dataoutbuffer[3][12] ), .B1(
        n4701), .Y(n3285) );
  CLKBUFX2TS U4027 ( .A(dataIn_WEST[12]), .Y(n3279) );
  CLKBUFX2TS U4028 ( .A(dataIn_NORTH[12]), .Y(n3281) );
  INVX2TS U4029 ( .A(n3281), .Y(n4044) );
  CLKBUFX2TS U4030 ( .A(dataIn_SOUTH[12]), .Y(n3282) );
  INVX2TS U4031 ( .A(n3282), .Y(n4161) );
  OAI22X1TS U4032 ( .A0(n3579), .A1(n4044), .B0(n3567), .B1(n4161), .Y(n3283)
         );
  AOI21X1TS U4033 ( .A0(n4687), .A1(n3279), .B0(n3283), .Y(n3284) );
  CLKBUFX2TS U4034 ( .A(dataIn_EAST[21]), .Y(n3286) );
  INVX2TS U4035 ( .A(n3286), .Y(n4043) );
  CLKBUFX2TS U4036 ( .A(cacheDataOut[21]), .Y(n3287) );
  AOI22X1TS U4037 ( .A0(n3287), .A1(n3232), .B0(\dataoutbuffer[3][21] ), .B1(
        n4701), .Y(n3295) );
  CLKBUFX2TS U4038 ( .A(dataIn_WEST[21]), .Y(n3288) );
  CLKBUFX2TS U4039 ( .A(dataIn_NORTH[21]), .Y(n3290) );
  INVX2TS U4040 ( .A(n3290), .Y(n4039) );
  CLKBUFX2TS U4041 ( .A(dataIn_SOUTH[21]), .Y(n3291) );
  OAI22X1TS U4042 ( .A0(n3579), .A1(n4039), .B0(n3567), .B1(n3292), .Y(n3293)
         );
  AOI21X1TS U4043 ( .A0(n4687), .A1(n3288), .B0(n3293), .Y(n3294) );
  CLKBUFX2TS U4044 ( .A(dataIn_EAST[27]), .Y(n3296) );
  INVX2TS U4045 ( .A(n3296), .Y(n5259) );
  CLKBUFX2TS U4046 ( .A(cacheDataOut[27]), .Y(n3297) );
  AOI22X1TS U4047 ( .A0(n3297), .A1(n3232), .B0(\dataoutbuffer[3][27] ), .B1(
        n4701), .Y(n3304) );
  CLKBUFX2TS U4048 ( .A(dataIn_WEST[27]), .Y(n3298) );
  CLKBUFX2TS U4049 ( .A(dataIn_NORTH[27]), .Y(n3300) );
  INVX2TS U4050 ( .A(n3300), .Y(n4004) );
  CLKBUFX2TS U4051 ( .A(dataIn_SOUTH[27]), .Y(n3301) );
  INVX2TS U4052 ( .A(n3301), .Y(n5260) );
  OAI22X1TS U4053 ( .A0(n3579), .A1(n4004), .B0(n3567), .B1(n5260), .Y(n3302)
         );
  AOI21X1TS U4054 ( .A0(n4687), .A1(n3298), .B0(n3302), .Y(n3303) );
  AOI22X1TS U4055 ( .A0(n3005), .A1(n4616), .B0(
        \destinationAddressbuffer[6][6] ), .B1(n4612), .Y(n3306) );
  AOI22X1TS U4056 ( .A0(n4615), .A1(n3001), .B0(n4614), .B1(n3004), .Y(n3305)
         );
  AOI22X1TS U4057 ( .A0(n2980), .A1(n4607), .B0(writeOutbuffer[6]), .B1(n4612), 
        .Y(n3308) );
  AOI22X1TS U4058 ( .A0(n4616), .A1(n2983), .B0(n4614), .B1(n2982), .Y(n3307)
         );
  AOI22X1TS U4059 ( .A0(n2990), .A1(n4616), .B0(
        \destinationAddressbuffer[6][8] ), .B1(n4612), .Y(n3310) );
  AOI22X1TS U4060 ( .A0(n4607), .A1(n2988), .B0(n4614), .B1(n2989), .Y(n3309)
         );
  AOI22X1TS U4061 ( .A0(n3117), .A1(n4607), .B0(
        \destinationAddressbuffer[6][13] ), .B1(n4612), .Y(n3312) );
  AOI22X1TS U4062 ( .A0(n4616), .A1(n3115), .B0(n4613), .B1(n3116), .Y(n3311)
         );
  AOI22X1TS U4063 ( .A0(n3122), .A1(n4613), .B0(
        \destinationAddressbuffer[6][9] ), .B1(n4612), .Y(n3314) );
  AOI22X1TS U4064 ( .A0(n4615), .A1(n3121), .B0(n4616), .B1(n3123), .Y(n3313)
         );
  OAI32X1TS U4065 ( .A0(n3615), .A1(n3613), .A2(n3876), .B0(n4471), .B1(n3615), 
        .Y(n4473) );
  NAND2X1TS U4066 ( .A(n3319), .B(n4467), .Y(n4466) );
  NOR2X2TS U4067 ( .A(n4469), .B(n4466), .Y(n4583) );
  INVX2TS U4068 ( .A(n4473), .Y(n4579) );
  AOI22X1TS U4069 ( .A0(n3002), .A1(n4583), .B0(
        \destinationAddressbuffer[7][6] ), .B1(n4579), .Y(n3322) );
  NOR2X2TS U4070 ( .A(n4467), .B(n4469), .Y(n4580) );
  AOI22X1TS U4071 ( .A0(n3004), .A1(n4584), .B0(n3005), .B1(n4580), .Y(n3321)
         );
  AOI22X1TS U4072 ( .A0(n2976), .A1(n4580), .B0(
        \destinationAddressbuffer[7][7] ), .B1(n4579), .Y(n3324) );
  AOI22X1TS U4073 ( .A0(n2975), .A1(n4584), .B0(n2972), .B1(n4583), .Y(n3323)
         );
  INVX2TS U4074 ( .A(n4583), .Y(n3964) );
  NOR3XLTS U4075 ( .A(n3876), .B(n3615), .C(n3614), .Y(n3325) );
  BUFX3TS U4076 ( .A(n3325), .Y(n4323) );
  AOI22X1TS U4077 ( .A0(n3155), .A1(n4323), .B0(\dataoutbuffer[7][10] ), .B1(
        n4579), .Y(n3328) );
  INVX2TS U4078 ( .A(n4580), .Y(n3975) );
  OAI22X1TS U4079 ( .A0(n3157), .A1(n3975), .B0(n5086), .B1(n3969), .Y(n3326)
         );
  AOI21X1TS U4080 ( .A0(n3154), .A1(n4584), .B0(n3326), .Y(n3327) );
  AOI22X1TS U4081 ( .A0(n2964), .A1(n4323), .B0(\dataoutbuffer[7][13] ), .B1(
        n4579), .Y(n3331) );
  OAI22X1TS U4082 ( .A0(n2963), .A1(n3969), .B0(n4117), .B1(n3964), .Y(n3329)
         );
  AOI21X1TS U4083 ( .A0(n2965), .A1(n4584), .B0(n3329), .Y(n3330) );
  AOI22X1TS U4084 ( .A0(n3207), .A1(n4323), .B0(\dataoutbuffer[7][17] ), .B1(
        n4579), .Y(n3334) );
  OAI22X1TS U4085 ( .A0(n3209), .A1(n3964), .B0(n4207), .B1(n3969), .Y(n3332)
         );
  AOI21X1TS U4086 ( .A0(n3206), .A1(n4584), .B0(n3332), .Y(n3333) );
  AOI22X1TS U4087 ( .A0(n3061), .A1(n4323), .B0(\dataoutbuffer[7][9] ), .B1(
        n4579), .Y(n3337) );
  OAI22X1TS U4088 ( .A0(n5075), .A1(n3969), .B0(n5074), .B1(n3964), .Y(n3335)
         );
  AOI21X1TS U4089 ( .A0(n3062), .A1(n4584), .B0(n3335), .Y(n3336) );
  AOI22X1TS U4090 ( .A0(n3052), .A1(n4323), .B0(\dataoutbuffer[7][8] ), .B1(
        n4579), .Y(n3340) );
  OAI22X1TS U4091 ( .A0(n3056), .A1(n3969), .B0(n4166), .B1(n3964), .Y(n3338)
         );
  AOI21X1TS U4092 ( .A0(n3053), .A1(n4584), .B0(n3338), .Y(n3339) );
  CLKBUFX2TS U4093 ( .A(dataIn_EAST[15]), .Y(n3341) );
  INVX2TS U4094 ( .A(n3341), .Y(n5135) );
  CLKBUFX2TS U4095 ( .A(cacheDataOut[15]), .Y(n3342) );
  AOI22X1TS U4096 ( .A0(n3342), .A1(n4323), .B0(\dataoutbuffer[7][15] ), .B1(
        n4579), .Y(n3349) );
  CLKBUFX2TS U4097 ( .A(dataIn_SOUTH[15]), .Y(n3343) );
  CLKBUFX2TS U4098 ( .A(dataIn_WEST[15]), .Y(n3344) );
  INVX2TS U4099 ( .A(n3344), .Y(n4211) );
  CLKBUFX2TS U4100 ( .A(dataIn_NORTH[15]), .Y(n3345) );
  OAI22X1TS U4101 ( .A0(n4211), .A1(n3975), .B0(n3346), .B1(n3968), .Y(n3347)
         );
  AOI21X1TS U4102 ( .A0(n3343), .A1(n4586), .B0(n3347), .Y(n3348) );
  AOI22X1TS U4103 ( .A0(n3278), .A1(n4323), .B0(\dataoutbuffer[7][12] ), .B1(
        n4579), .Y(n3352) );
  OAI22X1TS U4104 ( .A0(n3280), .A1(n3975), .B0(n4044), .B1(n3968), .Y(n3350)
         );
  AOI21X1TS U4105 ( .A0(n3282), .A1(n4586), .B0(n3350), .Y(n3351) );
  CLKBUFX2TS U4106 ( .A(dataIn_EAST[14]), .Y(n3353) );
  CLKBUFX2TS U4107 ( .A(cacheDataOut[14]), .Y(n3354) );
  AOI22X1TS U4108 ( .A0(n3354), .A1(n4323), .B0(\dataoutbuffer[7][14] ), .B1(
        n4579), .Y(n3361) );
  CLKBUFX2TS U4109 ( .A(dataIn_SOUTH[14]), .Y(n3355) );
  CLKBUFX2TS U4110 ( .A(dataIn_WEST[14]), .Y(n3356) );
  CLKBUFX2TS U4111 ( .A(dataIn_NORTH[14]), .Y(n3358) );
  OAI22X1TS U4112 ( .A0(n3357), .A1(n3975), .B0(n5123), .B1(n3968), .Y(n3359)
         );
  AOI21X1TS U4113 ( .A0(n3355), .A1(n4586), .B0(n3359), .Y(n3360) );
  CLKBUFX2TS U4114 ( .A(dataIn_WEST[11]), .Y(n3362) );
  INVX2TS U4115 ( .A(n3362), .Y(n4102) );
  CLKBUFX2TS U4116 ( .A(cacheDataOut[11]), .Y(n3363) );
  AOI22X1TS U4117 ( .A0(n3363), .A1(n4323), .B0(\dataoutbuffer[7][11] ), .B1(
        n4579), .Y(n3370) );
  CLKBUFX2TS U4118 ( .A(dataIn_SOUTH[11]), .Y(n3364) );
  CLKBUFX2TS U4119 ( .A(dataIn_EAST[11]), .Y(n3366) );
  INVX2TS U4120 ( .A(n3366), .Y(n4106) );
  CLKBUFX2TS U4121 ( .A(dataIn_NORTH[11]), .Y(n3367) );
  INVX2TS U4122 ( .A(n3367), .Y(n4029) );
  OAI22X1TS U4123 ( .A0(n4106), .A1(n3964), .B0(n4029), .B1(n3968), .Y(n3368)
         );
  AOI21X1TS U4124 ( .A0(n3364), .A1(n4586), .B0(n3368), .Y(n3369) );
  AOI22X1TS U4125 ( .A0(n3043), .A1(n4323), .B0(\dataoutbuffer[7][16] ), .B1(
        n4579), .Y(n3373) );
  OAI22X1TS U4126 ( .A0(n3045), .A1(n3968), .B0(n5145), .B1(n3964), .Y(n3371)
         );
  AOI21X1TS U4127 ( .A0(n3047), .A1(n4586), .B0(n3371), .Y(n3372) );
  INVX2TS U4128 ( .A(n4615), .Y(n4064) );
  AOI22X1TS U4129 ( .A0(n2976), .A1(n4616), .B0(
        \destinationAddressbuffer[6][7] ), .B1(n4612), .Y(n3375) );
  AOI22X1TS U4130 ( .A0(n4613), .A1(n2972), .B0(n4614), .B1(n2975), .Y(n3374)
         );
  AOI22X1TS U4131 ( .A0(n3039), .A1(n4616), .B0(
        \destinationAddressbuffer[6][12] ), .B1(n4612), .Y(n3377) );
  AOI22X1TS U4132 ( .A0(n4613), .A1(n3035), .B0(n4614), .B1(n3038), .Y(n3376)
         );
  AOI22X1TS U4133 ( .A0(n3031), .A1(n4616), .B0(
        \destinationAddressbuffer[6][10] ), .B1(n4612), .Y(n3379) );
  AOI22X1TS U4134 ( .A0(n4613), .A1(n3028), .B0(n4614), .B1(n3030), .Y(n3378)
         );
  OAI32X1TS U4135 ( .A0(n3615), .A1(n3613), .A2(n3384), .B0(n4526), .B1(n3615), 
        .Y(n4528) );
  NOR2X2TS U4136 ( .A(n4522), .B(n4524), .Y(n4760) );
  INVX2TS U4137 ( .A(n4760), .Y(n4229) );
  NOR3XLTS U4138 ( .A(n3615), .B(n3614), .C(n3384), .Y(n3385) );
  BUFX3TS U4139 ( .A(n3385), .Y(n4436) );
  INVX2TS U4140 ( .A(n4528), .Y(n4744) );
  AOI22X1TS U4141 ( .A0(n3354), .A1(n4436), .B0(\dataoutbuffer[1][14] ), .B1(
        n4744), .Y(n3389) );
  NOR2X2TS U4142 ( .A(n4524), .B(n4521), .Y(n4758) );
  INVX2TS U4143 ( .A(n4758), .Y(n4240) );
  OAI22X1TS U4144 ( .A0(n5124), .A1(n4240), .B0(n5123), .B1(n3875), .Y(n3387)
         );
  AOI21X1TS U4145 ( .A0(n3355), .A1(n4759), .B0(n3387), .Y(n3388) );
  AOI22X1TS U4146 ( .A0(n3363), .A1(n4436), .B0(\dataoutbuffer[1][11] ), .B1(
        n4744), .Y(n3392) );
  OAI22X1TS U4147 ( .A0(n4106), .A1(n4240), .B0(n4029), .B1(n3875), .Y(n3390)
         );
  AOI21X1TS U4148 ( .A0(n3364), .A1(n4759), .B0(n3390), .Y(n3391) );
  AOI22X1TS U4149 ( .A0(n3137), .A1(n4436), .B0(\dataoutbuffer[1][31] ), .B1(
        n4744), .Y(n3395) );
  OAI22X1TS U4150 ( .A0(n3140), .A1(n4229), .B0(n5306), .B1(n3875), .Y(n3393)
         );
  AOI21X1TS U4151 ( .A0(n3138), .A1(n4759), .B0(n3393), .Y(n3394) );
  CLKBUFX2TS U4152 ( .A(dataIn_WEST[28]), .Y(n3396) );
  INVX2TS U4153 ( .A(n3396), .Y(n3951) );
  CLKBUFX2TS U4154 ( .A(cacheDataOut[28]), .Y(n3397) );
  AOI22X1TS U4155 ( .A0(n3397), .A1(n3232), .B0(\dataoutbuffer[3][28] ), .B1(
        n4701), .Y(n3404) );
  CLKBUFX2TS U4156 ( .A(dataIn_NORTH[28]), .Y(n3398) );
  CLKBUFX2TS U4157 ( .A(dataIn_EAST[28]), .Y(n3399) );
  INVX2TS U4158 ( .A(n3399), .Y(n5270) );
  CLKBUFX2TS U4159 ( .A(dataIn_SOUTH[28]), .Y(n3400) );
  OAI22X1TS U4160 ( .A0(n3575), .A1(n5270), .B0(n3567), .B1(n3401), .Y(n3402)
         );
  AOI21X1TS U4161 ( .A0(n4703), .A1(n3398), .B0(n3402), .Y(n3403) );
  CLKBUFX2TS U4162 ( .A(dataIn_WEST[18]), .Y(n3405) );
  CLKBUFX2TS U4163 ( .A(cacheDataOut[18]), .Y(n3407) );
  AOI22X1TS U4164 ( .A0(n3407), .A1(n3232), .B0(\dataoutbuffer[3][18] ), .B1(
        n4701), .Y(n3414) );
  CLKBUFX2TS U4165 ( .A(dataIn_NORTH[18]), .Y(n3408) );
  CLKBUFX2TS U4166 ( .A(dataIn_EAST[18]), .Y(n3410) );
  INVX2TS U4167 ( .A(n3410), .Y(n4205) );
  CLKBUFX2TS U4168 ( .A(dataIn_SOUTH[18]), .Y(n3411) );
  INVX2TS U4169 ( .A(n3411), .Y(n5166) );
  OAI22X1TS U4170 ( .A0(n3575), .A1(n4205), .B0(n3567), .B1(n5166), .Y(n3412)
         );
  AOI21X1TS U4171 ( .A0(n4703), .A1(n3408), .B0(n3412), .Y(n3413) );
  AOI22X1TS U4172 ( .A0(n3061), .A1(n3232), .B0(\dataoutbuffer[3][9] ), .B1(
        n4701), .Y(n3417) );
  OAI22X1TS U4173 ( .A0(n3575), .A1(n5074), .B0(n3567), .B1(n5075), .Y(n3415)
         );
  AOI21X1TS U4174 ( .A0(n4703), .A1(n3062), .B0(n3415), .Y(n3416) );
  AOI22X1TS U4175 ( .A0(n3342), .A1(n3232), .B0(\dataoutbuffer[3][15] ), .B1(
        n4701), .Y(n3420) );
  OAI22X1TS U4176 ( .A0(n3579), .A1(n3346), .B0(n3575), .B1(n5135), .Y(n3418)
         );
  AOI21X1TS U4177 ( .A0(n4702), .A1(n3343), .B0(n3418), .Y(n3419) );
  AOI22X1TS U4178 ( .A0(n3019), .A1(n3232), .B0(\dataoutbuffer[3][0] ), .B1(
        n4701), .Y(n3423) );
  INVX2TS U4179 ( .A(n3020), .Y(n4980) );
  OAI22X1TS U4180 ( .A0(n3579), .A1(n4980), .B0(n3575), .B1(n3023), .Y(n3421)
         );
  AOI21X1TS U4181 ( .A0(n4702), .A1(n3017), .B0(n3421), .Y(n3422) );
  AOI22X1TS U4182 ( .A0(n3010), .A1(n3232), .B0(\dataoutbuffer[3][1] ), .B1(
        n4701), .Y(n3426) );
  INVX2TS U4183 ( .A(n3011), .Y(n4991) );
  OAI22X1TS U4184 ( .A0(n3579), .A1(n4991), .B0(n3575), .B1(n4990), .Y(n3424)
         );
  AOI21X1TS U4185 ( .A0(n4702), .A1(n3008), .B0(n3424), .Y(n3425) );
  CLKBUFX2TS U4186 ( .A(dataIn_WEST[26]), .Y(n3427) );
  INVX2TS U4187 ( .A(n3427), .Y(n4089) );
  CLKBUFX2TS U4188 ( .A(cacheDataOut[26]), .Y(n3428) );
  AOI22X1TS U4189 ( .A0(n3428), .A1(n3232), .B0(\dataoutbuffer[3][26] ), .B1(
        n4701), .Y(n3435) );
  CLKBUFX2TS U4190 ( .A(dataIn_SOUTH[26]), .Y(n3429) );
  CLKBUFX2TS U4191 ( .A(dataIn_NORTH[26]), .Y(n3431) );
  INVX2TS U4192 ( .A(n3431), .Y(n4060) );
  CLKBUFX2TS U4193 ( .A(dataIn_EAST[26]), .Y(n3432) );
  INVX2TS U4194 ( .A(n3432), .Y(n4085) );
  OAI22X1TS U4195 ( .A0(n3579), .A1(n4060), .B0(n3575), .B1(n4085), .Y(n3433)
         );
  AOI21X1TS U4196 ( .A0(n4702), .A1(n3429), .B0(n3433), .Y(n3434) );
  AOI22X1TS U4197 ( .A0(n3164), .A1(n3232), .B0(\dataoutbuffer[3][4] ), .B1(
        n4701), .Y(n3438) );
  OAI22X1TS U4198 ( .A0(n3579), .A1(n5022), .B0(n3575), .B1(n5023), .Y(n3436)
         );
  AOI21X1TS U4199 ( .A0(n4702), .A1(n3165), .B0(n3436), .Y(n3437) );
  AOI22X1TS U4200 ( .A0(n3354), .A1(n3232), .B0(\dataoutbuffer[3][14] ), .B1(
        n4701), .Y(n3441) );
  OAI22X1TS U4201 ( .A0(n3579), .A1(n5123), .B0(n3575), .B1(n5124), .Y(n3439)
         );
  AOI21X1TS U4202 ( .A0(n4702), .A1(n3355), .B0(n3439), .Y(n3440) );
  CLKBUFX2TS U4203 ( .A(dataIn_WEST[3]), .Y(n3442) );
  INVX2TS U4204 ( .A(n3442), .Y(n3985) );
  CLKBUFX2TS U4205 ( .A(cacheDataOut[3]), .Y(n3443) );
  AOI22X1TS U4206 ( .A0(n3443), .A1(n3232), .B0(\dataoutbuffer[3][3] ), .B1(
        n4701), .Y(n3449) );
  CLKBUFX2TS U4207 ( .A(dataIn_SOUTH[3]), .Y(n3444) );
  CLKBUFX2TS U4208 ( .A(dataIn_NORTH[3]), .Y(n3445) );
  CLKBUFX2TS U4209 ( .A(dataIn_EAST[3]), .Y(n3446) );
  OAI22X1TS U4210 ( .A0(n3579), .A1(n5012), .B0(n3575), .B1(n5011), .Y(n3447)
         );
  AOI21X1TS U4211 ( .A0(n4702), .A1(n3444), .B0(n3447), .Y(n3448) );
  AOI22X1TS U4212 ( .A0(n3128), .A1(n3232), .B0(\dataoutbuffer[3][29] ), .B1(
        n4701), .Y(n3452) );
  OAI22X1TS U4213 ( .A0(n3579), .A1(n3127), .B0(n3575), .B1(n4171), .Y(n3450)
         );
  AOI21X1TS U4214 ( .A0(n4702), .A1(n3129), .B0(n3450), .Y(n3451) );
  AOI22X1TS U4215 ( .A0(n3198), .A1(n4417), .B0(\dataoutbuffer[2][7] ), .B1(
        n4728), .Y(n3455) );
  OAI22X1TS U4216 ( .A0(n3538), .A1(n5054), .B0(n3533), .B1(n3201), .Y(n3453)
         );
  AOI21X1TS U4217 ( .A0(n4729), .A1(n3199), .B0(n3453), .Y(n3454) );
  CLKBUFX2TS U4218 ( .A(dataIn_SOUTH[30]), .Y(n3456) );
  INVX2TS U4219 ( .A(n3456), .Y(n5292) );
  CLKBUFX2TS U4220 ( .A(cacheDataOut[30]), .Y(n3457) );
  AOI22X1TS U4221 ( .A0(n3457), .A1(n4417), .B0(\dataoutbuffer[2][30] ), .B1(
        n4728), .Y(n3464) );
  CLKBUFX2TS U4222 ( .A(dataIn_EAST[30]), .Y(n3458) );
  CLKBUFX2TS U4223 ( .A(dataIn_NORTH[30]), .Y(n3459) );
  CLKBUFX2TS U4224 ( .A(dataIn_WEST[30]), .Y(n3461) );
  INVX2TS U4225 ( .A(n3461), .Y(n4198) );
  OAI22X1TS U4226 ( .A0(n3538), .A1(n3460), .B0(n3533), .B1(n4198), .Y(n3462)
         );
  AOI21X1TS U4227 ( .A0(n4729), .A1(n3458), .B0(n3462), .Y(n3463) );
  AOI22X1TS U4228 ( .A0(n3207), .A1(n4417), .B0(\dataoutbuffer[2][17] ), .B1(
        n4728), .Y(n3467) );
  OAI22X1TS U4229 ( .A0(n3538), .A1(n5156), .B0(n3533), .B1(n4206), .Y(n3465)
         );
  AOI21X1TS U4230 ( .A0(n4729), .A1(n3208), .B0(n3465), .Y(n3466) );
  AOI22X1TS U4231 ( .A0(n3260), .A1(n4417), .B0(\dataoutbuffer[2][19] ), .B1(
        n4728), .Y(n3470) );
  OAI22X1TS U4232 ( .A0(n3538), .A1(n4014), .B0(n3542), .B1(n5177), .Y(n3468)
         );
  AOI21X1TS U4233 ( .A0(n4731), .A1(n3261), .B0(n3468), .Y(n3469) );
  AOI22X1TS U4234 ( .A0(n3244), .A1(n4417), .B0(\dataoutbuffer[2][20] ), .B1(
        n4728), .Y(n3473) );
  OAI22X1TS U4235 ( .A0(n3538), .A1(n3248), .B0(n3542), .B1(n5188), .Y(n3471)
         );
  AOI21X1TS U4236 ( .A0(n4731), .A1(n3245), .B0(n3471), .Y(n3472) );
  AOI22X1TS U4237 ( .A0(n3407), .A1(n4417), .B0(\dataoutbuffer[2][18] ), .B1(
        n4728), .Y(n3476) );
  OAI22X1TS U4238 ( .A0(n3538), .A1(n3409), .B0(n3542), .B1(n4205), .Y(n3474)
         );
  AOI21X1TS U4239 ( .A0(n4731), .A1(n3405), .B0(n3474), .Y(n3475) );
  AOI22X1TS U4240 ( .A0(n3363), .A1(n4417), .B0(\dataoutbuffer[2][11] ), .B1(
        n4728), .Y(n3479) );
  OAI22X1TS U4241 ( .A0(n3538), .A1(n4029), .B0(n3537), .B1(n3365), .Y(n3477)
         );
  AOI21X1TS U4242 ( .A0(n4729), .A1(n3366), .B0(n3477), .Y(n3478) );
  CLKBUFX2TS U4243 ( .A(dataIn_WEST[22]), .Y(n3480) );
  INVX2TS U4244 ( .A(n3480), .Y(n4223) );
  CLKBUFX2TS U4245 ( .A(cacheDataOut[22]), .Y(n3481) );
  AOI22X1TS U4246 ( .A0(n3481), .A1(n4417), .B0(\dataoutbuffer[2][22] ), .B1(
        n4728), .Y(n3488) );
  CLKBUFX2TS U4247 ( .A(dataIn_SOUTH[22]), .Y(n3482) );
  CLKBUFX2TS U4248 ( .A(dataIn_NORTH[22]), .Y(n3483) );
  CLKBUFX2TS U4249 ( .A(dataIn_EAST[22]), .Y(n3485) );
  INVX2TS U4250 ( .A(n3485), .Y(n4227) );
  OAI22X1TS U4251 ( .A0(n3538), .A1(n3484), .B0(n3542), .B1(n4227), .Y(n3486)
         );
  AOI21X1TS U4252 ( .A0(n4730), .A1(n3482), .B0(n3486), .Y(n3487) );
  CLKBUFX2TS U4253 ( .A(dataIn_WEST[2]), .Y(n3489) );
  INVX2TS U4254 ( .A(n3489), .Y(n4132) );
  CLKBUFX2TS U4255 ( .A(cacheDataOut[2]), .Y(n3490) );
  AOI22X1TS U4256 ( .A0(n3490), .A1(n4417), .B0(\dataoutbuffer[2][2] ), .B1(
        n4728), .Y(n3498) );
  CLKBUFX2TS U4257 ( .A(dataIn_SOUTH[2]), .Y(n3491) );
  CLKBUFX2TS U4258 ( .A(dataIn_NORTH[2]), .Y(n3493) );
  CLKBUFX2TS U4259 ( .A(dataIn_EAST[2]), .Y(n3495) );
  OAI22X1TS U4260 ( .A0(n3538), .A1(n3494), .B0(n3542), .B1(n5001), .Y(n3496)
         );
  AOI21X1TS U4261 ( .A0(n4730), .A1(n3491), .B0(n3496), .Y(n3497) );
  INVX2TS U4262 ( .A(n3343), .Y(n5134) );
  AOI22X1TS U4263 ( .A0(n3342), .A1(n4417), .B0(\dataoutbuffer[2][15] ), .B1(
        n4728), .Y(n3501) );
  OAI22X1TS U4264 ( .A0(n3538), .A1(n3346), .B0(n3542), .B1(n5135), .Y(n3499)
         );
  AOI21X1TS U4265 ( .A0(n4731), .A1(n3344), .B0(n3499), .Y(n3500) );
  AOI22X1TS U4266 ( .A0(n3428), .A1(n4417), .B0(\dataoutbuffer[2][26] ), .B1(
        n4728), .Y(n3504) );
  OAI22X1TS U4267 ( .A0(n3538), .A1(n4060), .B0(n3542), .B1(n4085), .Y(n3502)
         );
  AOI21X1TS U4268 ( .A0(n4730), .A1(n3429), .B0(n3502), .Y(n3503) );
  AOI22X1TS U4269 ( .A0(n3269), .A1(n4417), .B0(\dataoutbuffer[2][6] ), .B1(
        n4728), .Y(n3507) );
  OAI22X1TS U4270 ( .A0(n3538), .A1(n5044), .B0(n3533), .B1(n4018), .Y(n3505)
         );
  AOI21X1TS U4271 ( .A0(n4729), .A1(n3270), .B0(n3505), .Y(n3506) );
  AOI22X1TS U4272 ( .A0(n3278), .A1(n4417), .B0(\dataoutbuffer[2][12] ), .B1(
        n4728), .Y(n3510) );
  OAI22X1TS U4273 ( .A0(n3538), .A1(n4044), .B0(n3537), .B1(n4161), .Y(n3508)
         );
  AOI21X1TS U4274 ( .A0(n4731), .A1(n3279), .B0(n3508), .Y(n3509) );
  AOI22X1TS U4275 ( .A0(n3443), .A1(n4417), .B0(\dataoutbuffer[2][3] ), .B1(
        n4728), .Y(n3513) );
  OAI22X1TS U4276 ( .A0(n3538), .A1(n5012), .B0(n3533), .B1(n3985), .Y(n3511)
         );
  AOI21X1TS U4277 ( .A0(n4730), .A1(n3444), .B0(n3511), .Y(n3512) );
  AOI22X1TS U4278 ( .A0(n3287), .A1(n4417), .B0(\dataoutbuffer[2][21] ), .B1(
        n4728), .Y(n3516) );
  OAI22X1TS U4279 ( .A0(n3538), .A1(n4039), .B0(n3537), .B1(n3292), .Y(n3514)
         );
  AOI21X1TS U4280 ( .A0(n4731), .A1(n3288), .B0(n3514), .Y(n3515) );
  AOI22X1TS U4281 ( .A0(n3297), .A1(n4417), .B0(\dataoutbuffer[2][27] ), .B1(
        n4728), .Y(n3519) );
  OAI22X1TS U4282 ( .A0(n3538), .A1(n4004), .B0(n3537), .B1(n5260), .Y(n3517)
         );
  AOI21X1TS U4283 ( .A0(n4731), .A1(n3298), .B0(n3517), .Y(n3518) );
  AOI22X1TS U4284 ( .A0(n3397), .A1(n4417), .B0(\dataoutbuffer[2][28] ), .B1(
        n4728), .Y(n3522) );
  INVX2TS U4285 ( .A(n3398), .Y(n3947) );
  OAI22X1TS U4286 ( .A0(n3538), .A1(n3947), .B0(n3537), .B1(n3401), .Y(n3520)
         );
  AOI21X1TS U4287 ( .A0(n4731), .A1(n3396), .B0(n3520), .Y(n3521) );
  AOI22X1TS U4288 ( .A0(n3354), .A1(n4417), .B0(\dataoutbuffer[2][14] ), .B1(
        n4728), .Y(n3525) );
  OAI22X1TS U4289 ( .A0(n3538), .A1(n5123), .B0(n3533), .B1(n3357), .Y(n3523)
         );
  AOI21X1TS U4290 ( .A0(n4730), .A1(n3355), .B0(n3523), .Y(n3524) );
  CLKBUFX2TS U4291 ( .A(dataIn_EAST[5]), .Y(n3526) );
  CLKBUFX2TS U4292 ( .A(cacheDataOut[5]), .Y(n3527) );
  AOI22X1TS U4293 ( .A0(n3527), .A1(n4417), .B0(\dataoutbuffer[2][5] ), .B1(
        n4728), .Y(n3536) );
  CLKBUFX2TS U4294 ( .A(dataIn_SOUTH[5]), .Y(n3528) );
  CLKBUFX2TS U4295 ( .A(dataIn_NORTH[5]), .Y(n3530) );
  CLKBUFX2TS U4296 ( .A(dataIn_WEST[5]), .Y(n3532) );
  INVX2TS U4297 ( .A(n3532), .Y(n4141) );
  OAI22X1TS U4298 ( .A0(n3538), .A1(n3531), .B0(n3533), .B1(n4141), .Y(n3534)
         );
  AOI21X1TS U4299 ( .A0(n4730), .A1(n3528), .B0(n3534), .Y(n3535) );
  INVX2TS U4300 ( .A(n3233), .Y(n5239) );
  AOI22X1TS U4301 ( .A0(n3230), .A1(n4417), .B0(\dataoutbuffer[2][25] ), .B1(
        n4728), .Y(n3541) );
  OAI22X1TS U4302 ( .A0(n3538), .A1(n5238), .B0(n3537), .B1(n3236), .Y(n3539)
         );
  AOI21X1TS U4303 ( .A0(n4731), .A1(n3229), .B0(n3539), .Y(n3540) );
  AOI22X1TS U4304 ( .A0(n3198), .A1(n3232), .B0(\dataoutbuffer[3][7] ), .B1(
        n4701), .Y(n3545) );
  OAI22X1TS U4305 ( .A0(n3567), .A1(n5055), .B0(n3574), .B1(n3201), .Y(n3543)
         );
  AOI21X1TS U4306 ( .A0(n4696), .A1(n3199), .B0(n3543), .Y(n3544) );
  AOI22X1TS U4307 ( .A0(n3043), .A1(n3232), .B0(\dataoutbuffer[3][16] ), .B1(
        n4701), .Y(n3548) );
  OAI22X1TS U4308 ( .A0(n3567), .A1(n5146), .B0(n3574), .B1(n4219), .Y(n3546)
         );
  AOI21X1TS U4309 ( .A0(n4703), .A1(n3044), .B0(n3546), .Y(n3547) );
  AOI22X1TS U4310 ( .A0(n3052), .A1(n3232), .B0(\dataoutbuffer[3][8] ), .B1(
        n4701), .Y(n3551) );
  OAI22X1TS U4311 ( .A0(n3567), .A1(n3056), .B0(n3574), .B1(n4170), .Y(n3549)
         );
  AOI21X1TS U4312 ( .A0(n4703), .A1(n3053), .B0(n3549), .Y(n3550) );
  AOI22X1TS U4313 ( .A0(n3363), .A1(n3232), .B0(\dataoutbuffer[3][11] ), .B1(
        n4701), .Y(n3554) );
  OAI22X1TS U4314 ( .A0(n3579), .A1(n4029), .B0(n3574), .B1(n4102), .Y(n3552)
         );
  AOI21X1TS U4315 ( .A0(n4696), .A1(n3366), .B0(n3552), .Y(n3553) );
  INVX2TS U4316 ( .A(n3458), .Y(n5293) );
  AOI22X1TS U4317 ( .A0(n3457), .A1(n3232), .B0(\dataoutbuffer[3][30] ), .B1(
        n4701), .Y(n3557) );
  OAI22X1TS U4318 ( .A0(n3579), .A1(n3460), .B0(n3574), .B1(n4198), .Y(n3555)
         );
  AOI21X1TS U4319 ( .A0(n4702), .A1(n3456), .B0(n3555), .Y(n3556) );
  AOI22X1TS U4320 ( .A0(n3527), .A1(n3232), .B0(\dataoutbuffer[3][5] ), .B1(
        n4701), .Y(n3560) );
  OAI22X1TS U4321 ( .A0(n3579), .A1(n3531), .B0(n3574), .B1(n4141), .Y(n3558)
         );
  AOI21X1TS U4322 ( .A0(n4702), .A1(n3528), .B0(n3558), .Y(n3559) );
  AOI22X1TS U4323 ( .A0(n2964), .A1(n3232), .B0(\dataoutbuffer[3][13] ), .B1(
        n4701), .Y(n3563) );
  OAI22X1TS U4324 ( .A0(n3579), .A1(n2966), .B0(n3574), .B1(n4113), .Y(n3561)
         );
  AOI21X1TS U4325 ( .A0(n4702), .A1(n2962), .B0(n3561), .Y(n3562) );
  INVX2TS U4326 ( .A(n3482), .Y(n5207) );
  AOI22X1TS U4327 ( .A0(n3481), .A1(n3232), .B0(\dataoutbuffer[3][22] ), .B1(
        n4701), .Y(n3566) );
  OAI22X1TS U4328 ( .A0(n3575), .A1(n4227), .B0(n3574), .B1(n4223), .Y(n3564)
         );
  AOI21X1TS U4329 ( .A0(n4703), .A1(n3483), .B0(n3564), .Y(n3565) );
  AOI22X1TS U4330 ( .A0(n3490), .A1(n3232), .B0(\dataoutbuffer[3][2] ), .B1(
        n4701), .Y(n3570) );
  OAI22X1TS U4331 ( .A0(n3575), .A1(n5001), .B0(n3574), .B1(n4132), .Y(n3568)
         );
  AOI21X1TS U4332 ( .A0(n4702), .A1(n3491), .B0(n3568), .Y(n3569) );
  AOI22X1TS U4333 ( .A0(n3137), .A1(n3232), .B0(\dataoutbuffer[3][31] ), .B1(
        n4701), .Y(n3573) );
  OAI22X1TS U4334 ( .A0(n3575), .A1(n5308), .B0(n3574), .B1(n3140), .Y(n3571)
         );
  AOI21X1TS U4335 ( .A0(n4702), .A1(n3138), .B0(n3571), .Y(n3572) );
  AOI22X1TS U4336 ( .A0(n2950), .A1(n3232), .B0(\dataoutbuffer[3][23] ), .B1(
        n4701), .Y(n3578) );
  OAI22X1TS U4337 ( .A0(n3575), .A1(n5217), .B0(n3574), .B1(n4215), .Y(n3576)
         );
  AOI21X1TS U4338 ( .A0(n4702), .A1(n2957), .B0(n3576), .Y(n3577) );
  AOI22X1TS U4339 ( .A0(n3061), .A1(n4455), .B0(\dataoutbuffer[0][9] ), .B1(
        n4787), .Y(n3582) );
  OAI22X1TS U4340 ( .A0(n3704), .A1(n5074), .B0(n3698), .B1(n5075), .Y(n3580)
         );
  AOI21X1TS U4341 ( .A0(n4790), .A1(n3062), .B0(n3580), .Y(n3581) );
  AOI22X1TS U4342 ( .A0(n3155), .A1(n4455), .B0(\dataoutbuffer[0][10] ), .B1(
        n4787), .Y(n3585) );
  OAI22X1TS U4343 ( .A0(n3704), .A1(n5085), .B0(n3698), .B1(n5086), .Y(n3583)
         );
  AOI21X1TS U4344 ( .A0(n4788), .A1(n3156), .B0(n3583), .Y(n3584) );
  AOI22X1TS U4345 ( .A0(n3278), .A1(n4455), .B0(\dataoutbuffer[0][12] ), .B1(
        n4787), .Y(n3588) );
  OAI22X1TS U4346 ( .A0(n3704), .A1(n4162), .B0(n3698), .B1(n4161), .Y(n3586)
         );
  AOI21X1TS U4347 ( .A0(n4788), .A1(n3279), .B0(n3586), .Y(n3587) );
  AOI22X1TS U4348 ( .A0(n3342), .A1(n4455), .B0(\dataoutbuffer[0][15] ), .B1(
        n4787), .Y(n3591) );
  OAI22X1TS U4349 ( .A0(n3704), .A1(n5135), .B0(n3698), .B1(n5134), .Y(n3589)
         );
  AOI21X1TS U4350 ( .A0(n4788), .A1(n3344), .B0(n3589), .Y(n3590) );
  AOI22X1TS U4351 ( .A0(n3287), .A1(n4455), .B0(\dataoutbuffer[0][21] ), .B1(
        n4787), .Y(n3594) );
  OAI22X1TS U4352 ( .A0(n3704), .A1(n4043), .B0(n3698), .B1(n3292), .Y(n3592)
         );
  AOI21X1TS U4353 ( .A0(n4788), .A1(n3288), .B0(n3592), .Y(n3593) );
  AOI22X1TS U4354 ( .A0(n3363), .A1(n4455), .B0(\dataoutbuffer[0][11] ), .B1(
        n4787), .Y(n3597) );
  OAI22X1TS U4355 ( .A0(n3704), .A1(n4106), .B0(n3698), .B1(n3365), .Y(n3595)
         );
  AOI21X1TS U4356 ( .A0(n4788), .A1(n3362), .B0(n3595), .Y(n3596) );
  AOI22X1TS U4357 ( .A0(n3230), .A1(n4455), .B0(\dataoutbuffer[0][25] ), .B1(
        n4787), .Y(n3600) );
  OAI22X1TS U4358 ( .A0(n3699), .A1(n5238), .B0(n3698), .B1(n3236), .Y(n3598)
         );
  AOI21X1TS U4359 ( .A0(n4782), .A1(n3233), .B0(n3598), .Y(n3599) );
  AOI22X1TS U4360 ( .A0(n3407), .A1(n4455), .B0(\dataoutbuffer[0][18] ), .B1(
        n4787), .Y(n3603) );
  OAI22X1TS U4361 ( .A0(n3699), .A1(n3409), .B0(n3698), .B1(n5166), .Y(n3601)
         );
  AOI21X1TS U4362 ( .A0(n4788), .A1(n3405), .B0(n3601), .Y(n3602) );
  AOI22X1TS U4363 ( .A0(n3297), .A1(n4455), .B0(\dataoutbuffer[0][27] ), .B1(
        n4787), .Y(n3606) );
  OAI22X1TS U4364 ( .A0(n3699), .A1(n4004), .B0(n3698), .B1(n5260), .Y(n3604)
         );
  AOI21X1TS U4365 ( .A0(n4788), .A1(n3298), .B0(n3604), .Y(n3605) );
  OAI32X1TS U4366 ( .A0(n3615), .A1(n3613), .A2(n3708), .B0(n4489), .B1(n3615), 
        .Y(n4491) );
  NOR2X2TS U4367 ( .A(n4486), .B(n4488), .Y(n4642) );
  INVX2TS U4368 ( .A(n4642), .Y(n4140) );
  NOR3XLTS U4369 ( .A(n3615), .B(n3708), .C(n3614), .Y(n3616) );
  BUFX3TS U4370 ( .A(n3616), .Y(n4361) );
  INVX2TS U4371 ( .A(n4491), .Y(n4128) );
  AOI22X1TS U4372 ( .A0(n3407), .A1(n4361), .B0(\dataoutbuffer[5][18] ), .B1(
        n4128), .Y(n3622) );
  NOR2X2TS U4373 ( .A(n4488), .B(n4485), .Y(n4643) );
  INVX2TS U4374 ( .A(n4643), .Y(n4157) );
  OAI22X1TS U4375 ( .A0(n3409), .A1(n4077), .B0(n4205), .B1(n4157), .Y(n3620)
         );
  AOI21X1TS U4376 ( .A0(n3411), .A1(n4644), .B0(n3620), .Y(n3621) );
  AOI22X1TS U4377 ( .A0(n3244), .A1(n4361), .B0(\dataoutbuffer[5][20] ), .B1(
        n4128), .Y(n3625) );
  OAI22X1TS U4378 ( .A0(n3248), .A1(n4077), .B0(n5188), .B1(n4157), .Y(n3623)
         );
  AOI21X1TS U4379 ( .A0(n3249), .A1(n4644), .B0(n3623), .Y(n3624) );
  AOI22X1TS U4380 ( .A0(n3287), .A1(n4361), .B0(\dataoutbuffer[5][21] ), .B1(
        n4128), .Y(n3628) );
  OAI22X1TS U4381 ( .A0(n4043), .A1(n4157), .B0(n4039), .B1(n4077), .Y(n3626)
         );
  AOI21X1TS U4382 ( .A0(n3291), .A1(n4644), .B0(n3626), .Y(n3627) );
  AOI22X1TS U4383 ( .A0(n3155), .A1(n4361), .B0(\dataoutbuffer[5][10] ), .B1(
        n4128), .Y(n3631) );
  OAI22X1TS U4384 ( .A0(n3157), .A1(n4140), .B0(n4022), .B1(n4077), .Y(n3629)
         );
  AOI21X1TS U4385 ( .A0(n3159), .A1(n4644), .B0(n3629), .Y(n3630) );
  AOI22X1TS U4386 ( .A0(n3354), .A1(n4361), .B0(\dataoutbuffer[5][14] ), .B1(
        n4128), .Y(n3634) );
  OAI22X1TS U4387 ( .A0(n3357), .A1(n4140), .B0(n5123), .B1(n4077), .Y(n3632)
         );
  AOI21X1TS U4388 ( .A0(n3355), .A1(n4644), .B0(n3632), .Y(n3633) );
  AOI22X1TS U4389 ( .A0(n3207), .A1(n4361), .B0(\dataoutbuffer[5][17] ), .B1(
        n4128), .Y(n3637) );
  OAI22X1TS U4390 ( .A0(n4206), .A1(n4140), .B0(n5156), .B1(n4077), .Y(n3635)
         );
  AOI21X1TS U4391 ( .A0(n3211), .A1(n4644), .B0(n3635), .Y(n3636) );
  AOI22X1TS U4392 ( .A0(n3297), .A1(n4361), .B0(\dataoutbuffer[5][27] ), .B1(
        n4128), .Y(n3640) );
  OAI22X1TS U4393 ( .A0(n3299), .A1(n4140), .B0(n4004), .B1(n4077), .Y(n3638)
         );
  AOI21X1TS U4394 ( .A0(n3301), .A1(n4644), .B0(n3638), .Y(n3639) );
  AOI22X1TS U4395 ( .A0(n3043), .A1(n4361), .B0(\dataoutbuffer[5][16] ), .B1(
        n4128), .Y(n3643) );
  OAI22X1TS U4396 ( .A0(n3045), .A1(n4077), .B0(n4219), .B1(n4140), .Y(n3641)
         );
  AOI21X1TS U4397 ( .A0(n3047), .A1(n4644), .B0(n3641), .Y(n3642) );
  AOI22X1TS U4398 ( .A0(n3146), .A1(n4455), .B0(\dataoutbuffer[0][24] ), .B1(
        n4787), .Y(n3646) );
  OAI22X1TS U4399 ( .A0(n3700), .A1(n4179), .B0(n3704), .B1(n5227), .Y(n3644)
         );
  AOI21X1TS U4400 ( .A0(n4790), .A1(n3145), .B0(n3644), .Y(n3645) );
  AOI22X1TS U4401 ( .A0(n2964), .A1(n4455), .B0(\dataoutbuffer[0][13] ), .B1(
        n4787), .Y(n3649) );
  OAI22X1TS U4402 ( .A0(n3700), .A1(n4113), .B0(n3704), .B1(n4117), .Y(n3647)
         );
  AOI21X1TS U4403 ( .A0(n4789), .A1(n2962), .B0(n3647), .Y(n3648) );
  AOI22X1TS U4404 ( .A0(n3428), .A1(n4455), .B0(\dataoutbuffer[0][26] ), .B1(
        n4787), .Y(n3652) );
  OAI22X1TS U4405 ( .A0(n3700), .A1(n4089), .B0(n3704), .B1(n4085), .Y(n3650)
         );
  AOI21X1TS U4406 ( .A0(n4789), .A1(n3429), .B0(n3650), .Y(n3651) );
  AOI22X1TS U4407 ( .A0(n3137), .A1(n4455), .B0(\dataoutbuffer[0][31] ), .B1(
        n4787), .Y(n3655) );
  OAI22X1TS U4408 ( .A0(n3700), .A1(n3140), .B0(n3704), .B1(n5308), .Y(n3653)
         );
  AOI21X1TS U4409 ( .A0(n4789), .A1(n3138), .B0(n3653), .Y(n3654) );
  AOI22X1TS U4410 ( .A0(n3354), .A1(n4455), .B0(\dataoutbuffer[0][14] ), .B1(
        n4787), .Y(n3658) );
  OAI22X1TS U4411 ( .A0(n3700), .A1(n3357), .B0(n3704), .B1(n5124), .Y(n3656)
         );
  AOI21X1TS U4412 ( .A0(n4789), .A1(n3355), .B0(n3656), .Y(n3657) );
  AOI22X1TS U4413 ( .A0(n3527), .A1(n4455), .B0(\dataoutbuffer[0][5] ), .B1(
        n4787), .Y(n3661) );
  OAI22X1TS U4414 ( .A0(n3700), .A1(n4141), .B0(n3704), .B1(n5033), .Y(n3659)
         );
  AOI21X1TS U4415 ( .A0(n4789), .A1(n3528), .B0(n3659), .Y(n3660) );
  AOI22X1TS U4416 ( .A0(n2950), .A1(n4455), .B0(\dataoutbuffer[0][23] ), .B1(
        n4787), .Y(n3664) );
  OAI22X1TS U4417 ( .A0(n3699), .A1(n2954), .B0(n3704), .B1(n5217), .Y(n3662)
         );
  AOI21X1TS U4418 ( .A0(n4788), .A1(n2949), .B0(n3662), .Y(n3663) );
  AOI22X1TS U4419 ( .A0(n3481), .A1(n4455), .B0(\dataoutbuffer[0][22] ), .B1(
        n4787), .Y(n3667) );
  OAI22X1TS U4420 ( .A0(n3699), .A1(n3484), .B0(n3704), .B1(n4227), .Y(n3665)
         );
  AOI21X1TS U4421 ( .A0(n4789), .A1(n3482), .B0(n3665), .Y(n3666) );
  AOI22X1TS U4422 ( .A0(n3244), .A1(n4455), .B0(\dataoutbuffer[0][20] ), .B1(
        n4787), .Y(n3670) );
  OAI22X1TS U4423 ( .A0(n3699), .A1(n3248), .B0(n3704), .B1(n5188), .Y(n3668)
         );
  AOI21X1TS U4424 ( .A0(n4788), .A1(n3245), .B0(n3668), .Y(n3669) );
  AOI22X1TS U4425 ( .A0(n3260), .A1(n4455), .B0(\dataoutbuffer[0][19] ), .B1(
        n4787), .Y(n3673) );
  OAI22X1TS U4426 ( .A0(n3699), .A1(n4014), .B0(n3704), .B1(n5177), .Y(n3671)
         );
  AOI21X1TS U4427 ( .A0(n4788), .A1(n3261), .B0(n3671), .Y(n3672) );
  AOI22X1TS U4428 ( .A0(n3019), .A1(n4455), .B0(\dataoutbuffer[0][0] ), .B1(
        n4787), .Y(n3676) );
  OAI22X1TS U4429 ( .A0(n3699), .A1(n4980), .B0(n3704), .B1(n3023), .Y(n3674)
         );
  AOI21X1TS U4430 ( .A0(n4789), .A1(n3017), .B0(n3674), .Y(n3675) );
  AOI22X1TS U4431 ( .A0(n3490), .A1(n4455), .B0(\dataoutbuffer[0][2] ), .B1(
        n4787), .Y(n3679) );
  OAI22X1TS U4432 ( .A0(n3699), .A1(n3494), .B0(n3704), .B1(n5001), .Y(n3677)
         );
  AOI21X1TS U4433 ( .A0(n4789), .A1(n3491), .B0(n3677), .Y(n3678) );
  AOI22X1TS U4434 ( .A0(n3010), .A1(n4455), .B0(\dataoutbuffer[0][1] ), .B1(
        n4787), .Y(n3682) );
  OAI22X1TS U4435 ( .A0(n3699), .A1(n4991), .B0(n3704), .B1(n4990), .Y(n3680)
         );
  AOI21X1TS U4436 ( .A0(n4789), .A1(n3008), .B0(n3680), .Y(n3681) );
  AOI22X1TS U4437 ( .A0(n3164), .A1(n4455), .B0(\dataoutbuffer[0][4] ), .B1(
        n4787), .Y(n3685) );
  OAI22X1TS U4438 ( .A0(n3699), .A1(n5022), .B0(n3704), .B1(n5023), .Y(n3683)
         );
  AOI21X1TS U4439 ( .A0(n4789), .A1(n3165), .B0(n3683), .Y(n3684) );
  AOI22X1TS U4440 ( .A0(n3443), .A1(n4455), .B0(\dataoutbuffer[0][3] ), .B1(
        n4787), .Y(n3688) );
  OAI22X1TS U4441 ( .A0(n3699), .A1(n5012), .B0(n3704), .B1(n5011), .Y(n3686)
         );
  AOI21X1TS U4442 ( .A0(n4789), .A1(n3444), .B0(n3686), .Y(n3687) );
  AOI22X1TS U4443 ( .A0(n3397), .A1(n4455), .B0(\dataoutbuffer[0][28] ), .B1(
        n4787), .Y(n3691) );
  OAI22X1TS U4444 ( .A0(n3700), .A1(n3951), .B0(n3699), .B1(n3947), .Y(n3689)
         );
  AOI21X1TS U4445 ( .A0(n4782), .A1(n3399), .B0(n3689), .Y(n3690) );
  AOI22X1TS U4446 ( .A0(n3457), .A1(n4455), .B0(\dataoutbuffer[0][30] ), .B1(
        n4787), .Y(n3694) );
  OAI22X1TS U4447 ( .A0(n3700), .A1(n4198), .B0(n3699), .B1(n3460), .Y(n3692)
         );
  AOI21X1TS U4448 ( .A0(n4782), .A1(n3458), .B0(n3692), .Y(n3693) );
  AOI22X1TS U4449 ( .A0(n3269), .A1(n4455), .B0(\dataoutbuffer[0][6] ), .B1(
        n4787), .Y(n3697) );
  OAI22X1TS U4450 ( .A0(n3700), .A1(n4018), .B0(n3699), .B1(n5044), .Y(n3695)
         );
  AOI21X1TS U4451 ( .A0(n4782), .A1(n3270), .B0(n3695), .Y(n3696) );
  AOI22X1TS U4452 ( .A0(n3128), .A1(n4455), .B0(\dataoutbuffer[0][29] ), .B1(
        n4787), .Y(n3703) );
  OAI22X1TS U4453 ( .A0(n3700), .A1(n4175), .B0(n3699), .B1(n3127), .Y(n3701)
         );
  AOI21X1TS U4454 ( .A0(n4789), .A1(n3129), .B0(n3701), .Y(n3702) );
  AOI22X1TS U4455 ( .A0(n2964), .A1(n4436), .B0(\dataoutbuffer[1][13] ), .B1(
        n4744), .Y(n3707) );
  OAI22X1TS U4456 ( .A0(n4113), .A1(n4229), .B0(n2966), .B1(n3875), .Y(n3705)
         );
  AOI21X1TS U4457 ( .A0(n2962), .A1(n4759), .B0(n3705), .Y(n3706) );
  NOR3XLTS U4458 ( .A(n3877), .B(n3615), .C(n3708), .Y(n3709) );
  BUFX3TS U4459 ( .A(n3709), .Y(n4380) );
  AOI22X1TS U4460 ( .A0(n3043), .A1(n4380), .B0(\dataoutbuffer[4][16] ), .B1(
        n4671), .Y(n3712) );
  OAI22X1TS U4461 ( .A0(n3827), .A1(n5145), .B0(n3807), .B1(n5146), .Y(n3710)
         );
  AOI21X1TS U4462 ( .A0(n4674), .A1(n3044), .B0(n3710), .Y(n3711) );
  AOI22X1TS U4463 ( .A0(n3244), .A1(n4380), .B0(\dataoutbuffer[4][20] ), .B1(
        n4671), .Y(n3715) );
  OAI22X1TS U4464 ( .A0(n3827), .A1(n5188), .B0(n3807), .B1(n5187), .Y(n3713)
         );
  AOI21X1TS U4465 ( .A0(n4674), .A1(n3247), .B0(n3713), .Y(n3714) );
  AOI22X1TS U4466 ( .A0(n2964), .A1(n4380), .B0(\dataoutbuffer[4][13] ), .B1(
        n4671), .Y(n3718) );
  OAI22X1TS U4467 ( .A0(n3827), .A1(n4117), .B0(n3807), .B1(n2963), .Y(n3716)
         );
  AOI21X1TS U4468 ( .A0(n4674), .A1(n2965), .B0(n3716), .Y(n3717) );
  AOI22X1TS U4469 ( .A0(n3061), .A1(n4380), .B0(\dataoutbuffer[4][9] ), .B1(
        n4671), .Y(n3721) );
  OAI22X1TS U4470 ( .A0(n3827), .A1(n5074), .B0(n3807), .B1(n5075), .Y(n3719)
         );
  AOI21X1TS U4471 ( .A0(n4674), .A1(n3062), .B0(n3719), .Y(n3720) );
  AOI22X1TS U4472 ( .A0(n3198), .A1(n4380), .B0(\dataoutbuffer[4][7] ), .B1(
        n4671), .Y(n3724) );
  OAI22X1TS U4473 ( .A0(n3831), .A1(n3201), .B0(n3807), .B1(n5055), .Y(n3722)
         );
  AOI21X1TS U4474 ( .A0(n4672), .A1(n3199), .B0(n3722), .Y(n3723) );
  AOI22X1TS U4475 ( .A0(n3269), .A1(n4380), .B0(\dataoutbuffer[4][6] ), .B1(
        n4671), .Y(n3727) );
  OAI22X1TS U4476 ( .A0(n3831), .A1(n4018), .B0(n3807), .B1(n5043), .Y(n3725)
         );
  AOI21X1TS U4477 ( .A0(n4672), .A1(n3270), .B0(n3725), .Y(n3726) );
  AOI22X1TS U4478 ( .A0(n3207), .A1(n4380), .B0(\dataoutbuffer[4][17] ), .B1(
        n4671), .Y(n3730) );
  OAI22X1TS U4479 ( .A0(n3831), .A1(n4206), .B0(n3807), .B1(n4207), .Y(n3728)
         );
  AOI21X1TS U4480 ( .A0(n4672), .A1(n3208), .B0(n3728), .Y(n3729) );
  AOI22X1TS U4481 ( .A0(n3052), .A1(n4380), .B0(\dataoutbuffer[4][8] ), .B1(
        n4671), .Y(n3733) );
  OAI22X1TS U4482 ( .A0(n3831), .A1(n4170), .B0(n3807), .B1(n3056), .Y(n3731)
         );
  AOI21X1TS U4483 ( .A0(n4674), .A1(n3053), .B0(n3731), .Y(n3732) );
  AOI22X1TS U4484 ( .A0(n3269), .A1(n4361), .B0(\dataoutbuffer[5][6] ), .B1(
        n4641), .Y(n3736) );
  OAI22X1TS U4485 ( .A0(n5044), .A1(n4077), .B0(n5043), .B1(n4243), .Y(n3734)
         );
  AOI21X1TS U4486 ( .A0(n3270), .A1(n4643), .B0(n3734), .Y(n3735) );
  AOI22X1TS U4487 ( .A0(n3397), .A1(n4361), .B0(\dataoutbuffer[5][28] ), .B1(
        n4641), .Y(n3739) );
  OAI22X1TS U4488 ( .A0(n5270), .A1(n4157), .B0(n3947), .B1(n4077), .Y(n3737)
         );
  AOI21X1TS U4489 ( .A0(n3400), .A1(n4644), .B0(n3737), .Y(n3738) );
  AOI22X1TS U4490 ( .A0(n3198), .A1(n4361), .B0(\dataoutbuffer[5][7] ), .B1(
        n4641), .Y(n3742) );
  OAI22X1TS U4491 ( .A0(n5055), .A1(n4243), .B0(n5054), .B1(n4077), .Y(n3740)
         );
  AOI21X1TS U4492 ( .A0(n3199), .A1(n4643), .B0(n3740), .Y(n3741) );
  AOI22X1TS U4493 ( .A0(n3137), .A1(n4361), .B0(\dataoutbuffer[5][31] ), .B1(
        n4641), .Y(n3745) );
  OAI22X1TS U4494 ( .A0(n3140), .A1(n4140), .B0(n5306), .B1(n4077), .Y(n3743)
         );
  AOI21X1TS U4495 ( .A0(n3138), .A1(n4644), .B0(n3743), .Y(n3744) );
  AOI22X1TS U4496 ( .A0(n3260), .A1(n4361), .B0(\dataoutbuffer[5][19] ), .B1(
        n4641), .Y(n3748) );
  OAI22X1TS U4497 ( .A0(n3262), .A1(n4140), .B0(n4014), .B1(n4077), .Y(n3746)
         );
  AOI21X1TS U4498 ( .A0(n3264), .A1(n4644), .B0(n3746), .Y(n3747) );
  AOI22X1TS U4499 ( .A0(n3443), .A1(n4361), .B0(\dataoutbuffer[5][3] ), .B1(
        n4641), .Y(n3751) );
  OAI22X1TS U4500 ( .A0(n5012), .A1(n4077), .B0(n3985), .B1(n4140), .Y(n3749)
         );
  AOI21X1TS U4501 ( .A0(n3444), .A1(n4644), .B0(n3749), .Y(n3750) );
  AOI22X1TS U4502 ( .A0(n3115), .A1(n4642), .B0(
        \destinationAddressbuffer[5][13] ), .B1(n4641), .Y(n3753) );
  AOI22X1TS U4503 ( .A0(n3116), .A1(n4643), .B0(n3117), .B1(n4644), .Y(n3752)
         );
  AOI22X1TS U4504 ( .A0(n3122), .A1(n4643), .B0(
        \destinationAddressbuffer[5][9] ), .B1(n4641), .Y(n3755) );
  AOI22X1TS U4505 ( .A0(n3123), .A1(n4642), .B0(n3121), .B1(n4644), .Y(n3754)
         );
  AOI22X1TS U4506 ( .A0(n3527), .A1(n4380), .B0(\dataoutbuffer[4][5] ), .B1(
        n4671), .Y(n3758) );
  OAI22X1TS U4507 ( .A0(n3827), .A1(n5033), .B0(n3831), .B1(n4141), .Y(n3756)
         );
  AOI21X1TS U4508 ( .A0(n4674), .A1(n3530), .B0(n3756), .Y(n3757) );
  AOI22X1TS U4509 ( .A0(n3481), .A1(n4380), .B0(\dataoutbuffer[4][22] ), .B1(
        n4671), .Y(n3761) );
  OAI22X1TS U4510 ( .A0(n3827), .A1(n4227), .B0(n3831), .B1(n4223), .Y(n3759)
         );
  AOI21X1TS U4511 ( .A0(n4674), .A1(n3483), .B0(n3759), .Y(n3760) );
  AOI22X1TS U4512 ( .A0(n3397), .A1(n4380), .B0(\dataoutbuffer[4][28] ), .B1(
        n4671), .Y(n3764) );
  OAI22X1TS U4513 ( .A0(n3827), .A1(n5270), .B0(n3831), .B1(n3951), .Y(n3762)
         );
  AOI21X1TS U4514 ( .A0(n4673), .A1(n3400), .B0(n3762), .Y(n3763) );
  AOI22X1TS U4515 ( .A0(n3137), .A1(n4380), .B0(\dataoutbuffer[4][31] ), .B1(
        n4671), .Y(n3767) );
  OAI22X1TS U4516 ( .A0(n3827), .A1(n5308), .B0(n3831), .B1(n3140), .Y(n3765)
         );
  AOI21X1TS U4517 ( .A0(n4673), .A1(n3138), .B0(n3765), .Y(n3766) );
  AOI22X1TS U4518 ( .A0(n3443), .A1(n4380), .B0(\dataoutbuffer[4][3] ), .B1(
        n4671), .Y(n3770) );
  OAI22X1TS U4519 ( .A0(n3827), .A1(n5011), .B0(n3831), .B1(n3985), .Y(n3768)
         );
  AOI21X1TS U4520 ( .A0(n4673), .A1(n3444), .B0(n3768), .Y(n3769) );
  AOI22X1TS U4521 ( .A0(n3407), .A1(n4380), .B0(\dataoutbuffer[4][18] ), .B1(
        n4671), .Y(n3773) );
  OAI22X1TS U4522 ( .A0(n3827), .A1(n4205), .B0(n3831), .B1(n3406), .Y(n3771)
         );
  AOI21X1TS U4523 ( .A0(n4673), .A1(n3411), .B0(n3771), .Y(n3772) );
  AOI22X1TS U4524 ( .A0(n3128), .A1(n4380), .B0(\dataoutbuffer[4][29] ), .B1(
        n4671), .Y(n3776) );
  OAI22X1TS U4525 ( .A0(n3827), .A1(n4171), .B0(n3831), .B1(n4175), .Y(n3774)
         );
  AOI21X1TS U4526 ( .A0(n4673), .A1(n3129), .B0(n3774), .Y(n3775) );
  AOI22X1TS U4527 ( .A0(n3010), .A1(n4380), .B0(\dataoutbuffer[4][1] ), .B1(
        n4671), .Y(n3779) );
  OAI22X1TS U4528 ( .A0(n3826), .A1(n4991), .B0(n3831), .B1(n4084), .Y(n3777)
         );
  AOI21X1TS U4529 ( .A0(n4672), .A1(n3013), .B0(n3777), .Y(n3778) );
  AOI22X1TS U4530 ( .A0(n3019), .A1(n4380), .B0(\dataoutbuffer[4][0] ), .B1(
        n4671), .Y(n3782) );
  OAI22X1TS U4531 ( .A0(n3826), .A1(n4980), .B0(n3831), .B1(n4118), .Y(n3780)
         );
  AOI21X1TS U4532 ( .A0(n4672), .A1(n3022), .B0(n3780), .Y(n3781) );
  AOI22X1TS U4533 ( .A0(n3354), .A1(n4380), .B0(\dataoutbuffer[4][14] ), .B1(
        n4671), .Y(n3785) );
  OAI22X1TS U4534 ( .A0(n3826), .A1(n5123), .B0(n3831), .B1(n3357), .Y(n3783)
         );
  AOI21X1TS U4535 ( .A0(n4673), .A1(n3355), .B0(n3783), .Y(n3784) );
  AOI22X1TS U4536 ( .A0(n3230), .A1(n4380), .B0(\dataoutbuffer[4][25] ), .B1(
        n4671), .Y(n3788) );
  OAI22X1TS U4537 ( .A0(n3826), .A1(n5238), .B0(n3831), .B1(n4183), .Y(n3786)
         );
  AOI21X1TS U4538 ( .A0(n4672), .A1(n3233), .B0(n3786), .Y(n3787) );
  AOI22X1TS U4539 ( .A0(n3342), .A1(n4380), .B0(\dataoutbuffer[4][15] ), .B1(
        n4671), .Y(n3791) );
  OAI22X1TS U4540 ( .A0(n3826), .A1(n3346), .B0(n3831), .B1(n4211), .Y(n3789)
         );
  AOI21X1TS U4541 ( .A0(n4672), .A1(n3341), .B0(n3789), .Y(n3790) );
  AOI22X1TS U4542 ( .A0(n3278), .A1(n4380), .B0(\dataoutbuffer[4][12] ), .B1(
        n4671), .Y(n3794) );
  OAI22X1TS U4543 ( .A0(n3827), .A1(n4162), .B0(n3826), .B1(n4044), .Y(n3792)
         );
  AOI21X1TS U4544 ( .A0(n4666), .A1(n3279), .B0(n3792), .Y(n3793) );
  AOI22X1TS U4545 ( .A0(n2950), .A1(n4380), .B0(\dataoutbuffer[4][23] ), .B1(
        n4671), .Y(n3797) );
  OAI22X1TS U4546 ( .A0(n3827), .A1(n5217), .B0(n3826), .B1(n2954), .Y(n3795)
         );
  AOI21X1TS U4547 ( .A0(n4666), .A1(n2949), .B0(n3795), .Y(n3796) );
  AOI22X1TS U4548 ( .A0(n3287), .A1(n4380), .B0(\dataoutbuffer[4][21] ), .B1(
        n4671), .Y(n3800) );
  OAI22X1TS U4549 ( .A0(n3827), .A1(n4043), .B0(n3826), .B1(n4039), .Y(n3798)
         );
  AOI21X1TS U4550 ( .A0(n4666), .A1(n3288), .B0(n3798), .Y(n3799) );
  AOI22X1TS U4551 ( .A0(n3260), .A1(n4380), .B0(\dataoutbuffer[4][19] ), .B1(
        n4671), .Y(n3803) );
  OAI22X1TS U4552 ( .A0(n3827), .A1(n5177), .B0(n3826), .B1(n4014), .Y(n3801)
         );
  AOI21X1TS U4553 ( .A0(n4666), .A1(n3261), .B0(n3801), .Y(n3802) );
  AOI22X1TS U4554 ( .A0(n3155), .A1(n4380), .B0(\dataoutbuffer[4][10] ), .B1(
        n4671), .Y(n3806) );
  OAI22X1TS U4555 ( .A0(n3827), .A1(n5085), .B0(n3826), .B1(n4022), .Y(n3804)
         );
  AOI21X1TS U4556 ( .A0(n4666), .A1(n3156), .B0(n3804), .Y(n3805) );
  AOI22X1TS U4557 ( .A0(n3146), .A1(n4380), .B0(\dataoutbuffer[4][24] ), .B1(
        n4671), .Y(n3810) );
  OAI22X1TS U4558 ( .A0(n3827), .A1(n5227), .B0(n3826), .B1(n5228), .Y(n3808)
         );
  AOI21X1TS U4559 ( .A0(n4673), .A1(n3149), .B0(n3808), .Y(n3809) );
  AOI22X1TS U4560 ( .A0(n3457), .A1(n4380), .B0(\dataoutbuffer[4][30] ), .B1(
        n4671), .Y(n3813) );
  OAI22X1TS U4561 ( .A0(n3827), .A1(n5293), .B0(n3826), .B1(n3460), .Y(n3811)
         );
  AOI21X1TS U4562 ( .A0(n4673), .A1(n3456), .B0(n3811), .Y(n3812) );
  AOI22X1TS U4563 ( .A0(n3164), .A1(n4380), .B0(\dataoutbuffer[4][4] ), .B1(
        n4671), .Y(n3816) );
  OAI22X1TS U4564 ( .A0(n3827), .A1(n5023), .B0(n3826), .B1(n5022), .Y(n3814)
         );
  AOI21X1TS U4565 ( .A0(n4673), .A1(n3165), .B0(n3814), .Y(n3815) );
  AOI22X1TS U4566 ( .A0(n3297), .A1(n4380), .B0(\dataoutbuffer[4][27] ), .B1(
        n4671), .Y(n3819) );
  OAI22X1TS U4567 ( .A0(n3827), .A1(n5259), .B0(n3826), .B1(n4004), .Y(n3817)
         );
  AOI21X1TS U4568 ( .A0(n4673), .A1(n3301), .B0(n3817), .Y(n3818) );
  AOI22X1TS U4569 ( .A0(n3363), .A1(n4380), .B0(\dataoutbuffer[4][11] ), .B1(
        n4671), .Y(n3822) );
  OAI22X1TS U4570 ( .A0(n3827), .A1(n4106), .B0(n3826), .B1(n4029), .Y(n3820)
         );
  AOI21X1TS U4571 ( .A0(n4673), .A1(n3364), .B0(n3820), .Y(n3821) );
  AOI22X1TS U4572 ( .A0(n3490), .A1(n4380), .B0(\dataoutbuffer[4][2] ), .B1(
        n4671), .Y(n3825) );
  OAI22X1TS U4573 ( .A0(n3827), .A1(n5001), .B0(n3826), .B1(n3494), .Y(n3823)
         );
  AOI21X1TS U4574 ( .A0(n4673), .A1(n3491), .B0(n3823), .Y(n3824) );
  AOI22X1TS U4575 ( .A0(n3428), .A1(n4380), .B0(\dataoutbuffer[4][26] ), .B1(
        n4671), .Y(n3830) );
  OAI22X1TS U4576 ( .A0(n3827), .A1(n4085), .B0(n3826), .B1(n4060), .Y(n3828)
         );
  AOI21X1TS U4577 ( .A0(n4673), .A1(n3429), .B0(n3828), .Y(n3829) );
  AOI22X1TS U4578 ( .A0(n3397), .A1(n4436), .B0(\dataoutbuffer[1][28] ), .B1(
        n4757), .Y(n3834) );
  OAI22X1TS U4579 ( .A0(n5270), .A1(n4240), .B0(n3947), .B1(n3875), .Y(n3832)
         );
  AOI21X1TS U4580 ( .A0(n3400), .A1(n4759), .B0(n3832), .Y(n3833) );
  AOI22X1TS U4581 ( .A0(n3527), .A1(n4436), .B0(\dataoutbuffer[1][5] ), .B1(
        n4757), .Y(n3837) );
  OAI22X1TS U4582 ( .A0(n5033), .A1(n4240), .B0(n3531), .B1(n3875), .Y(n3835)
         );
  AOI21X1TS U4583 ( .A0(n3528), .A1(n4759), .B0(n3835), .Y(n3836) );
  AOI22X1TS U4584 ( .A0(n3198), .A1(n4436), .B0(\dataoutbuffer[1][7] ), .B1(
        n4757), .Y(n3840) );
  OAI22X1TS U4585 ( .A0(n5055), .A1(n4228), .B0(n5054), .B1(n3875), .Y(n3838)
         );
  AOI21X1TS U4586 ( .A0(n3199), .A1(n4758), .B0(n3838), .Y(n3839) );
  AOI22X1TS U4587 ( .A0(n3297), .A1(n4436), .B0(\dataoutbuffer[1][27] ), .B1(
        n4757), .Y(n3843) );
  OAI22X1TS U4588 ( .A0(n4004), .A1(n3875), .B0(n5259), .B1(n4240), .Y(n3841)
         );
  AOI21X1TS U4589 ( .A0(n3301), .A1(n4759), .B0(n3841), .Y(n3842) );
  AOI22X1TS U4590 ( .A0(n3269), .A1(n4436), .B0(\dataoutbuffer[1][6] ), .B1(
        n4757), .Y(n3846) );
  OAI22X1TS U4591 ( .A0(n5044), .A1(n3875), .B0(n5043), .B1(n4228), .Y(n3844)
         );
  AOI21X1TS U4592 ( .A0(n3270), .A1(n4758), .B0(n3844), .Y(n3845) );
  AOI22X1TS U4593 ( .A0(n3443), .A1(n4436), .B0(\dataoutbuffer[1][3] ), .B1(
        n4757), .Y(n3849) );
  OAI22X1TS U4594 ( .A0(n5012), .A1(n3875), .B0(n5011), .B1(n4240), .Y(n3847)
         );
  AOI21X1TS U4595 ( .A0(n3444), .A1(n4759), .B0(n3847), .Y(n3848) );
  AOI22X1TS U4596 ( .A0(n3428), .A1(n4436), .B0(\dataoutbuffer[1][26] ), .B1(
        n4757), .Y(n3852) );
  OAI22X1TS U4597 ( .A0(n4089), .A1(n4229), .B0(n4060), .B1(n3875), .Y(n3850)
         );
  AOI21X1TS U4598 ( .A0(n3429), .A1(n4759), .B0(n3850), .Y(n3851) );
  AOI22X1TS U4599 ( .A0(n3164), .A1(n4436), .B0(\dataoutbuffer[1][4] ), .B1(
        n4757), .Y(n3855) );
  OAI22X1TS U4600 ( .A0(n5022), .A1(n3875), .B0(n4136), .B1(n4229), .Y(n3853)
         );
  AOI21X1TS U4601 ( .A0(n3165), .A1(n4759), .B0(n3853), .Y(n3854) );
  AOI22X1TS U4602 ( .A0(n3490), .A1(n4436), .B0(\dataoutbuffer[1][2] ), .B1(
        n4757), .Y(n3858) );
  OAI22X1TS U4603 ( .A0(n3494), .A1(n3875), .B0(n4132), .B1(n4229), .Y(n3856)
         );
  AOI21X1TS U4604 ( .A0(n3491), .A1(n4759), .B0(n3856), .Y(n3857) );
  AOI22X1TS U4605 ( .A0(n3287), .A1(n4436), .B0(\dataoutbuffer[1][21] ), .B1(
        n4757), .Y(n3861) );
  OAI22X1TS U4606 ( .A0(n3292), .A1(n4228), .B0(n4039), .B1(n3875), .Y(n3859)
         );
  AOI21X1TS U4607 ( .A0(n3288), .A1(n4760), .B0(n3859), .Y(n3860) );
  AOI22X1TS U4608 ( .A0(n3010), .A1(n4436), .B0(\dataoutbuffer[1][1] ), .B1(
        n4757), .Y(n3864) );
  OAI22X1TS U4609 ( .A0(n4991), .A1(n3875), .B0(n4084), .B1(n4229), .Y(n3862)
         );
  AOI21X1TS U4610 ( .A0(n3008), .A1(n4759), .B0(n3862), .Y(n3863) );
  AOI22X1TS U4611 ( .A0(n3260), .A1(n4436), .B0(\dataoutbuffer[1][19] ), .B1(
        n4757), .Y(n3867) );
  OAI22X1TS U4612 ( .A0(n3262), .A1(n4229), .B0(n4014), .B1(n3875), .Y(n3865)
         );
  AOI21X1TS U4613 ( .A0(n3264), .A1(n4759), .B0(n3865), .Y(n3866) );
  AOI22X1TS U4614 ( .A0(n3019), .A1(n4436), .B0(\dataoutbuffer[1][0] ), .B1(
        n4757), .Y(n3870) );
  OAI22X1TS U4615 ( .A0(n4980), .A1(n3875), .B0(n4118), .B1(n4229), .Y(n3868)
         );
  AOI21X1TS U4616 ( .A0(n3017), .A1(n4759), .B0(n3868), .Y(n3869) );
  AOI22X1TS U4617 ( .A0(n3116), .A1(n4758), .B0(
        \destinationAddressbuffer[1][13] ), .B1(n4757), .Y(n3872) );
  AOI22X1TS U4618 ( .A0(n3115), .A1(n4760), .B0(n3117), .B1(n4759), .Y(n3871)
         );
  AOI22X1TS U4619 ( .A0(n3123), .A1(n4760), .B0(
        \destinationAddressbuffer[1][9] ), .B1(n4757), .Y(n3874) );
  AOI22X1TS U4620 ( .A0(n3121), .A1(n4759), .B0(n3122), .B1(n4758), .Y(n3873)
         );
  NOR3XLTS U4621 ( .A(n3877), .B(n3876), .C(n3615), .Y(n3878) );
  BUFX3TS U4622 ( .A(n3878), .Y(n4342) );
  AOI22X1TS U4623 ( .A0(n3397), .A1(n4342), .B0(\dataoutbuffer[6][28] ), .B1(
        n4612), .Y(n3881) );
  OAI22X1TS U4624 ( .A0(n4064), .A1(n3401), .B0(n4076), .B1(n3951), .Y(n3879)
         );
  AOI21X1TS U4625 ( .A0(n4614), .A1(n3398), .B0(n3879), .Y(n3880) );
  AOI22X1TS U4626 ( .A0(n3407), .A1(n4342), .B0(\dataoutbuffer[6][18] ), .B1(
        n4612), .Y(n3884) );
  OAI22X1TS U4627 ( .A0(n4064), .A1(n5166), .B0(n4076), .B1(n3406), .Y(n3882)
         );
  AOI21X1TS U4628 ( .A0(n4614), .A1(n3408), .B0(n3882), .Y(n3883) );
  AOI22X1TS U4629 ( .A0(n3198), .A1(n4342), .B0(\dataoutbuffer[6][7] ), .B1(
        n4612), .Y(n3887) );
  OAI22X1TS U4630 ( .A0(n4064), .A1(n5055), .B0(n4076), .B1(n3201), .Y(n3885)
         );
  AOI21X1TS U4631 ( .A0(n4613), .A1(n3199), .B0(n3885), .Y(n3886) );
  AOI22X1TS U4632 ( .A0(n3122), .A1(n4583), .B0(
        \destinationAddressbuffer[7][9] ), .B1(n4318), .Y(n3889) );
  AOI22X1TS U4633 ( .A0(n3123), .A1(n4580), .B0(n3121), .B1(n4586), .Y(n3888)
         );
  AOI22X1TS U4634 ( .A0(n3115), .A1(n4580), .B0(
        \destinationAddressbuffer[7][13] ), .B1(n4318), .Y(n3892) );
  AOI22X1TS U4635 ( .A0(n3116), .A1(n4583), .B0(n3117), .B1(n4586), .Y(n3891)
         );
  AOI22X1TS U4636 ( .A0(n3035), .A1(n4583), .B0(
        \destinationAddressbuffer[7][12] ), .B1(n4318), .Y(n3895) );
  AOI22X1TS U4637 ( .A0(n3038), .A1(n4584), .B0(n3039), .B1(n4580), .Y(n3894)
         );
  AOI22X1TS U4638 ( .A0(n3031), .A1(n4580), .B0(
        \destinationAddressbuffer[7][10] ), .B1(n4318), .Y(n3897) );
  AOI22X1TS U4639 ( .A0(n3030), .A1(n4584), .B0(n3028), .B1(n4583), .Y(n3896)
         );
  AOI22X1TS U4640 ( .A0(n3137), .A1(n4323), .B0(\dataoutbuffer[7][31] ), .B1(
        n4318), .Y(n3900) );
  OAI22X1TS U4641 ( .A0(n3140), .A1(n3975), .B0(n5306), .B1(n3968), .Y(n3898)
         );
  AOI21X1TS U4642 ( .A0(n3138), .A1(n4586), .B0(n3898), .Y(n3899) );
  AOI22X1TS U4643 ( .A0(n3230), .A1(n4323), .B0(\dataoutbuffer[7][25] ), .B1(
        n4318), .Y(n3903) );
  OAI22X1TS U4644 ( .A0(n3236), .A1(n3969), .B0(n4183), .B1(n3975), .Y(n3901)
         );
  AOI21X1TS U4645 ( .A0(n3234), .A1(n4584), .B0(n3901), .Y(n3902) );
  AOI22X1TS U4646 ( .A0(n3481), .A1(n4323), .B0(\dataoutbuffer[7][22] ), .B1(
        n4318), .Y(n3906) );
  OAI22X1TS U4647 ( .A0(n3484), .A1(n3968), .B0(n4223), .B1(n3975), .Y(n3904)
         );
  AOI21X1TS U4648 ( .A0(n3482), .A1(n4586), .B0(n3904), .Y(n3905) );
  AOI22X1TS U4649 ( .A0(n3269), .A1(n4323), .B0(\dataoutbuffer[7][6] ), .B1(
        n4318), .Y(n3909) );
  OAI22X1TS U4650 ( .A0(n5044), .A1(n3968), .B0(n4018), .B1(n3975), .Y(n3907)
         );
  AOI21X1TS U4651 ( .A0(n3273), .A1(n4586), .B0(n3907), .Y(n3908) );
  AOI22X1TS U4652 ( .A0(n3244), .A1(n4323), .B0(\dataoutbuffer[7][20] ), .B1(
        n4318), .Y(n3912) );
  OAI22X1TS U4653 ( .A0(n3246), .A1(n3975), .B0(n5187), .B1(n3969), .Y(n3910)
         );
  AOI21X1TS U4654 ( .A0(n3247), .A1(n4584), .B0(n3910), .Y(n3911) );
  AOI22X1TS U4655 ( .A0(n3073), .A1(n4580), .B0(
        \destinationAddressbuffer[7][11] ), .B1(n4318), .Y(n3914) );
  AOI22X1TS U4656 ( .A0(n3077), .A1(n4584), .B0(n3078), .B1(n4586), .Y(n3913)
         );
  AOI22X1TS U4657 ( .A0(n3128), .A1(n4323), .B0(\dataoutbuffer[7][29] ), .B1(
        n4318), .Y(n3917) );
  OAI22X1TS U4658 ( .A0(n3130), .A1(n3969), .B0(n4175), .B1(n3975), .Y(n3915)
         );
  AOI21X1TS U4659 ( .A0(n3126), .A1(n4584), .B0(n3915), .Y(n3916) );
  AOI22X1TS U4660 ( .A0(n3260), .A1(n4323), .B0(\dataoutbuffer[7][19] ), .B1(
        n4318), .Y(n3920) );
  OAI22X1TS U4661 ( .A0(n3262), .A1(n3975), .B0(n5176), .B1(n3969), .Y(n3918)
         );
  AOI21X1TS U4662 ( .A0(n3263), .A1(n4584), .B0(n3918), .Y(n3919) );
  AOI22X1TS U4663 ( .A0(n2990), .A1(n4580), .B0(
        \destinationAddressbuffer[7][8] ), .B1(n4318), .Y(n3922) );
  AOI22X1TS U4664 ( .A0(n2989), .A1(n4584), .B0(n2988), .B1(n4586), .Y(n3921)
         );
  AOI22X1TS U4665 ( .A0(n3428), .A1(n4323), .B0(\dataoutbuffer[7][26] ), .B1(
        n4318), .Y(n3925) );
  OAI22X1TS U4666 ( .A0(n3430), .A1(n3969), .B0(n4089), .B1(n3975), .Y(n3923)
         );
  AOI21X1TS U4667 ( .A0(n3431), .A1(n4584), .B0(n3923), .Y(n3924) );
  AOI22X1TS U4668 ( .A0(n3146), .A1(n4323), .B0(\dataoutbuffer[7][24] ), .B1(
        n4318), .Y(n3928) );
  OAI22X1TS U4669 ( .A0(n5228), .A1(n3968), .B0(n5227), .B1(n3964), .Y(n3926)
         );
  AOI21X1TS U4670 ( .A0(n3149), .A1(n4586), .B0(n3926), .Y(n3927) );
  AOI22X1TS U4671 ( .A0(n2950), .A1(n4323), .B0(\dataoutbuffer[7][23] ), .B1(
        n4318), .Y(n3931) );
  OAI22X1TS U4672 ( .A0(n5217), .A1(n3964), .B0(n2958), .B1(n3969), .Y(n3929)
         );
  AOI21X1TS U4673 ( .A0(n2953), .A1(n4584), .B0(n3929), .Y(n3930) );
  AOI22X1TS U4674 ( .A0(n3407), .A1(n4323), .B0(\dataoutbuffer[7][18] ), .B1(
        n4318), .Y(n3934) );
  OAI22X1TS U4675 ( .A0(n5166), .A1(n3969), .B0(n4205), .B1(n3964), .Y(n3932)
         );
  AOI21X1TS U4676 ( .A0(n3408), .A1(n4584), .B0(n3932), .Y(n3933) );
  AOI22X1TS U4677 ( .A0(n3019), .A1(n4323), .B0(\dataoutbuffer[7][0] ), .B1(
        n4318), .Y(n3937) );
  OAI22X1TS U4678 ( .A0(n3023), .A1(n3964), .B0(n4980), .B1(n3968), .Y(n3935)
         );
  AOI21X1TS U4679 ( .A0(n3017), .A1(n4586), .B0(n3935), .Y(n3936) );
  AOI22X1TS U4680 ( .A0(n3490), .A1(n4323), .B0(\dataoutbuffer[7][2] ), .B1(
        n4318), .Y(n3940) );
  OAI22X1TS U4681 ( .A0(n5001), .A1(n3964), .B0(n3494), .B1(n3968), .Y(n3938)
         );
  AOI21X1TS U4682 ( .A0(n3491), .A1(n4586), .B0(n3938), .Y(n3939) );
  AOI22X1TS U4683 ( .A0(n3457), .A1(n4323), .B0(\dataoutbuffer[7][30] ), .B1(
        n4318), .Y(n3943) );
  OAI22X1TS U4684 ( .A0(n5293), .A1(n3964), .B0(n5292), .B1(n3969), .Y(n3941)
         );
  AOI21X1TS U4685 ( .A0(n3459), .A1(n4584), .B0(n3941), .Y(n3942) );
  AOI22X1TS U4686 ( .A0(n3297), .A1(n4323), .B0(\dataoutbuffer[7][27] ), .B1(
        n4318), .Y(n3946) );
  OAI22X1TS U4687 ( .A0(n5260), .A1(n3969), .B0(n5259), .B1(n3964), .Y(n3944)
         );
  AOI21X1TS U4688 ( .A0(n3300), .A1(n4584), .B0(n3944), .Y(n3945) );
  AOI22X1TS U4689 ( .A0(n3397), .A1(n4323), .B0(\dataoutbuffer[7][28] ), .B1(
        n4318), .Y(n3950) );
  OAI22X1TS U4690 ( .A0(n5270), .A1(n3964), .B0(n3947), .B1(n3968), .Y(n3948)
         );
  AOI21X1TS U4691 ( .A0(n3400), .A1(n4586), .B0(n3948), .Y(n3949) );
  AOI22X1TS U4692 ( .A0(n3287), .A1(n4323), .B0(\dataoutbuffer[7][21] ), .B1(
        n4318), .Y(n3954) );
  OAI22X1TS U4693 ( .A0(n3292), .A1(n3969), .B0(n4043), .B1(n3964), .Y(n3952)
         );
  AOI21X1TS U4694 ( .A0(n3290), .A1(n4584), .B0(n3952), .Y(n3953) );
  AOI22X1TS U4695 ( .A0(n3527), .A1(n4323), .B0(\dataoutbuffer[7][5] ), .B1(
        n4318), .Y(n3957) );
  OAI22X1TS U4696 ( .A0(n5033), .A1(n3964), .B0(n3531), .B1(n3968), .Y(n3955)
         );
  AOI21X1TS U4697 ( .A0(n3528), .A1(n4586), .B0(n3955), .Y(n3956) );
  AOI22X1TS U4698 ( .A0(n3010), .A1(n4323), .B0(\dataoutbuffer[7][1] ), .B1(
        n4318), .Y(n3960) );
  OAI22X1TS U4699 ( .A0(n4991), .A1(n3968), .B0(n4990), .B1(n3964), .Y(n3958)
         );
  AOI21X1TS U4700 ( .A0(n3008), .A1(n4586), .B0(n3958), .Y(n3959) );
  AOI22X1TS U4701 ( .A0(n3443), .A1(n4323), .B0(\dataoutbuffer[7][3] ), .B1(
        n4318), .Y(n3963) );
  OAI22X1TS U4702 ( .A0(n5012), .A1(n3968), .B0(n5011), .B1(n3964), .Y(n3961)
         );
  AOI21X1TS U4703 ( .A0(n3444), .A1(n4586), .B0(n3961), .Y(n3962) );
  AOI22X1TS U4704 ( .A0(n3164), .A1(n4323), .B0(\dataoutbuffer[7][4] ), .B1(
        n4318), .Y(n3967) );
  OAI22X1TS U4705 ( .A0(n5023), .A1(n3964), .B0(n5022), .B1(n3968), .Y(n3965)
         );
  AOI21X1TS U4706 ( .A0(n3165), .A1(n4586), .B0(n3965), .Y(n3966) );
  AOI22X1TS U4707 ( .A0(n3198), .A1(n4323), .B0(\dataoutbuffer[7][7] ), .B1(
        n4318), .Y(n3972) );
  OAI22X1TS U4708 ( .A0(n5055), .A1(n3969), .B0(n5054), .B1(n3968), .Y(n3970)
         );
  AOI21X1TS U4709 ( .A0(n3199), .A1(n4583), .B0(n3970), .Y(n3971) );
  AOI22X1TS U4710 ( .A0(n2979), .A1(n4583), .B0(writeOutbuffer[7]), .B1(n4318), 
        .Y(n3974) );
  AOI22X1TS U4711 ( .A0(n2982), .A1(n4584), .B0(n2980), .B1(n4586), .Y(n3973)
         );
  AOI22X1TS U4712 ( .A0(n3061), .A1(n4342), .B0(\dataoutbuffer[6][9] ), .B1(
        n4612), .Y(n3978) );
  OAI22X1TS U4713 ( .A0(n4076), .A1(n3064), .B0(n4072), .B1(n5074), .Y(n3976)
         );
  AOI21X1TS U4714 ( .A0(n4614), .A1(n3062), .B0(n3976), .Y(n3977) );
  AOI22X1TS U4715 ( .A0(n3137), .A1(n4342), .B0(\dataoutbuffer[6][31] ), .B1(
        n4612), .Y(n3981) );
  OAI22X1TS U4716 ( .A0(n4076), .A1(n3140), .B0(n4072), .B1(n5308), .Y(n3979)
         );
  AOI21X1TS U4717 ( .A0(n4615), .A1(n3138), .B0(n3979), .Y(n3980) );
  AOI22X1TS U4718 ( .A0(n3230), .A1(n4342), .B0(\dataoutbuffer[6][25] ), .B1(
        n4612), .Y(n3984) );
  OAI22X1TS U4719 ( .A0(n4076), .A1(n4183), .B0(n4072), .B1(n5239), .Y(n3982)
         );
  AOI21X1TS U4720 ( .A0(n4615), .A1(n3235), .B0(n3982), .Y(n3983) );
  AOI22X1TS U4721 ( .A0(n3443), .A1(n4342), .B0(\dataoutbuffer[6][3] ), .B1(
        n4612), .Y(n3988) );
  OAI22X1TS U4722 ( .A0(n4076), .A1(n3985), .B0(n4072), .B1(n5011), .Y(n3986)
         );
  AOI21X1TS U4723 ( .A0(n4615), .A1(n3444), .B0(n3986), .Y(n3987) );
  AOI22X1TS U4724 ( .A0(n3527), .A1(n4342), .B0(\dataoutbuffer[6][5] ), .B1(
        n4612), .Y(n3991) );
  OAI22X1TS U4725 ( .A0(n4064), .A1(n3529), .B0(n4072), .B1(n5033), .Y(n3989)
         );
  AOI21X1TS U4726 ( .A0(n4614), .A1(n3530), .B0(n3989), .Y(n3990) );
  AOI22X1TS U4727 ( .A0(n3052), .A1(n4342), .B0(\dataoutbuffer[6][8] ), .B1(
        n4612), .Y(n3994) );
  OAI22X1TS U4728 ( .A0(n4064), .A1(n3056), .B0(n4072), .B1(n4166), .Y(n3992)
         );
  AOI21X1TS U4729 ( .A0(n4614), .A1(n3053), .B0(n3992), .Y(n3993) );
  AOI22X1TS U4730 ( .A0(n3146), .A1(n4342), .B0(\dataoutbuffer[6][24] ), .B1(
        n4612), .Y(n3997) );
  OAI22X1TS U4731 ( .A0(n4064), .A1(n3150), .B0(n4072), .B1(n5227), .Y(n3995)
         );
  AOI21X1TS U4732 ( .A0(n4616), .A1(n3147), .B0(n3995), .Y(n3996) );
  AOI22X1TS U4733 ( .A0(n3043), .A1(n4342), .B0(\dataoutbuffer[6][16] ), .B1(
        n4612), .Y(n4000) );
  OAI22X1TS U4734 ( .A0(n4064), .A1(n5146), .B0(n4072), .B1(n5145), .Y(n3998)
         );
  AOI21X1TS U4735 ( .A0(n4616), .A1(n3046), .B0(n3998), .Y(n3999) );
  AOI22X1TS U4736 ( .A0(n3128), .A1(n4342), .B0(\dataoutbuffer[6][29] ), .B1(
        n4612), .Y(n4003) );
  OAI22X1TS U4737 ( .A0(n4076), .A1(n4175), .B0(n4071), .B1(n3127), .Y(n4001)
         );
  AOI21X1TS U4738 ( .A0(n4613), .A1(n3132), .B0(n4001), .Y(n4002) );
  AOI22X1TS U4739 ( .A0(n3297), .A1(n4342), .B0(\dataoutbuffer[6][27] ), .B1(
        n4612), .Y(n4007) );
  OAI22X1TS U4740 ( .A0(n4076), .A1(n3299), .B0(n4071), .B1(n4004), .Y(n4005)
         );
  AOI21X1TS U4741 ( .A0(n4613), .A1(n3296), .B0(n4005), .Y(n4006) );
  AOI22X1TS U4742 ( .A0(n3342), .A1(n4342), .B0(\dataoutbuffer[6][15] ), .B1(
        n4612), .Y(n4010) );
  OAI22X1TS U4743 ( .A0(n4076), .A1(n4211), .B0(n4071), .B1(n3346), .Y(n4008)
         );
  AOI21X1TS U4744 ( .A0(n4613), .A1(n3341), .B0(n4008), .Y(n4009) );
  AOI22X1TS U4745 ( .A0(n3457), .A1(n4342), .B0(\dataoutbuffer[6][30] ), .B1(
        n4612), .Y(n4013) );
  OAI22X1TS U4746 ( .A0(n4076), .A1(n4198), .B0(n4071), .B1(n3460), .Y(n4011)
         );
  AOI21X1TS U4747 ( .A0(n4615), .A1(n3456), .B0(n4011), .Y(n4012) );
  AOI22X1TS U4748 ( .A0(n3260), .A1(n4342), .B0(\dataoutbuffer[6][19] ), .B1(
        n4612), .Y(n4017) );
  OAI22X1TS U4749 ( .A0(n4064), .A1(n5176), .B0(n4071), .B1(n4014), .Y(n4015)
         );
  AOI21X1TS U4750 ( .A0(n4613), .A1(n3259), .B0(n4015), .Y(n4016) );
  AOI22X1TS U4751 ( .A0(n3269), .A1(n4342), .B0(\dataoutbuffer[6][6] ), .B1(
        n4612), .Y(n4021) );
  OAI22X1TS U4752 ( .A0(n4076), .A1(n4018), .B0(n4071), .B1(n5044), .Y(n4019)
         );
  AOI21X1TS U4753 ( .A0(n4613), .A1(n3270), .B0(n4019), .Y(n4020) );
  AOI22X1TS U4754 ( .A0(n3155), .A1(n4342), .B0(\dataoutbuffer[6][10] ), .B1(
        n4612), .Y(n4025) );
  OAI22X1TS U4755 ( .A0(n4064), .A1(n5086), .B0(n4071), .B1(n4022), .Y(n4023)
         );
  AOI21X1TS U4756 ( .A0(n4616), .A1(n3156), .B0(n4023), .Y(n4024) );
  AOI22X1TS U4757 ( .A0(n3019), .A1(n4342), .B0(\dataoutbuffer[6][0] ), .B1(
        n4612), .Y(n4028) );
  OAI22X1TS U4758 ( .A0(n4064), .A1(n3018), .B0(n4071), .B1(n4980), .Y(n4026)
         );
  AOI21X1TS U4759 ( .A0(n4616), .A1(n3021), .B0(n4026), .Y(n4027) );
  AOI22X1TS U4760 ( .A0(n3363), .A1(n4342), .B0(\dataoutbuffer[6][11] ), .B1(
        n4612), .Y(n4032) );
  OAI22X1TS U4761 ( .A0(n4064), .A1(n3365), .B0(n4071), .B1(n4029), .Y(n4030)
         );
  AOI21X1TS U4762 ( .A0(n4613), .A1(n3366), .B0(n4030), .Y(n4031) );
  AOI22X1TS U4763 ( .A0(n3207), .A1(n4342), .B0(\dataoutbuffer[6][17] ), .B1(
        n4612), .Y(n4035) );
  OAI22X1TS U4764 ( .A0(n4064), .A1(n4207), .B0(n4071), .B1(n5156), .Y(n4033)
         );
  AOI21X1TS U4765 ( .A0(n4613), .A1(n3208), .B0(n4033), .Y(n4034) );
  AOI22X1TS U4766 ( .A0(n3481), .A1(n4342), .B0(\dataoutbuffer[6][22] ), .B1(
        n4612), .Y(n4038) );
  OAI22X1TS U4767 ( .A0(n4064), .A1(n5207), .B0(n4071), .B1(n3484), .Y(n4036)
         );
  AOI21X1TS U4768 ( .A0(n4616), .A1(n3480), .B0(n4036), .Y(n4037) );
  AOI22X1TS U4769 ( .A0(n3287), .A1(n4342), .B0(\dataoutbuffer[6][21] ), .B1(
        n4612), .Y(n4042) );
  OAI22X1TS U4770 ( .A0(n4064), .A1(n3292), .B0(n4071), .B1(n4039), .Y(n4040)
         );
  AOI21X1TS U4771 ( .A0(n4616), .A1(n3288), .B0(n4040), .Y(n4041) );
  AOI22X1TS U4772 ( .A0(n3278), .A1(n4342), .B0(\dataoutbuffer[6][12] ), .B1(
        n4612), .Y(n4047) );
  OAI22X1TS U4773 ( .A0(n4072), .A1(n4162), .B0(n4071), .B1(n4044), .Y(n4045)
         );
  AOI21X1TS U4774 ( .A0(n4615), .A1(n3282), .B0(n4045), .Y(n4046) );
  AOI22X1TS U4775 ( .A0(n3244), .A1(n4342), .B0(\dataoutbuffer[6][20] ), .B1(
        n4612), .Y(n4050) );
  OAI22X1TS U4776 ( .A0(n4072), .A1(n5188), .B0(n4071), .B1(n3248), .Y(n4048)
         );
  AOI21X1TS U4777 ( .A0(n4615), .A1(n3249), .B0(n4048), .Y(n4049) );
  AOI22X1TS U4778 ( .A0(n3164), .A1(n4342), .B0(\dataoutbuffer[6][4] ), .B1(
        n4612), .Y(n4053) );
  OAI22X1TS U4779 ( .A0(n4072), .A1(n5023), .B0(n4071), .B1(n5022), .Y(n4051)
         );
  AOI21X1TS U4780 ( .A0(n4616), .A1(n3167), .B0(n4051), .Y(n4052) );
  AOI22X1TS U4781 ( .A0(n3490), .A1(n4342), .B0(\dataoutbuffer[6][2] ), .B1(
        n4612), .Y(n4056) );
  OAI22X1TS U4782 ( .A0(n4072), .A1(n5001), .B0(n4071), .B1(n3494), .Y(n4054)
         );
  AOI21X1TS U4783 ( .A0(n4616), .A1(n3489), .B0(n4054), .Y(n4055) );
  AOI22X1TS U4784 ( .A0(n3010), .A1(n4342), .B0(\dataoutbuffer[6][1] ), .B1(
        n4612), .Y(n4059) );
  OAI22X1TS U4785 ( .A0(n4072), .A1(n4990), .B0(n4071), .B1(n4991), .Y(n4057)
         );
  AOI21X1TS U4786 ( .A0(n4616), .A1(n3012), .B0(n4057), .Y(n4058) );
  AOI22X1TS U4787 ( .A0(n3428), .A1(n4342), .B0(\dataoutbuffer[6][26] ), .B1(
        n4612), .Y(n4063) );
  OAI22X1TS U4788 ( .A0(n4072), .A1(n4085), .B0(n4071), .B1(n4060), .Y(n4061)
         );
  AOI21X1TS U4789 ( .A0(n4616), .A1(n3427), .B0(n4061), .Y(n4062) );
  AOI22X1TS U4790 ( .A0(n2950), .A1(n4342), .B0(\dataoutbuffer[6][23] ), .B1(
        n4612), .Y(n4067) );
  OAI22X1TS U4791 ( .A0(n4072), .A1(n5217), .B0(n4071), .B1(n2954), .Y(n4065)
         );
  AOI21X1TS U4792 ( .A0(n4615), .A1(n2957), .B0(n4065), .Y(n4066) );
  AOI22X1TS U4793 ( .A0(n3354), .A1(n4342), .B0(\dataoutbuffer[6][14] ), .B1(
        n4612), .Y(n4070) );
  OAI22X1TS U4794 ( .A0(n4072), .A1(n5124), .B0(n4071), .B1(n5123), .Y(n4068)
         );
  AOI21X1TS U4795 ( .A0(n4615), .A1(n3355), .B0(n4068), .Y(n4069) );
  AOI22X1TS U4796 ( .A0(n2964), .A1(n4342), .B0(\dataoutbuffer[6][13] ), .B1(
        n4612), .Y(n4075) );
  OAI22X1TS U4797 ( .A0(n4072), .A1(n4117), .B0(n4071), .B1(n2966), .Y(n4073)
         );
  AOI21X1TS U4798 ( .A0(n4615), .A1(n2962), .B0(n4073), .Y(n4074) );
  AOI22X1TS U4799 ( .A0(n3128), .A1(n4361), .B0(\dataoutbuffer[5][29] ), .B1(
        n4641), .Y(n4080) );
  OAI22X1TS U4800 ( .A0(n3130), .A1(n4243), .B0(n4171), .B1(n4157), .Y(n4078)
         );
  AOI21X1TS U4801 ( .A0(n3126), .A1(n4645), .B0(n4078), .Y(n4079) );
  AOI22X1TS U4802 ( .A0(n3010), .A1(n4361), .B0(\dataoutbuffer[5][1] ), .B1(
        n4641), .Y(n4083) );
  OAI22X1TS U4803 ( .A0(n3009), .A1(n4243), .B0(n4990), .B1(n4157), .Y(n4081)
         );
  AOI21X1TS U4804 ( .A0(n3011), .A1(n4645), .B0(n4081), .Y(n4082) );
  AOI22X1TS U4805 ( .A0(n3428), .A1(n4361), .B0(\dataoutbuffer[5][26] ), .B1(
        n4641), .Y(n4088) );
  OAI22X1TS U4806 ( .A0(n3430), .A1(n4243), .B0(n4085), .B1(n4157), .Y(n4086)
         );
  AOI21X1TS U4807 ( .A0(n3431), .A1(n4645), .B0(n4086), .Y(n4087) );
  AOI22X1TS U4808 ( .A0(n3061), .A1(n4361), .B0(\dataoutbuffer[5][9] ), .B1(
        n4128), .Y(n4092) );
  OAI22X1TS U4809 ( .A0(n5075), .A1(n4243), .B0(n5074), .B1(n4157), .Y(n4090)
         );
  AOI21X1TS U4810 ( .A0(n3062), .A1(n4645), .B0(n4090), .Y(n4091) );
  AOI22X1TS U4811 ( .A0(n3457), .A1(n4361), .B0(\dataoutbuffer[5][30] ), .B1(
        n4641), .Y(n4095) );
  OAI22X1TS U4812 ( .A0(n5293), .A1(n4157), .B0(n5292), .B1(n4243), .Y(n4093)
         );
  AOI21X1TS U4813 ( .A0(n3459), .A1(n4645), .B0(n4093), .Y(n4094) );
  AOI22X1TS U4814 ( .A0(n3481), .A1(n4361), .B0(\dataoutbuffer[5][22] ), .B1(
        n4128), .Y(n4098) );
  OAI22X1TS U4815 ( .A0(n5207), .A1(n4243), .B0(n4227), .B1(n4157), .Y(n4096)
         );
  AOI21X1TS U4816 ( .A0(n3483), .A1(n4645), .B0(n4096), .Y(n4097) );
  AOI22X1TS U4817 ( .A0(n3052), .A1(n4361), .B0(\dataoutbuffer[5][8] ), .B1(
        n4128), .Y(n4101) );
  OAI22X1TS U4818 ( .A0(n3056), .A1(n4243), .B0(n4166), .B1(n4157), .Y(n4099)
         );
  AOI21X1TS U4819 ( .A0(n3053), .A1(n4645), .B0(n4099), .Y(n4100) );
  AOI22X1TS U4820 ( .A0(n3363), .A1(n4361), .B0(\dataoutbuffer[5][11] ), .B1(
        n4128), .Y(n4105) );
  OAI22X1TS U4821 ( .A0(n4102), .A1(n4140), .B0(n3365), .B1(n4243), .Y(n4103)
         );
  AOI21X1TS U4822 ( .A0(n3367), .A1(n4645), .B0(n4103), .Y(n4104) );
  AOI22X1TS U4823 ( .A0(n3342), .A1(n4361), .B0(\dataoutbuffer[5][15] ), .B1(
        n4128), .Y(n4109) );
  OAI22X1TS U4824 ( .A0(n4211), .A1(n4140), .B0(n5134), .B1(n4243), .Y(n4107)
         );
  AOI21X1TS U4825 ( .A0(n3345), .A1(n4645), .B0(n4107), .Y(n4108) );
  AOI22X1TS U4826 ( .A0(n3278), .A1(n4361), .B0(\dataoutbuffer[5][12] ), .B1(
        n4128), .Y(n4112) );
  OAI22X1TS U4827 ( .A0(n3280), .A1(n4140), .B0(n4161), .B1(n4243), .Y(n4110)
         );
  AOI21X1TS U4828 ( .A0(n3281), .A1(n4645), .B0(n4110), .Y(n4111) );
  AOI22X1TS U4829 ( .A0(n2964), .A1(n4361), .B0(\dataoutbuffer[5][13] ), .B1(
        n4128), .Y(n4116) );
  OAI22X1TS U4830 ( .A0(n2963), .A1(n4243), .B0(n4113), .B1(n4140), .Y(n4114)
         );
  AOI21X1TS U4831 ( .A0(n2965), .A1(n4645), .B0(n4114), .Y(n4115) );
  AOI22X1TS U4832 ( .A0(n3019), .A1(n4361), .B0(\dataoutbuffer[5][0] ), .B1(
        n4641), .Y(n4121) );
  OAI22X1TS U4833 ( .A0(n3018), .A1(n4243), .B0(n4118), .B1(n4140), .Y(n4119)
         );
  AOI21X1TS U4834 ( .A0(n3020), .A1(n4645), .B0(n4119), .Y(n4120) );
  AOI22X1TS U4835 ( .A0(n2950), .A1(n4361), .B0(\dataoutbuffer[5][23] ), .B1(
        n4128), .Y(n4124) );
  OAI22X1TS U4836 ( .A0(n4215), .A1(n4140), .B0(n2958), .B1(n4243), .Y(n4122)
         );
  AOI21X1TS U4837 ( .A0(n2953), .A1(n4645), .B0(n4122), .Y(n4123) );
  AOI22X1TS U4838 ( .A0(n3146), .A1(n4361), .B0(\dataoutbuffer[5][24] ), .B1(
        n4128), .Y(n4127) );
  OAI22X1TS U4839 ( .A0(n4179), .A1(n4140), .B0(n3150), .B1(n4243), .Y(n4125)
         );
  AOI21X1TS U4840 ( .A0(n3145), .A1(n4645), .B0(n4125), .Y(n4126) );
  AOI22X1TS U4841 ( .A0(n3230), .A1(n4361), .B0(\dataoutbuffer[5][25] ), .B1(
        n4128), .Y(n4131) );
  OAI22X1TS U4842 ( .A0(n3236), .A1(n4243), .B0(n4183), .B1(n4140), .Y(n4129)
         );
  AOI21X1TS U4843 ( .A0(n3234), .A1(n4645), .B0(n4129), .Y(n4130) );
  AOI22X1TS U4844 ( .A0(n3490), .A1(n4361), .B0(\dataoutbuffer[5][2] ), .B1(
        n4641), .Y(n4135) );
  OAI22X1TS U4845 ( .A0(n3492), .A1(n4243), .B0(n4132), .B1(n4140), .Y(n4133)
         );
  AOI21X1TS U4846 ( .A0(n3493), .A1(n4645), .B0(n4133), .Y(n4134) );
  AOI22X1TS U4847 ( .A0(n3164), .A1(n4361), .B0(\dataoutbuffer[5][4] ), .B1(
        n4641), .Y(n4139) );
  OAI22X1TS U4848 ( .A0(n3166), .A1(n4243), .B0(n4136), .B1(n4140), .Y(n4137)
         );
  AOI21X1TS U4849 ( .A0(n3163), .A1(n4645), .B0(n4137), .Y(n4138) );
  AOI22X1TS U4850 ( .A0(n3527), .A1(n4361), .B0(\dataoutbuffer[5][5] ), .B1(
        n4641), .Y(n4144) );
  OAI22X1TS U4851 ( .A0(n4141), .A1(n4140), .B0(n3529), .B1(n4243), .Y(n4142)
         );
  AOI21X1TS U4852 ( .A0(n3530), .A1(n4645), .B0(n4142), .Y(n4143) );
  AOI22X1TS U4853 ( .A0(n3031), .A1(n4642), .B0(
        \destinationAddressbuffer[5][10] ), .B1(n4641), .Y(n4146) );
  AOI22X1TS U4854 ( .A0(n3030), .A1(n4645), .B0(n3028), .B1(n4643), .Y(n4145)
         );
  AOI22X1TS U4855 ( .A0(n2972), .A1(n4643), .B0(
        \destinationAddressbuffer[5][7] ), .B1(n4641), .Y(n4148) );
  AOI22X1TS U4856 ( .A0(n2975), .A1(n4645), .B0(n2976), .B1(n4642), .Y(n4147)
         );
  AOI22X1TS U4857 ( .A0(n3039), .A1(n4642), .B0(
        \destinationAddressbuffer[5][12] ), .B1(n4641), .Y(n4150) );
  AOI22X1TS U4858 ( .A0(n3038), .A1(n4645), .B0(n3035), .B1(n4643), .Y(n4149)
         );
  AOI22X1TS U4859 ( .A0(n2983), .A1(n4642), .B0(writeOutbuffer[5]), .B1(n4641), 
        .Y(n4152) );
  AOI22X1TS U4860 ( .A0(n2982), .A1(n4645), .B0(n2980), .B1(n4644), .Y(n4151)
         );
  AOI22X1TS U4861 ( .A0(n3073), .A1(n4642), .B0(
        \destinationAddressbuffer[5][11] ), .B1(n4641), .Y(n4154) );
  AOI22X1TS U4862 ( .A0(n3077), .A1(n4645), .B0(n3078), .B1(n4644), .Y(n4153)
         );
  AOI22X1TS U4863 ( .A0(n2990), .A1(n4642), .B0(
        \destinationAddressbuffer[5][8] ), .B1(n4641), .Y(n4156) );
  AOI22X1TS U4864 ( .A0(n2989), .A1(n4645), .B0(n2988), .B1(n4644), .Y(n4155)
         );
  AOI22X1TS U4865 ( .A0(n3155), .A1(n4436), .B0(\dataoutbuffer[1][10] ), .B1(
        n4744), .Y(n4160) );
  OAI22X1TS U4866 ( .A0(n5086), .A1(n4228), .B0(n5085), .B1(n4240), .Y(n4158)
         );
  AOI21X1TS U4867 ( .A0(n3154), .A1(n4761), .B0(n4158), .Y(n4159) );
  AOI22X1TS U4868 ( .A0(n3278), .A1(n4436), .B0(\dataoutbuffer[1][12] ), .B1(
        n4744), .Y(n4165) );
  OAI22X1TS U4869 ( .A0(n4162), .A1(n4240), .B0(n4161), .B1(n4228), .Y(n4163)
         );
  AOI21X1TS U4870 ( .A0(n3281), .A1(n4761), .B0(n4163), .Y(n4164) );
  AOI22X1TS U4871 ( .A0(n3052), .A1(n4436), .B0(\dataoutbuffer[1][8] ), .B1(
        n4744), .Y(n4169) );
  OAI22X1TS U4872 ( .A0(n3056), .A1(n4228), .B0(n4166), .B1(n4240), .Y(n4167)
         );
  AOI21X1TS U4873 ( .A0(n3053), .A1(n4761), .B0(n4167), .Y(n4168) );
  AOI22X1TS U4874 ( .A0(n3128), .A1(n4436), .B0(\dataoutbuffer[1][29] ), .B1(
        n4757), .Y(n4174) );
  OAI22X1TS U4875 ( .A0(n3130), .A1(n4228), .B0(n4171), .B1(n4240), .Y(n4172)
         );
  AOI21X1TS U4876 ( .A0(n3126), .A1(n4761), .B0(n4172), .Y(n4173) );
  AOI22X1TS U4877 ( .A0(n3146), .A1(n4436), .B0(\dataoutbuffer[1][24] ), .B1(
        n4757), .Y(n4178) );
  OAI22X1TS U4878 ( .A0(n5227), .A1(n4240), .B0(n3150), .B1(n4228), .Y(n4176)
         );
  AOI21X1TS U4879 ( .A0(n3145), .A1(n4761), .B0(n4176), .Y(n4177) );
  AOI22X1TS U4880 ( .A0(n3230), .A1(n4436), .B0(\dataoutbuffer[1][25] ), .B1(
        n4757), .Y(n4182) );
  OAI22X1TS U4881 ( .A0(n5239), .A1(n4240), .B0(n3236), .B1(n4228), .Y(n4180)
         );
  AOI21X1TS U4882 ( .A0(n3234), .A1(n4761), .B0(n4180), .Y(n4181) );
  AOI22X1TS U4883 ( .A0(n3061), .A1(n4436), .B0(\dataoutbuffer[1][9] ), .B1(
        n4744), .Y(n4186) );
  OAI22X1TS U4884 ( .A0(n5075), .A1(n4228), .B0(n5074), .B1(n4240), .Y(n4184)
         );
  AOI21X1TS U4885 ( .A0(n3062), .A1(n4761), .B0(n4184), .Y(n4185) );
  AOI22X1TS U4886 ( .A0(n3039), .A1(n4760), .B0(
        \destinationAddressbuffer[1][12] ), .B1(n4757), .Y(n4188) );
  AOI22X1TS U4887 ( .A0(n3038), .A1(n4761), .B0(n3035), .B1(n4758), .Y(n4187)
         );
  AOI22X1TS U4888 ( .A0(n2976), .A1(n4760), .B0(
        \destinationAddressbuffer[1][7] ), .B1(n4744), .Y(n4191) );
  AOI22X1TS U4889 ( .A0(n2975), .A1(n4761), .B0(n2972), .B1(n4758), .Y(n4190)
         );
  AOI22X1TS U4890 ( .A0(n3031), .A1(n4760), .B0(
        \destinationAddressbuffer[1][10] ), .B1(n4757), .Y(n4194) );
  AOI22X1TS U4891 ( .A0(n3030), .A1(n4761), .B0(n3028), .B1(n4758), .Y(n4193)
         );
  AOI22X1TS U4892 ( .A0(n3002), .A1(n4758), .B0(
        \destinationAddressbuffer[1][6] ), .B1(n4744), .Y(n4197) );
  AOI22X1TS U4893 ( .A0(n3004), .A1(n4761), .B0(n3005), .B1(n4760), .Y(n4196)
         );
  AOI22X1TS U4894 ( .A0(n3457), .A1(n4436), .B0(\dataoutbuffer[1][30] ), .B1(
        n4757), .Y(n4201) );
  OAI22X1TS U4895 ( .A0(n4198), .A1(n4229), .B0(n5292), .B1(n4228), .Y(n4199)
         );
  AOI21X1TS U4896 ( .A0(n3459), .A1(n4761), .B0(n4199), .Y(n4200) );
  AOI22X1TS U4897 ( .A0(n3407), .A1(n4436), .B0(\dataoutbuffer[1][18] ), .B1(
        n4757), .Y(n4204) );
  OAI22X1TS U4898 ( .A0(n3406), .A1(n4229), .B0(n5166), .B1(n4228), .Y(n4202)
         );
  AOI21X1TS U4899 ( .A0(n3408), .A1(n4761), .B0(n4202), .Y(n4203) );
  AOI22X1TS U4900 ( .A0(n3207), .A1(n4436), .B0(\dataoutbuffer[1][17] ), .B1(
        n4744), .Y(n4210) );
  OAI22X1TS U4901 ( .A0(n4207), .A1(n4228), .B0(n4206), .B1(n4229), .Y(n4208)
         );
  AOI21X1TS U4902 ( .A0(n3206), .A1(n4761), .B0(n4208), .Y(n4209) );
  AOI22X1TS U4903 ( .A0(n3342), .A1(n4436), .B0(\dataoutbuffer[1][15] ), .B1(
        n4744), .Y(n4214) );
  OAI22X1TS U4904 ( .A0(n4211), .A1(n4229), .B0(n5134), .B1(n4228), .Y(n4212)
         );
  AOI21X1TS U4905 ( .A0(n3345), .A1(n4761), .B0(n4212), .Y(n4213) );
  AOI22X1TS U4906 ( .A0(n2950), .A1(n4436), .B0(\dataoutbuffer[1][23] ), .B1(
        n4757), .Y(n4218) );
  OAI22X1TS U4907 ( .A0(n4215), .A1(n4229), .B0(n2958), .B1(n4228), .Y(n4216)
         );
  AOI21X1TS U4908 ( .A0(n2953), .A1(n4761), .B0(n4216), .Y(n4217) );
  AOI22X1TS U4909 ( .A0(n3043), .A1(n4436), .B0(\dataoutbuffer[1][16] ), .B1(
        n4744), .Y(n4222) );
  OAI22X1TS U4910 ( .A0(n4219), .A1(n4229), .B0(n5146), .B1(n4228), .Y(n4220)
         );
  AOI21X1TS U4911 ( .A0(n3044), .A1(n4761), .B0(n4220), .Y(n4221) );
  AOI22X1TS U4912 ( .A0(n3481), .A1(n4436), .B0(\dataoutbuffer[1][22] ), .B1(
        n4757), .Y(n4226) );
  OAI22X1TS U4913 ( .A0(n5207), .A1(n4228), .B0(n4223), .B1(n4229), .Y(n4224)
         );
  AOI21X1TS U4914 ( .A0(n3483), .A1(n4761), .B0(n4224), .Y(n4225) );
  AOI22X1TS U4915 ( .A0(n3244), .A1(n4436), .B0(\dataoutbuffer[1][20] ), .B1(
        n4757), .Y(n4232) );
  OAI22X1TS U4916 ( .A0(n3246), .A1(n4229), .B0(n5187), .B1(n4228), .Y(n4230)
         );
  AOI21X1TS U4917 ( .A0(n3247), .A1(n4761), .B0(n4230), .Y(n4231) );
  AOI22X1TS U4918 ( .A0(n2990), .A1(n4760), .B0(
        \destinationAddressbuffer[1][8] ), .B1(n4744), .Y(n4234) );
  AOI22X1TS U4919 ( .A0(n2989), .A1(n4761), .B0(n2988), .B1(n4759), .Y(n4233)
         );
  AOI22X1TS U4920 ( .A0(n3073), .A1(n4760), .B0(
        \destinationAddressbuffer[1][11] ), .B1(n4757), .Y(n4237) );
  AOI22X1TS U4921 ( .A0(n3077), .A1(n4761), .B0(n3078), .B1(n4759), .Y(n4236)
         );
  AOI22X1TS U4922 ( .A0(n2983), .A1(n4760), .B0(writeOutbuffer[1]), .B1(n4744), 
        .Y(n4239) );
  AOI22X1TS U4923 ( .A0(n2982), .A1(n4761), .B0(n2980), .B1(n4759), .Y(n4238)
         );
  AOI22X1TS U4924 ( .A0(n3005), .A1(n4642), .B0(
        \destinationAddressbuffer[5][6] ), .B1(n4641), .Y(n4242) );
  AOI22X1TS U4925 ( .A0(n3002), .A1(n4643), .B0(n3004), .B1(n4645), .Y(n4241)
         );
  AOI22X1TS U4926 ( .A0(N375), .A1(read_reg[2]), .B0(n5329), .B1(n5326), .Y(
        n4282) );
  NAND2X1TS U4927 ( .A(N373), .B(n5325), .Y(n4246) );
  XNOR2X1TS U4928 ( .A(n4282), .B(n4245), .Y(n4256) );
  INVX2TS U4929 ( .A(n4258), .Y(n4255) );
  OAI21XLTS U4930 ( .A0(N373), .A1(n5325), .B0(n4246), .Y(n4279) );
  ADDHXLTS U4931 ( .A(n4249), .B(n4248), .CO(n4258), .S(n4260) );
  INVX2TS U4932 ( .A(n4260), .Y(n4250) );
  AOI21X1TS U4933 ( .A0(n4280), .A1(n4250), .B0(n4279), .Y(n4252) );
  OAI22X1TS U4934 ( .A0(n4280), .A1(n4250), .B0(n4256), .B1(n4255), .Y(n4251)
         );
  AOI21X1TS U4935 ( .A0(n4259), .A1(n4252), .B0(n4251), .Y(n4253) );
  INVX2TS U4936 ( .A(n4257), .Y(n4261) );
  NAND2X1TS U4937 ( .A(n4261), .B(n4258), .Y(n4264) );
  XNOR2X1TS U4938 ( .A(N375), .B(n4262), .Y(n4263) );
  INVX2TS U4939 ( .A(n4276), .Y(n4271) );
  ADDHXLTS U4940 ( .A(N373), .B(n4265), .CO(n4267), .S(n4274) );
  XNOR2X1TS U4941 ( .A(read_reg[1]), .B(n4275), .Y(n4268) );
  OAI2BB2XLTS U4942 ( .B0(n5328), .B1(n4273), .A0N(n4284), .A1N(n4272), .Y(
        N4718) );
  AOI22X1TS U4943 ( .A0(read_reg[0]), .A1(n4273), .B0(n4278), .B1(n5325), .Y(
        n2889) );
  OAI2BB2XLTS U4944 ( .B0(n5327), .B1(n4277), .A0N(n4284), .A1N(n4274), .Y(
        n2888) );
  OAI2BB2XLTS U4945 ( .B0(n5323), .B1(n4277), .A0N(n4284), .A1N(n4275), .Y(
        n2887) );
  OAI2BB2XLTS U4946 ( .B0(n5326), .B1(n4277), .A0N(n4284), .A1N(n4276), .Y(
        n2886) );
  OAI211XLTS U4947 ( .A0(n4283), .A1(n4282), .B0(n4280), .C0(n4279), .Y(n4281)
         );
  AO21XLTS U4948 ( .A0(n4283), .A1(n4282), .B0(n4281), .Y(n4285) );
  AOI21X1TS U4949 ( .A0(n2890), .A1(n4285), .B0(n4284), .Y(n2885) );
  OAI2BB2XLTS U4950 ( .B0(n4286), .B1(n5329), .A0N(n2891), .A1N(n2890), .Y(
        n2884) );
  AOI22X1TS U4951 ( .A0(n2907), .A1(n4580), .B0(\requesterAddressbuffer[7][0] ), .B1(n4318), .Y(n4289) );
  AOI22X1TS U4952 ( .A0(n2905), .A1(n4586), .B0(n2909), .B1(n4583), .Y(n4288)
         );
  NAND2X1TS U4953 ( .A(n2910), .B(n4584), .Y(n4287) );
  NAND2X1TS U4954 ( .A(n2921), .B(n4323), .Y(n4543) );
  CLKBUFX2TS U4955 ( .A(requesterAddressIn_EAST[1]), .Y(n4290) );
  AOI22X1TS U4956 ( .A0(n4290), .A1(n4583), .B0(\requesterAddressbuffer[7][1] ), .B1(n4318), .Y(n4297) );
  CLKBUFX2TS U4957 ( .A(requesterAddressIn_WEST[1]), .Y(n4291) );
  CLKBUFX2TS U4958 ( .A(requesterAddressIn_NORTH[1]), .Y(n4292) );
  AOI22X1TS U4959 ( .A0(n4291), .A1(n4580), .B0(n4292), .B1(n4584), .Y(n4296)
         );
  CLKBUFX2TS U4960 ( .A(requesterAddressIn_SOUTH[1]), .Y(n4293) );
  NAND2X1TS U4961 ( .A(n4293), .B(n4586), .Y(n4295) );
  CLKBUFX2TS U4962 ( .A(readRequesterAddress[1]), .Y(n4294) );
  NAND2X1TS U4963 ( .A(n4294), .B(n4323), .Y(n4551) );
  CLKBUFX2TS U4964 ( .A(requesterAddressIn_WEST[2]), .Y(n4298) );
  AOI22X1TS U4965 ( .A0(n4298), .A1(n4580), .B0(\requesterAddressbuffer[7][2] ), .B1(n4318), .Y(n4305) );
  CLKBUFX2TS U4966 ( .A(requesterAddressIn_EAST[2]), .Y(n4299) );
  CLKBUFX2TS U4967 ( .A(requesterAddressIn_SOUTH[2]), .Y(n4300) );
  AOI22X1TS U4968 ( .A0(n4299), .A1(n4583), .B0(n4300), .B1(n4586), .Y(n4304)
         );
  CLKBUFX2TS U4969 ( .A(requesterAddressIn_NORTH[2]), .Y(n4301) );
  NAND2X1TS U4970 ( .A(n4301), .B(n4584), .Y(n4303) );
  CLKBUFX2TS U4971 ( .A(readRequesterAddress[2]), .Y(n4302) );
  NAND2X1TS U4972 ( .A(n4302), .B(n4323), .Y(n4559) );
  AOI22X1TS U4973 ( .A0(n2926), .A1(n4580), .B0(\requesterAddressbuffer[7][3] ), .B1(n4318), .Y(n4308) );
  AOI22X1TS U4974 ( .A0(n2924), .A1(n4584), .B0(n2928), .B1(n4583), .Y(n4307)
         );
  NAND2X1TS U4975 ( .A(n2927), .B(n4586), .Y(n4306) );
  NAND2X1TS U4976 ( .A(n2936), .B(n4323), .Y(n4567) );
  CLKBUFX2TS U4977 ( .A(requesterAddressIn_WEST[4]), .Y(n4309) );
  AOI22X1TS U4978 ( .A0(n4309), .A1(n4580), .B0(\requesterAddressbuffer[7][4] ), .B1(n4318), .Y(n4316) );
  CLKBUFX2TS U4979 ( .A(requesterAddressIn_EAST[4]), .Y(n4310) );
  CLKBUFX2TS U4980 ( .A(requesterAddressIn_NORTH[4]), .Y(n4311) );
  AOI22X1TS U4981 ( .A0(n4310), .A1(n4583), .B0(n4311), .B1(n4584), .Y(n4315)
         );
  CLKBUFX2TS U4982 ( .A(requesterAddressIn_SOUTH[4]), .Y(n4312) );
  NAND2X1TS U4983 ( .A(n4312), .B(n4586), .Y(n4314) );
  CLKBUFX2TS U4984 ( .A(readRequesterAddress[4]), .Y(n4313) );
  NAND2X1TS U4985 ( .A(n4313), .B(n4323), .Y(n4575) );
  CLKBUFX2TS U4986 ( .A(requesterAddressIn_WEST[5]), .Y(n4317) );
  AOI22X1TS U4987 ( .A0(n4317), .A1(n4580), .B0(\requesterAddressbuffer[7][5] ), .B1(n4318), .Y(n4326) );
  CLKBUFX2TS U4988 ( .A(requesterAddressIn_EAST[5]), .Y(n4319) );
  CLKBUFX2TS U4989 ( .A(requesterAddressIn_NORTH[5]), .Y(n4320) );
  AOI22X1TS U4990 ( .A0(n4319), .A1(n4583), .B0(n4320), .B1(n4584), .Y(n4325)
         );
  CLKBUFX2TS U4991 ( .A(requesterAddressIn_SOUTH[5]), .Y(n4321) );
  NAND2X1TS U4992 ( .A(n4321), .B(n4586), .Y(n4324) );
  CLKBUFX2TS U4993 ( .A(readRequesterAddress[5]), .Y(n4322) );
  NAND2X1TS U4994 ( .A(n4322), .B(n4323), .Y(n4588) );
  AOI22X1TS U4995 ( .A0(n4614), .A1(n2910), .B0(\requesterAddressbuffer[6][0] ), .B1(n4612), .Y(n4329) );
  AOI22X1TS U4996 ( .A0(n2907), .A1(n4616), .B0(n2909), .B1(n4613), .Y(n4328)
         );
  NAND2X1TS U4997 ( .A(n2905), .B(n4607), .Y(n4327) );
  NAND2X1TS U4998 ( .A(n2921), .B(n4342), .Y(n4592) );
  AOI22X1TS U4999 ( .A0(n4293), .A1(n4607), .B0(\requesterAddressbuffer[6][1] ), .B1(n4612), .Y(n4332) );
  AOI22X1TS U5000 ( .A0(n4616), .A1(n4291), .B0(n4614), .B1(n4292), .Y(n4331)
         );
  NAND2X1TS U5001 ( .A(n4613), .B(n4290), .Y(n4330) );
  NAND2X1TS U5002 ( .A(n4342), .B(n4294), .Y(n4596) );
  AOI22X1TS U5003 ( .A0(n4300), .A1(n4607), .B0(\requesterAddressbuffer[6][2] ), .B1(n4612), .Y(n4335) );
  AOI22X1TS U5004 ( .A0(n4616), .A1(n4298), .B0(n4614), .B1(n4301), .Y(n4334)
         );
  NAND2X1TS U5005 ( .A(n4613), .B(n4299), .Y(n4333) );
  NAND2X1TS U5006 ( .A(n4342), .B(n4302), .Y(n4600) );
  AOI22X1TS U5007 ( .A0(n2928), .A1(n4613), .B0(\requesterAddressbuffer[6][3] ), .B1(n4612), .Y(n4338) );
  AOI22X1TS U5008 ( .A0(n4615), .A1(n2927), .B0(n4616), .B1(n2926), .Y(n4337)
         );
  NAND2X1TS U5009 ( .A(n4614), .B(n2924), .Y(n4336) );
  NAND2X1TS U5010 ( .A(n4342), .B(n2936), .Y(n4604) );
  AOI22X1TS U5011 ( .A0(n4311), .A1(n4614), .B0(\requesterAddressbuffer[6][4] ), .B1(n4612), .Y(n4341) );
  AOI22X1TS U5012 ( .A0(n4607), .A1(n4312), .B0(n4616), .B1(n4309), .Y(n4340)
         );
  NAND2X1TS U5013 ( .A(n4613), .B(n4310), .Y(n4339) );
  NAND2X1TS U5014 ( .A(n4342), .B(n4313), .Y(n4609) );
  AOI22X1TS U5015 ( .A0(n4320), .A1(n4614), .B0(\requesterAddressbuffer[6][5] ), .B1(n4612), .Y(n4345) );
  AOI22X1TS U5016 ( .A0(n4616), .A1(n4317), .B0(n4613), .B1(n4319), .Y(n4344)
         );
  NAND2X1TS U5017 ( .A(n4615), .B(n4321), .Y(n4343) );
  NAND2X1TS U5018 ( .A(n4342), .B(n4322), .Y(n4618) );
  AOI22X1TS U5019 ( .A0(n2907), .A1(n4642), .B0(\requesterAddressbuffer[5][0] ), .B1(n4641), .Y(n4348) );
  AOI22X1TS U5020 ( .A0(n2909), .A1(n4643), .B0(n2910), .B1(n4645), .Y(n4347)
         );
  NAND2X1TS U5021 ( .A(n2905), .B(n4644), .Y(n4346) );
  NAND2X1TS U5022 ( .A(n2921), .B(n4361), .Y(n4622) );
  AOI22X1TS U5023 ( .A0(n4291), .A1(n4642), .B0(\requesterAddressbuffer[5][1] ), .B1(n4641), .Y(n4351) );
  AOI22X1TS U5024 ( .A0(n4290), .A1(n4643), .B0(n4292), .B1(n4645), .Y(n4350)
         );
  NAND2X1TS U5025 ( .A(n4293), .B(n4644), .Y(n4349) );
  NAND2X1TS U5026 ( .A(n4294), .B(n4361), .Y(n4626) );
  AOI22X1TS U5027 ( .A0(n4298), .A1(n4642), .B0(\requesterAddressbuffer[5][2] ), .B1(n4641), .Y(n4354) );
  AOI22X1TS U5028 ( .A0(n4299), .A1(n4643), .B0(n4301), .B1(n4645), .Y(n4353)
         );
  NAND2X1TS U5029 ( .A(n4300), .B(n4644), .Y(n4352) );
  NAND2X1TS U5030 ( .A(n4302), .B(n4361), .Y(n4630) );
  AOI22X1TS U5031 ( .A0(n2928), .A1(n4643), .B0(\requesterAddressbuffer[5][3] ), .B1(n4641), .Y(n4357) );
  AOI22X1TS U5032 ( .A0(n2924), .A1(n4645), .B0(n2926), .B1(n4642), .Y(n4356)
         );
  NAND2X1TS U5033 ( .A(n2927), .B(n4644), .Y(n4355) );
  NAND2X1TS U5034 ( .A(n2936), .B(n4361), .Y(n4634) );
  AOI22X1TS U5035 ( .A0(n4310), .A1(n4643), .B0(\requesterAddressbuffer[5][4] ), .B1(n4641), .Y(n4360) );
  AOI22X1TS U5036 ( .A0(n4309), .A1(n4642), .B0(n4311), .B1(n4645), .Y(n4359)
         );
  NAND2X1TS U5037 ( .A(n4312), .B(n4644), .Y(n4358) );
  NAND2X1TS U5038 ( .A(n4313), .B(n4361), .Y(n4638) );
  AOI22X1TS U5039 ( .A0(n4319), .A1(n4643), .B0(\requesterAddressbuffer[5][5] ), .B1(n4641), .Y(n4364) );
  AOI22X1TS U5040 ( .A0(n4321), .A1(n4644), .B0(n4317), .B1(n4642), .Y(n4363)
         );
  NAND2X1TS U5041 ( .A(n4320), .B(n4645), .Y(n4362) );
  NAND2X1TS U5042 ( .A(n4322), .B(n4361), .Y(n4647) );
  AOI22X1TS U5043 ( .A0(n2905), .A1(n4673), .B0(\requesterAddressbuffer[4][0] ), .B1(n4671), .Y(n4367) );
  AOI22X1TS U5044 ( .A0(n2907), .A1(n4666), .B0(n2910), .B1(n4674), .Y(n4366)
         );
  NAND2X1TS U5045 ( .A(n2909), .B(n4672), .Y(n4365) );
  NAND2X1TS U5046 ( .A(n2921), .B(n4380), .Y(n4651) );
  AOI22X1TS U5047 ( .A0(n4290), .A1(n4672), .B0(\requesterAddressbuffer[4][1] ), .B1(n4671), .Y(n4370) );
  AOI22X1TS U5048 ( .A0(n4291), .A1(n4666), .B0(n4293), .B1(n4673), .Y(n4369)
         );
  NAND2X1TS U5049 ( .A(n4292), .B(n4674), .Y(n4368) );
  NAND2X1TS U5050 ( .A(n4294), .B(n4380), .Y(n4655) );
  AOI22X1TS U5051 ( .A0(n4300), .A1(n4673), .B0(\requesterAddressbuffer[4][2] ), .B1(n4671), .Y(n4373) );
  AOI22X1TS U5052 ( .A0(n4298), .A1(n4666), .B0(n4301), .B1(n4674), .Y(n4372)
         );
  NAND2X1TS U5053 ( .A(n4299), .B(n4672), .Y(n4371) );
  NAND2X1TS U5054 ( .A(n4302), .B(n4380), .Y(n4659) );
  AOI22X1TS U5055 ( .A0(n2924), .A1(n4674), .B0(\requesterAddressbuffer[4][3] ), .B1(n4671), .Y(n4376) );
  AOI22X1TS U5056 ( .A0(n2927), .A1(n4673), .B0(n2928), .B1(n4672), .Y(n4375)
         );
  NAND2X1TS U5057 ( .A(n2926), .B(n4666), .Y(n4374) );
  NAND2X1TS U5058 ( .A(n2936), .B(n4380), .Y(n4663) );
  AOI22X1TS U5059 ( .A0(n4310), .A1(n4672), .B0(\requesterAddressbuffer[4][4] ), .B1(n4671), .Y(n4379) );
  AOI22X1TS U5060 ( .A0(n4312), .A1(n4673), .B0(n4309), .B1(n4666), .Y(n4378)
         );
  NAND2X1TS U5061 ( .A(n4311), .B(n4674), .Y(n4377) );
  NAND2X1TS U5062 ( .A(n4313), .B(n4380), .Y(n4668) );
  AOI22X1TS U5063 ( .A0(n4319), .A1(n4672), .B0(\requesterAddressbuffer[4][5] ), .B1(n4671), .Y(n4383) );
  AOI22X1TS U5064 ( .A0(n4317), .A1(n4666), .B0(n4320), .B1(n4674), .Y(n4382)
         );
  NAND2X1TS U5065 ( .A(n4321), .B(n4673), .Y(n4381) );
  NAND2X1TS U5066 ( .A(n4322), .B(n4380), .Y(n4676) );
  AOI22X1TS U5067 ( .A0(n2907), .A1(n4687), .B0(\requesterAddressbuffer[3][0] ), .B1(n4701), .Y(n4386) );
  AOI22X1TS U5068 ( .A0(n2905), .A1(n4702), .B0(n2909), .B1(n4696), .Y(n4385)
         );
  NAND2X1TS U5069 ( .A(n2910), .B(n4703), .Y(n4384) );
  NAND2X1TS U5070 ( .A(n2921), .B(n3232), .Y(n4680) );
  AOI22X1TS U5071 ( .A0(n4290), .A1(n4696), .B0(\requesterAddressbuffer[3][1] ), .B1(n4701), .Y(n4389) );
  AOI22X1TS U5072 ( .A0(n4291), .A1(n4687), .B0(n4292), .B1(n4703), .Y(n4388)
         );
  NAND2X1TS U5073 ( .A(n4293), .B(n4702), .Y(n4387) );
  NAND2X1TS U5074 ( .A(n4294), .B(n3232), .Y(n4684) );
  AOI22X1TS U5075 ( .A0(n4298), .A1(n4687), .B0(\requesterAddressbuffer[3][2] ), .B1(n4701), .Y(n4392) );
  AOI22X1TS U5076 ( .A0(n4299), .A1(n4696), .B0(n4300), .B1(n4702), .Y(n4391)
         );
  NAND2X1TS U5077 ( .A(n4301), .B(n4703), .Y(n4390) );
  NAND2X1TS U5078 ( .A(n4302), .B(n3232), .Y(n4689) );
  AOI22X1TS U5079 ( .A0(n2928), .A1(n4696), .B0(\requesterAddressbuffer[3][3] ), .B1(n4701), .Y(n4395) );
  AOI22X1TS U5080 ( .A0(n2924), .A1(n4703), .B0(n2926), .B1(n4687), .Y(n4394)
         );
  NAND2X1TS U5081 ( .A(n2927), .B(n4702), .Y(n4393) );
  NAND2X1TS U5082 ( .A(n2936), .B(n3232), .Y(n4693) );
  AOI22X1TS U5083 ( .A0(n4309), .A1(n4687), .B0(\requesterAddressbuffer[3][4] ), .B1(n4701), .Y(n4398) );
  AOI22X1TS U5084 ( .A0(n4310), .A1(n4696), .B0(n4311), .B1(n4703), .Y(n4397)
         );
  NAND2X1TS U5085 ( .A(n4312), .B(n4702), .Y(n4396) );
  NAND2X1TS U5086 ( .A(n4313), .B(n3232), .Y(n4698) );
  AOI22X1TS U5087 ( .A0(n4319), .A1(n4696), .B0(\requesterAddressbuffer[3][5] ), .B1(n4701), .Y(n4401) );
  AOI22X1TS U5088 ( .A0(n4317), .A1(n4687), .B0(n4320), .B1(n4703), .Y(n4400)
         );
  NAND2X1TS U5089 ( .A(n4321), .B(n4702), .Y(n4399) );
  NAND2X1TS U5090 ( .A(n4322), .B(n3232), .Y(n4705) );
  AOI22X1TS U5091 ( .A0(n2905), .A1(n4730), .B0(\requesterAddressbuffer[2][0] ), .B1(n4728), .Y(n4404) );
  AOI22X1TS U5092 ( .A0(n2907), .A1(n4731), .B0(n2909), .B1(n4729), .Y(n4403)
         );
  NAND2X1TS U5093 ( .A(n2910), .B(n2952), .Y(n4402) );
  NAND2X1TS U5094 ( .A(n2921), .B(n4417), .Y(n4709) );
  AOI22X1TS U5095 ( .A0(n4293), .A1(n4730), .B0(\requesterAddressbuffer[2][1] ), .B1(n4728), .Y(n4407) );
  AOI22X1TS U5096 ( .A0(n4291), .A1(n4731), .B0(n4292), .B1(n2952), .Y(n4406)
         );
  NAND2X1TS U5097 ( .A(n4290), .B(n4729), .Y(n4405) );
  NAND2X1TS U5098 ( .A(n4294), .B(n4417), .Y(n4713) );
  AOI22X1TS U5099 ( .A0(n4298), .A1(n4731), .B0(\requesterAddressbuffer[2][2] ), .B1(n4728), .Y(n4410) );
  AOI22X1TS U5100 ( .A0(n4301), .A1(n2952), .B0(n4300), .B1(n4730), .Y(n4409)
         );
  NAND2X1TS U5101 ( .A(n4299), .B(n4729), .Y(n4408) );
  NAND2X1TS U5102 ( .A(n4302), .B(n4417), .Y(n4717) );
  AOI22X1TS U5103 ( .A0(n2924), .A1(n2952), .B0(\requesterAddressbuffer[2][3] ), .B1(n4728), .Y(n4413) );
  AOI22X1TS U5104 ( .A0(n2927), .A1(n4730), .B0(n2928), .B1(n4729), .Y(n4412)
         );
  NAND2X1TS U5105 ( .A(n2926), .B(n4731), .Y(n4411) );
  NAND2X1TS U5106 ( .A(n2936), .B(n4417), .Y(n4721) );
  AOI22X1TS U5107 ( .A0(n4309), .A1(n4731), .B0(\requesterAddressbuffer[2][4] ), .B1(n4728), .Y(n4416) );
  AOI22X1TS U5108 ( .A0(n4310), .A1(n4729), .B0(n4312), .B1(n4730), .Y(n4415)
         );
  NAND2X1TS U5109 ( .A(n4311), .B(n2952), .Y(n4414) );
  NAND2X1TS U5110 ( .A(n4313), .B(n4417), .Y(n4725) );
  AOI22X1TS U5111 ( .A0(n4317), .A1(n4731), .B0(\requesterAddressbuffer[2][5] ), .B1(n4728), .Y(n4420) );
  AOI22X1TS U5112 ( .A0(n4321), .A1(n4730), .B0(n4319), .B1(n4729), .Y(n4419)
         );
  NAND2X1TS U5113 ( .A(n4320), .B(n2952), .Y(n4418) );
  NAND2X1TS U5114 ( .A(n4322), .B(n4417), .Y(n4733) );
  AOI22X1TS U5115 ( .A0(n2909), .A1(n4758), .B0(\requesterAddressbuffer[1][0] ), .B1(n4757), .Y(n4423) );
  AOI22X1TS U5116 ( .A0(n2905), .A1(n4759), .B0(n2907), .B1(n4760), .Y(n4422)
         );
  NAND2X1TS U5117 ( .A(n2910), .B(n4761), .Y(n4421) );
  NAND2X1TS U5118 ( .A(n2921), .B(n4436), .Y(n4737) );
  AOI22X1TS U5119 ( .A0(n4291), .A1(n4760), .B0(\requesterAddressbuffer[1][1] ), .B1(n4757), .Y(n4426) );
  AOI22X1TS U5120 ( .A0(n4290), .A1(n4758), .B0(n4292), .B1(n4761), .Y(n4425)
         );
  NAND2X1TS U5121 ( .A(n4293), .B(n4759), .Y(n4424) );
  NAND2X1TS U5122 ( .A(n4294), .B(n4436), .Y(n4741) );
  AOI22X1TS U5123 ( .A0(n4298), .A1(n4760), .B0(\requesterAddressbuffer[1][2] ), .B1(n4757), .Y(n4429) );
  AOI22X1TS U5124 ( .A0(n4299), .A1(n4758), .B0(n4300), .B1(n4759), .Y(n4428)
         );
  NAND2X1TS U5125 ( .A(n4301), .B(n4761), .Y(n4427) );
  NAND2X1TS U5126 ( .A(n4302), .B(n4436), .Y(n4746) );
  AOI22X1TS U5127 ( .A0(n2928), .A1(n4758), .B0(\requesterAddressbuffer[1][3] ), .B1(n4757), .Y(n4432) );
  AOI22X1TS U5128 ( .A0(n2926), .A1(n4760), .B0(n2927), .B1(n4759), .Y(n4431)
         );
  NAND2X1TS U5129 ( .A(n2924), .B(n4761), .Y(n4430) );
  NAND2X1TS U5130 ( .A(n2936), .B(n4436), .Y(n4750) );
  AOI22X1TS U5131 ( .A0(n4309), .A1(n4760), .B0(\requesterAddressbuffer[1][4] ), .B1(n4757), .Y(n4435) );
  AOI22X1TS U5132 ( .A0(n4310), .A1(n4758), .B0(n4312), .B1(n4759), .Y(n4434)
         );
  NAND2X1TS U5133 ( .A(n4311), .B(n4761), .Y(n4433) );
  NAND2X1TS U5134 ( .A(n4313), .B(n4436), .Y(n4754) );
  AOI22X1TS U5135 ( .A0(n4317), .A1(n4760), .B0(\requesterAddressbuffer[1][5] ), .B1(n4757), .Y(n4439) );
  AOI22X1TS U5136 ( .A0(n4319), .A1(n4758), .B0(n4320), .B1(n4761), .Y(n4438)
         );
  NAND2X1TS U5137 ( .A(n4321), .B(n4759), .Y(n4437) );
  NAND2X1TS U5138 ( .A(n4322), .B(n4436), .Y(n4763) );
  AOI22X1TS U5139 ( .A0(n2905), .A1(n4789), .B0(\requesterAddressbuffer[0][0] ), .B1(n4787), .Y(n4442) );
  AOI22X1TS U5140 ( .A0(n2909), .A1(n4782), .B0(n2910), .B1(n4790), .Y(n4441)
         );
  NAND2X1TS U5141 ( .A(n2907), .B(n4788), .Y(n4440) );
  NAND2X1TS U5142 ( .A(n2921), .B(n4455), .Y(n4767) );
  AOI22X1TS U5143 ( .A0(n4292), .A1(n4790), .B0(\requesterAddressbuffer[0][1] ), .B1(n4787), .Y(n4445) );
  AOI22X1TS U5144 ( .A0(n4290), .A1(n4782), .B0(n4291), .B1(n4788), .Y(n4444)
         );
  NAND2X1TS U5145 ( .A(n4293), .B(n4789), .Y(n4443) );
  NAND2X1TS U5146 ( .A(n4294), .B(n4455), .Y(n4771) );
  AOI22X1TS U5147 ( .A0(n4299), .A1(n4782), .B0(\requesterAddressbuffer[0][2] ), .B1(n4787), .Y(n4448) );
  AOI22X1TS U5148 ( .A0(n4301), .A1(n4790), .B0(n4300), .B1(n4789), .Y(n4447)
         );
  NAND2X1TS U5149 ( .A(n4298), .B(n4788), .Y(n4446) );
  NAND2X1TS U5150 ( .A(n4302), .B(n4455), .Y(n4775) );
  AOI22X1TS U5151 ( .A0(n2924), .A1(n4790), .B0(\requesterAddressbuffer[0][3] ), .B1(n4787), .Y(n4451) );
  AOI22X1TS U5152 ( .A0(n2926), .A1(n4788), .B0(n2927), .B1(n4789), .Y(n4450)
         );
  NAND2X1TS U5153 ( .A(n2928), .B(n4782), .Y(n4449) );
  NAND2X1TS U5154 ( .A(n2936), .B(n4455), .Y(n4779) );
  AOI22X1TS U5155 ( .A0(n4312), .A1(n4789), .B0(\requesterAddressbuffer[0][4] ), .B1(n4787), .Y(n4454) );
  AOI22X1TS U5156 ( .A0(n4310), .A1(n4782), .B0(n4311), .B1(n4790), .Y(n4453)
         );
  NAND2X1TS U5157 ( .A(n4309), .B(n4788), .Y(n4452) );
  NAND2X1TS U5158 ( .A(n4313), .B(n4455), .Y(n4784) );
  AOI22X1TS U5159 ( .A0(n4317), .A1(n4788), .B0(\requesterAddressbuffer[0][5] ), .B1(n4787), .Y(n4458) );
  AOI22X1TS U5160 ( .A0(n4319), .A1(n4782), .B0(n4320), .B1(n4790), .Y(n4457)
         );
  NAND2X1TS U5161 ( .A(n4321), .B(n4789), .Y(n4456) );
  NAND2X1TS U5162 ( .A(n4322), .B(n4455), .Y(n4792) );
  CLKBUFX2TS U5163 ( .A(readIn_SOUTH), .Y(n4459) );
  INVX2TS U5164 ( .A(n4459), .Y(n4797) );
  CLKBUFX2TS U5165 ( .A(readIn_NORTH), .Y(n4460) );
  AOI22X1TS U5166 ( .A0(n4463), .A1(n4797), .B0(n4461), .B1(n4462), .Y(n4470)
         );
  CLKBUFX2TS U5167 ( .A(readIn_WEST), .Y(n4464) );
  INVX2TS U5168 ( .A(n4464), .Y(n4799) );
  CLKBUFX2TS U5169 ( .A(readIn_EAST), .Y(n4465) );
  OAI22X1TS U5170 ( .A0(n4467), .A1(n4799), .B0(n4466), .B1(n4796), .Y(n4468)
         );
  AOI211XLTS U5171 ( .A0(n4471), .A1(n4470), .B0(n4469), .C0(n4468), .Y(n4472)
         );
  OAI22X1TS U5172 ( .A0(n4475), .A1(n4799), .B0(n4474), .B1(n4796), .Y(n4476)
         );
  AOI211XLTS U5173 ( .A0(n4478), .A1(n4460), .B0(n4477), .C0(n4476), .Y(n4479)
         );
  OA21XLTS U5174 ( .A0(n4482), .A1(readOutbuffer[6]), .B0(n4481), .Y(n2569) );
  AOI22X1TS U5175 ( .A0(n4484), .A1(n4797), .B0(n4461), .B1(n4483), .Y(n4525)
         );
  OAI22X1TS U5176 ( .A0(n4486), .A1(n4799), .B0(n4485), .B1(n4796), .Y(n4487)
         );
  AOI211XLTS U5177 ( .A0(n4489), .A1(n4525), .B0(n4488), .C0(n4487), .Y(n4490)
         );
  OAI22X1TS U5178 ( .A0(n4493), .A1(n4799), .B0(n4492), .B1(n4796), .Y(n4494)
         );
  AOI211XLTS U5179 ( .A0(n4496), .A1(n4460), .B0(n4495), .C0(n4494), .Y(n4497)
         );
  OA21XLTS U5180 ( .A0(n4500), .A1(readOutbuffer[4]), .B0(n4499), .Y(n2567) );
  AOI22X1TS U5181 ( .A0(n4503), .A1(n4460), .B0(n4459), .B1(n4502), .Y(n4505)
         );
  OAI22X1TS U5182 ( .A0(n4506), .A1(n4505), .B0(n4504), .B1(n4796), .Y(n4507)
         );
  AOI211XLTS U5183 ( .A0(n4509), .A1(n4464), .B0(n4508), .C0(n4507), .Y(n4510)
         );
  NOR3XLTS U5184 ( .A(n4796), .B(n4517), .C(n4512), .Y(n4516) );
  OAI2BB2XLTS U5185 ( .B0(n4514), .B1(n4797), .A0N(n4513), .A1N(n4460), .Y(
        n4515) );
  OAI22X1TS U5186 ( .A0(n4522), .A1(n4799), .B0(n4521), .B1(n4796), .Y(n4523)
         );
  AOI211XLTS U5187 ( .A0(n4526), .A1(n4525), .B0(n4524), .C0(n4523), .Y(n4527)
         );
  OAI22X1TS U5188 ( .A0(n4530), .A1(n4799), .B0(n4529), .B1(n4796), .Y(n4534)
         );
  OAI22X1TS U5189 ( .A0(n4532), .A1(n4461), .B0(n4531), .B1(n4797), .Y(n4533)
         );
  NOR3XLTS U5190 ( .A(n4535), .B(n4534), .C(n4533), .Y(n4536) );
  CLKBUFX2TS U5191 ( .A(destinationAddressIn_EAST[0]), .Y(n4538) );
  AOI22X1TS U5192 ( .A0(n4538), .A1(n4583), .B0(
        \destinationAddressbuffer[7][0] ), .B1(n4579), .Y(n4545) );
  CLKBUFX2TS U5193 ( .A(destinationAddressIn_SOUTH[0]), .Y(n4539) );
  CLKBUFX2TS U5194 ( .A(destinationAddressIn_WEST[0]), .Y(n4540) );
  AOI22X1TS U5195 ( .A0(n4539), .A1(n4586), .B0(n4540), .B1(n4580), .Y(n4544)
         );
  CLKBUFX2TS U5196 ( .A(destinationAddressIn_NORTH[0]), .Y(n4541) );
  NAND2X1TS U5197 ( .A(n4541), .B(n4584), .Y(n4542) );
  CLKBUFX2TS U5198 ( .A(destinationAddressIn_WEST[1]), .Y(n4546) );
  AOI22X1TS U5199 ( .A0(n4546), .A1(n4580), .B0(
        \destinationAddressbuffer[7][1] ), .B1(n4579), .Y(n4553) );
  CLKBUFX2TS U5200 ( .A(destinationAddressIn_EAST[1]), .Y(n4547) );
  CLKBUFX2TS U5201 ( .A(destinationAddressIn_NORTH[1]), .Y(n4548) );
  AOI22X1TS U5202 ( .A0(n4547), .A1(n4583), .B0(n4548), .B1(n4584), .Y(n4552)
         );
  CLKBUFX2TS U5203 ( .A(destinationAddressIn_SOUTH[1]), .Y(n4549) );
  NAND2X1TS U5204 ( .A(n4549), .B(n4586), .Y(n4550) );
  CLKBUFX2TS U5205 ( .A(destinationAddressIn_WEST[2]), .Y(n4554) );
  AOI22X1TS U5206 ( .A0(n4554), .A1(n4580), .B0(
        \destinationAddressbuffer[7][2] ), .B1(n4579), .Y(n4561) );
  CLKBUFX2TS U5207 ( .A(destinationAddressIn_EAST[2]), .Y(n4555) );
  CLKBUFX2TS U5208 ( .A(destinationAddressIn_SOUTH[2]), .Y(n4556) );
  AOI22X1TS U5209 ( .A0(n4555), .A1(n4583), .B0(n4556), .B1(n4586), .Y(n4560)
         );
  CLKBUFX2TS U5210 ( .A(destinationAddressIn_NORTH[2]), .Y(n4557) );
  NAND2X1TS U5211 ( .A(n4557), .B(n4584), .Y(n4558) );
  CLKBUFX2TS U5212 ( .A(destinationAddressIn_EAST[3]), .Y(n4562) );
  AOI22X1TS U5213 ( .A0(n4562), .A1(n4583), .B0(
        \destinationAddressbuffer[7][3] ), .B1(n4579), .Y(n4569) );
  CLKBUFX2TS U5214 ( .A(destinationAddressIn_NORTH[3]), .Y(n4563) );
  CLKBUFX2TS U5215 ( .A(destinationAddressIn_WEST[3]), .Y(n4564) );
  AOI22X1TS U5216 ( .A0(n4563), .A1(n4584), .B0(n4564), .B1(n4580), .Y(n4568)
         );
  CLKBUFX2TS U5217 ( .A(destinationAddressIn_SOUTH[3]), .Y(n4565) );
  NAND2X1TS U5218 ( .A(n4565), .B(n4586), .Y(n4566) );
  CLKBUFX2TS U5219 ( .A(destinationAddressIn_WEST[4]), .Y(n4570) );
  AOI22X1TS U5220 ( .A0(n4570), .A1(n4580), .B0(
        \destinationAddressbuffer[7][4] ), .B1(n4579), .Y(n4577) );
  CLKBUFX2TS U5221 ( .A(destinationAddressIn_EAST[4]), .Y(n4571) );
  CLKBUFX2TS U5222 ( .A(destinationAddressIn_NORTH[4]), .Y(n4572) );
  AOI22X1TS U5223 ( .A0(n4571), .A1(n4583), .B0(n4572), .B1(n4584), .Y(n4576)
         );
  CLKBUFX2TS U5224 ( .A(destinationAddressIn_SOUTH[4]), .Y(n4573) );
  NAND2X1TS U5225 ( .A(n4573), .B(n4586), .Y(n4574) );
  CLKBUFX2TS U5226 ( .A(destinationAddressIn_WEST[5]), .Y(n4578) );
  AOI22X1TS U5227 ( .A0(n4578), .A1(n4580), .B0(
        \destinationAddressbuffer[7][5] ), .B1(n4579), .Y(n4590) );
  CLKBUFX2TS U5228 ( .A(destinationAddressIn_NORTH[5]), .Y(n4581) );
  CLKBUFX2TS U5229 ( .A(destinationAddressIn_EAST[5]), .Y(n4582) );
  AOI22X1TS U5230 ( .A0(n4581), .A1(n4584), .B0(n4582), .B1(n4583), .Y(n4589)
         );
  CLKBUFX2TS U5231 ( .A(destinationAddressIn_SOUTH[5]), .Y(n4585) );
  NAND2X1TS U5232 ( .A(n4585), .B(n4586), .Y(n4587) );
  AOI22X1TS U5233 ( .A0(n4540), .A1(n4616), .B0(
        \destinationAddressbuffer[6][0] ), .B1(n4612), .Y(n4594) );
  AOI22X1TS U5234 ( .A0(n4607), .A1(n4539), .B0(n4614), .B1(n4541), .Y(n4593)
         );
  NAND2X1TS U5235 ( .A(n4613), .B(n4538), .Y(n4591) );
  AOI22X1TS U5236 ( .A0(n4548), .A1(n4614), .B0(
        \destinationAddressbuffer[6][1] ), .B1(n4612), .Y(n4598) );
  AOI22X1TS U5237 ( .A0(n4607), .A1(n4549), .B0(n4613), .B1(n4547), .Y(n4597)
         );
  NAND2X1TS U5238 ( .A(n4616), .B(n4546), .Y(n4595) );
  AOI22X1TS U5239 ( .A0(n4556), .A1(n4607), .B0(
        \destinationAddressbuffer[6][2] ), .B1(n4612), .Y(n4602) );
  AOI22X1TS U5240 ( .A0(n4613), .A1(n4555), .B0(n4614), .B1(n4557), .Y(n4601)
         );
  NAND2X1TS U5241 ( .A(n4616), .B(n4554), .Y(n4599) );
  AOI22X1TS U5242 ( .A0(n4562), .A1(n4613), .B0(
        \destinationAddressbuffer[6][3] ), .B1(n4612), .Y(n4606) );
  AOI22X1TS U5243 ( .A0(n4607), .A1(n4565), .B0(n4616), .B1(n4564), .Y(n4605)
         );
  NAND2X1TS U5244 ( .A(n4614), .B(n4563), .Y(n4603) );
  AOI22X1TS U5245 ( .A0(n4573), .A1(n4607), .B0(
        \destinationAddressbuffer[6][4] ), .B1(n4612), .Y(n4611) );
  AOI22X1TS U5246 ( .A0(n4613), .A1(n4571), .B0(n4614), .B1(n4572), .Y(n4610)
         );
  NAND2X1TS U5247 ( .A(n4616), .B(n4570), .Y(n4608) );
  AOI22X1TS U5248 ( .A0(n4582), .A1(n4613), .B0(
        \destinationAddressbuffer[6][5] ), .B1(n4612), .Y(n4620) );
  AOI22X1TS U5249 ( .A0(n4615), .A1(n4585), .B0(n4614), .B1(n4581), .Y(n4619)
         );
  NAND2X1TS U5250 ( .A(n4616), .B(n4578), .Y(n4617) );
  AOI22X1TS U5251 ( .A0(n4538), .A1(n4643), .B0(
        \destinationAddressbuffer[5][0] ), .B1(n4641), .Y(n4624) );
  AOI22X1TS U5252 ( .A0(n4539), .A1(n4644), .B0(n4540), .B1(n4642), .Y(n4623)
         );
  NAND2X1TS U5253 ( .A(n4541), .B(n4645), .Y(n4621) );
  AOI22X1TS U5254 ( .A0(n4546), .A1(n4642), .B0(
        \destinationAddressbuffer[5][1] ), .B1(n4641), .Y(n4628) );
  AOI22X1TS U5255 ( .A0(n4547), .A1(n4643), .B0(n4549), .B1(n4644), .Y(n4627)
         );
  NAND2X1TS U5256 ( .A(n4548), .B(n4645), .Y(n4625) );
  AOI22X1TS U5257 ( .A0(n4555), .A1(n4643), .B0(
        \destinationAddressbuffer[5][2] ), .B1(n4641), .Y(n4632) );
  AOI22X1TS U5258 ( .A0(n4554), .A1(n4642), .B0(n4556), .B1(n4644), .Y(n4631)
         );
  NAND2X1TS U5259 ( .A(n4557), .B(n4645), .Y(n4629) );
  AOI22X1TS U5260 ( .A0(n4562), .A1(n4643), .B0(
        \destinationAddressbuffer[5][3] ), .B1(n4641), .Y(n4636) );
  AOI22X1TS U5261 ( .A0(n4563), .A1(n4645), .B0(n4564), .B1(n4642), .Y(n4635)
         );
  NAND2X1TS U5262 ( .A(n4565), .B(n4644), .Y(n4633) );
  AOI22X1TS U5263 ( .A0(n4571), .A1(n4643), .B0(
        \destinationAddressbuffer[5][4] ), .B1(n4641), .Y(n4640) );
  AOI22X1TS U5264 ( .A0(n4570), .A1(n4642), .B0(n4573), .B1(n4644), .Y(n4639)
         );
  NAND2X1TS U5265 ( .A(n4572), .B(n4645), .Y(n4637) );
  AOI22X1TS U5266 ( .A0(n4578), .A1(n4642), .B0(
        \destinationAddressbuffer[5][5] ), .B1(n4641), .Y(n4649) );
  AOI22X1TS U5267 ( .A0(n4585), .A1(n4644), .B0(n4582), .B1(n4643), .Y(n4648)
         );
  NAND2X1TS U5268 ( .A(n4581), .B(n4645), .Y(n4646) );
  AOI22X1TS U5269 ( .A0(n4541), .A1(n4674), .B0(
        \destinationAddressbuffer[4][0] ), .B1(n4671), .Y(n4653) );
  AOI22X1TS U5270 ( .A0(n4672), .A1(n4538), .B0(n4673), .B1(n4539), .Y(n4652)
         );
  NAND2X1TS U5271 ( .A(n4666), .B(n4540), .Y(n4650) );
  AOI22X1TS U5272 ( .A0(n4547), .A1(n4672), .B0(
        \destinationAddressbuffer[4][1] ), .B1(n4671), .Y(n4657) );
  AOI22X1TS U5273 ( .A0(n4674), .A1(n4548), .B0(n4666), .B1(n4546), .Y(n4656)
         );
  NAND2X1TS U5274 ( .A(n4673), .B(n4549), .Y(n4654) );
  AOI22X1TS U5275 ( .A0(n4554), .A1(n4666), .B0(
        \destinationAddressbuffer[4][2] ), .B1(n4671), .Y(n4661) );
  AOI22X1TS U5276 ( .A0(n4672), .A1(n4555), .B0(n4674), .B1(n4557), .Y(n4660)
         );
  NAND2X1TS U5277 ( .A(n4673), .B(n4556), .Y(n4658) );
  AOI22X1TS U5278 ( .A0(n4563), .A1(n4674), .B0(
        \destinationAddressbuffer[4][3] ), .B1(n4671), .Y(n4665) );
  AOI22X1TS U5279 ( .A0(n4666), .A1(n4564), .B0(n4673), .B1(n4565), .Y(n4664)
         );
  NAND2X1TS U5280 ( .A(n4672), .B(n4562), .Y(n4662) );
  AOI22X1TS U5281 ( .A0(n4573), .A1(n4673), .B0(
        \destinationAddressbuffer[4][4] ), .B1(n4671), .Y(n4670) );
  AOI22X1TS U5282 ( .A0(n4672), .A1(n4571), .B0(n4666), .B1(n4570), .Y(n4669)
         );
  NAND2X1TS U5283 ( .A(n4674), .B(n4572), .Y(n4667) );
  AOI22X1TS U5284 ( .A0(n4582), .A1(n4672), .B0(
        \destinationAddressbuffer[4][5] ), .B1(n4671), .Y(n4678) );
  AOI22X1TS U5285 ( .A0(n4674), .A1(n4581), .B0(n4673), .B1(n4585), .Y(n4677)
         );
  NAND2X1TS U5286 ( .A(n4666), .B(n4578), .Y(n4675) );
  AOI22X1TS U5287 ( .A0(n4538), .A1(n4696), .B0(
        \destinationAddressbuffer[3][0] ), .B1(n4701), .Y(n4682) );
  AOI22X1TS U5288 ( .A0(n4703), .A1(n4541), .B0(n4702), .B1(n4539), .Y(n4681)
         );
  NAND2X1TS U5289 ( .A(n4687), .B(n4540), .Y(n4679) );
  AOI22X1TS U5290 ( .A0(n4547), .A1(n4696), .B0(
        \destinationAddressbuffer[3][1] ), .B1(n4701), .Y(n4686) );
  AOI22X1TS U5291 ( .A0(n4703), .A1(n4548), .B0(n4687), .B1(n4546), .Y(n4685)
         );
  NAND2X1TS U5292 ( .A(n4702), .B(n4549), .Y(n4683) );
  AOI22X1TS U5293 ( .A0(n4556), .A1(n4702), .B0(
        \destinationAddressbuffer[3][2] ), .B1(n4701), .Y(n4691) );
  AOI22X1TS U5294 ( .A0(n4703), .A1(n4557), .B0(n4687), .B1(n4554), .Y(n4690)
         );
  NAND2X1TS U5295 ( .A(n4696), .B(n4555), .Y(n4688) );
  AOI22X1TS U5296 ( .A0(n4563), .A1(n4703), .B0(
        \destinationAddressbuffer[3][3] ), .B1(n4701), .Y(n4695) );
  AOI22X1TS U5297 ( .A0(n4696), .A1(n4562), .B0(n4702), .B1(n4565), .Y(n4694)
         );
  NAND2X1TS U5298 ( .A(n4687), .B(n4564), .Y(n4692) );
  AOI22X1TS U5299 ( .A0(n4571), .A1(n4696), .B0(
        \destinationAddressbuffer[3][4] ), .B1(n4701), .Y(n4700) );
  AOI22X1TS U5300 ( .A0(n4703), .A1(n4572), .B0(n4702), .B1(n4573), .Y(n4699)
         );
  NAND2X1TS U5301 ( .A(n4687), .B(n4570), .Y(n4697) );
  AOI22X1TS U5302 ( .A0(n4582), .A1(n4696), .B0(
        \destinationAddressbuffer[3][5] ), .B1(n4701), .Y(n4707) );
  AOI22X1TS U5303 ( .A0(n4703), .A1(n4581), .B0(n4702), .B1(n4585), .Y(n4706)
         );
  NAND2X1TS U5304 ( .A(n4687), .B(n4578), .Y(n4704) );
  AOI22X1TS U5305 ( .A0(n4540), .A1(n4731), .B0(
        \destinationAddressbuffer[2][0] ), .B1(n4728), .Y(n4711) );
  AOI22X1TS U5306 ( .A0(n4729), .A1(n4538), .B0(n4730), .B1(n4539), .Y(n4710)
         );
  NAND2X1TS U5307 ( .A(n2952), .B(n4541), .Y(n4708) );
  AOI22X1TS U5308 ( .A0(n4548), .A1(n2952), .B0(
        \destinationAddressbuffer[2][1] ), .B1(n4728), .Y(n4715) );
  AOI22X1TS U5309 ( .A0(n4729), .A1(n4547), .B0(n4730), .B1(n4549), .Y(n4714)
         );
  NAND2X1TS U5310 ( .A(n4731), .B(n4546), .Y(n4712) );
  AOI22X1TS U5311 ( .A0(n4557), .A1(n2952), .B0(
        \destinationAddressbuffer[2][2] ), .B1(n4728), .Y(n4719) );
  AOI22X1TS U5312 ( .A0(n4729), .A1(n4555), .B0(n4730), .B1(n4556), .Y(n4718)
         );
  NAND2X1TS U5313 ( .A(n4731), .B(n4554), .Y(n4716) );
  AOI22X1TS U5314 ( .A0(n4564), .A1(n4731), .B0(
        \destinationAddressbuffer[2][3] ), .B1(n4728), .Y(n4723) );
  AOI22X1TS U5315 ( .A0(n2952), .A1(n4563), .B0(n4729), .B1(n4562), .Y(n4722)
         );
  NAND2X1TS U5316 ( .A(n4730), .B(n4565), .Y(n4720) );
  AOI22X1TS U5317 ( .A0(n4570), .A1(n4731), .B0(
        \destinationAddressbuffer[2][4] ), .B1(n4728), .Y(n4727) );
  AOI22X1TS U5318 ( .A0(n4729), .A1(n4571), .B0(n4730), .B1(n4573), .Y(n4726)
         );
  NAND2X1TS U5319 ( .A(n2952), .B(n4572), .Y(n4724) );
  AOI22X1TS U5320 ( .A0(n4582), .A1(n4729), .B0(
        \destinationAddressbuffer[2][5] ), .B1(n4728), .Y(n4735) );
  AOI22X1TS U5321 ( .A0(n4731), .A1(n4578), .B0(n4730), .B1(n4585), .Y(n4734)
         );
  NAND2X1TS U5322 ( .A(n2952), .B(n4581), .Y(n4732) );
  AOI22X1TS U5323 ( .A0(n4538), .A1(n4758), .B0(
        \destinationAddressbuffer[1][0] ), .B1(n4744), .Y(n4739) );
  AOI22X1TS U5324 ( .A0(n4541), .A1(n4761), .B0(n4540), .B1(n4760), .Y(n4738)
         );
  NAND2X1TS U5325 ( .A(n4539), .B(n4759), .Y(n4736) );
  AOI22X1TS U5326 ( .A0(n4547), .A1(n4758), .B0(
        \destinationAddressbuffer[1][1] ), .B1(n4744), .Y(n4743) );
  AOI22X1TS U5327 ( .A0(n4546), .A1(n4760), .B0(n4549), .B1(n4759), .Y(n4742)
         );
  NAND2X1TS U5328 ( .A(n4548), .B(n4761), .Y(n4740) );
  AOI22X1TS U5329 ( .A0(n4554), .A1(n4760), .B0(
        \destinationAddressbuffer[1][2] ), .B1(n4744), .Y(n4748) );
  AOI22X1TS U5330 ( .A0(n4557), .A1(n4761), .B0(n4555), .B1(n4758), .Y(n4747)
         );
  NAND2X1TS U5331 ( .A(n4556), .B(n4759), .Y(n4745) );
  AOI22X1TS U5332 ( .A0(n4564), .A1(n4760), .B0(
        \destinationAddressbuffer[1][3] ), .B1(n4757), .Y(n4752) );
  AOI22X1TS U5333 ( .A0(n4563), .A1(n4761), .B0(n4562), .B1(n4758), .Y(n4751)
         );
  NAND2X1TS U5334 ( .A(n4565), .B(n4759), .Y(n4749) );
  AOI22X1TS U5335 ( .A0(n4570), .A1(n4760), .B0(
        \destinationAddressbuffer[1][4] ), .B1(n4757), .Y(n4756) );
  AOI22X1TS U5336 ( .A0(n4571), .A1(n4758), .B0(n4573), .B1(n4759), .Y(n4755)
         );
  NAND2X1TS U5337 ( .A(n4572), .B(n4761), .Y(n4753) );
  AOI22X1TS U5338 ( .A0(n4582), .A1(n4758), .B0(
        \destinationAddressbuffer[1][5] ), .B1(n4757), .Y(n4765) );
  AOI22X1TS U5339 ( .A0(n4578), .A1(n4760), .B0(n4585), .B1(n4759), .Y(n4764)
         );
  NAND2X1TS U5340 ( .A(n4581), .B(n4761), .Y(n4762) );
  AOI22X1TS U5341 ( .A0(n4541), .A1(n4790), .B0(
        \destinationAddressbuffer[0][0] ), .B1(n4787), .Y(n4769) );
  AOI22X1TS U5342 ( .A0(n4788), .A1(n4540), .B0(n4782), .B1(n4538), .Y(n4768)
         );
  NAND2X1TS U5343 ( .A(n4789), .B(n4539), .Y(n4766) );
  AOI22X1TS U5344 ( .A0(n4548), .A1(n4790), .B0(
        \destinationAddressbuffer[0][1] ), .B1(n4787), .Y(n4773) );
  AOI22X1TS U5345 ( .A0(n4782), .A1(n4547), .B0(n4789), .B1(n4549), .Y(n4772)
         );
  NAND2X1TS U5346 ( .A(n4788), .B(n4546), .Y(n4770) );
  AOI22X1TS U5347 ( .A0(n4557), .A1(n4790), .B0(
        \destinationAddressbuffer[0][2] ), .B1(n4787), .Y(n4777) );
  AOI22X1TS U5348 ( .A0(n4788), .A1(n4554), .B0(n4789), .B1(n4556), .Y(n4776)
         );
  NAND2X1TS U5349 ( .A(n4782), .B(n4555), .Y(n4774) );
  AOI22X1TS U5350 ( .A0(n4562), .A1(n4782), .B0(
        \destinationAddressbuffer[0][3] ), .B1(n4787), .Y(n4781) );
  AOI22X1TS U5351 ( .A0(n4790), .A1(n4563), .B0(n4789), .B1(n4565), .Y(n4780)
         );
  NAND2X1TS U5352 ( .A(n4788), .B(n4564), .Y(n4778) );
  AOI22X1TS U5353 ( .A0(n4571), .A1(n4782), .B0(
        \destinationAddressbuffer[0][4] ), .B1(n4787), .Y(n4786) );
  AOI22X1TS U5354 ( .A0(n4790), .A1(n4572), .B0(n4789), .B1(n4573), .Y(n4785)
         );
  NAND2X1TS U5355 ( .A(n4788), .B(n4570), .Y(n4783) );
  AOI22X1TS U5356 ( .A0(n4578), .A1(n4788), .B0(
        \destinationAddressbuffer[0][5] ), .B1(n4787), .Y(n4794) );
  AOI22X1TS U5357 ( .A0(n4790), .A1(n4581), .B0(n4789), .B1(n4585), .Y(n4793)
         );
  NAND2X1TS U5358 ( .A(n4782), .B(n4582), .Y(n4791) );
  INVX2TS U5359 ( .A(n4795), .Y(n4819) );
  OAI22X1TS U5360 ( .A0(n4797), .A1(n4815), .B0(n4796), .B1(n4816), .Y(n4801)
         );
  OAI211XLTS U5361 ( .A0(n4799), .A1(n4821), .B0(empty_reg), .C0(n4798), .Y(
        n4800) );
  AOI211XLTS U5362 ( .A0(n4460), .A1(n4819), .B0(n4801), .C0(n4800), .Y(n4811)
         );
  AO22XLTS U5363 ( .A0(readOutbuffer[2]), .A1(n5310), .B0(readOutbuffer[7]), 
        .B1(n2895), .Y(n4808) );
  AOI22X1TS U5364 ( .A0(readOutbuffer[3]), .A1(n2891), .B0(readOutbuffer[5]), 
        .B1(n2892), .Y(n4806) );
  AOI22X1TS U5365 ( .A0(readOutbuffer[4]), .A1(n5295), .B0(readOutbuffer[1]), 
        .B1(n2894), .Y(n4805) );
  AOI22X1TS U5366 ( .A0(readOutbuffer[6]), .A1(n2893), .B0(readOutbuffer[0]), 
        .B1(n5312), .Y(n4804) );
  NAND3XLTS U5367 ( .A(n4806), .B(n4805), .C(n4804), .Y(n4807) );
  CLKAND2X2TS U5368 ( .A(n4932), .B(n4809), .Y(n4825) );
  OAI2BB2XLTS U5369 ( .B0(n4811), .B1(n4810), .A0N(n4825), .A1N(readOut), .Y(
        n2450) );
  AO22XLTS U5370 ( .A0(writeOutbuffer[4]), .A1(n5249), .B0(writeOutbuffer[2]), 
        .B1(n5310), .Y(n4824) );
  AOI22X1TS U5371 ( .A0(writeOutbuffer[3]), .A1(n2891), .B0(writeOutbuffer[0]), 
        .B1(n5312), .Y(n4814) );
  AOI22X1TS U5372 ( .A0(writeOutbuffer[6]), .A1(n2893), .B0(writeOutbuffer[5]), 
        .B1(n2892), .Y(n4813) );
  AOI22X1TS U5373 ( .A0(writeOutbuffer[7]), .A1(n2895), .B0(writeOutbuffer[1]), 
        .B1(n2894), .Y(n4812) );
  NAND3XLTS U5374 ( .A(n4814), .B(n4813), .C(n4812), .Y(n4823) );
  OAI22X1TS U5375 ( .A0(n4817), .A1(n4816), .B0(n2981), .B1(n4815), .Y(n4818)
         );
  AOI21X1TS U5376 ( .A0(n2982), .A1(n4819), .B0(n4818), .Y(n4820) );
  OAI211XLTS U5377 ( .A0(n2984), .A1(n4821), .B0(empty_reg), .C0(n4820), .Y(
        n4822) );
  OAI2BB2XLTS U5378 ( .B0(n2896), .B1(n4826), .A0N(writeOut), .A1N(n4825), .Y(
        n2449) );
  AOI22X1TS U5379 ( .A0(n3002), .A1(n5280), .B0(n3004), .B1(n5290), .Y(n4834)
         );
  AOI22X1TS U5380 ( .A0(n3001), .A1(n5304), .B0(n3005), .B1(n2908), .Y(n4833)
         );
  AOI22X1TS U5381 ( .A0(\destinationAddressbuffer[2][6] ), .A1(n5310), .B0(
        \destinationAddressbuffer[0][6] ), .B1(n5312), .Y(n4830) );
  AOI22X1TS U5382 ( .A0(\destinationAddressbuffer[4][6] ), .A1(n5295), .B0(
        \destinationAddressbuffer[1][6] ), .B1(n2894), .Y(n4829) );
  AOI22X1TS U5383 ( .A0(\destinationAddressbuffer[3][6] ), .A1(n2891), .B0(
        \destinationAddressbuffer[7][6] ), .B1(n2895), .Y(n4828) );
  AOI22X1TS U5384 ( .A0(\destinationAddressbuffer[6][6] ), .A1(n2893), .B0(
        \destinationAddressbuffer[5][6] ), .B1(n2892), .Y(n4827) );
  NAND4XLTS U5385 ( .A(n4830), .B(n4829), .C(n4828), .D(n4827), .Y(n4831) );
  AOI22X1TS U5386 ( .A0(n5318), .A1(destinationAddressOut[6]), .B0(n2890), 
        .B1(n4831), .Y(n4832) );
  AOI22X1TS U5387 ( .A0(n2974), .A1(n5304), .B0(n2972), .B1(n5280), .Y(n4842)
         );
  AOI22X1TS U5388 ( .A0(n2975), .A1(n5290), .B0(n2976), .B1(n2908), .Y(n4841)
         );
  AOI22X1TS U5389 ( .A0(\destinationAddressbuffer[3][7] ), .A1(n2891), .B0(
        \destinationAddressbuffer[2][7] ), .B1(n5310), .Y(n4838) );
  AOI22X1TS U5390 ( .A0(\destinationAddressbuffer[6][7] ), .A1(n2893), .B0(
        \destinationAddressbuffer[7][7] ), .B1(n2895), .Y(n4837) );
  AOI22X1TS U5391 ( .A0(\destinationAddressbuffer[0][7] ), .A1(n5312), .B0(
        \destinationAddressbuffer[5][7] ), .B1(n2892), .Y(n4836) );
  AOI22X1TS U5392 ( .A0(\destinationAddressbuffer[4][7] ), .A1(n5295), .B0(
        \destinationAddressbuffer[1][7] ), .B1(n2894), .Y(n4835) );
  NAND4XLTS U5393 ( .A(n4838), .B(n4837), .C(n4836), .D(n4835), .Y(n4839) );
  AOI22X1TS U5394 ( .A0(n4932), .A1(destinationAddressOut[7]), .B0(n2890), 
        .B1(n4839), .Y(n4840) );
  AOI22X1TS U5395 ( .A0(n2989), .A1(n5290), .B0(n2990), .B1(n2908), .Y(n4850)
         );
  AOI22X1TS U5396 ( .A0(n2987), .A1(n5280), .B0(n2988), .B1(n5304), .Y(n4849)
         );
  AOI22X1TS U5397 ( .A0(\destinationAddressbuffer[6][8] ), .A1(n2893), .B0(
        \destinationAddressbuffer[3][8] ), .B1(n2891), .Y(n4846) );
  AOI22X1TS U5398 ( .A0(\destinationAddressbuffer[4][8] ), .A1(n5295), .B0(
        \destinationAddressbuffer[5][8] ), .B1(n2892), .Y(n4845) );
  AOI22X1TS U5399 ( .A0(\destinationAddressbuffer[2][8] ), .A1(n5310), .B0(
        \destinationAddressbuffer[7][8] ), .B1(n4884), .Y(n4844) );
  AOI22X1TS U5400 ( .A0(\destinationAddressbuffer[0][8] ), .A1(n5312), .B0(
        \destinationAddressbuffer[1][8] ), .B1(n2894), .Y(n4843) );
  NAND4XLTS U5401 ( .A(n4846), .B(n4845), .C(n4844), .D(n4843), .Y(n4847) );
  AOI22X1TS U5402 ( .A0(n5318), .A1(destinationAddressOut[8]), .B0(n2890), 
        .B1(n4847), .Y(n4848) );
  AOI22X1TS U5403 ( .A0(n3121), .A1(n5304), .B0(n3122), .B1(n5280), .Y(n4858)
         );
  AOI22X1TS U5404 ( .A0(n3120), .A1(n5290), .B0(n3123), .B1(n2908), .Y(n4857)
         );
  AOI22X1TS U5405 ( .A0(\destinationAddressbuffer[4][9] ), .A1(n5295), .B0(
        \destinationAddressbuffer[2][9] ), .B1(n5310), .Y(n4854) );
  AOI22X1TS U5406 ( .A0(\destinationAddressbuffer[7][9] ), .A1(n2895), .B0(
        \destinationAddressbuffer[1][9] ), .B1(n2894), .Y(n4853) );
  AOI22X1TS U5407 ( .A0(\destinationAddressbuffer[0][9] ), .A1(n5312), .B0(
        \destinationAddressbuffer[5][9] ), .B1(n2892), .Y(n4852) );
  AOI22X1TS U5408 ( .A0(\destinationAddressbuffer[6][9] ), .A1(n2893), .B0(
        \destinationAddressbuffer[3][9] ), .B1(n2891), .Y(n4851) );
  NAND4XLTS U5409 ( .A(n4854), .B(n4853), .C(n4852), .D(n4851), .Y(n4855) );
  AOI22X1TS U5410 ( .A0(n4932), .A1(destinationAddressOut[9]), .B0(n2890), 
        .B1(n4855), .Y(n4856) );
  AOI22X1TS U5411 ( .A0(n3027), .A1(n5304), .B0(n3030), .B1(n5290), .Y(n4866)
         );
  AOI22X1TS U5412 ( .A0(n3028), .A1(n5280), .B0(n3031), .B1(n2908), .Y(n4865)
         );
  AOI22X1TS U5413 ( .A0(\destinationAddressbuffer[3][10] ), .A1(n2891), .B0(
        \destinationAddressbuffer[5][10] ), .B1(n2892), .Y(n4862) );
  AOI22X1TS U5414 ( .A0(\destinationAddressbuffer[2][10] ), .A1(n5310), .B0(
        \destinationAddressbuffer[0][10] ), .B1(n5312), .Y(n4861) );
  AOI22X1TS U5415 ( .A0(\destinationAddressbuffer[4][10] ), .A1(n5295), .B0(
        \destinationAddressbuffer[7][10] ), .B1(n2895), .Y(n4860) );
  AOI22X1TS U5416 ( .A0(\destinationAddressbuffer[6][10] ), .A1(n2893), .B0(
        \destinationAddressbuffer[1][10] ), .B1(n2894), .Y(n4859) );
  NAND4XLTS U5417 ( .A(n4862), .B(n4861), .C(n4860), .D(n4859), .Y(n4863) );
  AOI22X1TS U5418 ( .A0(n4932), .A1(destinationAddressOut[10]), .B0(n2890), 
        .B1(n4863), .Y(n4864) );
  AOI22X1TS U5419 ( .A0(n3075), .A1(n5280), .B0(n3077), .B1(n5290), .Y(n4874)
         );
  AOI22X1TS U5420 ( .A0(n3073), .A1(n2908), .B0(n3078), .B1(n5304), .Y(n4873)
         );
  AOI22X1TS U5421 ( .A0(\destinationAddressbuffer[6][11] ), .A1(n2893), .B0(
        \destinationAddressbuffer[2][11] ), .B1(n5310), .Y(n4870) );
  AOI22X1TS U5422 ( .A0(\destinationAddressbuffer[0][11] ), .A1(n5312), .B0(
        \destinationAddressbuffer[5][11] ), .B1(n2892), .Y(n4869) );
  AOI22X1TS U5423 ( .A0(\destinationAddressbuffer[3][11] ), .A1(n2891), .B0(
        \destinationAddressbuffer[1][11] ), .B1(n2894), .Y(n4868) );
  AOI22X1TS U5424 ( .A0(\destinationAddressbuffer[4][11] ), .A1(n5295), .B0(
        \destinationAddressbuffer[7][11] ), .B1(n2895), .Y(n4867) );
  NAND4XLTS U5425 ( .A(n4870), .B(n4869), .C(n4868), .D(n4867), .Y(n4871) );
  AOI22X1TS U5426 ( .A0(n5318), .A1(destinationAddressOut[11]), .B0(n2890), 
        .B1(n4871), .Y(n4872) );
  AOI22X1TS U5427 ( .A0(n3038), .A1(n5290), .B0(n3039), .B1(n2908), .Y(n4883)
         );
  AOI22X1TS U5428 ( .A0(n3037), .A1(n5304), .B0(n3035), .B1(n5280), .Y(n4882)
         );
  AOI22X1TS U5429 ( .A0(\destinationAddressbuffer[2][12] ), .A1(n5310), .B0(
        \destinationAddressbuffer[5][12] ), .B1(n2892), .Y(n4879) );
  AOI22X1TS U5430 ( .A0(\destinationAddressbuffer[6][12] ), .A1(n2893), .B0(
        \destinationAddressbuffer[7][12] ), .B1(n4884), .Y(n4878) );
  AOI22X1TS U5431 ( .A0(\destinationAddressbuffer[4][12] ), .A1(n5295), .B0(
        \destinationAddressbuffer[3][12] ), .B1(n4875), .Y(n4877) );
  AOI22X1TS U5432 ( .A0(\destinationAddressbuffer[0][12] ), .A1(n5312), .B0(
        \destinationAddressbuffer[1][12] ), .B1(n2894), .Y(n4876) );
  NAND4XLTS U5433 ( .A(n4879), .B(n4878), .C(n4877), .D(n4876), .Y(n4880) );
  AOI22X1TS U5434 ( .A0(n5318), .A1(destinationAddressOut[12]), .B0(n2890), 
        .B1(n4880), .Y(n4881) );
  AOI22X1TS U5435 ( .A0(n3114), .A1(n5290), .B0(n3116), .B1(n5280), .Y(n4892)
         );
  AOI22X1TS U5436 ( .A0(n3115), .A1(n2908), .B0(n3117), .B1(n5304), .Y(n4891)
         );
  AOI22X1TS U5437 ( .A0(\destinationAddressbuffer[4][13] ), .A1(n5295), .B0(
        \destinationAddressbuffer[0][13] ), .B1(n5312), .Y(n4888) );
  AOI22X1TS U5438 ( .A0(\destinationAddressbuffer[3][13] ), .A1(n2891), .B0(
        \destinationAddressbuffer[5][13] ), .B1(n2892), .Y(n4887) );
  AOI22X1TS U5439 ( .A0(\destinationAddressbuffer[6][13] ), .A1(n5311), .B0(
        \destinationAddressbuffer[7][13] ), .B1(n4884), .Y(n4886) );
  AOI22X1TS U5440 ( .A0(\destinationAddressbuffer[2][13] ), .A1(n5310), .B0(
        \destinationAddressbuffer[1][13] ), .B1(n2894), .Y(n4885) );
  NAND4XLTS U5441 ( .A(n4888), .B(n4887), .C(n4886), .D(n4885), .Y(n4889) );
  AOI22X1TS U5442 ( .A0(n4932), .A1(destinationAddressOut[13]), .B0(n2890), 
        .B1(n4889), .Y(n4890) );
  AOI22X1TS U5443 ( .A0(n4539), .A1(n5304), .B0(n4541), .B1(n5290), .Y(n4901)
         );
  AOI22X1TS U5444 ( .A0(n4538), .A1(n5280), .B0(n4540), .B1(n2908), .Y(n4900)
         );
  AOI22X1TS U5445 ( .A0(\destinationAddressbuffer[7][0] ), .A1(n2895), .B0(
        \destinationAddressbuffer[1][0] ), .B1(n2894), .Y(n4896) );
  AOI22X1TS U5446 ( .A0(\destinationAddressbuffer[3][0] ), .A1(n2891), .B0(
        \destinationAddressbuffer[0][0] ), .B1(n5312), .Y(n4895) );
  AOI22X1TS U5447 ( .A0(\destinationAddressbuffer[6][0] ), .A1(n2893), .B0(
        \destinationAddressbuffer[5][0] ), .B1(n2892), .Y(n4894) );
  AOI22X1TS U5448 ( .A0(\destinationAddressbuffer[4][0] ), .A1(n5295), .B0(
        \destinationAddressbuffer[2][0] ), .B1(n5310), .Y(n4893) );
  NAND4XLTS U5449 ( .A(n4896), .B(n4895), .C(n4894), .D(n4893), .Y(n4897) );
  AOI22X1TS U5450 ( .A0(n4932), .A1(destinationAddressOut[0]), .B0(n2890), 
        .B1(n4897), .Y(n4899) );
  AOI22X1TS U5451 ( .A0(n4546), .A1(n2908), .B0(n4547), .B1(n5280), .Y(n4909)
         );
  AOI22X1TS U5452 ( .A0(n4549), .A1(n5304), .B0(n4548), .B1(n5290), .Y(n4908)
         );
  AOI22X1TS U5453 ( .A0(\destinationAddressbuffer[3][1] ), .A1(n2891), .B0(
        \destinationAddressbuffer[1][1] ), .B1(n2894), .Y(n4905) );
  AOI22X1TS U5454 ( .A0(\destinationAddressbuffer[4][1] ), .A1(n5295), .B0(
        \destinationAddressbuffer[5][1] ), .B1(n2892), .Y(n4904) );
  AOI22X1TS U5455 ( .A0(\destinationAddressbuffer[6][1] ), .A1(n2893), .B0(
        \destinationAddressbuffer[2][1] ), .B1(n5310), .Y(n4903) );
  AOI22X1TS U5456 ( .A0(\destinationAddressbuffer[0][1] ), .A1(n5312), .B0(
        \destinationAddressbuffer[7][1] ), .B1(n2895), .Y(n4902) );
  NAND4XLTS U5457 ( .A(n4905), .B(n4904), .C(n4903), .D(n4902), .Y(n4906) );
  AOI22X1TS U5458 ( .A0(n5318), .A1(destinationAddressOut[1]), .B0(n2890), 
        .B1(n4906), .Y(n4907) );
  NAND2X1TS U5459 ( .A(n4294), .B(n2922), .Y(n4949) );
  AOI22X1TS U5460 ( .A0(n4554), .A1(n2908), .B0(n4556), .B1(n5304), .Y(n4917)
         );
  AOI22X1TS U5461 ( .A0(n4557), .A1(n5290), .B0(n4555), .B1(n5280), .Y(n4916)
         );
  AOI22X1TS U5462 ( .A0(\destinationAddressbuffer[2][2] ), .A1(n5310), .B0(
        \destinationAddressbuffer[1][2] ), .B1(n2894), .Y(n4913) );
  AOI22X1TS U5463 ( .A0(\destinationAddressbuffer[0][2] ), .A1(n5312), .B0(
        \destinationAddressbuffer[5][2] ), .B1(n2892), .Y(n4912) );
  AOI22X1TS U5464 ( .A0(\destinationAddressbuffer[6][2] ), .A1(n5311), .B0(
        \destinationAddressbuffer[7][2] ), .B1(n2895), .Y(n4911) );
  AOI22X1TS U5465 ( .A0(\destinationAddressbuffer[4][2] ), .A1(n5249), .B0(
        \destinationAddressbuffer[3][2] ), .B1(n2891), .Y(n4910) );
  NAND4XLTS U5466 ( .A(n4913), .B(n4912), .C(n4911), .D(n4910), .Y(n4914) );
  AOI22X1TS U5467 ( .A0(n4932), .A1(destinationAddressOut[2]), .B0(n2890), 
        .B1(n4914), .Y(n4915) );
  NAND2X1TS U5468 ( .A(n4302), .B(n2922), .Y(n4958) );
  AOI22X1TS U5469 ( .A0(n4565), .A1(n5304), .B0(n4562), .B1(n5280), .Y(n4926)
         );
  AOI22X1TS U5470 ( .A0(n4563), .A1(n5290), .B0(n4564), .B1(n2908), .Y(n4925)
         );
  AOI22X1TS U5471 ( .A0(\destinationAddressbuffer[3][3] ), .A1(n2891), .B0(
        \destinationAddressbuffer[2][3] ), .B1(n5310), .Y(n4921) );
  AOI22X1TS U5472 ( .A0(\destinationAddressbuffer[4][3] ), .A1(n5249), .B0(
        \destinationAddressbuffer[5][3] ), .B1(n2892), .Y(n4920) );
  AOI22X1TS U5473 ( .A0(\destinationAddressbuffer[0][3] ), .A1(n5312), .B0(
        \destinationAddressbuffer[1][3] ), .B1(n2894), .Y(n4919) );
  AOI22X1TS U5474 ( .A0(\destinationAddressbuffer[6][3] ), .A1(n2893), .B0(
        \destinationAddressbuffer[7][3] ), .B1(n2895), .Y(n4918) );
  NAND4XLTS U5475 ( .A(n4921), .B(n4920), .C(n4919), .D(n4918), .Y(n4922) );
  AOI22X1TS U5476 ( .A0(n5318), .A1(destinationAddressOut[3]), .B0(n2890), 
        .B1(n4922), .Y(n4924) );
  AOI22X1TS U5477 ( .A0(n4572), .A1(n5290), .B0(n4573), .B1(n5304), .Y(n4935)
         );
  AOI22X1TS U5478 ( .A0(n4570), .A1(n2908), .B0(n4571), .B1(n5280), .Y(n4934)
         );
  AOI22X1TS U5479 ( .A0(\destinationAddressbuffer[6][4] ), .A1(n5311), .B0(
        \destinationAddressbuffer[2][4] ), .B1(n5310), .Y(n4930) );
  AOI22X1TS U5480 ( .A0(\destinationAddressbuffer[4][4] ), .A1(n5295), .B0(
        \destinationAddressbuffer[5][4] ), .B1(n2892), .Y(n4929) );
  AOI22X1TS U5481 ( .A0(\destinationAddressbuffer[3][4] ), .A1(n2891), .B0(
        \destinationAddressbuffer[0][4] ), .B1(n5312), .Y(n4928) );
  AOI22X1TS U5482 ( .A0(\destinationAddressbuffer[7][4] ), .A1(n2895), .B0(
        \destinationAddressbuffer[1][4] ), .B1(n2894), .Y(n4927) );
  NAND4XLTS U5483 ( .A(n4930), .B(n4929), .C(n4928), .D(n4927), .Y(n4931) );
  AOI22X1TS U5484 ( .A0(n4932), .A1(destinationAddressOut[4]), .B0(n2890), 
        .B1(n4931), .Y(n4933) );
  NAND2X1TS U5485 ( .A(n4313), .B(n2922), .Y(n4967) );
  AOI22X1TS U5486 ( .A0(n4578), .A1(n2908), .B0(n4581), .B1(n5290), .Y(n4943)
         );
  AOI22X1TS U5487 ( .A0(n4585), .A1(n5304), .B0(n4582), .B1(n5280), .Y(n4942)
         );
  AOI22X1TS U5488 ( .A0(\destinationAddressbuffer[3][5] ), .A1(n2891), .B0(
        \destinationAddressbuffer[7][5] ), .B1(n2895), .Y(n4939) );
  AOI22X1TS U5489 ( .A0(\destinationAddressbuffer[6][5] ), .A1(n5311), .B0(
        \destinationAddressbuffer[5][5] ), .B1(n2892), .Y(n4938) );
  AOI22X1TS U5490 ( .A0(\destinationAddressbuffer[4][5] ), .A1(n5249), .B0(
        \destinationAddressbuffer[2][5] ), .B1(n5310), .Y(n4937) );
  AOI22X1TS U5491 ( .A0(\destinationAddressbuffer[0][5] ), .A1(n5312), .B0(
        \destinationAddressbuffer[1][5] ), .B1(n2894), .Y(n4936) );
  NAND4XLTS U5492 ( .A(n4939), .B(n4938), .C(n4937), .D(n4936), .Y(n4940) );
  AOI22X1TS U5493 ( .A0(n5318), .A1(destinationAddressOut[5]), .B0(n2890), 
        .B1(n4940), .Y(n4941) );
  NAND2X1TS U5494 ( .A(n4322), .B(n2922), .Y(n4976) );
  AOI22X1TS U5495 ( .A0(n4291), .A1(n2908), .B0(n4292), .B1(n5290), .Y(n4952)
         );
  AOI22X1TS U5496 ( .A0(n4290), .A1(n5280), .B0(n4293), .B1(n5304), .Y(n4951)
         );
  AOI22X1TS U5497 ( .A0(\requesterAddressbuffer[6][1] ), .A1(n5311), .B0(
        \requesterAddressbuffer[7][1] ), .B1(n2895), .Y(n4947) );
  AOI22X1TS U5498 ( .A0(\requesterAddressbuffer[4][1] ), .A1(n5295), .B0(
        \requesterAddressbuffer[0][1] ), .B1(n5312), .Y(n4946) );
  AOI22X1TS U5499 ( .A0(\requesterAddressbuffer[2][1] ), .A1(n5310), .B0(
        \requesterAddressbuffer[1][1] ), .B1(n2894), .Y(n4945) );
  AOI22X1TS U5500 ( .A0(\requesterAddressbuffer[3][1] ), .A1(n2891), .B0(
        \requesterAddressbuffer[5][1] ), .B1(n2892), .Y(n4944) );
  NAND4XLTS U5501 ( .A(n4947), .B(n4946), .C(n4945), .D(n4944), .Y(n4948) );
  AOI22X1TS U5502 ( .A0(n5318), .A1(requesterAddressOut[1]), .B0(n2890), .B1(
        n4948), .Y(n4950) );
  AOI22X1TS U5503 ( .A0(n4298), .A1(n2908), .B0(n4300), .B1(n5304), .Y(n4961)
         );
  AOI22X1TS U5504 ( .A0(n4299), .A1(n5280), .B0(n4301), .B1(n5290), .Y(n4960)
         );
  AOI22X1TS U5505 ( .A0(\requesterAddressbuffer[3][2] ), .A1(n2891), .B0(
        \requesterAddressbuffer[2][2] ), .B1(n5310), .Y(n4956) );
  AOI22X1TS U5506 ( .A0(\requesterAddressbuffer[6][2] ), .A1(n2893), .B0(
        \requesterAddressbuffer[5][2] ), .B1(n2892), .Y(n4955) );
  AOI22X1TS U5507 ( .A0(\requesterAddressbuffer[4][2] ), .A1(n5249), .B0(
        \requesterAddressbuffer[0][2] ), .B1(n5312), .Y(n4954) );
  AOI22X1TS U5508 ( .A0(\requesterAddressbuffer[7][2] ), .A1(n2895), .B0(
        \requesterAddressbuffer[1][2] ), .B1(n2894), .Y(n4953) );
  NAND4XLTS U5509 ( .A(n4956), .B(n4955), .C(n4954), .D(n4953), .Y(n4957) );
  AOI22X1TS U5510 ( .A0(n5318), .A1(requesterAddressOut[2]), .B0(n2890), .B1(
        n4957), .Y(n4959) );
  AOI22X1TS U5511 ( .A0(n4312), .A1(n5304), .B0(n4311), .B1(n5290), .Y(n4970)
         );
  AOI22X1TS U5512 ( .A0(n4310), .A1(n5280), .B0(n4309), .B1(n2908), .Y(n4969)
         );
  AOI22X1TS U5513 ( .A0(\requesterAddressbuffer[2][4] ), .A1(n5310), .B0(
        \requesterAddressbuffer[1][4] ), .B1(n2894), .Y(n4965) );
  AOI22X1TS U5514 ( .A0(\requesterAddressbuffer[6][4] ), .A1(n2893), .B0(
        \requesterAddressbuffer[4][4] ), .B1(n5249), .Y(n4964) );
  AOI22X1TS U5515 ( .A0(\requesterAddressbuffer[3][4] ), .A1(n2891), .B0(
        \requesterAddressbuffer[0][4] ), .B1(n5312), .Y(n4963) );
  AOI22X1TS U5516 ( .A0(\requesterAddressbuffer[7][4] ), .A1(n2895), .B0(
        \requesterAddressbuffer[5][4] ), .B1(n2892), .Y(n4962) );
  NAND4XLTS U5517 ( .A(n4965), .B(n4964), .C(n4963), .D(n4962), .Y(n4966) );
  AOI22X1TS U5518 ( .A0(n5318), .A1(requesterAddressOut[4]), .B0(n2890), .B1(
        n4966), .Y(n4968) );
  AOI22X1TS U5519 ( .A0(n4321), .A1(n5304), .B0(n4320), .B1(n5290), .Y(n4979)
         );
  AOI22X1TS U5520 ( .A0(n4317), .A1(n2908), .B0(n4319), .B1(n5280), .Y(n4978)
         );
  AOI22X1TS U5521 ( .A0(\requesterAddressbuffer[0][5] ), .A1(n5312), .B0(
        \requesterAddressbuffer[5][5] ), .B1(n2892), .Y(n4974) );
  AOI22X1TS U5522 ( .A0(\requesterAddressbuffer[3][5] ), .A1(n2891), .B0(
        \requesterAddressbuffer[2][5] ), .B1(n5310), .Y(n4973) );
  AOI22X1TS U5523 ( .A0(\requesterAddressbuffer[7][5] ), .A1(n2895), .B0(
        \requesterAddressbuffer[1][5] ), .B1(n2894), .Y(n4972) );
  AOI22X1TS U5524 ( .A0(\requesterAddressbuffer[6][5] ), .A1(n2893), .B0(
        \requesterAddressbuffer[4][5] ), .B1(n5295), .Y(n4971) );
  NAND4XLTS U5525 ( .A(n4974), .B(n4973), .C(n4972), .D(n4971), .Y(n4975) );
  AOI22X1TS U5526 ( .A0(n5318), .A1(requesterAddressOut[5]), .B0(n2890), .B1(
        n4975), .Y(n4977) );
  AOI22X1TS U5527 ( .A0(n3022), .A1(n5280), .B0(n3019), .B1(n2922), .Y(n4989)
         );
  OAI22X1TS U5528 ( .A0(n3018), .A1(n5291), .B0(n4980), .B1(n5305), .Y(n4981)
         );
  AOI21X1TS U5529 ( .A0(n3021), .A1(n2908), .B0(n4981), .Y(n4988) );
  AOI22X1TS U5530 ( .A0(\dataoutbuffer[1][0] ), .A1(n2894), .B0(
        \dataoutbuffer[5][0] ), .B1(n2892), .Y(n4985) );
  AOI22X1TS U5531 ( .A0(\dataoutbuffer[0][0] ), .A1(n5312), .B0(
        \dataoutbuffer[6][0] ), .B1(n2893), .Y(n4984) );
  AOI22X1TS U5532 ( .A0(\dataoutbuffer[2][0] ), .A1(n5310), .B0(
        \dataoutbuffer[4][0] ), .B1(n5249), .Y(n4983) );
  AOI22X1TS U5533 ( .A0(\dataoutbuffer[3][0] ), .A1(n2891), .B0(
        \dataoutbuffer[7][0] ), .B1(n2895), .Y(n4982) );
  NAND4XLTS U5534 ( .A(n4985), .B(n4984), .C(n4983), .D(n4982), .Y(n4986) );
  AOI22X1TS U5535 ( .A0(n5318), .A1(dataOut[0]), .B0(n2890), .B1(n4986), .Y(
        n4987) );
  AOI22X1TS U5536 ( .A0(n3008), .A1(n5304), .B0(n3012), .B1(n2908), .Y(n5000)
         );
  OAI22X1TS U5537 ( .A0(n4991), .A1(n5305), .B0(n4990), .B1(n5307), .Y(n4992)
         );
  AOI21X1TS U5538 ( .A0(n3010), .A1(n2922), .B0(n4992), .Y(n4999) );
  AOI22X1TS U5539 ( .A0(\dataoutbuffer[0][1] ), .A1(n5312), .B0(
        \dataoutbuffer[2][1] ), .B1(n5310), .Y(n4996) );
  AOI22X1TS U5540 ( .A0(\dataoutbuffer[5][1] ), .A1(n2892), .B0(
        \dataoutbuffer[7][1] ), .B1(n2895), .Y(n4995) );
  AOI22X1TS U5541 ( .A0(\dataoutbuffer[6][1] ), .A1(n2893), .B0(
        \dataoutbuffer[1][1] ), .B1(n2894), .Y(n4994) );
  AOI22X1TS U5542 ( .A0(\dataoutbuffer[3][1] ), .A1(n2891), .B0(
        \dataoutbuffer[4][1] ), .B1(n5249), .Y(n4993) );
  NAND4XLTS U5543 ( .A(n4996), .B(n4995), .C(n4994), .D(n4993), .Y(n4997) );
  AOI22X1TS U5544 ( .A0(n5318), .A1(dataOut[1]), .B0(n2890), .B1(n4997), .Y(
        n4998) );
  AOI22X1TS U5545 ( .A0(n3493), .A1(n5290), .B0(n3490), .B1(n2922), .Y(n5010)
         );
  OAI22X1TS U5546 ( .A0(n5001), .A1(n5307), .B0(n3492), .B1(n5291), .Y(n5002)
         );
  AOI21X1TS U5547 ( .A0(n3489), .A1(n2908), .B0(n5002), .Y(n5009) );
  AOI22X1TS U5548 ( .A0(\dataoutbuffer[0][2] ), .A1(n5312), .B0(
        \dataoutbuffer[6][2] ), .B1(n2893), .Y(n5006) );
  AOI22X1TS U5549 ( .A0(\dataoutbuffer[2][2] ), .A1(n5310), .B0(
        \dataoutbuffer[3][2] ), .B1(n2891), .Y(n5005) );
  AOI22X1TS U5550 ( .A0(\dataoutbuffer[4][2] ), .A1(n5295), .B0(
        \dataoutbuffer[5][2] ), .B1(n2892), .Y(n5004) );
  AOI22X1TS U5551 ( .A0(\dataoutbuffer[1][2] ), .A1(n2894), .B0(
        \dataoutbuffer[7][2] ), .B1(n2895), .Y(n5003) );
  NAND4XLTS U5552 ( .A(n5006), .B(n5005), .C(n5004), .D(n5003), .Y(n5007) );
  AOI22X1TS U5553 ( .A0(n5318), .A1(dataOut[2]), .B0(n2890), .B1(n5007), .Y(
        n5008) );
  AOI22X1TS U5554 ( .A0(n3444), .A1(n5304), .B0(n3443), .B1(n2922), .Y(n5021)
         );
  OAI22X1TS U5555 ( .A0(n5012), .A1(n5305), .B0(n5011), .B1(n5307), .Y(n5013)
         );
  AOI21X1TS U5556 ( .A0(n3442), .A1(n2908), .B0(n5013), .Y(n5020) );
  AOI22X1TS U5557 ( .A0(\dataoutbuffer[4][3] ), .A1(n5295), .B0(
        \dataoutbuffer[5][3] ), .B1(n2892), .Y(n5017) );
  AOI22X1TS U5558 ( .A0(\dataoutbuffer[3][3] ), .A1(n2891), .B0(
        \dataoutbuffer[7][3] ), .B1(n2895), .Y(n5016) );
  AOI22X1TS U5559 ( .A0(\dataoutbuffer[0][3] ), .A1(n5312), .B0(
        \dataoutbuffer[1][3] ), .B1(n2894), .Y(n5015) );
  AOI22X1TS U5560 ( .A0(\dataoutbuffer[2][3] ), .A1(n5310), .B0(
        \dataoutbuffer[6][3] ), .B1(n2893), .Y(n5014) );
  NAND4XLTS U5561 ( .A(n5017), .B(n5016), .C(n5015), .D(n5014), .Y(n5018) );
  AOI22X1TS U5562 ( .A0(n5318), .A1(dataOut[3]), .B0(n2890), .B1(n5018), .Y(
        n5019) );
  AOI22X1TS U5563 ( .A0(n3165), .A1(n5304), .B0(n3164), .B1(n2922), .Y(n5032)
         );
  OAI22X1TS U5564 ( .A0(n5023), .A1(n5307), .B0(n5022), .B1(n5305), .Y(n5024)
         );
  AOI21X1TS U5565 ( .A0(n3167), .A1(n2908), .B0(n5024), .Y(n5031) );
  AOI22X1TS U5566 ( .A0(\dataoutbuffer[6][4] ), .A1(n2893), .B0(
        \dataoutbuffer[1][4] ), .B1(n2894), .Y(n5028) );
  AOI22X1TS U5567 ( .A0(\dataoutbuffer[4][4] ), .A1(n5295), .B0(
        \dataoutbuffer[5][4] ), .B1(n2892), .Y(n5027) );
  AOI22X1TS U5568 ( .A0(\dataoutbuffer[2][4] ), .A1(n5310), .B0(
        \dataoutbuffer[3][4] ), .B1(n2891), .Y(n5026) );
  AOI22X1TS U5569 ( .A0(\dataoutbuffer[0][4] ), .A1(n5312), .B0(
        \dataoutbuffer[7][4] ), .B1(n2895), .Y(n5025) );
  NAND4XLTS U5570 ( .A(n5028), .B(n5027), .C(n5026), .D(n5025), .Y(n5029) );
  AOI22X1TS U5571 ( .A0(n5318), .A1(dataOut[4]), .B0(n2890), .B1(n5029), .Y(
        n5030) );
  AOI22X1TS U5572 ( .A0(n3532), .A1(n2908), .B0(n3530), .B1(n5290), .Y(n5042)
         );
  OAI22X1TS U5573 ( .A0(n5033), .A1(n5307), .B0(n3529), .B1(n5291), .Y(n5034)
         );
  AOI21X1TS U5574 ( .A0(n3527), .A1(n2922), .B0(n5034), .Y(n5041) );
  AOI22X1TS U5575 ( .A0(\dataoutbuffer[0][5] ), .A1(n5312), .B0(
        \dataoutbuffer[5][5] ), .B1(n2892), .Y(n5038) );
  AOI22X1TS U5576 ( .A0(\dataoutbuffer[2][5] ), .A1(n5310), .B0(
        \dataoutbuffer[3][5] ), .B1(n2891), .Y(n5037) );
  AOI22X1TS U5577 ( .A0(\dataoutbuffer[4][5] ), .A1(n5295), .B0(
        \dataoutbuffer[6][5] ), .B1(n2893), .Y(n5036) );
  AOI22X1TS U5578 ( .A0(\dataoutbuffer[1][5] ), .A1(n2894), .B0(
        \dataoutbuffer[7][5] ), .B1(n2895), .Y(n5035) );
  NAND4XLTS U5579 ( .A(n5038), .B(n5037), .C(n5036), .D(n5035), .Y(n5039) );
  AOI22X1TS U5580 ( .A0(n5318), .A1(dataOut[5]), .B0(n2890), .B1(n5039), .Y(
        n5040) );
  AOI22X1TS U5581 ( .A0(n3270), .A1(n5280), .B0(n3269), .B1(n2922), .Y(n5053)
         );
  OAI22X1TS U5582 ( .A0(n5044), .A1(n5305), .B0(n5043), .B1(n5291), .Y(n5045)
         );
  AOI21X1TS U5583 ( .A0(n3268), .A1(n2908), .B0(n5045), .Y(n5052) );
  AOI22X1TS U5584 ( .A0(\dataoutbuffer[2][6] ), .A1(n5310), .B0(
        \dataoutbuffer[7][6] ), .B1(n2895), .Y(n5049) );
  AOI22X1TS U5585 ( .A0(\dataoutbuffer[3][6] ), .A1(n2891), .B0(
        \dataoutbuffer[4][6] ), .B1(n5295), .Y(n5048) );
  AOI22X1TS U5586 ( .A0(\dataoutbuffer[0][6] ), .A1(n5312), .B0(
        \dataoutbuffer[5][6] ), .B1(n2892), .Y(n5047) );
  AOI22X1TS U5587 ( .A0(\dataoutbuffer[6][6] ), .A1(n2893), .B0(
        \dataoutbuffer[1][6] ), .B1(n2894), .Y(n5046) );
  NAND4XLTS U5588 ( .A(n5049), .B(n5048), .C(n5047), .D(n5046), .Y(n5050) );
  AOI22X1TS U5589 ( .A0(n5318), .A1(dataOut[6]), .B0(n2890), .B1(n5050), .Y(
        n5051) );
  AOI22X1TS U5590 ( .A0(n3200), .A1(n2908), .B0(n3198), .B1(n2922), .Y(n5064)
         );
  OAI22X1TS U5591 ( .A0(n5055), .A1(n5291), .B0(n5054), .B1(n5305), .Y(n5056)
         );
  AOI21X1TS U5592 ( .A0(n3199), .A1(n5280), .B0(n5056), .Y(n5063) );
  AOI22X1TS U5593 ( .A0(\dataoutbuffer[3][7] ), .A1(n2891), .B0(
        \dataoutbuffer[1][7] ), .B1(n2894), .Y(n5060) );
  AOI22X1TS U5594 ( .A0(\dataoutbuffer[4][7] ), .A1(n5295), .B0(
        \dataoutbuffer[5][7] ), .B1(n2892), .Y(n5059) );
  AOI22X1TS U5595 ( .A0(\dataoutbuffer[0][7] ), .A1(n5312), .B0(
        \dataoutbuffer[6][7] ), .B1(n2893), .Y(n5058) );
  AOI22X1TS U5596 ( .A0(\dataoutbuffer[2][7] ), .A1(n5310), .B0(
        \dataoutbuffer[7][7] ), .B1(n2895), .Y(n5057) );
  NAND4XLTS U5597 ( .A(n5060), .B(n5059), .C(n5058), .D(n5057), .Y(n5061) );
  AOI22X1TS U5598 ( .A0(n5318), .A1(dataOut[7]), .B0(n2890), .B1(n5061), .Y(
        n5062) );
  AOI22X1TS U5599 ( .A0(n3053), .A1(n5290), .B0(n3051), .B1(n5280), .Y(n5073)
         );
  AOI22X1TS U5600 ( .A0(n3055), .A1(n5304), .B0(n3052), .B1(n2922), .Y(n5072)
         );
  AOI22X1TS U5601 ( .A0(\dataoutbuffer[0][8] ), .A1(n5312), .B0(
        \dataoutbuffer[6][8] ), .B1(n2893), .Y(n5068) );
  AOI22X1TS U5602 ( .A0(\dataoutbuffer[2][8] ), .A1(n5310), .B0(
        \dataoutbuffer[5][8] ), .B1(n2892), .Y(n5067) );
  AOI22X1TS U5603 ( .A0(\dataoutbuffer[1][8] ), .A1(n2894), .B0(
        \dataoutbuffer[7][8] ), .B1(n2895), .Y(n5066) );
  AOI22X1TS U5604 ( .A0(\dataoutbuffer[3][8] ), .A1(n2891), .B0(
        \dataoutbuffer[4][8] ), .B1(n5295), .Y(n5065) );
  NAND4XLTS U5605 ( .A(n5068), .B(n5067), .C(n5066), .D(n5065), .Y(n5069) );
  AOI22X1TS U5606 ( .A0(n5318), .A1(dataOut[8]), .B0(n2890), .B1(n5069), .Y(
        n5071) );
  NAND2X1TS U5607 ( .A(n3054), .B(n2908), .Y(n5070) );
  AOI22X1TS U5608 ( .A0(n3062), .A1(n5290), .B0(n3063), .B1(n2908), .Y(n5084)
         );
  OAI22X1TS U5609 ( .A0(n5075), .A1(n5291), .B0(n5074), .B1(n5307), .Y(n5076)
         );
  AOI21X1TS U5610 ( .A0(n3061), .A1(n2922), .B0(n5076), .Y(n5083) );
  AOI22X1TS U5611 ( .A0(\dataoutbuffer[0][9] ), .A1(n5312), .B0(
        \dataoutbuffer[7][9] ), .B1(n2895), .Y(n5080) );
  AOI22X1TS U5612 ( .A0(\dataoutbuffer[4][9] ), .A1(n5295), .B0(
        \dataoutbuffer[6][9] ), .B1(n2893), .Y(n5079) );
  AOI22X1TS U5613 ( .A0(\dataoutbuffer[3][9] ), .A1(n2891), .B0(
        \dataoutbuffer[5][9] ), .B1(n2892), .Y(n5078) );
  AOI22X1TS U5614 ( .A0(\dataoutbuffer[2][9] ), .A1(n5310), .B0(
        \dataoutbuffer[1][9] ), .B1(n2894), .Y(n5077) );
  NAND4XLTS U5615 ( .A(n5080), .B(n5079), .C(n5078), .D(n5077), .Y(n5081) );
  AOI22X1TS U5616 ( .A0(n5318), .A1(dataOut[9]), .B0(n2890), .B1(n5081), .Y(
        n5082) );
  AOI22X1TS U5617 ( .A0(n3154), .A1(n5290), .B0(n3155), .B1(n2922), .Y(n5095)
         );
  OAI22X1TS U5618 ( .A0(n5086), .A1(n5291), .B0(n5085), .B1(n5307), .Y(n5087)
         );
  AOI21X1TS U5619 ( .A0(n3156), .A1(n2908), .B0(n5087), .Y(n5094) );
  AOI22X1TS U5620 ( .A0(\dataoutbuffer[1][10] ), .A1(n2894), .B0(
        \dataoutbuffer[7][10] ), .B1(n2895), .Y(n5091) );
  AOI22X1TS U5621 ( .A0(\dataoutbuffer[0][10] ), .A1(n5312), .B0(
        \dataoutbuffer[2][10] ), .B1(n5310), .Y(n5090) );
  AOI22X1TS U5622 ( .A0(\dataoutbuffer[3][10] ), .A1(n2891), .B0(
        \dataoutbuffer[4][10] ), .B1(n5295), .Y(n5089) );
  AOI22X1TS U5623 ( .A0(\dataoutbuffer[6][10] ), .A1(n2893), .B0(
        \dataoutbuffer[5][10] ), .B1(n2892), .Y(n5088) );
  NAND4XLTS U5624 ( .A(n5091), .B(n5090), .C(n5089), .D(n5088), .Y(n5092) );
  AOI22X1TS U5625 ( .A0(n5318), .A1(dataOut[10]), .B0(n2890), .B1(n5092), .Y(
        n5093) );
  AOI22X1TS U5626 ( .A0(n3366), .A1(n5280), .B0(n3364), .B1(n5304), .Y(n5104)
         );
  AOI22X1TS U5627 ( .A0(n3367), .A1(n5290), .B0(n3363), .B1(n2922), .Y(n5103)
         );
  AOI22X1TS U5628 ( .A0(\dataoutbuffer[2][11] ), .A1(n5310), .B0(
        \dataoutbuffer[6][11] ), .B1(n2893), .Y(n5099) );
  AOI22X1TS U5629 ( .A0(\dataoutbuffer[3][11] ), .A1(n2891), .B0(
        \dataoutbuffer[4][11] ), .B1(n5295), .Y(n5098) );
  AOI22X1TS U5630 ( .A0(\dataoutbuffer[5][11] ), .A1(n2892), .B0(
        \dataoutbuffer[7][11] ), .B1(n2895), .Y(n5097) );
  AOI22X1TS U5631 ( .A0(\dataoutbuffer[0][11] ), .A1(n5312), .B0(
        \dataoutbuffer[1][11] ), .B1(n2894), .Y(n5096) );
  NAND4XLTS U5632 ( .A(n5099), .B(n5098), .C(n5097), .D(n5096), .Y(n5100) );
  AOI22X1TS U5633 ( .A0(n5318), .A1(dataOut[11]), .B0(n2890), .B1(n5100), .Y(
        n5102) );
  NAND2X1TS U5634 ( .A(n3362), .B(n2908), .Y(n5101) );
  AOI22X1TS U5635 ( .A0(n3277), .A1(n5280), .B0(n3282), .B1(n5304), .Y(n5113)
         );
  AOI22X1TS U5636 ( .A0(n3281), .A1(n5290), .B0(n3278), .B1(n2922), .Y(n5112)
         );
  AOI22X1TS U5637 ( .A0(\dataoutbuffer[6][12] ), .A1(n2893), .B0(
        \dataoutbuffer[1][12] ), .B1(n2894), .Y(n5108) );
  AOI22X1TS U5638 ( .A0(\dataoutbuffer[0][12] ), .A1(n5312), .B0(
        \dataoutbuffer[5][12] ), .B1(n2892), .Y(n5107) );
  AOI22X1TS U5639 ( .A0(\dataoutbuffer[3][12] ), .A1(n2891), .B0(
        \dataoutbuffer[4][12] ), .B1(n5295), .Y(n5106) );
  AOI22X1TS U5640 ( .A0(\dataoutbuffer[2][12] ), .A1(n5310), .B0(
        \dataoutbuffer[7][12] ), .B1(n2895), .Y(n5105) );
  NAND4XLTS U5641 ( .A(n5108), .B(n5107), .C(n5106), .D(n5105), .Y(n5109) );
  AOI22X1TS U5642 ( .A0(n5318), .A1(dataOut[12]), .B0(n2890), .B1(n5109), .Y(
        n5111) );
  NAND2X1TS U5643 ( .A(n3279), .B(n2908), .Y(n5110) );
  AOI22X1TS U5644 ( .A0(n2962), .A1(n5304), .B0(n2965), .B1(n5290), .Y(n5122)
         );
  AOI22X1TS U5645 ( .A0(n2967), .A1(n2908), .B0(n2964), .B1(n2922), .Y(n5121)
         );
  AOI22X1TS U5646 ( .A0(\dataoutbuffer[0][13] ), .A1(n5312), .B0(
        \dataoutbuffer[1][13] ), .B1(n2894), .Y(n5117) );
  AOI22X1TS U5647 ( .A0(\dataoutbuffer[6][13] ), .A1(n2893), .B0(
        \dataoutbuffer[5][13] ), .B1(n2892), .Y(n5116) );
  AOI22X1TS U5648 ( .A0(\dataoutbuffer[2][13] ), .A1(n5310), .B0(
        \dataoutbuffer[3][13] ), .B1(n2891), .Y(n5115) );
  AOI22X1TS U5649 ( .A0(\dataoutbuffer[4][13] ), .A1(n5295), .B0(
        \dataoutbuffer[7][13] ), .B1(n2895), .Y(n5114) );
  NAND4XLTS U5650 ( .A(n5117), .B(n5116), .C(n5115), .D(n5114), .Y(n5118) );
  AOI22X1TS U5651 ( .A0(n5318), .A1(dataOut[13]), .B0(n2890), .B1(n5118), .Y(
        n5120) );
  NAND2X1TS U5652 ( .A(n2968), .B(n5280), .Y(n5119) );
  AOI22X1TS U5653 ( .A0(n3356), .A1(n2908), .B0(n3354), .B1(n2922), .Y(n5133)
         );
  OAI22X1TS U5654 ( .A0(n5124), .A1(n5307), .B0(n5123), .B1(n5305), .Y(n5125)
         );
  AOI21X1TS U5655 ( .A0(n3355), .A1(n5304), .B0(n5125), .Y(n5132) );
  AOI22X1TS U5656 ( .A0(\dataoutbuffer[4][14] ), .A1(n5295), .B0(
        \dataoutbuffer[7][14] ), .B1(n2895), .Y(n5129) );
  AOI22X1TS U5657 ( .A0(\dataoutbuffer[3][14] ), .A1(n2891), .B0(
        \dataoutbuffer[6][14] ), .B1(n2893), .Y(n5128) );
  AOI22X1TS U5658 ( .A0(\dataoutbuffer[0][14] ), .A1(n5312), .B0(
        \dataoutbuffer[1][14] ), .B1(n2894), .Y(n5127) );
  AOI22X1TS U5659 ( .A0(\dataoutbuffer[2][14] ), .A1(n5310), .B0(
        \dataoutbuffer[5][14] ), .B1(n2892), .Y(n5126) );
  NAND4XLTS U5660 ( .A(n5129), .B(n5128), .C(n5127), .D(n5126), .Y(n5130) );
  AOI22X1TS U5661 ( .A0(n5318), .A1(dataOut[14]), .B0(n2890), .B1(n5130), .Y(
        n5131) );
  AOI22X1TS U5662 ( .A0(n3345), .A1(n5290), .B0(n3342), .B1(n2922), .Y(n5144)
         );
  OAI22X1TS U5663 ( .A0(n5135), .A1(n5307), .B0(n5134), .B1(n5291), .Y(n5136)
         );
  AOI21X1TS U5664 ( .A0(n3344), .A1(n2908), .B0(n5136), .Y(n5143) );
  AOI22X1TS U5665 ( .A0(\dataoutbuffer[4][15] ), .A1(n5295), .B0(
        \dataoutbuffer[6][15] ), .B1(n2893), .Y(n5140) );
  AOI22X1TS U5666 ( .A0(\dataoutbuffer[0][15] ), .A1(n5312), .B0(
        \dataoutbuffer[1][15] ), .B1(n2894), .Y(n5139) );
  AOI22X1TS U5667 ( .A0(\dataoutbuffer[2][15] ), .A1(n5310), .B0(
        \dataoutbuffer[3][15] ), .B1(n2891), .Y(n5138) );
  AOI22X1TS U5668 ( .A0(\dataoutbuffer[5][15] ), .A1(n2892), .B0(
        \dataoutbuffer[7][15] ), .B1(n2895), .Y(n5137) );
  NAND4XLTS U5669 ( .A(n5140), .B(n5139), .C(n5138), .D(n5137), .Y(n5141) );
  AOI22X1TS U5670 ( .A0(n5318), .A1(dataOut[15]), .B0(n2890), .B1(n5141), .Y(
        n5142) );
  AOI22X1TS U5671 ( .A0(n3044), .A1(n5290), .B0(n3043), .B1(n2922), .Y(n5155)
         );
  OAI22X1TS U5672 ( .A0(n5146), .A1(n5291), .B0(n5145), .B1(n5307), .Y(n5147)
         );
  AOI21X1TS U5673 ( .A0(n3046), .A1(n2908), .B0(n5147), .Y(n5154) );
  AOI22X1TS U5674 ( .A0(\dataoutbuffer[2][16] ), .A1(n5310), .B0(
        \dataoutbuffer[1][16] ), .B1(n2894), .Y(n5151) );
  AOI22X1TS U5675 ( .A0(\dataoutbuffer[5][16] ), .A1(n2892), .B0(
        \dataoutbuffer[7][16] ), .B1(n2895), .Y(n5150) );
  AOI22X1TS U5676 ( .A0(\dataoutbuffer[0][16] ), .A1(n5312), .B0(
        \dataoutbuffer[6][16] ), .B1(n2893), .Y(n5149) );
  AOI22X1TS U5677 ( .A0(\dataoutbuffer[3][16] ), .A1(n2891), .B0(
        \dataoutbuffer[4][16] ), .B1(n5295), .Y(n5148) );
  NAND4XLTS U5678 ( .A(n5151), .B(n5150), .C(n5149), .D(n5148), .Y(n5152) );
  AOI22X1TS U5679 ( .A0(n5318), .A1(dataOut[16]), .B0(n2890), .B1(n5152), .Y(
        n5153) );
  AOI22X1TS U5680 ( .A0(n3211), .A1(n5304), .B0(n3207), .B1(n2922), .Y(n5165)
         );
  OAI22X1TS U5681 ( .A0(n3209), .A1(n5307), .B0(n5156), .B1(n5305), .Y(n5157)
         );
  AOI21X1TS U5682 ( .A0(n3210), .A1(n2908), .B0(n5157), .Y(n5164) );
  AOI22X1TS U5683 ( .A0(\dataoutbuffer[4][17] ), .A1(n5295), .B0(
        \dataoutbuffer[6][17] ), .B1(n2893), .Y(n5161) );
  AOI22X1TS U5684 ( .A0(\dataoutbuffer[2][17] ), .A1(n5310), .B0(
        \dataoutbuffer[5][17] ), .B1(n2892), .Y(n5160) );
  AOI22X1TS U5685 ( .A0(\dataoutbuffer[0][17] ), .A1(n5312), .B0(
        \dataoutbuffer[7][17] ), .B1(n2895), .Y(n5159) );
  AOI22X1TS U5686 ( .A0(\dataoutbuffer[3][17] ), .A1(n2891), .B0(
        \dataoutbuffer[1][17] ), .B1(n2894), .Y(n5158) );
  NAND4XLTS U5687 ( .A(n5161), .B(n5160), .C(n5159), .D(n5158), .Y(n5162) );
  AOI22X1TS U5688 ( .A0(n5318), .A1(dataOut[17]), .B0(n2890), .B1(n5162), .Y(
        n5163) );
  AOI22X1TS U5689 ( .A0(n3405), .A1(n2908), .B0(n3407), .B1(n2922), .Y(n5175)
         );
  OAI22X1TS U5690 ( .A0(n3409), .A1(n5305), .B0(n5166), .B1(n5291), .Y(n5167)
         );
  AOI21X1TS U5691 ( .A0(n3410), .A1(n5280), .B0(n5167), .Y(n5174) );
  AOI22X1TS U5692 ( .A0(\dataoutbuffer[6][18] ), .A1(n2893), .B0(
        \dataoutbuffer[1][18] ), .B1(n2894), .Y(n5171) );
  AOI22X1TS U5693 ( .A0(\dataoutbuffer[2][18] ), .A1(n5310), .B0(
        \dataoutbuffer[3][18] ), .B1(n2891), .Y(n5170) );
  AOI22X1TS U5694 ( .A0(\dataoutbuffer[0][18] ), .A1(n5312), .B0(
        \dataoutbuffer[5][18] ), .B1(n2892), .Y(n5169) );
  AOI22X1TS U5695 ( .A0(\dataoutbuffer[4][18] ), .A1(n5295), .B0(
        \dataoutbuffer[7][18] ), .B1(n2895), .Y(n5168) );
  NAND4XLTS U5696 ( .A(n5171), .B(n5170), .C(n5169), .D(n5168), .Y(n5172) );
  AOI22X1TS U5697 ( .A0(n5318), .A1(dataOut[18]), .B0(n2890), .B1(n5172), .Y(
        n5173) );
  AOI22X1TS U5698 ( .A0(n3261), .A1(n2908), .B0(n3263), .B1(n5290), .Y(n5186)
         );
  OAI22X1TS U5699 ( .A0(n5177), .A1(n5307), .B0(n5176), .B1(n5291), .Y(n5178)
         );
  AOI21X1TS U5700 ( .A0(n3260), .A1(n2922), .B0(n5178), .Y(n5185) );
  AOI22X1TS U5701 ( .A0(\dataoutbuffer[3][19] ), .A1(n2891), .B0(
        \dataoutbuffer[7][19] ), .B1(n2895), .Y(n5182) );
  AOI22X1TS U5702 ( .A0(\dataoutbuffer[1][19] ), .A1(n2894), .B0(
        \dataoutbuffer[5][19] ), .B1(n2892), .Y(n5181) );
  AOI22X1TS U5703 ( .A0(\dataoutbuffer[0][19] ), .A1(n5312), .B0(
        \dataoutbuffer[6][19] ), .B1(n2893), .Y(n5180) );
  AOI22X1TS U5704 ( .A0(\dataoutbuffer[2][19] ), .A1(n5310), .B0(
        \dataoutbuffer[4][19] ), .B1(n5295), .Y(n5179) );
  NAND4XLTS U5705 ( .A(n5182), .B(n5181), .C(n5180), .D(n5179), .Y(n5183) );
  AOI22X1TS U5706 ( .A0(n5318), .A1(dataOut[19]), .B0(n2890), .B1(n5183), .Y(
        n5184) );
  AOI22X1TS U5707 ( .A0(n3247), .A1(n5290), .B0(n3244), .B1(n2922), .Y(n5197)
         );
  OAI22X1TS U5708 ( .A0(n5188), .A1(n5307), .B0(n5187), .B1(n5291), .Y(n5189)
         );
  AOI21X1TS U5709 ( .A0(n3245), .A1(n2908), .B0(n5189), .Y(n5196) );
  AOI22X1TS U5710 ( .A0(\dataoutbuffer[0][20] ), .A1(n5312), .B0(
        \dataoutbuffer[3][20] ), .B1(n2891), .Y(n5193) );
  AOI22X1TS U5711 ( .A0(\dataoutbuffer[2][20] ), .A1(n5310), .B0(
        \dataoutbuffer[4][20] ), .B1(n5295), .Y(n5192) );
  AOI22X1TS U5712 ( .A0(\dataoutbuffer[1][20] ), .A1(n2894), .B0(
        \dataoutbuffer[7][20] ), .B1(n2895), .Y(n5191) );
  AOI22X1TS U5713 ( .A0(\dataoutbuffer[6][20] ), .A1(n2893), .B0(
        \dataoutbuffer[5][20] ), .B1(n2892), .Y(n5190) );
  NAND4XLTS U5714 ( .A(n5193), .B(n5192), .C(n5191), .D(n5190), .Y(n5194) );
  AOI22X1TS U5715 ( .A0(n5318), .A1(dataOut[20]), .B0(n2890), .B1(n5194), .Y(
        n5195) );
  AOI22X1TS U5716 ( .A0(n3291), .A1(n5304), .B0(n3290), .B1(n5290), .Y(n5206)
         );
  AOI22X1TS U5717 ( .A0(n3286), .A1(n5280), .B0(n3287), .B1(n2922), .Y(n5205)
         );
  AOI22X1TS U5718 ( .A0(\dataoutbuffer[0][21] ), .A1(n5312), .B0(
        \dataoutbuffer[7][21] ), .B1(n2895), .Y(n5201) );
  AOI22X1TS U5719 ( .A0(\dataoutbuffer[3][21] ), .A1(n2891), .B0(
        \dataoutbuffer[4][21] ), .B1(n5295), .Y(n5200) );
  AOI22X1TS U5720 ( .A0(\dataoutbuffer[6][21] ), .A1(n2893), .B0(
        \dataoutbuffer[5][21] ), .B1(n2892), .Y(n5199) );
  AOI22X1TS U5721 ( .A0(\dataoutbuffer[2][21] ), .A1(n5310), .B0(
        \dataoutbuffer[1][21] ), .B1(n2894), .Y(n5198) );
  NAND4XLTS U5722 ( .A(n5201), .B(n5200), .C(n5199), .D(n5198), .Y(n5202) );
  AOI22X1TS U5723 ( .A0(n5318), .A1(dataOut[21]), .B0(n2890), .B1(n5202), .Y(
        n5204) );
  NAND2X1TS U5724 ( .A(n3288), .B(n2908), .Y(n5203) );
  AOI22X1TS U5725 ( .A0(n3480), .A1(n2908), .B0(n3481), .B1(n2922), .Y(n5216)
         );
  OAI22X1TS U5726 ( .A0(n5207), .A1(n5291), .B0(n3484), .B1(n5305), .Y(n5208)
         );
  AOI21X1TS U5727 ( .A0(n3485), .A1(n5280), .B0(n5208), .Y(n5215) );
  AOI22X1TS U5728 ( .A0(\dataoutbuffer[2][22] ), .A1(n5310), .B0(
        \dataoutbuffer[6][22] ), .B1(n5311), .Y(n5212) );
  AOI22X1TS U5729 ( .A0(\dataoutbuffer[1][22] ), .A1(n2894), .B0(
        \dataoutbuffer[5][22] ), .B1(n2892), .Y(n5211) );
  AOI22X1TS U5730 ( .A0(\dataoutbuffer[3][22] ), .A1(n2891), .B0(
        \dataoutbuffer[4][22] ), .B1(n5295), .Y(n5210) );
  AOI22X1TS U5731 ( .A0(\dataoutbuffer[0][22] ), .A1(n5312), .B0(
        \dataoutbuffer[7][22] ), .B1(n2895), .Y(n5209) );
  NAND4XLTS U5732 ( .A(n5212), .B(n5211), .C(n5210), .D(n5209), .Y(n5213) );
  AOI22X1TS U5733 ( .A0(n5318), .A1(dataOut[22]), .B0(n2890), .B1(n5213), .Y(
        n5214) );
  AOI22X1TS U5734 ( .A0(n2957), .A1(n5304), .B0(n2950), .B1(n2922), .Y(n5226)
         );
  OAI22X1TS U5735 ( .A0(n2954), .A1(n5305), .B0(n5217), .B1(n5307), .Y(n5218)
         );
  AOI21X1TS U5736 ( .A0(n2949), .A1(n2908), .B0(n5218), .Y(n5225) );
  AOI22X1TS U5737 ( .A0(\dataoutbuffer[0][23] ), .A1(n5312), .B0(
        \dataoutbuffer[3][23] ), .B1(n2891), .Y(n5222) );
  AOI22X1TS U5738 ( .A0(\dataoutbuffer[2][23] ), .A1(n5310), .B0(
        \dataoutbuffer[7][23] ), .B1(n2895), .Y(n5221) );
  AOI22X1TS U5739 ( .A0(\dataoutbuffer[4][23] ), .A1(n5295), .B0(
        \dataoutbuffer[5][23] ), .B1(n2892), .Y(n5220) );
  AOI22X1TS U5740 ( .A0(\dataoutbuffer[6][23] ), .A1(n2893), .B0(
        \dataoutbuffer[1][23] ), .B1(n2894), .Y(n5219) );
  NAND4XLTS U5741 ( .A(n5222), .B(n5221), .C(n5220), .D(n5219), .Y(n5223) );
  AOI22X1TS U5742 ( .A0(n5318), .A1(dataOut[23]), .B0(n2890), .B1(n5223), .Y(
        n5224) );
  AOI22X1TS U5743 ( .A0(n3149), .A1(n5304), .B0(n3146), .B1(n2922), .Y(n5237)
         );
  OAI22X1TS U5744 ( .A0(n5228), .A1(n5305), .B0(n5227), .B1(n5307), .Y(n5229)
         );
  AOI21X1TS U5745 ( .A0(n3147), .A1(n2908), .B0(n5229), .Y(n5236) );
  AOI22X1TS U5746 ( .A0(\dataoutbuffer[2][24] ), .A1(n5310), .B0(
        \dataoutbuffer[6][24] ), .B1(n5311), .Y(n5233) );
  AOI22X1TS U5747 ( .A0(\dataoutbuffer[3][24] ), .A1(n2891), .B0(
        \dataoutbuffer[5][24] ), .B1(n2892), .Y(n5232) );
  AOI22X1TS U5748 ( .A0(\dataoutbuffer[0][24] ), .A1(n5312), .B0(
        \dataoutbuffer[7][24] ), .B1(n2895), .Y(n5231) );
  AOI22X1TS U5749 ( .A0(\dataoutbuffer[4][24] ), .A1(n5295), .B0(
        \dataoutbuffer[1][24] ), .B1(n2894), .Y(n5230) );
  NAND4XLTS U5750 ( .A(n5233), .B(n5232), .C(n5231), .D(n5230), .Y(n5234) );
  AOI22X1TS U5751 ( .A0(n5318), .A1(dataOut[24]), .B0(n2890), .B1(n5234), .Y(
        n5235) );
  AOI22X1TS U5752 ( .A0(n3235), .A1(n5304), .B0(n3230), .B1(n2922), .Y(n5248)
         );
  OAI22X1TS U5753 ( .A0(n5239), .A1(n5307), .B0(n5238), .B1(n5305), .Y(n5240)
         );
  AOI21X1TS U5754 ( .A0(n3229), .A1(n2908), .B0(n5240), .Y(n5247) );
  AOI22X1TS U5755 ( .A0(\dataoutbuffer[6][25] ), .A1(n2893), .B0(
        \dataoutbuffer[5][25] ), .B1(n2892), .Y(n5244) );
  AOI22X1TS U5756 ( .A0(\dataoutbuffer[4][25] ), .A1(n5295), .B0(
        \dataoutbuffer[1][25] ), .B1(n2894), .Y(n5243) );
  AOI22X1TS U5757 ( .A0(\dataoutbuffer[0][25] ), .A1(n5312), .B0(
        \dataoutbuffer[7][25] ), .B1(n2895), .Y(n5242) );
  AOI22X1TS U5758 ( .A0(\dataoutbuffer[2][25] ), .A1(n5310), .B0(
        \dataoutbuffer[3][25] ), .B1(n2891), .Y(n5241) );
  NAND4XLTS U5759 ( .A(n5244), .B(n5243), .C(n5242), .D(n5241), .Y(n5245) );
  AOI22X1TS U5760 ( .A0(n5318), .A1(dataOut[25]), .B0(n2890), .B1(n5245), .Y(
        n5246) );
  AOI22X1TS U5761 ( .A0(n3429), .A1(n5304), .B0(n3431), .B1(n5290), .Y(n5258)
         );
  AOI22X1TS U5762 ( .A0(n3427), .A1(n2908), .B0(n3428), .B1(n2922), .Y(n5257)
         );
  AOI22X1TS U5763 ( .A0(\dataoutbuffer[3][26] ), .A1(n2891), .B0(
        \dataoutbuffer[1][26] ), .B1(n2894), .Y(n5253) );
  AOI22X1TS U5764 ( .A0(\dataoutbuffer[0][26] ), .A1(n5312), .B0(
        \dataoutbuffer[6][26] ), .B1(n2893), .Y(n5252) );
  AOI22X1TS U5765 ( .A0(\dataoutbuffer[2][26] ), .A1(n5310), .B0(
        \dataoutbuffer[7][26] ), .B1(n2895), .Y(n5251) );
  AOI22X1TS U5766 ( .A0(\dataoutbuffer[4][26] ), .A1(n5249), .B0(
        \dataoutbuffer[5][26] ), .B1(n2892), .Y(n5250) );
  NAND4XLTS U5767 ( .A(n5253), .B(n5252), .C(n5251), .D(n5250), .Y(n5254) );
  AOI22X1TS U5768 ( .A0(n5318), .A1(dataOut[26]), .B0(n2890), .B1(n5254), .Y(
        n5256) );
  NAND2X1TS U5769 ( .A(n3432), .B(n5280), .Y(n5255) );
  AOI22X1TS U5770 ( .A0(n3300), .A1(n5290), .B0(n3297), .B1(n2922), .Y(n5269)
         );
  OAI22X1TS U5771 ( .A0(n5260), .A1(n5291), .B0(n5259), .B1(n5307), .Y(n5261)
         );
  AOI21X1TS U5772 ( .A0(n3298), .A1(n2908), .B0(n5261), .Y(n5268) );
  AOI22X1TS U5773 ( .A0(\dataoutbuffer[0][27] ), .A1(n5312), .B0(
        \dataoutbuffer[2][27] ), .B1(n5310), .Y(n5265) );
  AOI22X1TS U5774 ( .A0(\dataoutbuffer[3][27] ), .A1(n2891), .B0(
        \dataoutbuffer[7][27] ), .B1(n2895), .Y(n5264) );
  AOI22X1TS U5775 ( .A0(\dataoutbuffer[4][27] ), .A1(n5295), .B0(
        \dataoutbuffer[6][27] ), .B1(n2893), .Y(n5263) );
  AOI22X1TS U5776 ( .A0(\dataoutbuffer[1][27] ), .A1(n2894), .B0(
        \dataoutbuffer[5][27] ), .B1(n2892), .Y(n5262) );
  NAND4XLTS U5777 ( .A(n5265), .B(n5264), .C(n5263), .D(n5262), .Y(n5266) );
  AOI22X1TS U5778 ( .A0(n5318), .A1(dataOut[27]), .B0(n2890), .B1(n5266), .Y(
        n5267) );
  AOI22X1TS U5779 ( .A0(n3398), .A1(n5290), .B0(n3397), .B1(n2922), .Y(n5279)
         );
  OAI22X1TS U5780 ( .A0(n5270), .A1(n5307), .B0(n3401), .B1(n5291), .Y(n5271)
         );
  AOI21X1TS U5781 ( .A0(n3396), .A1(n2908), .B0(n5271), .Y(n5278) );
  AOI22X1TS U5782 ( .A0(\dataoutbuffer[0][28] ), .A1(n5312), .B0(
        \dataoutbuffer[5][28] ), .B1(n2892), .Y(n5275) );
  AOI22X1TS U5783 ( .A0(\dataoutbuffer[3][28] ), .A1(n2891), .B0(
        \dataoutbuffer[7][28] ), .B1(n2895), .Y(n5274) );
  AOI22X1TS U5784 ( .A0(\dataoutbuffer[2][28] ), .A1(n5310), .B0(
        \dataoutbuffer[6][28] ), .B1(n2893), .Y(n5273) );
  AOI22X1TS U5785 ( .A0(\dataoutbuffer[4][28] ), .A1(n5295), .B0(
        \dataoutbuffer[1][28] ), .B1(n2894), .Y(n5272) );
  NAND4XLTS U5786 ( .A(n5275), .B(n5274), .C(n5273), .D(n5272), .Y(n5276) );
  AOI22X1TS U5787 ( .A0(n5318), .A1(dataOut[28]), .B0(n2890), .B1(n5276), .Y(
        n5277) );
  AOI22X1TS U5788 ( .A0(n3126), .A1(n5290), .B0(n3132), .B1(n5280), .Y(n5289)
         );
  AOI22X1TS U5789 ( .A0(n3129), .A1(n5304), .B0(n3128), .B1(n2922), .Y(n5288)
         );
  AOI22X1TS U5790 ( .A0(\dataoutbuffer[0][29] ), .A1(n5312), .B0(
        \dataoutbuffer[4][29] ), .B1(n5295), .Y(n5284) );
  AOI22X1TS U5791 ( .A0(\dataoutbuffer[6][29] ), .A1(n2893), .B0(
        \dataoutbuffer[5][29] ), .B1(n2892), .Y(n5283) );
  AOI22X1TS U5792 ( .A0(\dataoutbuffer[3][29] ), .A1(n2891), .B0(
        \dataoutbuffer[1][29] ), .B1(n2894), .Y(n5282) );
  AOI22X1TS U5793 ( .A0(\dataoutbuffer[2][29] ), .A1(n5310), .B0(
        \dataoutbuffer[7][29] ), .B1(n2895), .Y(n5281) );
  NAND4XLTS U5794 ( .A(n5284), .B(n5283), .C(n5282), .D(n5281), .Y(n5285) );
  AOI22X1TS U5795 ( .A0(n5318), .A1(dataOut[29]), .B0(n2890), .B1(n5285), .Y(
        n5287) );
  NAND2X1TS U5796 ( .A(n3131), .B(n2908), .Y(n5286) );
  AOI22X1TS U5797 ( .A0(n3461), .A1(n2908), .B0(n3459), .B1(n5290), .Y(n5303)
         );
  OAI22X1TS U5798 ( .A0(n5293), .A1(n5307), .B0(n5292), .B1(n5291), .Y(n5294)
         );
  AOI21X1TS U5799 ( .A0(n3457), .A1(n2922), .B0(n5294), .Y(n5302) );
  AOI22X1TS U5800 ( .A0(\dataoutbuffer[3][30] ), .A1(n2891), .B0(
        \dataoutbuffer[1][30] ), .B1(n2894), .Y(n5299) );
  AOI22X1TS U5801 ( .A0(\dataoutbuffer[0][30] ), .A1(n5312), .B0(
        \dataoutbuffer[6][30] ), .B1(n5311), .Y(n5298) );
  AOI22X1TS U5802 ( .A0(\dataoutbuffer[2][30] ), .A1(n5310), .B0(
        \dataoutbuffer[5][30] ), .B1(n2892), .Y(n5297) );
  AOI22X1TS U5803 ( .A0(\dataoutbuffer[4][30] ), .A1(n5295), .B0(
        \dataoutbuffer[7][30] ), .B1(n2895), .Y(n5296) );
  NAND4XLTS U5804 ( .A(n5299), .B(n5298), .C(n5297), .D(n5296), .Y(n5300) );
  AOI22X1TS U5805 ( .A0(n5318), .A1(dataOut[30]), .B0(n2890), .B1(n5300), .Y(
        n5301) );
  AOI22X1TS U5806 ( .A0(n3138), .A1(n5304), .B0(n3139), .B1(n2908), .Y(n5321)
         );
  OAI22X1TS U5807 ( .A0(n5308), .A1(n5307), .B0(n5306), .B1(n5305), .Y(n5309)
         );
  AOI21X1TS U5808 ( .A0(n3137), .A1(n2922), .B0(n5309), .Y(n5320) );
  AOI22X1TS U5809 ( .A0(\dataoutbuffer[2][31] ), .A1(n5310), .B0(
        \dataoutbuffer[1][31] ), .B1(n2894), .Y(n5316) );
  AOI22X1TS U5810 ( .A0(\dataoutbuffer[5][31] ), .A1(n2892), .B0(
        \dataoutbuffer[7][31] ), .B1(n2895), .Y(n5315) );
  AOI22X1TS U5811 ( .A0(\dataoutbuffer[3][31] ), .A1(n2891), .B0(
        \dataoutbuffer[6][31] ), .B1(n5311), .Y(n5314) );
  AOI22X1TS U5812 ( .A0(\dataoutbuffer[0][31] ), .A1(n5312), .B0(
        \dataoutbuffer[4][31] ), .B1(n5295), .Y(n5313) );
  NAND4XLTS U5813 ( .A(n5316), .B(n5315), .C(n5314), .D(n5313), .Y(n5317) );
  AOI22X1TS U5814 ( .A0(n5318), .A1(dataOut[31]), .B0(n2890), .B1(n5317), .Y(
        n5319) );
endmodule

