
module incomingPortHandler_0 ( clk, reset, localRouterAddress, 
        destinationAddressIn, requesterAddressIn, readIn, writeIn, 
        outputPortSelect, memRead, memWrite );
  input [5:0] localRouterAddress;
  input [13:0] destinationAddressIn;
  input [5:0] requesterAddressIn;
  output [3:0] outputPortSelect;
  input clk, reset, readIn, writeIn;
  output memRead, memWrite;
  wire   n45, n44, n43, n42, n1, n2, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n3;

  DFFQX1TS memWrite_reg ( .D(n1), .CK(clk), .Q(memWrite) );
  DFFQX1TS memRead_reg ( .D(n2), .CK(clk), .Q(memRead) );
  DFFHQX4TS \outputPortSelect_reg[2]  ( .D(n44), .CK(clk), .Q(
        outputPortSelect[2]) );
  DFFQX1TS \outputPortSelect_reg[0]  ( .D(n42), .CK(clk), .Q(
        outputPortSelect[0]) );
  DFFQX1TS \outputPortSelect_reg[3]  ( .D(n45), .CK(clk), .Q(
        outputPortSelect[3]) );
  DFFHQX1TS \outputPortSelect_reg[1]  ( .D(n43), .CK(clk), .Q(
        outputPortSelect[1]) );
  OAI211X1TS U1 ( .A0(localRouterAddress[4]), .A1(n9), .B0(n10), .C0(
        localRouterAddress[3]), .Y(n28) );
  INVXLTS U2 ( .A(destinationAddressIn[13]), .Y(n8) );
  NOR3BXLTS U3 ( .AN(n3), .B(writeIn), .C(readIn), .Y(n14) );
  NAND2XLTS U4 ( .A(localRouterAddress[2]), .B(n11), .Y(n19) );
  AOI2BB2XLTS U5 ( .B0(n12), .B1(localRouterAddress[1]), .A0N(
        destinationAddressIn[8]), .A1N(n7), .Y(n17) );
  INVX2TS U6 ( .A(reset), .Y(n3) );
  NOR2BX1TS U7 ( .AN(n15), .B(n16), .Y(n45) );
  NOR2X1TS U8 ( .A(n16), .B(n15), .Y(n44) );
  INVX2TS U9 ( .A(n22), .Y(n4) );
  OAI21X1TS U10 ( .A0(n17), .A1(n18), .B0(n19), .Y(n15) );
  NAND3BX1TS U11 ( .AN(n20), .B(n21), .C(n22), .Y(n16) );
  OAI22XLTS U12 ( .A0(localRouterAddress[1]), .A1(n12), .B0(
        localRouterAddress[2]), .B1(n11), .Y(n18) );
  AOI2BB1XLTS U13 ( .A0N(localRouterAddress[4]), .A1N(n9), .B0(n29), .Y(n23)
         );
  NAND3X1TS U14 ( .A(n17), .B(n21), .C(n31), .Y(n22) );
  AOI211XLTS U15 ( .A0(destinationAddressIn[8]), .A1(n7), .B0(n18), .C0(n6), 
        .Y(n31) );
  INVX2TS U16 ( .A(n19), .Y(n6) );
  AND4X1TS U17 ( .A(n32), .B(n23), .C(n26), .D(n25), .Y(n21) );
  XNOR2XLTS U18 ( .A(destinationAddressIn[11]), .B(localRouterAddress[3]), .Y(
        n32) );
  INVXLTS U19 ( .A(destinationAddressIn[10]), .Y(n11) );
  INVXLTS U20 ( .A(destinationAddressIn[12]), .Y(n9) );
  INVX2TS U21 ( .A(n13), .Y(n2) );
  AOI32XLTS U22 ( .A0(n4), .A1(n3), .A2(readIn), .B0(memRead), .B1(n14), .Y(
        n13) );
  INVX2TS U23 ( .A(n30), .Y(n1) );
  AOI32XLTS U24 ( .A0(n4), .A1(n3), .A2(writeIn), .B0(memWrite), .B1(n14), .Y(
        n30) );
  OAI21XLTS U25 ( .A0(readIn), .A1(writeIn), .B0(n3), .Y(n20) );
  NAND2XLTS U26 ( .A(localRouterAddress[5]), .B(n8), .Y(n25) );
  NAND2XLTS U27 ( .A(localRouterAddress[4]), .B(n9), .Y(n26) );
  NOR2XLTS U28 ( .A(n8), .B(localRouterAddress[5]), .Y(n29) );
  AOI211X1TS U29 ( .A0(n27), .A1(n28), .B0(n20), .C0(n29), .Y(n42) );
  AND2X2TS U30 ( .A(n26), .B(n25), .Y(n27) );
  INVXLTS U31 ( .A(destinationAddressIn[11]), .Y(n10) );
  AOI211X1TS U32 ( .A0(n23), .A1(n24), .B0(n20), .C0(n5), .Y(n43) );
  INVX2TS U33 ( .A(n25), .Y(n5) );
  NAND3BXLTS U34 ( .AN(localRouterAddress[3]), .B(n26), .C(
        destinationAddressIn[11]), .Y(n24) );
  INVXLTS U35 ( .A(destinationAddressIn[9]), .Y(n12) );
  INVXLTS U36 ( .A(localRouterAddress[0]), .Y(n7) );
endmodule


module cacheAccessArbiter ( clk, reset, cacheAddressIn_NORTH, 
        requesterAddressIn_NORTH, memRead_NORTH, memWrite_NORTH, dataIn_NORTH, 
        readReady_NORTH, requesterAddressOut_NORTH, cacheDataOut_NORTH, 
        cacheAddressIn_SOUTH, requesterAddressIn_SOUTH, memRead_SOUTH, 
        memWrite_SOUTH, dataIn_SOUTH, readReady_SOUTH, 
        requesterAddressOut_SOUTH, cacheDataOut_SOUTH, cacheAddressIn_EAST, 
        requesterAddressIn_EAST, memRead_EAST, memWrite_EAST, dataIn_EAST, 
        readReady_EAST, requesterAddressOut_EAST, cacheDataOut_EAST, 
        cacheAddressIn_WEST, requesterAddressIn_WEST, memRead_WEST, 
        memWrite_WEST, dataIn_WEST, readReady_WEST, requesterAddressOut_WEST, 
        cacheDataOut_WEST, cacheDataIn_A, cacheAddressIn_A, cacheDataOut_A, 
        memWrite_A, cacheDataIn_B, cacheAddressIn_B, cacheDataOut_B, 
        memWrite_B );
  input [7:0] cacheAddressIn_NORTH;
  input [5:0] requesterAddressIn_NORTH;
  input [31:0] dataIn_NORTH;
  output [5:0] requesterAddressOut_NORTH;
  output [31:0] cacheDataOut_NORTH;
  input [7:0] cacheAddressIn_SOUTH;
  input [5:0] requesterAddressIn_SOUTH;
  input [31:0] dataIn_SOUTH;
  output [5:0] requesterAddressOut_SOUTH;
  output [31:0] cacheDataOut_SOUTH;
  input [7:0] cacheAddressIn_EAST;
  input [5:0] requesterAddressIn_EAST;
  input [31:0] dataIn_EAST;
  output [5:0] requesterAddressOut_EAST;
  output [31:0] cacheDataOut_EAST;
  input [7:0] cacheAddressIn_WEST;
  input [5:0] requesterAddressIn_WEST;
  input [31:0] dataIn_WEST;
  output [5:0] requesterAddressOut_WEST;
  output [31:0] cacheDataOut_WEST;
  output [31:0] cacheDataIn_A;
  output [7:0] cacheAddressIn_A;
  input [31:0] cacheDataOut_A;
  output [31:0] cacheDataIn_B;
  output [7:0] cacheAddressIn_B;
  input [31:0] cacheDataOut_B;
  input clk, reset, memRead_NORTH, memWrite_NORTH, memRead_SOUTH,
         memWrite_SOUTH, memRead_EAST, memWrite_EAST, memRead_WEST,
         memWrite_WEST;
  output readReady_NORTH, readReady_SOUTH, readReady_EAST, readReady_WEST,
         memWrite_A, memWrite_B;
  wire   n3345, n3343, n3546, n1072, n3547, n1073, n3548, n1074, n3549, n1075,
         n3550, n1076, n3551, n1077, n3552, n1078, n3553, n1079, n3554, n1080,
         n3555, n1081, n3556, n1082, n3557, n1083, n3558, n1084, n3559, n1085,
         n3560, n1086, n3561, n1087, n3562, n1088, n3563, n1089, n3564, n1090,
         n3565, n1091, n3566, n1092, n3567, n1093, n3568, n1094, n3569, n1095,
         n3570, n1096, n3571, n1097, n3572, n1098, n3573, n1099, n3574, n1100,
         n3575, n1101, n3576, n1102, n3577, n1103, n3253,
         \requesterPortBuffer[7][0] , n3266, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3208, n3207, n3206, n3205, n3204,
         n3203, \requesterPortBuffer[0][0] , n3268,
         \requesterPortBuffer[0][1] , n3382, n1172, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3378, n3267, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3418, n3482, n3419, n3483, n3420, n3484, n3421, n3485, n3422, n3486,
         n3423, n3487, n3424, n3488, n3425, n3489, n3426, n3490, n3427, n3491,
         n3428, n3492, n3429, n3493, n3430, n3494, n3431, n3495, n3432, n3496,
         n3433, n3497, n3434, n3498, n3435, n3499, n3436, n3500, n3437, n3501,
         n3438, n3502, n3439, n3503, n3440, n3504, n3441, n3505, n3442, n3506,
         n3443, n3507, n3444, n3508, n3445, n3509, n3446, n3510, n3447, n3511,
         n3448, n3512, n3449, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3286, n3302, n3287, n3303, n3288, n3304, n3289, n3305,
         n3290, n3306, n3291, n3307, n3292, n3308, n3293, n3309, n3621, n1147,
         n3622, n1148, n3623, n1149, n3624, n1150, n3625, n1151, n3626, n1152,
         n3627, n1153, n3628, n1154, n3629, n1155, n3630, n1156, n3631, n1157,
         n3632, n1158, n3633, n1159, n3634, n1160, n3635, n1161, n3636, n1162,
         n3637, n1163, n3638, n1164, n3639, n1165, n3640, n1166, n3641, n1167,
         n3165, n3164, n3163, n3162, n3161, n3160, n3183, n3182, n3181, n3180,
         n3179, n3178, n3177, n3176, n3175, n3174, n3173, n3172, n3171, n3170,
         n3169, n3168, n3167, n3166, n3344, n3250, n3677, n3251, n3678, n3277,
         n3276, n3275, n3274, n3273, n3272, n3271, n3270, n3249, n3248, n3247,
         n3246, n3245, n3244, n3243, n3242, n3241, n3240, n3239, n3238, n3237,
         n3236, n3235, n3234, n3233, n3232, n3231, n3230, n3229, n3228, n3227,
         n3226, n3225, n3224, n3223, n3222, n3221, n3220, n3219, n3218, n3184,
         n3217, n3377, n3376, n3375, n3374, n3373, n3372, n3371, n3370, n3369,
         n3368, n3367, n3366, n3365, n3364, n3363, n3362, n3361, n3360, n3359,
         n3358, n3357, n3356, n3355, n3354, n3353, n3352, n3351, n3350, n3349,
         n3348, n3347, n3346, n3216, n3215, n3214, n3213, n3212, n3211, n3210,
         n3209, N10040, N10030, N10020, N10010, N10216, N10215, N10214, N10213,
         N10212, N10211, N10210, N10209, N10208, N10207, N10206, N10205,
         N10204, N10203, N10202, N10201, N10200, N10199, N10198, N10197,
         N10196, N10195, N10194, N10193, N10192, N10191, N10190, N10189,
         N10188, N10187, N10186, N10185, N10182, N10181, N10180, N10179,
         N10178, N10177, N10176, N10175, N10174, N10173, N10172, N10171,
         N10170, N10169, N10168, N10167, N10166, N10165, N10164, N10163,
         N10162, N10161, N10160, N10159, N10158, N10157, N10156, N10155,
         N10154, N10153, N10152, N10151, N10148, N10147, N10146, N10145,
         N10144, N10143, N10142, N10141, N10140, N10139, N10138, N10137,
         N10136, N10135, N10134, N10133, N10132, N10131, N10130, N10129,
         N10128, N10127, N10126, N10125, N10124, N10123, N10122, N10121,
         N10120, N10119, N10118, N10117, N10114, N10113, N10112, N10111,
         N10110, N10109, N10108, N10107, N10106, N10105, N10104, N10103,
         N10102, N10101, N10100, N10099, N10098, N10097, N10096, N10095,
         N10094, N10093, N10092, N10091, N10090, N10089, N10088, N10087,
         N10086, N10085, N10084, N10083, n3264, n3265, n3197, n3198, n3199,
         n3200, n3201, n3202, n3185, n3186, n3187, n3188, n3189, n3190,
         \requesterPortBuffer[4][1] , \requesterPortBuffer[4][0] ,
         \requesterPortBuffer[2][0] , \requesterPortBuffer[5][1] ,
         \requesterPortBuffer[5][0] , \requesterPortBuffer[6][1] ,
         \requesterPortBuffer[6][0] , n3252, \requesterPortBuffer[7][1] ,
         n3379, n1169, n3318, n1219, n3319, n1220, n3320, n1221, n3321, n1222,
         n3322, n1223, n3323, n1224, n3324, n1225, n3325, n1226, n3384, n1174,
         n3383, n1173, n3381, n1171, n3196, \requesterAddressBuffer[0][5] ,
         n3195, \requesterAddressBuffer[0][4] , n3193,
         \requesterAddressBuffer[0][2] , n3194, \requesterAddressBuffer[0][3] ,
         n3192, \requesterAddressBuffer[0][1] , n3191,
         \requesterAddressBuffer[0][0] , n3334, n1235, n3335, n1236, n3336,
         n1237, n3337, n1238, n3338, n1239, n3339, n1240, n3340, n1241, n3341,
         n1242, n3380, n1170, n3385, n1175, n3610, n1136, n3611, n1137, n3612,
         n1138, n3613, n1139, n3614, n1140, n3615, n1141, n3616, n1142, n3617,
         n1143, n3618, n1144, n3619, n1145, n3620, n1146, n3643, n910, n3644,
         n4621, n3642, n880, n596, n597, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n645, n646, n647, n648, n649, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n739, n740,
         n741, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n806, n807, n810, n811, n812, n813, n814,
         n816, n818, n819, n820, n821, n822, n824, n825, n827, n828, n830,
         n831, n832, n833, n835, n837, n844, n885, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n994, n996, n997, n998, n999, n1000, n1001,
         n1003, n1004, n1005, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1168, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1369, n1370, n1371, n1372, n1373, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1473, n1474, n1475, n1476, n1477, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1503, n1504, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1516, n1517, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
         n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
         n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
         n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
         n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
         n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
         n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
         n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2014,
         n2016, n2018, n2020, n2022, n2024, n2026, n2028, n2030, n2032, n2034,
         n2036, n2038, n2040, n2042, n2044, n2046, n2048, n2050, n2052, n2054,
         n2056, n2058, n2060, n2062, n2064, n2066, n2068, n2070, n2072, n2074,
         n2076, n2078, n2080, n2082, n2084, n2086, n2088, n2090, n2092, n2095,
         n2096, n2097, n2098, n2100, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n598, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n737, n738, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n803, n804,
         n805, n808, n809, n815, n817, n823, n826, n829, n834, n836, n838,
         n839, n840, n841, n842, n843, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n881, n882, n883, n884,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n911, n912, n913, n914, n915, n916, n917, n918, n993,
         n995, n1002, n1006, n1187, n1188, n1283, n1324, n1325, n1368, n1374,
         n1472, n1478, n1492, n1502, n1505, n1515, n1518, n1589, n1660, n1717,
         n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2015, n2017, n2019,
         n2021, n2023, n2025, n2027, n2029, n2031, n2033, n2035, n2037, n2039,
         n2041, n2043, n2045, n2047, n2049, n2051, n2053, n2055, n2057, n2059,
         n2061, n2063, n2065, n2067, n2069, n2071, n2073, n2075, n2077, n2079,
         n2081, n2083, n2085, n2087, n2089, n2091, n2093, n2094, n2099, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386;
  wire   [1:0] prevRequesterPort_B;
  wire   [5:0] prevRequesterAddress_B;
  wire   [5:0] prevRequesterAddress_A;

  DFFNSRX2TS \requesterPortBuffer_reg[4][1]  ( .D(n756), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[4][1] ) );
  DFFNSRX2TS \requesterPortBuffer_reg[4][0]  ( .D(n758), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[4][0] ) );
  DFFNSRX2TS \requesterPortBuffer_reg[5][1]  ( .D(n759), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[5][1] ) );
  DFFNSRX2TS \requesterPortBuffer_reg[5][0]  ( .D(n597), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[5][0] ) );
  DFFNSRX2TS \requesterPortBuffer_reg[6][1]  ( .D(n647), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[6][1] ) );
  DFFNSRX2TS \requesterPortBuffer_reg[6][0]  ( .D(n646), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[6][0] ) );
  DFFNSRX2TS \requesterPortBuffer_reg[2][0]  ( .D(n757), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[2][0] ) );
  DFFNSRX2TS \requesterPortBuffer_reg[7][0]  ( .D(n3253), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[7][0] ) );
  DFFNSRX2TS \requesterPortBuffer_reg[7][1]  ( .D(n3252), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[7][1] ) );
  DFFNSRX2TS \addressToWriteBuffer_reg[7][7]  ( .D(n3278), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1930) );
  DFFNSRX2TS \addressToWriteBuffer_reg[7][6]  ( .D(n3279), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1929) );
  DFFNSRX2TS \addressToWriteBuffer_reg[7][5]  ( .D(n3280), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1928) );
  DFFNSRX2TS \addressToWriteBuffer_reg[7][4]  ( .D(n3281), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1927) );
  DFFNSRX2TS \addressToWriteBuffer_reg[7][3]  ( .D(n3282), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1926) );
  DFFNSRX2TS \addressToWriteBuffer_reg[7][2]  ( .D(n3283), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1925) );
  DFFNSRX2TS \addressToWriteBuffer_reg[7][1]  ( .D(n3284), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1924) );
  DFFNSRX2TS \addressToWriteBuffer_reg[7][0]  ( .D(n3285), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1923) );
  DFFNSRX2TS \requesterPortBuffer_reg[3][0]  ( .D(n648), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1963) );
  DFFNSRX2TS \requesterPortBuffer_reg[3][1]  ( .D(n715), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1964) );
  DFFNSRX2TS \requesterPortBuffer_reg[2][1]  ( .D(n649), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1966) );
  DFFNSRX2TS \requesterPortBuffer_reg[0][0]  ( .D(n645), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[0][0] ) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][31]  ( .D(n3386), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1962) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][30]  ( .D(n3387), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1961) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][29]  ( .D(n3388), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1960) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][28]  ( .D(n3389), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1959) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][27]  ( .D(n3390), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1958) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][26]  ( .D(n3391), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1957) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][25]  ( .D(n3392), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1956) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][24]  ( .D(n3393), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1955) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][23]  ( .D(n3394), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1954) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][22]  ( .D(n3395), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1953) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][21]  ( .D(n3396), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1952) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][20]  ( .D(n3397), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1951) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][19]  ( .D(n3398), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1950) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][18]  ( .D(n3399), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1949) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][17]  ( .D(n3400), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1948) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][16]  ( .D(n3401), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1947) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][15]  ( .D(n3402), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1946) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][14]  ( .D(n3403), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1945) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][13]  ( .D(n3404), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1944) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][12]  ( .D(n3405), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1943) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][11]  ( .D(n3406), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1942) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][10]  ( .D(n3407), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1941) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][9]  ( .D(n3408), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1940) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][8]  ( .D(n3409), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1939) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][7]  ( .D(n3410), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1938) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][6]  ( .D(n3411), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1937) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][5]  ( .D(n3412), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1936) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][4]  ( .D(n3413), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1935) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][3]  ( .D(n3414), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1934) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][2]  ( .D(n3415), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1933) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][1]  ( .D(n3416), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1932) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][0]  ( .D(n3417), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1931) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][31]  ( .D(n3450), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1858) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][30]  ( .D(n3451), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1857) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][29]  ( .D(n3452), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1856) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][28]  ( .D(n3453), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1855) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][27]  ( .D(n3454), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1854) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][26]  ( .D(n3455), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1853) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][25]  ( .D(n3456), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1852) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][24]  ( .D(n3457), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1851) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][23]  ( .D(n3458), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1850) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][22]  ( .D(n3459), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1849) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][21]  ( .D(n3460), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1848) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][20]  ( .D(n3461), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1847) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][19]  ( .D(n3462), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1846) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][18]  ( .D(n3463), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1845) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][17]  ( .D(n3464), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1844) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][16]  ( .D(n3465), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1843) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][15]  ( .D(n3466), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1842) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][14]  ( .D(n3467), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1841) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][13]  ( .D(n3468), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1840) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][12]  ( .D(n3469), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1839) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][11]  ( .D(n3470), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1838) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][10]  ( .D(n3471), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1837) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][9]  ( .D(n3472), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1836) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][8]  ( .D(n3473), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1835) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][7]  ( .D(n3474), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1834) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][6]  ( .D(n3475), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1833) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][5]  ( .D(n3476), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1832) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][4]  ( .D(n3477), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1831) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][3]  ( .D(n3478), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1830) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][2]  ( .D(n3479), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1829) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][1]  ( .D(n3480), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1828) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][0]  ( .D(n3481), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1827) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][31]  ( .D(n3418), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1826) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][30]  ( .D(n3419), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1824) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][29]  ( .D(n3420), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1822) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][28]  ( .D(n3421), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1820) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][27]  ( .D(n3422), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1818) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][26]  ( .D(n3423), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1816) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][25]  ( .D(n3424), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1814) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][24]  ( .D(n3425), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1812) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][23]  ( .D(n3426), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1810) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][22]  ( .D(n3427), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1808) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][21]  ( .D(n3428), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1806) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][20]  ( .D(n3429), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1804) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][19]  ( .D(n3430), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1802) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][18]  ( .D(n3431), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1800) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][17]  ( .D(n3432), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1798) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][16]  ( .D(n3433), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1796) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][15]  ( .D(n3434), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1794) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][14]  ( .D(n3435), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1792) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][13]  ( .D(n3436), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1790) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][12]  ( .D(n3437), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1788) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][11]  ( .D(n3438), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1786) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][10]  ( .D(n3439), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1784) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][9]  ( .D(n3440), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1782) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][8]  ( .D(n3441), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1780) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][7]  ( .D(n3442), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1778) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][6]  ( .D(n3443), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1776) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][5]  ( .D(n3444), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1774) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][4]  ( .D(n3445), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1772) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][3]  ( .D(n3446), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1770) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][2]  ( .D(n3447), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1768) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][1]  ( .D(n3448), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1766) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][0]  ( .D(n3449), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1764) );
  DFFNSRX2TS \isRead_reg[1]  ( .D(n3345), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .QN(n30) );
  DFFNSRX2TS \addressToWriteBuffer_reg[1][7]  ( .D(n3326), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n43) );
  DFFNSRX2TS \addressToWriteBuffer_reg[1][6]  ( .D(n3327), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n42) );
  DFFNSRX2TS \addressToWriteBuffer_reg[1][5]  ( .D(n3328), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n41) );
  DFFNSRX2TS \addressToWriteBuffer_reg[1][4]  ( .D(n3329), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n40) );
  DFFNSRX2TS \addressToWriteBuffer_reg[1][3]  ( .D(n3330), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n39) );
  DFFNSRX2TS \addressToWriteBuffer_reg[1][2]  ( .D(n3331), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n38) );
  DFFNSRX2TS \addressToWriteBuffer_reg[1][1]  ( .D(n3332), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n37) );
  DFFNSRX2TS \addressToWriteBuffer_reg[1][0]  ( .D(n3333), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n44) );
  DFFNSRX2TS \requesterAddressBuffer_reg[1][5]  ( .D(n3208), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n36) );
  DFFNSRX2TS \requesterAddressBuffer_reg[1][4]  ( .D(n3207), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n35) );
  DFFNSRX2TS \requesterAddressBuffer_reg[1][3]  ( .D(n3206), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n34) );
  DFFNSRX2TS \requesterAddressBuffer_reg[1][2]  ( .D(n3205), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n33) );
  DFFNSRX2TS \requesterAddressBuffer_reg[1][1]  ( .D(n3204), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n32) );
  DFFNSRX2TS \requesterAddressBuffer_reg[1][0]  ( .D(n3203), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n31) );
  DFFNSRX2TS \requesterPortBuffer_reg[0][1]  ( .D(n3268), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[0][1] ) );
  DFFNSRX2TS \isRead_reg[0]  ( .D(n3343), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        n2098), .QN(n45) );
  DFFNSRX2TS \addressToWriteBuffer_reg[5][7]  ( .D(n3294), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1890), .QN(n71) );
  DFFNSRX2TS \addressToWriteBuffer_reg[5][6]  ( .D(n3295), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1889), .QN(n70) );
  DFFNSRX2TS \addressToWriteBuffer_reg[5][5]  ( .D(n3296), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1888), .QN(n69) );
  DFFNSRX2TS \addressToWriteBuffer_reg[5][4]  ( .D(n3297), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1887), .QN(n68) );
  DFFNSRX2TS \addressToWriteBuffer_reg[5][3]  ( .D(n3298), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1886), .QN(n67) );
  DFFNSRX2TS \addressToWriteBuffer_reg[5][2]  ( .D(n3299), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1885), .QN(n66) );
  DFFNSRX2TS \addressToWriteBuffer_reg[5][1]  ( .D(n3300), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1884), .QN(n65) );
  DFFNSRX2TS \addressToWriteBuffer_reg[5][0]  ( .D(n3301), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1883), .QN(n64) );
  DFFNSRX2TS \addressToWriteBuffer_reg[3][7]  ( .D(n3310), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1882), .QN(n79) );
  DFFNSRX2TS \addressToWriteBuffer_reg[3][6]  ( .D(n3311), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1881), .QN(n78) );
  DFFNSRX2TS \addressToWriteBuffer_reg[3][5]  ( .D(n3312), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1880), .QN(n77) );
  DFFNSRX2TS \addressToWriteBuffer_reg[3][4]  ( .D(n3313), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1879), .QN(n76) );
  DFFNSRX2TS \addressToWriteBuffer_reg[3][3]  ( .D(n3314), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1878), .QN(n75) );
  DFFNSRX2TS \addressToWriteBuffer_reg[3][2]  ( .D(n3315), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1877), .QN(n74) );
  DFFNSRX2TS \addressToWriteBuffer_reg[3][1]  ( .D(n3316), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1876), .QN(n73) );
  DFFNSRX2TS \addressToWriteBuffer_reg[3][0]  ( .D(n3317), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1875), .QN(n72) );
  DFFNSRX2TS \addressToWriteBuffer_reg[6][7]  ( .D(n3286), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1874), .QN(n63) );
  DFFNSRX2TS \addressToWriteBuffer_reg[4][7]  ( .D(n3302), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1873), .QN(n62) );
  DFFNSRX2TS \addressToWriteBuffer_reg[6][6]  ( .D(n3287), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1872), .QN(n61) );
  DFFNSRX2TS \addressToWriteBuffer_reg[4][6]  ( .D(n3303), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1871), .QN(n60) );
  DFFNSRX2TS \addressToWriteBuffer_reg[6][5]  ( .D(n3288), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1870), .QN(n59) );
  DFFNSRX2TS \addressToWriteBuffer_reg[4][5]  ( .D(n3304), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1869), .QN(n58) );
  DFFNSRX2TS \addressToWriteBuffer_reg[6][4]  ( .D(n3289), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1868), .QN(n57) );
  DFFNSRX2TS \addressToWriteBuffer_reg[4][4]  ( .D(n3305), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1867), .QN(n56) );
  DFFNSRX2TS \addressToWriteBuffer_reg[6][3]  ( .D(n3290), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1866), .QN(n55) );
  DFFNSRX2TS \addressToWriteBuffer_reg[4][3]  ( .D(n3306), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1865), .QN(n54) );
  DFFNSRX2TS \addressToWriteBuffer_reg[6][2]  ( .D(n3291), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1864), .QN(n53) );
  DFFNSRX2TS \addressToWriteBuffer_reg[4][2]  ( .D(n3307), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1863), .QN(n52) );
  DFFNSRX2TS \addressToWriteBuffer_reg[6][1]  ( .D(n3292), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1862), .QN(n51) );
  DFFNSRX2TS \addressToWriteBuffer_reg[4][1]  ( .D(n3308), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1861), .QN(n50) );
  DFFNSRX2TS \addressToWriteBuffer_reg[6][0]  ( .D(n3293), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1860), .QN(n49) );
  DFFNSRX2TS \addressToWriteBuffer_reg[4][0]  ( .D(n3309), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1859), .QN(n48) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][31]  ( .D(n3514), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1922), .QN(n111) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][30]  ( .D(n3515), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1921), .QN(n110) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][29]  ( .D(n3516), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1920), .QN(n109) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][28]  ( .D(n3517), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1919), .QN(n108) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][27]  ( .D(n3518), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1918), .QN(n107) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][26]  ( .D(n3519), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1917), .QN(n106) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][25]  ( .D(n3520), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1916), .QN(n105) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][24]  ( .D(n3521), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1915), .QN(n104) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][23]  ( .D(n3522), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1914), .QN(n103) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][22]  ( .D(n3523), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1913), .QN(n102) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][21]  ( .D(n3524), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1912), .QN(n101) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][20]  ( .D(n3525), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1911), .QN(n100) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][19]  ( .D(n3526), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1910), .QN(n99) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][18]  ( .D(n3527), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1909), .QN(n98) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][17]  ( .D(n3528), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1908), .QN(n97) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][16]  ( .D(n3529), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1907), .QN(n96) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][15]  ( .D(n3530), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1906), .QN(n95) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][14]  ( .D(n3531), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1905), .QN(n94) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][13]  ( .D(n3532), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1904), .QN(n93) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][12]  ( .D(n3533), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1903), .QN(n92) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][11]  ( .D(n3534), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1902), .QN(n91) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][10]  ( .D(n3535), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1901), .QN(n90) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][9]  ( .D(n3536), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1900), .QN(n89) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][8]  ( .D(n3537), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1899), .QN(n88) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][7]  ( .D(n3538), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1898), .QN(n87) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][6]  ( .D(n3539), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1897), .QN(n86) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][5]  ( .D(n3540), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1896), .QN(n85) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][4]  ( .D(n3541), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1895), .QN(n84) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][3]  ( .D(n3542), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1894), .QN(n83) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][2]  ( .D(n3543), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1893), .QN(n82) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][1]  ( .D(n3544), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1892), .QN(n81) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][0]  ( .D(n3545), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1891), .QN(n80) );
  DFFNSRX2TS \requesterPortBuffer_reg[1][1]  ( .D(n3266), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2100), .QN(n47) );
  DFFNSRX2TS \requesterPortBuffer_reg[1][0]  ( .D(n3267), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2096), .QN(n46) );
  DFFNSRX2TS \nextEmptyBuffer_reg[1]  ( .D(n3643), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n318), .QN(n910) );
  DFFNSRX2TS \nextEmptyBuffer_reg[2]  ( .D(n3642), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n328), .QN(n880) );
  DFFNSRX2TS prevMemRead_B_reg ( .D(n3344), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .QN(n27) );
  DFFNSRX2TS prevMemRead_A_reg ( .D(n596), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .QN(n2) );
  DFFNSRX2TS \prevRequesterAddress_B_reg[5]  ( .D(n3197), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_B[5]), .QN(n8) );
  DFFNSRX2TS \prevRequesterAddress_B_reg[4]  ( .D(n3198), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_B[4]), .QN(n7) );
  DFFNSRX2TS \prevRequesterAddress_B_reg[3]  ( .D(n3199), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_B[3]), .QN(n6) );
  DFFNSRX2TS \prevRequesterAddress_B_reg[2]  ( .D(n3200), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_B[2]), .QN(n5) );
  DFFNSRX2TS \prevRequesterAddress_B_reg[1]  ( .D(n3201), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_B[1]), .QN(n4) );
  DFFNSRX2TS \prevRequesterAddress_B_reg[0]  ( .D(n3202), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_B[0]), .QN(n3) );
  DFFNSRX2TS \prevRequesterAddress_A_reg[5]  ( .D(n3185), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_A[5]), .QN(n251) );
  DFFNSRX2TS \prevRequesterAddress_A_reg[4]  ( .D(n3186), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_A[4]), .QN(n252) );
  DFFNSRX2TS \prevRequesterAddress_A_reg[3]  ( .D(n3187), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_A[3]), .QN(n253) );
  DFFNSRX2TS \prevRequesterAddress_A_reg[2]  ( .D(n3188), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_A[2]), .QN(n254) );
  DFFNSRX2TS \prevRequesterAddress_A_reg[1]  ( .D(n3189), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_A[1]), .QN(n255) );
  DFFNSRX2TS \prevRequesterAddress_A_reg[0]  ( .D(n3190), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_A[0]), .QN(n256) );
  DFFNSRX2TS \prevRequesterPort_B_reg[0]  ( .D(n3265), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterPort_B[0]), .QN(n26) );
  DFFNSRX2TS \prevRequesterPort_B_reg[1]  ( .D(n3264), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterPort_B[1]), .QN(n1) );
  DFFNSRX2TS \cacheAddressIn_A_reg[7]  ( .D(n3277), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_A[7]), .QN(n1974) );
  DFFNSRX2TS \cacheAddressIn_A_reg[6]  ( .D(n3276), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_A[6]), .QN(n1973) );
  DFFNSRX2TS \cacheAddressIn_A_reg[5]  ( .D(n3275), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_A[5]), .QN(n1972) );
  DFFNSRX2TS \cacheAddressIn_A_reg[4]  ( .D(n3274), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_A[4]), .QN(n1971) );
  DFFNSRX2TS \cacheAddressIn_A_reg[3]  ( .D(n3273), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_A[3]), .QN(n1970) );
  DFFNSRX2TS \cacheAddressIn_A_reg[2]  ( .D(n3272), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_A[2]), .QN(n1969) );
  DFFNSRX2TS \cacheAddressIn_A_reg[1]  ( .D(n3271), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_A[1]), .QN(n1968) );
  DFFNSRX2TS \cacheAddressIn_A_reg[0]  ( .D(n3270), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_A[0]), .QN(n1967) );
  DFFNSRX2TS \cacheDataIn_A_reg[31]  ( .D(n3249), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[31]), .QN(n2006) );
  DFFNSRX2TS \cacheDataIn_A_reg[30]  ( .D(n3248), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[30]), .QN(n2005) );
  DFFNSRX2TS \cacheDataIn_A_reg[29]  ( .D(n3247), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[29]), .QN(n2004) );
  DFFNSRX2TS \cacheDataIn_A_reg[28]  ( .D(n3246), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[28]), .QN(n2003) );
  DFFNSRX2TS \cacheDataIn_A_reg[27]  ( .D(n3245), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[27]), .QN(n2002) );
  DFFNSRX2TS \cacheDataIn_A_reg[26]  ( .D(n3244), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[26]), .QN(n2001) );
  DFFNSRX2TS \cacheDataIn_A_reg[25]  ( .D(n3243), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[25]), .QN(n2000) );
  DFFNSRX2TS \cacheDataIn_A_reg[24]  ( .D(n3242), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[24]), .QN(n1999) );
  DFFNSRX2TS \cacheDataIn_A_reg[23]  ( .D(n3241), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[23]), .QN(n1998) );
  DFFNSRX2TS \cacheDataIn_A_reg[22]  ( .D(n3240), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[22]), .QN(n1997) );
  DFFNSRX2TS \cacheDataIn_A_reg[21]  ( .D(n3239), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[21]), .QN(n1996) );
  DFFNSRX2TS \cacheDataIn_A_reg[20]  ( .D(n3238), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[20]), .QN(n1995) );
  DFFNSRX2TS \cacheDataIn_A_reg[19]  ( .D(n3237), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[19]), .QN(n1994) );
  DFFNSRX2TS \cacheDataIn_A_reg[18]  ( .D(n3236), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[18]), .QN(n1993) );
  DFFNSRX2TS \cacheDataIn_A_reg[17]  ( .D(n3235), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[17]), .QN(n1992) );
  DFFNSRX2TS \cacheDataIn_A_reg[16]  ( .D(n3234), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[16]), .QN(n1991) );
  DFFNSRX2TS \cacheDataIn_A_reg[15]  ( .D(n3233), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[15]), .QN(n1990) );
  DFFNSRX2TS \cacheDataIn_A_reg[14]  ( .D(n3232), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[14]), .QN(n1989) );
  DFFNSRX2TS \cacheDataIn_A_reg[13]  ( .D(n3231), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[13]), .QN(n1988) );
  DFFNSRX2TS \cacheDataIn_A_reg[12]  ( .D(n3230), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[12]), .QN(n1987) );
  DFFNSRX2TS \cacheDataIn_A_reg[11]  ( .D(n3229), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[11]), .QN(n1986) );
  DFFNSRX2TS \cacheDataIn_A_reg[10]  ( .D(n3228), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[10]), .QN(n1985) );
  DFFNSRX2TS \cacheDataIn_A_reg[9]  ( .D(n3227), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[9]), .QN(n1984) );
  DFFNSRX2TS \cacheDataIn_A_reg[8]  ( .D(n3226), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[8]), .QN(n1983) );
  DFFNSRX2TS \cacheDataIn_A_reg[7]  ( .D(n3225), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[7]), .QN(n1982) );
  DFFNSRX2TS \cacheDataIn_A_reg[6]  ( .D(n3224), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[6]), .QN(n1981) );
  DFFNSRX2TS \cacheDataIn_A_reg[5]  ( .D(n3223), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[5]), .QN(n1980) );
  DFFNSRX2TS \cacheDataIn_A_reg[4]  ( .D(n3222), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[4]), .QN(n1979) );
  DFFNSRX2TS \cacheDataIn_A_reg[3]  ( .D(n3221), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[3]), .QN(n1978) );
  DFFNSRX2TS \cacheDataIn_A_reg[2]  ( .D(n3220), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[2]), .QN(n1977) );
  DFFNSRX2TS \cacheDataIn_A_reg[1]  ( .D(n3219), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[1]), .QN(n1976) );
  DFFNSRX2TS \cacheDataIn_A_reg[0]  ( .D(n3218), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[0]), .QN(n1975) );
  DFFNSRX2TS memWrite_A_reg ( .D(n3184), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        memWrite_A), .QN(n2095) );
  DFFNSRX2TS memWrite_B_reg ( .D(n3217), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        memWrite_B), .QN(n2097) );
  DFFNSRX2TS \cacheDataIn_B_reg[31]  ( .D(n3377), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[31]), .QN(n2092) );
  DFFNSRX2TS \cacheDataIn_B_reg[30]  ( .D(n3376), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[30]), .QN(n2090) );
  DFFNSRX2TS \cacheDataIn_B_reg[29]  ( .D(n3375), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[29]), .QN(n2088) );
  DFFNSRX2TS \cacheDataIn_B_reg[28]  ( .D(n3374), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[28]), .QN(n2086) );
  DFFNSRX2TS \cacheDataIn_B_reg[27]  ( .D(n3373), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[27]), .QN(n2084) );
  DFFNSRX2TS \cacheDataIn_B_reg[26]  ( .D(n3372), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[26]), .QN(n2082) );
  DFFNSRX2TS \cacheDataIn_B_reg[25]  ( .D(n3371), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[25]), .QN(n2080) );
  DFFNSRX2TS \cacheDataIn_B_reg[24]  ( .D(n3370), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[24]), .QN(n2078) );
  DFFNSRX2TS \cacheDataIn_B_reg[23]  ( .D(n3369), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[23]), .QN(n2076) );
  DFFNSRX2TS \cacheDataIn_B_reg[22]  ( .D(n3368), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[22]), .QN(n2074) );
  DFFNSRX2TS \cacheDataIn_B_reg[21]  ( .D(n3367), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[21]), .QN(n2072) );
  DFFNSRX2TS \cacheDataIn_B_reg[20]  ( .D(n3366), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[20]), .QN(n2070) );
  DFFNSRX2TS \cacheDataIn_B_reg[19]  ( .D(n3365), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[19]), .QN(n2068) );
  DFFNSRX2TS \cacheDataIn_B_reg[18]  ( .D(n3364), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[18]), .QN(n2066) );
  DFFNSRX2TS \cacheDataIn_B_reg[17]  ( .D(n3363), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[17]), .QN(n2064) );
  DFFNSRX2TS \cacheDataIn_B_reg[16]  ( .D(n3362), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[16]), .QN(n2062) );
  DFFNSRX2TS \cacheDataIn_B_reg[15]  ( .D(n3361), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[15]), .QN(n2060) );
  DFFNSRX2TS \cacheDataIn_B_reg[14]  ( .D(n3360), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[14]), .QN(n2058) );
  DFFNSRX2TS \cacheDataIn_B_reg[13]  ( .D(n3359), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[13]), .QN(n2056) );
  DFFNSRX2TS \cacheDataIn_B_reg[12]  ( .D(n3358), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[12]), .QN(n2054) );
  DFFNSRX2TS \cacheDataIn_B_reg[11]  ( .D(n3357), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[11]), .QN(n2052) );
  DFFNSRX2TS \cacheDataIn_B_reg[10]  ( .D(n3356), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[10]), .QN(n2050) );
  DFFNSRX2TS \cacheDataIn_B_reg[9]  ( .D(n3355), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[9]), .QN(n2048) );
  DFFNSRX2TS \cacheDataIn_B_reg[8]  ( .D(n3354), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[8]), .QN(n2046) );
  DFFNSRX2TS \cacheDataIn_B_reg[7]  ( .D(n3353), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[7]), .QN(n2044) );
  DFFNSRX2TS \cacheDataIn_B_reg[6]  ( .D(n3352), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[6]), .QN(n2042) );
  DFFNSRX2TS \cacheDataIn_B_reg[5]  ( .D(n3351), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[5]), .QN(n2040) );
  DFFNSRX2TS \cacheDataIn_B_reg[4]  ( .D(n3350), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[4]), .QN(n2038) );
  DFFNSRX2TS \cacheDataIn_B_reg[3]  ( .D(n3349), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[3]), .QN(n2036) );
  DFFNSRX2TS \cacheDataIn_B_reg[2]  ( .D(n3348), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[2]), .QN(n2034) );
  DFFNSRX2TS \cacheDataIn_B_reg[1]  ( .D(n3347), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[1]), .QN(n2032) );
  DFFNSRX2TS \cacheDataIn_B_reg[0]  ( .D(n3346), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[0]), .QN(n2030) );
  DFFNSRX2TS \cacheAddressIn_B_reg[7]  ( .D(n3216), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_B[7]), .QN(n2028) );
  DFFNSRX2TS \cacheAddressIn_B_reg[6]  ( .D(n3215), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_B[6]), .QN(n2026) );
  DFFNSRX2TS \cacheAddressIn_B_reg[5]  ( .D(n3214), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_B[5]), .QN(n2024) );
  DFFNSRX2TS \cacheAddressIn_B_reg[4]  ( .D(n3213), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_B[4]), .QN(n2022) );
  DFFNSRX2TS \cacheAddressIn_B_reg[3]  ( .D(n3212), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_B[3]), .QN(n2020) );
  DFFNSRX2TS \cacheAddressIn_B_reg[2]  ( .D(n3211), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_B[2]), .QN(n2018) );
  DFFNSRX2TS \cacheAddressIn_B_reg[1]  ( .D(n3210), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_B[1]), .QN(n2016) );
  DFFNSRX2TS \cacheAddressIn_B_reg[0]  ( .D(n3209), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_B[0]), .QN(n2014) );
  EDFFX2TS \readReady_Concatenated_reg[3]  ( .D(N10040), .E(n2374), .CK(clk), 
        .Q(readReady_WEST) );
  EDFFX2TS \readReady_Concatenated_reg[2]  ( .D(N10030), .E(n2375), .CK(clk), 
        .Q(readReady_EAST) );
  EDFFX2TS \readReady_Concatenated_reg[1]  ( .D(N10020), .E(n2374), .CK(clk), 
        .Q(readReady_SOUTH) );
  EDFFX2TS \readReady_Concatenated_reg[0]  ( .D(N10010), .E(n2375), .CK(clk), 
        .Q(readReady_NORTH) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[0][5]  ( .D(n3165), .CK(clk), 
        .Q(requesterAddressOut_NORTH[5]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[0][4]  ( .D(n3164), .CK(clk), 
        .Q(requesterAddressOut_NORTH[4]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[0][3]  ( .D(n3163), .CK(clk), 
        .Q(requesterAddressOut_NORTH[3]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[0][2]  ( .D(n3162), .CK(clk), 
        .Q(requesterAddressOut_NORTH[2]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[0][1]  ( .D(n3161), .CK(clk), 
        .Q(requesterAddressOut_NORTH[1]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[0][0]  ( .D(n3160), .CK(clk), 
        .Q(requesterAddressOut_NORTH[0]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[2][5]  ( .D(n3177), .CK(clk), 
        .Q(requesterAddressOut_EAST[5]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[2][4]  ( .D(n3176), .CK(clk), 
        .Q(requesterAddressOut_EAST[4]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[2][3]  ( .D(n3175), .CK(clk), 
        .Q(requesterAddressOut_EAST[3]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[2][2]  ( .D(n3174), .CK(clk), 
        .Q(requesterAddressOut_EAST[2]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[2][1]  ( .D(n3173), .CK(clk), 
        .Q(requesterAddressOut_EAST[1]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[2][0]  ( .D(n3172), .CK(clk), 
        .Q(requesterAddressOut_EAST[0]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[1][5]  ( .D(n3171), .CK(clk), 
        .Q(requesterAddressOut_SOUTH[5]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[1][4]  ( .D(n3170), .CK(clk), 
        .Q(requesterAddressOut_SOUTH[4]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[1][3]  ( .D(n3169), .CK(clk), 
        .Q(requesterAddressOut_SOUTH[3]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[1][2]  ( .D(n3168), .CK(clk), 
        .Q(requesterAddressOut_SOUTH[2]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[1][1]  ( .D(n3167), .CK(clk), 
        .Q(requesterAddressOut_SOUTH[1]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[1][0]  ( .D(n3166), .CK(clk), 
        .Q(requesterAddressOut_SOUTH[0]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[3][5]  ( .D(n3183), .CK(clk), 
        .Q(requesterAddressOut_WEST[5]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[3][4]  ( .D(n3182), .CK(clk), 
        .Q(requesterAddressOut_WEST[4]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[3][3]  ( .D(n3181), .CK(clk), 
        .Q(requesterAddressOut_WEST[3]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[3][2]  ( .D(n3180), .CK(clk), 
        .Q(requesterAddressOut_WEST[2]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[3][1]  ( .D(n3179), .CK(clk), 
        .Q(requesterAddressOut_WEST[1]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[3][0]  ( .D(n3178), .CK(clk), 
        .Q(requesterAddressOut_WEST[0]) );
  TLATXLTS \dataOut_Concatenated_reg[3][31]  ( .G(clk), .D(N10216), .Q(
        cacheDataOut_WEST[31]) );
  TLATXLTS \dataOut_Concatenated_reg[3][30]  ( .G(clk), .D(N10215), .Q(
        cacheDataOut_WEST[30]) );
  TLATXLTS \dataOut_Concatenated_reg[3][29]  ( .G(clk), .D(N10214), .Q(
        cacheDataOut_WEST[29]) );
  TLATXLTS \dataOut_Concatenated_reg[3][28]  ( .G(clk), .D(N10213), .Q(
        cacheDataOut_WEST[28]) );
  TLATXLTS \dataOut_Concatenated_reg[3][27]  ( .G(clk), .D(N10212), .Q(
        cacheDataOut_WEST[27]) );
  TLATXLTS \dataOut_Concatenated_reg[3][26]  ( .G(clk), .D(N10211), .Q(
        cacheDataOut_WEST[26]) );
  TLATXLTS \dataOut_Concatenated_reg[3][25]  ( .G(clk), .D(N10210), .Q(
        cacheDataOut_WEST[25]) );
  TLATXLTS \dataOut_Concatenated_reg[3][24]  ( .G(clk), .D(N10209), .Q(
        cacheDataOut_WEST[24]) );
  TLATXLTS \dataOut_Concatenated_reg[3][23]  ( .G(clk), .D(N10208), .Q(
        cacheDataOut_WEST[23]) );
  TLATXLTS \dataOut_Concatenated_reg[3][22]  ( .G(clk), .D(N10207), .Q(
        cacheDataOut_WEST[22]) );
  TLATXLTS \dataOut_Concatenated_reg[3][21]  ( .G(clk), .D(N10206), .Q(
        cacheDataOut_WEST[21]) );
  TLATXLTS \dataOut_Concatenated_reg[3][20]  ( .G(clk), .D(N10205), .Q(
        cacheDataOut_WEST[20]) );
  TLATXLTS \dataOut_Concatenated_reg[3][19]  ( .G(clk), .D(N10204), .Q(
        cacheDataOut_WEST[19]) );
  TLATXLTS \dataOut_Concatenated_reg[3][18]  ( .G(clk), .D(N10203), .Q(
        cacheDataOut_WEST[18]) );
  TLATXLTS \dataOut_Concatenated_reg[3][17]  ( .G(clk), .D(N10202), .Q(
        cacheDataOut_WEST[17]) );
  TLATXLTS \dataOut_Concatenated_reg[3][16]  ( .G(clk), .D(N10201), .Q(
        cacheDataOut_WEST[16]) );
  TLATXLTS \dataOut_Concatenated_reg[3][15]  ( .G(clk), .D(N10200), .Q(
        cacheDataOut_WEST[15]) );
  TLATXLTS \dataOut_Concatenated_reg[3][14]  ( .G(clk), .D(N10199), .Q(
        cacheDataOut_WEST[14]) );
  TLATXLTS \dataOut_Concatenated_reg[3][13]  ( .G(clk), .D(N10198), .Q(
        cacheDataOut_WEST[13]) );
  TLATXLTS \dataOut_Concatenated_reg[3][12]  ( .G(clk), .D(N10197), .Q(
        cacheDataOut_WEST[12]) );
  TLATXLTS \dataOut_Concatenated_reg[3][11]  ( .G(clk), .D(N10196), .Q(
        cacheDataOut_WEST[11]) );
  TLATXLTS \dataOut_Concatenated_reg[3][10]  ( .G(clk), .D(N10195), .Q(
        cacheDataOut_WEST[10]) );
  TLATXLTS \dataOut_Concatenated_reg[3][9]  ( .G(clk), .D(N10194), .Q(
        cacheDataOut_WEST[9]) );
  TLATXLTS \dataOut_Concatenated_reg[3][8]  ( .G(clk), .D(N10193), .Q(
        cacheDataOut_WEST[8]) );
  TLATXLTS \dataOut_Concatenated_reg[3][7]  ( .G(clk), .D(N10192), .Q(
        cacheDataOut_WEST[7]) );
  TLATXLTS \dataOut_Concatenated_reg[3][6]  ( .G(clk), .D(N10191), .Q(
        cacheDataOut_WEST[6]) );
  TLATXLTS \dataOut_Concatenated_reg[3][5]  ( .G(clk), .D(N10190), .Q(
        cacheDataOut_WEST[5]) );
  TLATXLTS \dataOut_Concatenated_reg[3][4]  ( .G(clk), .D(N10189), .Q(
        cacheDataOut_WEST[4]) );
  TLATXLTS \dataOut_Concatenated_reg[3][3]  ( .G(clk), .D(N10188), .Q(
        cacheDataOut_WEST[3]) );
  TLATXLTS \dataOut_Concatenated_reg[3][2]  ( .G(clk), .D(N10187), .Q(
        cacheDataOut_WEST[2]) );
  TLATXLTS \dataOut_Concatenated_reg[3][1]  ( .G(clk), .D(N10186), .Q(
        cacheDataOut_WEST[1]) );
  TLATXLTS \dataOut_Concatenated_reg[3][0]  ( .G(clk), .D(N10185), .Q(
        cacheDataOut_WEST[0]) );
  TLATXLTS \dataOut_Concatenated_reg[2][31]  ( .G(clk), .D(N10182), .Q(
        cacheDataOut_EAST[31]) );
  TLATXLTS \dataOut_Concatenated_reg[2][30]  ( .G(clk), .D(N10181), .Q(
        cacheDataOut_EAST[30]) );
  TLATXLTS \dataOut_Concatenated_reg[2][29]  ( .G(clk), .D(N10180), .Q(
        cacheDataOut_EAST[29]) );
  TLATXLTS \dataOut_Concatenated_reg[2][28]  ( .G(clk), .D(N10179), .Q(
        cacheDataOut_EAST[28]) );
  TLATXLTS \dataOut_Concatenated_reg[2][27]  ( .G(clk), .D(N10178), .Q(
        cacheDataOut_EAST[27]) );
  TLATXLTS \dataOut_Concatenated_reg[2][26]  ( .G(clk), .D(N10177), .Q(
        cacheDataOut_EAST[26]) );
  TLATXLTS \dataOut_Concatenated_reg[2][25]  ( .G(clk), .D(N10176), .Q(
        cacheDataOut_EAST[25]) );
  TLATXLTS \dataOut_Concatenated_reg[2][24]  ( .G(clk), .D(N10175), .Q(
        cacheDataOut_EAST[24]) );
  TLATXLTS \dataOut_Concatenated_reg[2][23]  ( .G(clk), .D(N10174), .Q(
        cacheDataOut_EAST[23]) );
  TLATXLTS \dataOut_Concatenated_reg[2][22]  ( .G(clk), .D(N10173), .Q(
        cacheDataOut_EAST[22]) );
  TLATXLTS \dataOut_Concatenated_reg[2][21]  ( .G(clk), .D(N10172), .Q(
        cacheDataOut_EAST[21]) );
  TLATXLTS \dataOut_Concatenated_reg[2][20]  ( .G(clk), .D(N10171), .Q(
        cacheDataOut_EAST[20]) );
  TLATXLTS \dataOut_Concatenated_reg[2][19]  ( .G(clk), .D(N10170), .Q(
        cacheDataOut_EAST[19]) );
  TLATXLTS \dataOut_Concatenated_reg[2][18]  ( .G(clk), .D(N10169), .Q(
        cacheDataOut_EAST[18]) );
  TLATXLTS \dataOut_Concatenated_reg[2][17]  ( .G(clk), .D(N10168), .Q(
        cacheDataOut_EAST[17]) );
  TLATXLTS \dataOut_Concatenated_reg[2][16]  ( .G(clk), .D(N10167), .Q(
        cacheDataOut_EAST[16]) );
  TLATXLTS \dataOut_Concatenated_reg[2][15]  ( .G(clk), .D(N10166), .Q(
        cacheDataOut_EAST[15]) );
  TLATXLTS \dataOut_Concatenated_reg[2][14]  ( .G(clk), .D(N10165), .Q(
        cacheDataOut_EAST[14]) );
  TLATXLTS \dataOut_Concatenated_reg[2][13]  ( .G(clk), .D(N10164), .Q(
        cacheDataOut_EAST[13]) );
  TLATXLTS \dataOut_Concatenated_reg[2][12]  ( .G(clk), .D(N10163), .Q(
        cacheDataOut_EAST[12]) );
  TLATXLTS \dataOut_Concatenated_reg[2][11]  ( .G(clk), .D(N10162), .Q(
        cacheDataOut_EAST[11]) );
  TLATXLTS \dataOut_Concatenated_reg[2][10]  ( .G(clk), .D(N10161), .Q(
        cacheDataOut_EAST[10]) );
  TLATXLTS \dataOut_Concatenated_reg[2][9]  ( .G(clk), .D(N10160), .Q(
        cacheDataOut_EAST[9]) );
  TLATXLTS \dataOut_Concatenated_reg[2][8]  ( .G(clk), .D(N10159), .Q(
        cacheDataOut_EAST[8]) );
  TLATXLTS \dataOut_Concatenated_reg[2][7]  ( .G(clk), .D(N10158), .Q(
        cacheDataOut_EAST[7]) );
  TLATXLTS \dataOut_Concatenated_reg[2][6]  ( .G(clk), .D(N10157), .Q(
        cacheDataOut_EAST[6]) );
  TLATXLTS \dataOut_Concatenated_reg[2][5]  ( .G(clk), .D(N10156), .Q(
        cacheDataOut_EAST[5]) );
  TLATXLTS \dataOut_Concatenated_reg[2][4]  ( .G(clk), .D(N10155), .Q(
        cacheDataOut_EAST[4]) );
  TLATXLTS \dataOut_Concatenated_reg[2][3]  ( .G(clk), .D(N10154), .Q(
        cacheDataOut_EAST[3]) );
  TLATXLTS \dataOut_Concatenated_reg[2][2]  ( .G(clk), .D(N10153), .Q(
        cacheDataOut_EAST[2]) );
  TLATXLTS \dataOut_Concatenated_reg[2][1]  ( .G(clk), .D(N10152), .Q(
        cacheDataOut_EAST[1]) );
  TLATXLTS \dataOut_Concatenated_reg[2][0]  ( .G(clk), .D(N10151), .Q(
        cacheDataOut_EAST[0]) );
  TLATXLTS \dataOut_Concatenated_reg[1][31]  ( .G(clk), .D(N10148), .Q(
        cacheDataOut_SOUTH[31]) );
  TLATXLTS \dataOut_Concatenated_reg[1][30]  ( .G(clk), .D(N10147), .Q(
        cacheDataOut_SOUTH[30]) );
  TLATXLTS \dataOut_Concatenated_reg[1][29]  ( .G(clk), .D(N10146), .Q(
        cacheDataOut_SOUTH[29]) );
  TLATXLTS \dataOut_Concatenated_reg[1][28]  ( .G(clk), .D(N10145), .Q(
        cacheDataOut_SOUTH[28]) );
  TLATXLTS \dataOut_Concatenated_reg[1][27]  ( .G(clk), .D(N10144), .Q(
        cacheDataOut_SOUTH[27]) );
  TLATXLTS \dataOut_Concatenated_reg[1][26]  ( .G(clk), .D(N10143), .Q(
        cacheDataOut_SOUTH[26]) );
  TLATXLTS \dataOut_Concatenated_reg[1][25]  ( .G(clk), .D(N10142), .Q(
        cacheDataOut_SOUTH[25]) );
  TLATXLTS \dataOut_Concatenated_reg[1][24]  ( .G(clk), .D(N10141), .Q(
        cacheDataOut_SOUTH[24]) );
  TLATXLTS \dataOut_Concatenated_reg[1][23]  ( .G(clk), .D(N10140), .Q(
        cacheDataOut_SOUTH[23]) );
  TLATXLTS \dataOut_Concatenated_reg[1][22]  ( .G(clk), .D(N10139), .Q(
        cacheDataOut_SOUTH[22]) );
  TLATXLTS \dataOut_Concatenated_reg[1][21]  ( .G(clk), .D(N10138), .Q(
        cacheDataOut_SOUTH[21]) );
  TLATXLTS \dataOut_Concatenated_reg[1][20]  ( .G(clk), .D(N10137), .Q(
        cacheDataOut_SOUTH[20]) );
  TLATXLTS \dataOut_Concatenated_reg[1][19]  ( .G(clk), .D(N10136), .Q(
        cacheDataOut_SOUTH[19]) );
  TLATXLTS \dataOut_Concatenated_reg[1][18]  ( .G(clk), .D(N10135), .Q(
        cacheDataOut_SOUTH[18]) );
  TLATXLTS \dataOut_Concatenated_reg[1][17]  ( .G(clk), .D(N10134), .Q(
        cacheDataOut_SOUTH[17]) );
  TLATXLTS \dataOut_Concatenated_reg[1][16]  ( .G(clk), .D(N10133), .Q(
        cacheDataOut_SOUTH[16]) );
  TLATXLTS \dataOut_Concatenated_reg[1][15]  ( .G(clk), .D(N10132), .Q(
        cacheDataOut_SOUTH[15]) );
  TLATXLTS \dataOut_Concatenated_reg[1][14]  ( .G(clk), .D(N10131), .Q(
        cacheDataOut_SOUTH[14]) );
  TLATXLTS \dataOut_Concatenated_reg[1][13]  ( .G(clk), .D(N10130), .Q(
        cacheDataOut_SOUTH[13]) );
  TLATXLTS \dataOut_Concatenated_reg[1][12]  ( .G(clk), .D(N10129), .Q(
        cacheDataOut_SOUTH[12]) );
  TLATXLTS \dataOut_Concatenated_reg[1][11]  ( .G(clk), .D(N10128), .Q(
        cacheDataOut_SOUTH[11]) );
  TLATXLTS \dataOut_Concatenated_reg[1][10]  ( .G(clk), .D(N10127), .Q(
        cacheDataOut_SOUTH[10]) );
  TLATXLTS \dataOut_Concatenated_reg[1][9]  ( .G(clk), .D(N10126), .Q(
        cacheDataOut_SOUTH[9]) );
  TLATXLTS \dataOut_Concatenated_reg[1][8]  ( .G(clk), .D(N10125), .Q(
        cacheDataOut_SOUTH[8]) );
  TLATXLTS \dataOut_Concatenated_reg[1][7]  ( .G(clk), .D(N10124), .Q(
        cacheDataOut_SOUTH[7]) );
  TLATXLTS \dataOut_Concatenated_reg[1][6]  ( .G(clk), .D(N10123), .Q(
        cacheDataOut_SOUTH[6]) );
  TLATXLTS \dataOut_Concatenated_reg[1][5]  ( .G(clk), .D(N10122), .Q(
        cacheDataOut_SOUTH[5]) );
  TLATXLTS \dataOut_Concatenated_reg[1][4]  ( .G(clk), .D(N10121), .Q(
        cacheDataOut_SOUTH[4]) );
  TLATXLTS \dataOut_Concatenated_reg[1][3]  ( .G(clk), .D(N10120), .Q(
        cacheDataOut_SOUTH[3]) );
  TLATXLTS \dataOut_Concatenated_reg[1][2]  ( .G(clk), .D(N10119), .Q(
        cacheDataOut_SOUTH[2]) );
  TLATXLTS \dataOut_Concatenated_reg[1][1]  ( .G(clk), .D(N10118), .Q(
        cacheDataOut_SOUTH[1]) );
  TLATXLTS \dataOut_Concatenated_reg[1][0]  ( .G(clk), .D(N10117), .Q(
        cacheDataOut_SOUTH[0]) );
  TLATXLTS \dataOut_Concatenated_reg[0][31]  ( .G(clk), .D(N10114), .Q(
        cacheDataOut_NORTH[31]) );
  TLATXLTS \dataOut_Concatenated_reg[0][30]  ( .G(clk), .D(N10113), .Q(
        cacheDataOut_NORTH[30]) );
  TLATXLTS \dataOut_Concatenated_reg[0][29]  ( .G(clk), .D(N10112), .Q(
        cacheDataOut_NORTH[29]) );
  TLATXLTS \dataOut_Concatenated_reg[0][28]  ( .G(clk), .D(N10111), .Q(
        cacheDataOut_NORTH[28]) );
  TLATXLTS \dataOut_Concatenated_reg[0][27]  ( .G(clk), .D(N10110), .Q(
        cacheDataOut_NORTH[27]) );
  TLATXLTS \dataOut_Concatenated_reg[0][26]  ( .G(clk), .D(N10109), .Q(
        cacheDataOut_NORTH[26]) );
  TLATXLTS \dataOut_Concatenated_reg[0][25]  ( .G(clk), .D(N10108), .Q(
        cacheDataOut_NORTH[25]) );
  TLATXLTS \dataOut_Concatenated_reg[0][24]  ( .G(clk), .D(N10107), .Q(
        cacheDataOut_NORTH[24]) );
  TLATXLTS \dataOut_Concatenated_reg[0][23]  ( .G(clk), .D(N10106), .Q(
        cacheDataOut_NORTH[23]) );
  TLATXLTS \dataOut_Concatenated_reg[0][22]  ( .G(clk), .D(N10105), .Q(
        cacheDataOut_NORTH[22]) );
  TLATXLTS \dataOut_Concatenated_reg[0][21]  ( .G(clk), .D(N10104), .Q(
        cacheDataOut_NORTH[21]) );
  TLATXLTS \dataOut_Concatenated_reg[0][20]  ( .G(clk), .D(N10103), .Q(
        cacheDataOut_NORTH[20]) );
  TLATXLTS \dataOut_Concatenated_reg[0][19]  ( .G(clk), .D(N10102), .Q(
        cacheDataOut_NORTH[19]) );
  TLATXLTS \dataOut_Concatenated_reg[0][18]  ( .G(clk), .D(N10101), .Q(
        cacheDataOut_NORTH[18]) );
  TLATXLTS \dataOut_Concatenated_reg[0][17]  ( .G(clk), .D(N10100), .Q(
        cacheDataOut_NORTH[17]) );
  TLATXLTS \dataOut_Concatenated_reg[0][16]  ( .G(clk), .D(N10099), .Q(
        cacheDataOut_NORTH[16]) );
  TLATXLTS \dataOut_Concatenated_reg[0][15]  ( .G(clk), .D(N10098), .Q(
        cacheDataOut_NORTH[15]) );
  TLATXLTS \dataOut_Concatenated_reg[0][14]  ( .G(clk), .D(N10097), .Q(
        cacheDataOut_NORTH[14]) );
  TLATXLTS \dataOut_Concatenated_reg[0][13]  ( .G(clk), .D(N10096), .Q(
        cacheDataOut_NORTH[13]) );
  TLATXLTS \dataOut_Concatenated_reg[0][12]  ( .G(clk), .D(N10095), .Q(
        cacheDataOut_NORTH[12]) );
  TLATXLTS \dataOut_Concatenated_reg[0][11]  ( .G(clk), .D(N10094), .Q(
        cacheDataOut_NORTH[11]) );
  TLATXLTS \dataOut_Concatenated_reg[0][10]  ( .G(clk), .D(N10093), .Q(
        cacheDataOut_NORTH[10]) );
  TLATXLTS \dataOut_Concatenated_reg[0][9]  ( .G(clk), .D(N10092), .Q(
        cacheDataOut_NORTH[9]) );
  TLATXLTS \dataOut_Concatenated_reg[0][8]  ( .G(clk), .D(N10091), .Q(
        cacheDataOut_NORTH[8]) );
  TLATXLTS \dataOut_Concatenated_reg[0][7]  ( .G(clk), .D(N10090), .Q(
        cacheDataOut_NORTH[7]) );
  TLATXLTS \dataOut_Concatenated_reg[0][6]  ( .G(clk), .D(N10089), .Q(
        cacheDataOut_NORTH[6]) );
  TLATXLTS \dataOut_Concatenated_reg[0][5]  ( .G(clk), .D(N10088), .Q(
        cacheDataOut_NORTH[5]) );
  TLATXLTS \dataOut_Concatenated_reg[0][4]  ( .G(clk), .D(N10087), .Q(
        cacheDataOut_NORTH[4]) );
  TLATXLTS \dataOut_Concatenated_reg[0][3]  ( .G(clk), .D(N10086), .Q(
        cacheDataOut_NORTH[3]) );
  TLATXLTS \dataOut_Concatenated_reg[0][2]  ( .G(clk), .D(N10085), .Q(
        cacheDataOut_NORTH[2]) );
  TLATXLTS \dataOut_Concatenated_reg[0][1]  ( .G(clk), .D(N10084), .Q(
        cacheDataOut_NORTH[1]) );
  TLATXLTS \dataOut_Concatenated_reg[0][0]  ( .G(clk), .D(N10083), .Q(
        cacheDataOut_NORTH[0]) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][31]  ( .D(n3546), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1072) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][30]  ( .D(n3547), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1073) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][29]  ( .D(n3548), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1074) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][28]  ( .D(n3549), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1075) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][27]  ( .D(n3550), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1076) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][26]  ( .D(n3551), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1077) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][25]  ( .D(n3552), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1078) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][24]  ( .D(n3553), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1079) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][23]  ( .D(n3554), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1080) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][22]  ( .D(n3555), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1081) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][21]  ( .D(n3556), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1082) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][20]  ( .D(n3557), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1083) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][19]  ( .D(n3558), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1084) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][18]  ( .D(n3559), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1085) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][17]  ( .D(n3560), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1086) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][16]  ( .D(n3561), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1087) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][15]  ( .D(n3562), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1088) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][14]  ( .D(n3563), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1089) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][13]  ( .D(n3564), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1090) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][12]  ( .D(n3565), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1091) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][11]  ( .D(n3566), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1092) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][10]  ( .D(n3567), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1093) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][9]  ( .D(n3568), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1094) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][8]  ( .D(n3569), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1095) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][7]  ( .D(n3570), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1096) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][6]  ( .D(n3571), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1097) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][5]  ( .D(n3572), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1098) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][4]  ( .D(n3573), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1099) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][3]  ( .D(n3574), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1100) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][2]  ( .D(n3575), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1101) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][1]  ( .D(n3576), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1102) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][0]  ( .D(n3577), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1103) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][31]  ( .D(n3578), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n599) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][30]  ( .D(n3579), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n600) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][29]  ( .D(n3580), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n601) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][28]  ( .D(n3581), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n602) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][27]  ( .D(n3582), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n603) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][26]  ( .D(n3583), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n604) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][25]  ( .D(n3584), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n605) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][24]  ( .D(n3585), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n606) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][23]  ( .D(n3586), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n607) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][22]  ( .D(n3587), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n608) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][21]  ( .D(n3588), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n609) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][20]  ( .D(n3589), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n610) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][19]  ( .D(n3590), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n611) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][18]  ( .D(n3591), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n612) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][17]  ( .D(n3592), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n613) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][16]  ( .D(n3593), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n614) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][15]  ( .D(n3594), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n615) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][14]  ( .D(n3595), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n616) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][13]  ( .D(n3596), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n617) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][12]  ( .D(n3597), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n618) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][11]  ( .D(n3598), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n619) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][10]  ( .D(n3599), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n620) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][9]  ( .D(n3600), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n621) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][8]  ( .D(n3601), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n622) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][7]  ( .D(n3602), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n623) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][6]  ( .D(n3603), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n624) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][5]  ( .D(n3604), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n625) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][4]  ( .D(n3605), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n626) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][3]  ( .D(n3606), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n627) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][2]  ( .D(n3607), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n628) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][1]  ( .D(n3608), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n629) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][0]  ( .D(n3609), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n630) );
  DFFNSRXLTS \dataToWriteBuffer_reg[4][31]  ( .D(n3482), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1825) );
  DFFNSRXLTS \dataToWriteBuffer_reg[4][30]  ( .D(n3483), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1823) );
  DFFNSRXLTS \dataToWriteBuffer_reg[4][29]  ( .D(n3484), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1821) );
  DFFNSRXLTS \dataToWriteBuffer_reg[4][28]  ( .D(n3485), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1819) );
  DFFNSRXLTS \dataToWriteBuffer_reg[4][27]  ( .D(n3486), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1817) );
  DFFNSRXLTS \dataToWriteBuffer_reg[4][26]  ( .D(n3487), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1815) );
  DFFNSRXLTS \dataToWriteBuffer_reg[4][25]  ( .D(n3488), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1813) );
  DFFNSRXLTS \dataToWriteBuffer_reg[4][24]  ( .D(n3489), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1811) );
  DFFNSRXLTS \dataToWriteBuffer_reg[4][23]  ( .D(n3490), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1809) );
  DFFNSRXLTS \dataToWriteBuffer_reg[4][22]  ( .D(n3491), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1807) );
  DFFNSRXLTS \dataToWriteBuffer_reg[4][21]  ( .D(n3492), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1805) );
  DFFNSRXLTS \dataToWriteBuffer_reg[4][20]  ( .D(n3493), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1803) );
  DFFNSRXLTS \dataToWriteBuffer_reg[4][19]  ( .D(n3494), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1801) );
  DFFNSRXLTS \dataToWriteBuffer_reg[4][18]  ( .D(n3495), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1799) );
  DFFNSRXLTS \dataToWriteBuffer_reg[4][17]  ( .D(n3496), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1797) );
  DFFNSRXLTS \dataToWriteBuffer_reg[4][16]  ( .D(n3497), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1795) );
  DFFNSRXLTS \dataToWriteBuffer_reg[4][15]  ( .D(n3498), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1793) );
  DFFNSRXLTS \dataToWriteBuffer_reg[4][14]  ( .D(n3499), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1791) );
  DFFNSRXLTS \dataToWriteBuffer_reg[4][13]  ( .D(n3500), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1789) );
  DFFNSRXLTS \dataToWriteBuffer_reg[4][12]  ( .D(n3501), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1787) );
  DFFNSRXLTS \dataToWriteBuffer_reg[4][11]  ( .D(n3502), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1785) );
  DFFNSRXLTS \dataToWriteBuffer_reg[4][10]  ( .D(n3503), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1783) );
  DFFNSRXLTS \dataToWriteBuffer_reg[4][9]  ( .D(n3504), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1781) );
  DFFNSRXLTS \dataToWriteBuffer_reg[4][8]  ( .D(n3505), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1779) );
  DFFNSRXLTS \dataToWriteBuffer_reg[4][7]  ( .D(n3506), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1777) );
  DFFNSRXLTS \dataToWriteBuffer_reg[4][6]  ( .D(n3507), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1775) );
  DFFNSRXLTS \dataToWriteBuffer_reg[4][5]  ( .D(n3508), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1773) );
  DFFNSRXLTS \dataToWriteBuffer_reg[4][4]  ( .D(n3509), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1771) );
  DFFNSRXLTS \dataToWriteBuffer_reg[4][3]  ( .D(n3510), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1769) );
  DFFNSRXLTS \dataToWriteBuffer_reg[4][2]  ( .D(n3511), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1767) );
  DFFNSRXLTS \dataToWriteBuffer_reg[4][1]  ( .D(n3512), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1765) );
  DFFNSRXLTS \dataToWriteBuffer_reg[4][0]  ( .D(n3513), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1763) );
  DFFNSRXLTS \requesterAddressBuffer_reg[0][5]  ( .D(n3196), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressBuffer[0][5] ), .QN(n769) );
  DFFNSRXLTS \requesterAddressBuffer_reg[0][4]  ( .D(n3195), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressBuffer[0][4] ), .QN(n770) );
  DFFNSRXLTS \requesterAddressBuffer_reg[0][2]  ( .D(n3193), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressBuffer[0][2] ), .QN(n771) );
  DFFNSRXLTS \requesterAddressBuffer_reg[0][3]  ( .D(n3194), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressBuffer[0][3] ), .QN(n772) );
  DFFNSRXLTS \requesterAddressBuffer_reg[0][1]  ( .D(n3192), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressBuffer[0][1] ), .QN(n773) );
  DFFNSRXLTS \requesterAddressBuffer_reg[0][0]  ( .D(n3191), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressBuffer[0][0] ), .QN(n774) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][31]  ( .D(n3610), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n783), .QN(n1136) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][24]  ( .D(n3617), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n790), .QN(n1143) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][21]  ( .D(n3620), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n793), .QN(n1146) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][16]  ( .D(n3625), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n720), .QN(n1151) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][12]  ( .D(n3629), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n724), .QN(n1155) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][8]  ( .D(n3633), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n728), .QN(n1159) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][4]  ( .D(n3637), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n732), .QN(n1163) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][0]  ( .D(n3641), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n736), .QN(n1167) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][30]  ( .D(n3611), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n784), .QN(n1137) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][29]  ( .D(n3612), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n785), .QN(n1138) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][28]  ( .D(n3613), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n786), .QN(n1139) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][27]  ( .D(n3614), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n787), .QN(n1140) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][26]  ( .D(n3615), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n788), .QN(n1141) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][25]  ( .D(n3616), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n789), .QN(n1142) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][23]  ( .D(n3618), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n791), .QN(n1144) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][22]  ( .D(n3619), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n792), .QN(n1145) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][20]  ( .D(n3621), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n716), .QN(n1147) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][19]  ( .D(n3622), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n717), .QN(n1148) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][18]  ( .D(n3623), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n718), .QN(n1149) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][17]  ( .D(n3624), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n719), .QN(n1150) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][15]  ( .D(n3626), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n721), .QN(n1152) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][14]  ( .D(n3627), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n722), .QN(n1153) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][13]  ( .D(n3628), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n723), .QN(n1154) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][11]  ( .D(n3630), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n725), .QN(n1156) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][10]  ( .D(n3631), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n726), .QN(n1157) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][9]  ( .D(n3632), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n727), .QN(n1158) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][7]  ( .D(n3634), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n729), .QN(n1160) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][6]  ( .D(n3635), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n730), .QN(n1161) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][5]  ( .D(n3636), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n731), .QN(n1162) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][3]  ( .D(n3638), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n733), .QN(n1164) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][2]  ( .D(n3639), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n734), .QN(n1165) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][1]  ( .D(n3640), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n735), .QN(n1166) );
  DFFNSRXLTS \isWrite_reg[7]  ( .D(n3378), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .QN(n1965) );
  DFFNSRXLTS \isWrite_reg[6]  ( .D(n3379), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .QN(n1169) );
  DFFNSRXLTS \isWrite_reg[4]  ( .D(n3381), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .QN(n1171) );
  DFFNSRXLTS \isWrite_reg[2]  ( .D(n3383), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n768), .QN(n1173) );
  DFFNSRXLTS \isWrite_reg[5]  ( .D(n3380), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .QN(n1170) );
  DFFNSRXLTS \isWrite_reg[3]  ( .D(n3382), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .QN(n1172) );
  DFFNSRXLTS \isWrite_reg[0]  ( .D(n3385), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .QN(n1175) );
  DFFNSRXLTS \addressToWriteBuffer_reg[0][0]  ( .D(n3341), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n782), .QN(n1242) );
  DFFNSRXLTS \prevRequesterPort_A_reg[1]  ( .D(n3251), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n741), .QN(n3678) );
  DFFNSRXLTS \prevRequesterPort_A_reg[0]  ( .D(n3250), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n740), .QN(n3677) );
  DFFNSRXLTS \addressToWriteBuffer_reg[0][6]  ( .D(n3335), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n776), .QN(n1236) );
  DFFNSRXLTS \addressToWriteBuffer_reg[0][4]  ( .D(n3337), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n778), .QN(n1238) );
  DFFNSRXLTS \addressToWriteBuffer_reg[0][2]  ( .D(n3339), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n780), .QN(n1240) );
  DFFNSRXLTS \addressToWriteBuffer_reg[0][1]  ( .D(n3340), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n781), .QN(n1241) );
  DFFNSRXLTS \addressToWriteBuffer_reg[0][7]  ( .D(n3334), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n775), .QN(n1235) );
  DFFNSRXLTS \addressToWriteBuffer_reg[0][5]  ( .D(n3336), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n777), .QN(n1237) );
  DFFNSRXLTS \addressToWriteBuffer_reg[0][3]  ( .D(n3338), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n779), .QN(n1239) );
  DFFNSRXLTS \isWrite_reg[1]  ( .D(n3384), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .QN(n1174) );
  DFFNSRXLTS \addressToWriteBuffer_reg[2][7]  ( .D(n3318), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n760), .QN(n1219) );
  DFFNSRXLTS \addressToWriteBuffer_reg[2][6]  ( .D(n3319), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n761), .QN(n1220) );
  DFFNSRXLTS \addressToWriteBuffer_reg[2][5]  ( .D(n3320), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n762), .QN(n1221) );
  DFFNSRXLTS \addressToWriteBuffer_reg[2][4]  ( .D(n3321), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n763), .QN(n1222) );
  DFFNSRXLTS \addressToWriteBuffer_reg[2][3]  ( .D(n3322), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n764), .QN(n1223) );
  DFFNSRXLTS \addressToWriteBuffer_reg[2][2]  ( .D(n3323), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n765), .QN(n1224) );
  DFFNSRXLTS \addressToWriteBuffer_reg[2][1]  ( .D(n3324), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n766), .QN(n1225) );
  DFFNSRXLTS \addressToWriteBuffer_reg[2][0]  ( .D(n3325), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n767), .QN(n1226) );
  DFFNSRXLTS \nextEmptyBuffer_reg[0]  ( .D(n3644), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n9), .QN(n4621) );
  XNOR2X1TS U2 ( .A(n1443), .B(n298), .Y(n1448) );
  NOR2BX1TS U3 ( .AN(n1245), .B(n191), .Y(n1194) );
  NOR2BX1TS U4 ( .AN(n1367), .B(n330), .Y(n1332) );
  INVX2TS U5 ( .A(n1450), .Y(n144) );
  OR2X2TS U6 ( .A(memRead_SOUTH), .B(memWrite_SOUTH), .Y(n1442) );
  NAND2X1TS U7 ( .A(n1488), .B(n1461), .Y(n1189) );
  AND3X2TS U8 ( .A(n1038), .B(n341), .C(n806), .Y(n1005) );
  AND2X2TS U9 ( .A(n806), .B(n334), .Y(n340) );
  AND2X2TS U10 ( .A(n1282), .B(n801), .Y(n1249) );
  AND2X2TS U11 ( .A(n269), .B(n1109), .Y(n1044) );
  AND2X2TS U12 ( .A(n1186), .B(n10), .Y(n1114) );
  NAND2X1TS U13 ( .A(n259), .B(n1514), .Y(n1285) );
  OA21XLTS U14 ( .A0(n810), .A1(n1244), .B0(n1500), .Y(n1245) );
  NAND2X1TS U15 ( .A(n116), .B(n1514), .Y(n1326) );
  NOR2BX1TS U16 ( .AN(n1327), .B(n186), .Y(n1291) );
  OA21XLTS U17 ( .A0(n810), .A1(n1366), .B0(n1538), .Y(n1367) );
  AND2X2TS U18 ( .A(n1041), .B(n2373), .Y(n1109) );
  NAND2X1TS U19 ( .A(n1462), .B(n292), .Y(n1546) );
  CLKBUFX2TS U20 ( .A(n1373), .Y(n305) );
  CLKBUFX2TS U21 ( .A(n685), .Y(n684) );
  AOI222XLTS U22 ( .A0(memRead_EAST), .A1(n275), .B0(n1422), .B1(n1438), .C0(
        memRead_WEST), .C1(n1432), .Y(n1430) );
  INVX2TS U23 ( .A(n1442), .Y(n298) );
  AOI21X1TS U24 ( .A0(n342), .A1(n880), .B0(n818), .Y(n10) );
  AND2X2TS U25 ( .A(n1286), .B(n1284), .Y(n11) );
  AND2X2TS U26 ( .A(n1327), .B(n798), .Y(n12) );
  OR2X2TS U27 ( .A(n1461), .B(n145), .Y(n13) );
  NAND2X1TS U28 ( .A(n1326), .B(n798), .Y(n14) );
  NAND2X1TS U29 ( .A(n1244), .B(n329), .Y(n15) );
  OA21XLTS U30 ( .A0(n145), .A1(n1449), .B0(n1451), .Y(n16) );
  AND3X2TS U31 ( .A(n171), .B(n837), .C(n1691), .Y(n17) );
  AND3X2TS U32 ( .A(n1545), .B(n885), .C(n144), .Y(n18) );
  OR2X2TS U33 ( .A(n1189), .B(n182), .Y(n19) );
  OR2X2TS U34 ( .A(n178), .B(n1285), .Y(n20) );
  OR2X2TS U35 ( .A(n1326), .B(n187), .Y(n21) );
  AND3X2TS U36 ( .A(n1421), .B(n989), .C(n1420), .Y(n22) );
  OR2X2TS U37 ( .A(n183), .B(n795), .Y(n23) );
  OR2X2TS U38 ( .A(n179), .B(n822), .Y(n24) );
  OR3X1TS U39 ( .A(n1723), .B(n2362), .C(n1725), .Y(n25) );
  OR2X2TS U40 ( .A(n880), .B(n910), .Y(n28) );
  XOR2X1TS U41 ( .A(n123), .B(n329), .Y(n29) );
  CLKBUFX2TS U42 ( .A(memWrite_WEST), .Y(n112) );
  INVXLTS U43 ( .A(n18), .Y(n113) );
  INVXLTS U44 ( .A(n16), .Y(n114) );
  INVXLTS U45 ( .A(n16), .Y(n115) );
  INVXLTS U46 ( .A(n13), .Y(n116) );
  INVXLTS U47 ( .A(n13), .Y(n117) );
  INVX1TS U48 ( .A(n1443), .Y(n118) );
  INVXLTS U49 ( .A(n118), .Y(n119) );
  INVXLTS U50 ( .A(n166), .Y(n120) );
  INVXLTS U51 ( .A(n166), .Y(n121) );
  INVXLTS U52 ( .A(n318), .Y(n122) );
  INVXLTS U53 ( .A(n122), .Y(n123) );
  INVXLTS U54 ( .A(n17), .Y(n124) );
  INVXLTS U55 ( .A(n17), .Y(n125) );
  INVXLTS U56 ( .A(n1692), .Y(n126) );
  INVXLTS U57 ( .A(n126), .Y(n127) );
  INVXLTS U58 ( .A(n1750), .Y(n128) );
  INVXLTS U59 ( .A(n128), .Y(n129) );
  INVXLTS U60 ( .A(n1738), .Y(n130) );
  INVXLTS U61 ( .A(n130), .Y(n131) );
  INVXLTS U62 ( .A(n1726), .Y(n132) );
  INVXLTS U63 ( .A(n132), .Y(n133) );
  INVXLTS U64 ( .A(n29), .Y(n134) );
  INVXLTS U65 ( .A(n29), .Y(n135) );
  INVXLTS U66 ( .A(n989), .Y(n136) );
  INVXLTS U67 ( .A(n136), .Y(n137) );
  INVXLTS U68 ( .A(n25), .Y(n138) );
  INVXLTS U69 ( .A(n25), .Y(n139) );
  INVXLTS U70 ( .A(n1578), .Y(n140) );
  INVXLTS U71 ( .A(n140), .Y(n141) );
  INVXLTS U72 ( .A(n1595), .Y(n142) );
  INVXLTS U73 ( .A(n142), .Y(n143) );
  INVXLTS U74 ( .A(n1450), .Y(n145) );
  INVXLTS U75 ( .A(n15), .Y(n146) );
  INVXLTS U76 ( .A(n15), .Y(n147) );
  INVXLTS U77 ( .A(n14), .Y(n148) );
  INVXLTS U78 ( .A(n14), .Y(n149) );
  INVXLTS U79 ( .A(n24), .Y(n150) );
  INVXLTS U80 ( .A(n24), .Y(n151) );
  INVXLTS U81 ( .A(n23), .Y(n152) );
  INVXLTS U82 ( .A(n23), .Y(n153) );
  INVXLTS U83 ( .A(n12), .Y(n154) );
  INVXLTS U84 ( .A(n12), .Y(n155) );
  INVXLTS U85 ( .A(n12), .Y(n156) );
  INVXLTS U86 ( .A(n11), .Y(n157) );
  INVXLTS U87 ( .A(n11), .Y(n158) );
  INVXLTS U88 ( .A(n11), .Y(n159) );
  INVXLTS U89 ( .A(n20), .Y(n160) );
  INVXLTS U90 ( .A(n20), .Y(n161) );
  INVXLTS U91 ( .A(n20), .Y(n162) );
  INVXLTS U92 ( .A(n21), .Y(n163) );
  INVXLTS U93 ( .A(n21), .Y(n164) );
  INVXLTS U94 ( .A(n21), .Y(n165) );
  INVXLTS U95 ( .A(n1243), .Y(n166) );
  INVXLTS U96 ( .A(n19), .Y(n167) );
  INVXLTS U97 ( .A(n19), .Y(n168) );
  INVXLTS U98 ( .A(n19), .Y(n169) );
  INVXLTS U99 ( .A(n1443), .Y(n170) );
  INVXLTS U100 ( .A(n1443), .Y(n171) );
  INVXLTS U101 ( .A(n22), .Y(n172) );
  INVXLTS U102 ( .A(n22), .Y(n173) );
  INVXLTS U103 ( .A(n22), .Y(n174) );
  INVXLTS U104 ( .A(n9), .Y(n175) );
  INVXLTS U105 ( .A(n801), .Y(n176) );
  INVXLTS U106 ( .A(n176), .Y(n177) );
  INVXLTS U107 ( .A(n176), .Y(n178) );
  INVXLTS U108 ( .A(n176), .Y(n179) );
  INVXLTS U109 ( .A(n10), .Y(n180) );
  INVXLTS U110 ( .A(n180), .Y(n181) );
  INVXLTS U111 ( .A(n180), .Y(n182) );
  INVXLTS U112 ( .A(n180), .Y(n183) );
  INVXLTS U113 ( .A(n28), .Y(n184) );
  INVXLTS U114 ( .A(n28), .Y(n185) );
  INVXLTS U115 ( .A(n28), .Y(n186) );
  INVXLTS U116 ( .A(n28), .Y(n187) );
  INVXLTS U117 ( .A(n828), .Y(n188) );
  INVXLTS U118 ( .A(n188), .Y(n189) );
  INVXLTS U119 ( .A(n188), .Y(n190) );
  INVXLTS U120 ( .A(n188), .Y(n191) );
  XNOR2X1TS U180 ( .A(n1448), .B(n1447), .Y(n1545) );
  OR2XLTS U181 ( .A(n1691), .B(n119), .Y(n1666) );
  INVX2TS U182 ( .A(n1666), .Y(n257) );
  INVX2TS U183 ( .A(n1666), .Y(n258) );
  CLKBUFX2TS U184 ( .A(n1461), .Y(n259) );
  NAND3XLTS U185 ( .A(n259), .B(n1514), .C(n1488), .Y(n1366) );
  NAND2XLTS U186 ( .A(n259), .B(n1462), .Y(n1038) );
  XOR2XLTS U187 ( .A(n1448), .B(n998), .Y(n1461) );
  NAND2X1TS U188 ( .A(n1527), .B(n2385), .Y(n260) );
  OR2X2TS U189 ( .A(n272), .B(n292), .Y(n1592) );
  INVX2TS U190 ( .A(n1592), .Y(n261) );
  INVX2TS U191 ( .A(n1592), .Y(n262) );
  NAND2X1TS U192 ( .A(n289), .B(n2382), .Y(n263) );
  NAND2X1TS U193 ( .A(n289), .B(n2382), .Y(n264) );
  CLKBUFX2TS U194 ( .A(n1753), .Y(n265) );
  INVX2TS U195 ( .A(n1575), .Y(n266) );
  OR2X2TS U196 ( .A(n332), .B(n794), .Y(n1530) );
  INVX2TS U197 ( .A(n1530), .Y(n267) );
  INVX2TS U198 ( .A(n1530), .Y(n268) );
  OR2X2TS U199 ( .A(n824), .B(n308), .Y(n1108) );
  INVX2TS U200 ( .A(n1108), .Y(n269) );
  INVX2TS U201 ( .A(n1108), .Y(n270) );
  INVX2TS U202 ( .A(n1108), .Y(n271) );
  AOI21X1TS U203 ( .A0(n341), .A1(n1711), .B0(n2368), .Y(n1593) );
  INVX2TS U204 ( .A(n1593), .Y(n272) );
  INVX2TS U205 ( .A(n1593), .Y(n273) );
  INVX2TS U206 ( .A(n1593), .Y(n274) );
  OR2X2TS U207 ( .A(n337), .B(n259), .Y(n1372) );
  INVX2TS U208 ( .A(n1372), .Y(n275) );
  INVX2TS U209 ( .A(n1372), .Y(n276) );
  INVX2TS U210 ( .A(n1372), .Y(n277) );
  CLKBUFX2TS U211 ( .A(n1728), .Y(n278) );
  CLKBUFX2TS U212 ( .A(n1681), .Y(n279) );
  CLKBUFX2TS U213 ( .A(n1694), .Y(n280) );
  NOR2XLTS U214 ( .A(n1590), .B(n18), .Y(n1710) );
  CLKBUFX2TS U215 ( .A(n1662), .Y(n281) );
  AND2X2TS U216 ( .A(n300), .B(n2379), .Y(n1491) );
  INVX2TS U217 ( .A(n1491), .Y(n282) );
  INVX2TS U218 ( .A(n1491), .Y(n283) );
  OR2X2TS U219 ( .A(n310), .B(n116), .Y(n1110) );
  INVX2TS U220 ( .A(n1110), .Y(n284) );
  INVX2TS U221 ( .A(n1110), .Y(n285) );
  INVX2TS U222 ( .A(n1110), .Y(n286) );
  NAND2XLTS U223 ( .A(n1367), .B(n797), .Y(n287) );
  NAND2XLTS U224 ( .A(n1367), .B(n797), .Y(n288) );
  NAND2XLTS U225 ( .A(n1367), .B(n797), .Y(n1527) );
  AND2X2TS U226 ( .A(n1460), .B(n1038), .Y(n1369) );
  INVX2TS U227 ( .A(n1369), .Y(n289) );
  INVX2TS U228 ( .A(n1369), .Y(n290) );
  INVX2TS U229 ( .A(n1369), .Y(n291) );
  CLKBUFX2TS U230 ( .A(n1039), .Y(n292) );
  CLKBUFX2TS U231 ( .A(n1039), .Y(n293) );
  CLKBUFX2TS U232 ( .A(n1715), .Y(n294) );
  CLKBUFX2TS U233 ( .A(n1741), .Y(n295) );
  CLKBUFX2TS U234 ( .A(n1682), .Y(n296) );
  CLKBUFX2TS U235 ( .A(n1697), .Y(n297) );
  INVXLTS U236 ( .A(n1442), .Y(n299) );
  OAI22X1TS U237 ( .A0(n299), .A1(n119), .B0(n1447), .B1(n1448), .Y(n1450) );
  AND2XLTS U238 ( .A(n1245), .B(n329), .Y(n1489) );
  INVX2TS U239 ( .A(n1489), .Y(n300) );
  INVX2TS U240 ( .A(n1489), .Y(n301) );
  INVX2TS U241 ( .A(n1489), .Y(n302) );
  CLKBUFX2TS U242 ( .A(n794), .Y(n303) );
  CLKBUFX2TS U243 ( .A(n794), .Y(n304) );
  CLKBUFX2TS U244 ( .A(n1373), .Y(n306) );
  CLKBUFX2TS U245 ( .A(n1373), .Y(n307) );
  NOR2BXLTS U246 ( .AN(n1461), .B(n1546), .Y(n1373) );
  CLKBUFX2TS U247 ( .A(n137), .Y(n818) );
  INVX2TS U248 ( .A(n818), .Y(n308) );
  INVX2TS U249 ( .A(n818), .Y(n309) );
  INVX2TS U250 ( .A(n818), .Y(n310) );
  CLKBUFX2TS U251 ( .A(n1714), .Y(n311) );
  CLKBUFX2TS U252 ( .A(n1752), .Y(n312) );
  CLKBUFX2TS U253 ( .A(n1729), .Y(n313) );
  CLKBUFX2TS U254 ( .A(n1740), .Y(n314) );
  CLKBUFX2TS U255 ( .A(n1698), .Y(n315) );
  CLKBUFX2TS U256 ( .A(n835), .Y(n316) );
  CLKBUFX2TS U257 ( .A(n1447), .Y(n317) );
  NOR2XLTS U258 ( .A(n317), .B(n299), .Y(n1676) );
  CLKBUFX2TS U259 ( .A(n1376), .Y(n319) );
  CLKBUFX2TS U260 ( .A(n816), .Y(n320) );
  OAI31X1TS U261 ( .A0(n1689), .A1(n1676), .A2(n835), .B0(n2381), .Y(n1576) );
  INVXLTS U262 ( .A(n1109), .Y(n321) );
  AND2X2TS U263 ( .A(n154), .B(n2381), .Y(n1517) );
  INVX2TS U264 ( .A(n1517), .Y(n322) );
  INVX2TS U265 ( .A(n1517), .Y(n323) );
  AND2X2TS U266 ( .A(n157), .B(n2380), .Y(n1504) );
  INVX2TS U267 ( .A(n1504), .Y(n324) );
  INVX2TS U268 ( .A(n1504), .Y(n325) );
  AND2X2TS U269 ( .A(n853), .B(n2378), .Y(n1477) );
  INVX2TS U270 ( .A(n1477), .Y(n326) );
  INVX2TS U271 ( .A(n1477), .Y(n327) );
  INVX2TS U272 ( .A(n328), .Y(n329) );
  NAND3XLTS U273 ( .A(n329), .B(n1244), .C(n1234), .Y(n1190) );
  OR2X2TS U274 ( .A(n798), .B(n342), .Y(n1365) );
  INVX2TS U275 ( .A(n1365), .Y(n330) );
  INVX2TS U276 ( .A(n1365), .Y(n331) );
  INVX2TS U277 ( .A(n1365), .Y(n332) );
  INVX2TS U278 ( .A(n1365), .Y(n333) );
  AND2X1TS U279 ( .A(n1364), .B(n330), .Y(n1331) );
  CLKBUFX2TS U280 ( .A(n341), .Y(n812) );
  INVX2TS U281 ( .A(n812), .Y(n334) );
  INVX2TS U282 ( .A(n812), .Y(n335) );
  INVX2TS U283 ( .A(n812), .Y(n336) );
  INVX2TS U284 ( .A(n812), .Y(n337) );
  CLKAND2X2TS U285 ( .A(n1323), .B(n184), .Y(n1290) );
  AND2XLTS U286 ( .A(n1234), .B(n189), .Y(n1193) );
  INVX1TS U287 ( .A(n117), .Y(n824) );
  NAND2X1TS U288 ( .A(n2374), .B(n1003), .Y(n1693) );
  CLKBUFX2TS U289 ( .A(n1003), .Y(n2069) );
  CLKAND2X2TS U290 ( .A(n284), .B(n1109), .Y(n1043) );
  NAND2X1TS U291 ( .A(n1364), .B(n303), .Y(n1329) );
  NOR2X1TS U292 ( .A(n18), .B(n1690), .Y(n1462) );
  INVXLTS U293 ( .A(n2091), .Y(n2087) );
  OR2XLTS U294 ( .A(n813), .B(n1693), .Y(n338) );
  NAND2XLTS U295 ( .A(n1546), .B(n1439), .Y(n1475) );
  NAND2XLTS U296 ( .A(n1109), .B(n309), .Y(n1040) );
  NOR2XLTS U297 ( .A(n824), .B(n1546), .Y(n1377) );
  NAND2XLTS U298 ( .A(n145), .B(n1449), .Y(n1451) );
  NAND3XLTS U299 ( .A(n1284), .B(n1285), .C(n1282), .Y(n1246) );
  OA22XLTS U300 ( .A0(n1546), .A1(n824), .B0(n1679), .B1(n1439), .Y(n1421) );
  INVXLTS U301 ( .A(n1366), .Y(n794) );
  NAND2XLTS U302 ( .A(n1473), .B(n137), .Y(n1041) );
  OAI21XLTS U303 ( .A0(n1439), .A1(n1440), .B0(n813), .Y(n1432) );
  NOR2XLTS U304 ( .A(n1545), .B(n1690), .Y(n1449) );
  NOR2XLTS U305 ( .A(n1440), .B(n119), .Y(n1437) );
  AOI22XLTS U306 ( .A0(n1766), .A1(n695), .B0(n679), .B1(n1765), .Y(n1251) );
  AOI22XLTS U307 ( .A0(n1768), .A1(n696), .B0(n679), .B1(n1767), .Y(n1252) );
  AOI22XLTS U308 ( .A0(n1770), .A1(n696), .B0(n679), .B1(n1769), .Y(n1253) );
  AOI22XLTS U309 ( .A0(n1774), .A1(n693), .B0(n678), .B1(n1773), .Y(n1255) );
  AOI22XLTS U310 ( .A0(n1776), .A1(n693), .B0(n678), .B1(n1775), .Y(n1256) );
  AOI22XLTS U311 ( .A0(n1778), .A1(n693), .B0(n678), .B1(n1777), .Y(n1257) );
  AOI22XLTS U312 ( .A0(n1782), .A1(n692), .B0(n677), .B1(n1781), .Y(n1259) );
  AOI22XLTS U313 ( .A0(n1784), .A1(n692), .B0(n677), .B1(n1783), .Y(n1260) );
  AOI22XLTS U314 ( .A0(n1786), .A1(n692), .B0(n677), .B1(n1785), .Y(n1261) );
  AOI22XLTS U315 ( .A0(n1790), .A1(n691), .B0(n682), .B1(n1789), .Y(n1263) );
  AOI22XLTS U316 ( .A0(n1792), .A1(n691), .B0(n680), .B1(n1791), .Y(n1264) );
  AOI22XLTS U317 ( .A0(n1794), .A1(n691), .B0(n685), .B1(n1793), .Y(n1265) );
  AOI22XLTS U318 ( .A0(n1798), .A1(n690), .B0(n682), .B1(n1797), .Y(n1267) );
  AOI22XLTS U319 ( .A0(n1800), .A1(n690), .B0(n682), .B1(n1799), .Y(n1268) );
  AOI22XLTS U320 ( .A0(n1802), .A1(n690), .B0(n681), .B1(n1801), .Y(n1269) );
  AOI22XLTS U321 ( .A0(n1806), .A1(n689), .B0(n683), .B1(n1805), .Y(n1271) );
  AOI22XLTS U322 ( .A0(n1808), .A1(n689), .B0(n683), .B1(n1807), .Y(n1272) );
  AOI22XLTS U323 ( .A0(n1810), .A1(n689), .B0(n683), .B1(n1809), .Y(n1273) );
  AOI22XLTS U324 ( .A0(n1814), .A1(n688), .B0(n681), .B1(n1813), .Y(n1275) );
  AOI22XLTS U325 ( .A0(n1816), .A1(n688), .B0(n683), .B1(n1815), .Y(n1276) );
  AOI22XLTS U326 ( .A0(n1818), .A1(n688), .B0(n680), .B1(n1817), .Y(n1277) );
  AOI22XLTS U327 ( .A0(n1822), .A1(n687), .B0(n684), .B1(n1821), .Y(n1279) );
  AOI22XLTS U328 ( .A0(n1824), .A1(n687), .B0(n684), .B1(n1823), .Y(n1280) );
  AOI22XLTS U329 ( .A0(n1826), .A1(n687), .B0(n684), .B1(n1825), .Y(n1281) );
  AOI22XLTS U330 ( .A0(n2308), .A1(n2033), .B0(n2188), .B1(n2011), .Y(n1028)
         );
  AOI22XLTS U331 ( .A0(n2311), .A1(n2033), .B0(n2191), .B1(n2011), .Y(n1029)
         );
  AOI22XLTS U332 ( .A0(n2317), .A1(n2031), .B0(n2197), .B1(n2010), .Y(n1031)
         );
  AOI22XLTS U333 ( .A0(n2320), .A1(n2031), .B0(n2200), .B1(n2010), .Y(n1032)
         );
  AOI22XLTS U334 ( .A0(n2323), .A1(n2031), .B0(n2203), .B1(n2010), .Y(n1033)
         );
  AOI22XLTS U335 ( .A0(n2326), .A1(n2029), .B0(n2206), .B1(n2009), .Y(n1034)
         );
  AOI22XLTS U336 ( .A0(n2329), .A1(n2029), .B0(n2209), .B1(n2009), .Y(n1035)
         );
  AOI22XLTS U337 ( .A0(n2332), .A1(n2029), .B0(n2212), .B1(n2009), .Y(n1036)
         );
  AOI22XLTS U338 ( .A0(n914), .A1(n2257), .B0(n903), .B1(n2137), .Y(n1049) );
  AOI22XLTS U339 ( .A0(n914), .A1(n2260), .B0(n903), .B1(n2140), .Y(n1050) );
  AOI22XLTS U340 ( .A0(n914), .A1(n2263), .B0(n903), .B1(n2143), .Y(n1051) );
  AOI22XLTS U341 ( .A0(n2269), .A1(n2039), .B0(n2149), .B1(n2015), .Y(n1015)
         );
  AOI22XLTS U342 ( .A0(n2272), .A1(n2039), .B0(n2152), .B1(n2015), .Y(n1016)
         );
  AOI22XLTS U343 ( .A0(n2275), .A1(n2039), .B0(n2155), .B1(n2015), .Y(n1017)
         );
  AOI22XLTS U344 ( .A0(n2281), .A1(n2037), .B0(n2161), .B1(n2013), .Y(n1019)
         );
  AOI22XLTS U345 ( .A0(n2284), .A1(n2037), .B0(n2164), .B1(n2013), .Y(n1020)
         );
  AOI22XLTS U346 ( .A0(n2287), .A1(n2037), .B0(n2167), .B1(n2013), .Y(n1021)
         );
  AOI22XLTS U347 ( .A0(n2293), .A1(n2035), .B0(n2173), .B1(n2012), .Y(n1023)
         );
  AOI22XLTS U348 ( .A0(n2296), .A1(n2035), .B0(n2176), .B1(n2012), .Y(n1024)
         );
  AOI22XLTS U349 ( .A0(n2299), .A1(n2035), .B0(n2179), .B1(n2012), .Y(n1025)
         );
  AOI22XLTS U350 ( .A0(n2302), .A1(n2033), .B0(n2182), .B1(n2011), .Y(n1026)
         );
  AOI22XLTS U351 ( .A0(n915), .A1(n2242), .B0(n904), .B1(n2122), .Y(n1042) );
  AOI22XLTS U352 ( .A0(n915), .A1(n2245), .B0(n904), .B1(n2125), .Y(n1045) );
  AOI22XLTS U353 ( .A0(n915), .A1(n2248), .B0(n904), .B1(n2128), .Y(n1046) );
  AOI22XLTS U354 ( .A0(n913), .A1(n2269), .B0(n902), .B1(n2149), .Y(n1053) );
  AOI22XLTS U355 ( .A0(n913), .A1(n2272), .B0(n902), .B1(n2152), .Y(n1054) );
  AOI22XLTS U356 ( .A0(n913), .A1(n2275), .B0(n902), .B1(n2155), .Y(n1055) );
  AOI22XLTS U357 ( .A0(n917), .A1(n2281), .B0(n901), .B1(n2161), .Y(n1057) );
  AOI22XLTS U358 ( .A0(n917), .A1(n2284), .B0(n901), .B1(n2164), .Y(n1058) );
  AOI22XLTS U359 ( .A0(n918), .A1(n2287), .B0(n901), .B1(n2167), .Y(n1059) );
  AOI22XLTS U360 ( .A0(n912), .A1(n2293), .B0(n900), .B1(n2173), .Y(n1061) );
  AOI22XLTS U361 ( .A0(n912), .A1(n2296), .B0(n900), .B1(n2176), .Y(n1062) );
  AOI22XLTS U362 ( .A0(n912), .A1(n2299), .B0(n900), .B1(n2179), .Y(n1063) );
  AOI22XLTS U363 ( .A0(n911), .A1(n2305), .B0(n906), .B1(n2185), .Y(n1065) );
  AOI22XLTS U364 ( .A0(n911), .A1(n2308), .B0(n907), .B1(n2188), .Y(n1066) );
  AOI22XLTS U365 ( .A0(n911), .A1(n2311), .B0(n907), .B1(n2191), .Y(n1067) );
  AOI22XLTS U366 ( .A0(n909), .A1(n2317), .B0(n899), .B1(n2197), .Y(n1069) );
  AOI22XLTS U367 ( .A0(n909), .A1(n2323), .B0(n899), .B1(n2203), .Y(n1071) );
  AOI22XLTS U368 ( .A0(n908), .A1(n2326), .B0(n898), .B1(n2206), .Y(n1104) );
  AOI22XLTS U369 ( .A0(n908), .A1(n2329), .B0(n898), .B1(n2209), .Y(n1105) );
  AOI22XLTS U370 ( .A0(n908), .A1(n2332), .B0(n898), .B1(n2212), .Y(n1106) );
  AOI22XLTS U371 ( .A0(n2245), .A1(n2045), .B0(n2125), .B1(n2019), .Y(n1007)
         );
  AOI22XLTS U372 ( .A0(n2248), .A1(n2047), .B0(n2128), .B1(n2019), .Y(n1008)
         );
  AOI22XLTS U373 ( .A0(n2251), .A1(n2047), .B0(n2131), .B1(n2019), .Y(n1009)
         );
  AOI22XLTS U374 ( .A0(n2257), .A1(n2041), .B0(n2137), .B1(n2017), .Y(n1011)
         );
  AOI22XLTS U375 ( .A0(n2260), .A1(n2041), .B0(n2140), .B1(n2017), .Y(n1012)
         );
  AOI22XLTS U376 ( .A0(n2263), .A1(n2041), .B0(n2143), .B1(n2017), .Y(n1013)
         );
  AOI22XLTS U377 ( .A0(n909), .A1(n2320), .B0(n899), .B1(n2200), .Y(n1070) );
  AND2XLTS U378 ( .A(n1540), .B(n1450), .Y(n1488) );
  INVXLTS U379 ( .A(cacheDataOut_A[0]), .Y(n950) );
  INVXLTS U380 ( .A(cacheDataOut_A[1]), .Y(n949) );
  INVXLTS U381 ( .A(cacheDataOut_A[2]), .Y(n948) );
  INVXLTS U382 ( .A(cacheDataOut_A[3]), .Y(n947) );
  INVXLTS U383 ( .A(cacheDataOut_A[4]), .Y(n946) );
  INVXLTS U384 ( .A(cacheDataOut_A[5]), .Y(n945) );
  INVXLTS U385 ( .A(cacheDataOut_A[6]), .Y(n944) );
  INVXLTS U386 ( .A(cacheDataOut_A[7]), .Y(n943) );
  INVXLTS U387 ( .A(cacheDataOut_A[8]), .Y(n942) );
  INVXLTS U388 ( .A(cacheDataOut_A[9]), .Y(n941) );
  INVXLTS U389 ( .A(cacheDataOut_A[10]), .Y(n940) );
  INVXLTS U390 ( .A(cacheDataOut_A[11]), .Y(n939) );
  INVXLTS U391 ( .A(cacheDataOut_A[12]), .Y(n938) );
  INVXLTS U392 ( .A(cacheDataOut_A[13]), .Y(n937) );
  INVXLTS U393 ( .A(cacheDataOut_A[14]), .Y(n936) );
  INVXLTS U394 ( .A(cacheDataOut_A[15]), .Y(n935) );
  INVXLTS U395 ( .A(cacheDataOut_A[16]), .Y(n934) );
  INVXLTS U396 ( .A(cacheDataOut_A[17]), .Y(n933) );
  INVXLTS U397 ( .A(cacheDataOut_A[18]), .Y(n932) );
  INVXLTS U398 ( .A(cacheDataOut_A[19]), .Y(n931) );
  INVXLTS U399 ( .A(cacheDataOut_A[20]), .Y(n930) );
  INVXLTS U400 ( .A(cacheDataOut_A[21]), .Y(n929) );
  INVXLTS U401 ( .A(cacheDataOut_A[22]), .Y(n928) );
  INVXLTS U402 ( .A(cacheDataOut_A[23]), .Y(n927) );
  INVXLTS U403 ( .A(cacheDataOut_A[24]), .Y(n926) );
  INVXLTS U404 ( .A(cacheDataOut_A[25]), .Y(n925) );
  INVXLTS U405 ( .A(cacheDataOut_A[26]), .Y(n924) );
  INVXLTS U406 ( .A(cacheDataOut_A[27]), .Y(n923) );
  INVXLTS U407 ( .A(cacheDataOut_A[28]), .Y(n922) );
  INVXLTS U408 ( .A(cacheDataOut_A[29]), .Y(n921) );
  INVXLTS U409 ( .A(cacheDataOut_A[30]), .Y(n920) );
  INVXLTS U410 ( .A(cacheDataOut_A[31]), .Y(n919) );
  OAI222XLTS U411 ( .A0(n2021), .A1(n2218), .B0(n1692), .B1(n2338), .C0(n2069), 
        .C1(n774), .Y(n3191) );
  OAI222XLTS U412 ( .A0(n2021), .A1(n2219), .B0(n127), .B1(n2339), .C0(n2069), 
        .C1(n773), .Y(n3192) );
  OAI222XLTS U413 ( .A0(n2023), .A1(n2221), .B0(n1692), .B1(n2341), .C0(n2061), 
        .C1(n772), .Y(n3194) );
  OAI222XLTS U414 ( .A0(n2021), .A1(n2220), .B0(n127), .B1(n2340), .C0(n2063), 
        .C1(n771), .Y(n3193) );
  OAI222XLTS U415 ( .A0(n2023), .A1(n2222), .B0(n1692), .B1(n2342), .C0(n2067), 
        .C1(n770), .Y(n3195) );
  OAI222XLTS U416 ( .A0(n2023), .A1(n2223), .B0(n127), .B1(n2343), .C0(n2071), 
        .C1(n769), .Y(n3196) );
  OAI22XLTS U417 ( .A0(n1368), .A1(n44), .B0(n1463), .B1(n321), .Y(n3333) );
  INVXLTS U418 ( .A(memRead_EAST), .Y(n844) );
  CLKBUFX2TS U419 ( .A(n557), .Y(n552) );
  CLKBUFX2TS U420 ( .A(n557), .Y(n553) );
  CLKBUFX2TS U421 ( .A(n556), .Y(n554) );
  CLKBUFX2TS U422 ( .A(n477), .Y(n475) );
  NOR2X1TS U423 ( .A(n1573), .B(n1451), .Y(n1578) );
  NOR2X1TS U424 ( .A(n2363), .B(n293), .Y(n1446) );
  NOR4X1TS U425 ( .A(n556), .B(n258), .C(n835), .D(n1676), .Y(n1663) );
  INVX1TS U426 ( .A(n1189), .Y(n795) );
  NOR4XLTS U427 ( .A(n1661), .B(n339), .C(n476), .D(n281), .Y(n1553) );
  CLKBUFX2TS U428 ( .A(n1039), .Y(n341) );
  XNOR2X1TS U429 ( .A(n1542), .B(n1543), .Y(n1514) );
  OAI2BB1XLTS U430 ( .A0N(n145), .A1N(n1541), .B0(n1544), .Y(n1542) );
  OAI21XLTS U431 ( .A0(n1541), .A1(n144), .B0(n318), .Y(n1544) );
  NAND2XLTS U432 ( .A(n1486), .B(n820), .Y(n1115) );
  NOR2X1TS U433 ( .A(n833), .B(n299), .Y(n1662) );
  NOR2X1TS U434 ( .A(n1), .B(n26), .Y(n1725) );
  NOR2X1TS U435 ( .A(n828), .B(n123), .Y(n989) );
  AOI21X1TS U436 ( .A0(n190), .A1(n9), .B0(n184), .Y(n1284) );
  INVXLTS U437 ( .A(cacheDataOut_B[0]), .Y(n982) );
  INVXLTS U438 ( .A(cacheDataOut_B[1]), .Y(n981) );
  INVXLTS U439 ( .A(cacheDataOut_B[2]), .Y(n980) );
  INVXLTS U440 ( .A(cacheDataOut_B[3]), .Y(n979) );
  INVXLTS U441 ( .A(cacheDataOut_B[4]), .Y(n978) );
  INVXLTS U442 ( .A(cacheDataOut_B[5]), .Y(n977) );
  INVXLTS U443 ( .A(cacheDataOut_B[6]), .Y(n976) );
  INVXLTS U444 ( .A(cacheDataOut_B[7]), .Y(n975) );
  INVXLTS U445 ( .A(cacheDataOut_B[8]), .Y(n974) );
  INVXLTS U446 ( .A(cacheDataOut_B[9]), .Y(n973) );
  INVXLTS U447 ( .A(cacheDataOut_B[10]), .Y(n972) );
  INVXLTS U448 ( .A(cacheDataOut_B[11]), .Y(n971) );
  INVXLTS U449 ( .A(cacheDataOut_B[12]), .Y(n970) );
  INVXLTS U450 ( .A(cacheDataOut_B[13]), .Y(n969) );
  INVXLTS U451 ( .A(cacheDataOut_B[14]), .Y(n968) );
  INVXLTS U452 ( .A(cacheDataOut_B[15]), .Y(n967) );
  INVXLTS U453 ( .A(cacheDataOut_B[16]), .Y(n966) );
  INVXLTS U454 ( .A(cacheDataOut_B[17]), .Y(n965) );
  INVXLTS U455 ( .A(cacheDataOut_B[18]), .Y(n964) );
  INVXLTS U456 ( .A(cacheDataOut_B[19]), .Y(n963) );
  INVXLTS U457 ( .A(cacheDataOut_B[20]), .Y(n962) );
  INVXLTS U458 ( .A(cacheDataOut_B[21]), .Y(n961) );
  INVXLTS U459 ( .A(cacheDataOut_B[22]), .Y(n960) );
  INVXLTS U460 ( .A(cacheDataOut_B[23]), .Y(n959) );
  INVXLTS U461 ( .A(cacheDataOut_B[24]), .Y(n958) );
  INVXLTS U462 ( .A(cacheDataOut_B[25]), .Y(n957) );
  INVXLTS U463 ( .A(cacheDataOut_B[26]), .Y(n956) );
  INVXLTS U464 ( .A(cacheDataOut_B[27]), .Y(n955) );
  INVXLTS U465 ( .A(cacheDataOut_B[28]), .Y(n954) );
  INVXLTS U466 ( .A(cacheDataOut_B[29]), .Y(n953) );
  INVXLTS U467 ( .A(cacheDataOut_B[30]), .Y(n952) );
  INVXLTS U468 ( .A(cacheDataOut_B[31]), .Y(n951) );
  NOR2X1TS U469 ( .A(memRead_WEST), .B(memWrite_WEST), .Y(n1690) );
  NOR2X1TS U470 ( .A(memRead_EAST), .B(memWrite_EAST), .Y(n1443) );
  NOR2X1TS U471 ( .A(memRead_NORTH), .B(memWrite_NORTH), .Y(n1447) );
  AOI21XLTS U472 ( .A0(memRead_NORTH), .A1(n821), .B0(memRead_SOUTH), .Y(n1441) );
  OA22XLTS U473 ( .A0(n281), .A1(memWrite_NORTH), .B0(n832), .B1(
        memWrite_SOUTH), .Y(n1713) );
  AOI22XLTS U474 ( .A0(n258), .A1(memWrite_EAST), .B0(memWrite_SOUTH), .B1(
        n831), .Y(n1665) );
  NOR2X1TS U475 ( .A(n3677), .B(n3678), .Y(n1723) );
  AOI21XLTS U476 ( .A0(memRead_NORTH), .A1(n1426), .B0(memRead_SOUTH), .Y(
        n1425) );
  CLKBUFX2TS U477 ( .A(n4621), .Y(n342) );
  INVX2TS U478 ( .A(n1693), .Y(n806) );
  INVX2TS U479 ( .A(n2021), .Y(n2019) );
  INVX2TS U480 ( .A(n2023), .Y(n2017) );
  CLKBUFX2TS U481 ( .A(n2027), .Y(n2021) );
  CLKBUFX2TS U482 ( .A(n2027), .Y(n2023) );
  INVX2TS U483 ( .A(n2025), .Y(n2010) );
  INVX2TS U484 ( .A(n2027), .Y(n2009) );
  INVX2TS U485 ( .A(n2025), .Y(n2015) );
  CLKBUFX2TS U486 ( .A(n2027), .Y(n2025) );
  INVX2TS U487 ( .A(n2025), .Y(n2013) );
  INVX2TS U488 ( .A(n338), .Y(n2012) );
  INVX2TS U489 ( .A(n2025), .Y(n2011) );
  INVX2TS U490 ( .A(n2380), .Y(n2365) );
  CLKBUFX2TS U491 ( .A(n2067), .Y(n2051) );
  CLKBUFX2TS U492 ( .A(n2067), .Y(n2049) );
  CLKBUFX2TS U493 ( .A(n2061), .Y(n2057) );
  CLKBUFX2TS U494 ( .A(n2063), .Y(n2055) );
  CLKBUFX2TS U495 ( .A(n2063), .Y(n2053) );
  CLKBUFX2TS U496 ( .A(n2061), .Y(n2059) );
  INVX2TS U497 ( .A(n552), .Y(n541) );
  INVX2TS U498 ( .A(n2375), .Y(n2370) );
  INVX2TS U499 ( .A(n2374), .Y(n2371) );
  INVX2TS U500 ( .A(n2373), .Y(n2372) );
  INVX2TS U501 ( .A(n2373), .Y(n2362) );
  INVX2TS U502 ( .A(n2382), .Y(n2363) );
  INVX2TS U503 ( .A(n489), .Y(n486) );
  INVX2TS U504 ( .A(n490), .Y(n485) );
  INVX2TS U505 ( .A(n491), .Y(n484) );
  INVX2TS U506 ( .A(n492), .Y(n483) );
  INVX2TS U507 ( .A(n493), .Y(n482) );
  INVX2TS U508 ( .A(n494), .Y(n481) );
  INVX2TS U509 ( .A(n495), .Y(n480) );
  INVX2TS U510 ( .A(n497), .Y(n479) );
  INVX2TS U511 ( .A(n496), .Y(n478) );
  INVX2TS U512 ( .A(n552), .Y(n542) );
  INVX2TS U513 ( .A(n552), .Y(n543) );
  INVX2TS U514 ( .A(n553), .Y(n544) );
  INVX2TS U515 ( .A(n553), .Y(n545) );
  INVX2TS U516 ( .A(n554), .Y(n546) );
  INVX2TS U517 ( .A(n554), .Y(n547) );
  INVX2TS U518 ( .A(n554), .Y(n548) );
  INVX2TS U519 ( .A(n556), .Y(n550) );
  INVX2TS U520 ( .A(n556), .Y(n549) );
  INVX2TS U521 ( .A(n2377), .Y(n2368) );
  INVX2TS U522 ( .A(n553), .Y(n551) );
  INVX2TS U523 ( .A(n2379), .Y(n2366) );
  INVX2TS U524 ( .A(n2378), .Y(n2367) );
  INVX2TS U525 ( .A(n2376), .Y(n2369) );
  INVX2TS U526 ( .A(n2381), .Y(n2364) );
  NOR2X1TS U527 ( .A(n2362), .B(n1250), .Y(n1282) );
  CLKBUFX2TS U528 ( .A(n916), .Y(n915) );
  CLKBUFX2TS U529 ( .A(n916), .Y(n914) );
  CLKBUFX2TS U530 ( .A(n917), .Y(n913) );
  CLKBUFX2TS U531 ( .A(n1043), .Y(n912) );
  CLKBUFX2TS U532 ( .A(n916), .Y(n911) );
  CLKBUFX2TS U533 ( .A(n918), .Y(n909) );
  CLKBUFX2TS U534 ( .A(n918), .Y(n908) );
  CLKBUFX2TS U535 ( .A(n905), .Y(n904) );
  CLKBUFX2TS U536 ( .A(n905), .Y(n903) );
  CLKBUFX2TS U537 ( .A(n906), .Y(n902) );
  CLKBUFX2TS U538 ( .A(n906), .Y(n901) );
  CLKBUFX2TS U539 ( .A(n907), .Y(n900) );
  CLKBUFX2TS U540 ( .A(n1044), .Y(n899) );
  CLKBUFX2TS U541 ( .A(n905), .Y(n898) );
  CLKBUFX2TS U542 ( .A(n704), .Y(n703) );
  CLKBUFX2TS U543 ( .A(n704), .Y(n702) );
  CLKBUFX2TS U544 ( .A(n705), .Y(n701) );
  CLKBUFX2TS U545 ( .A(n705), .Y(n700) );
  CLKBUFX2TS U546 ( .A(n706), .Y(n699) );
  CLKBUFX2TS U547 ( .A(n706), .Y(n698) );
  CLKBUFX2TS U548 ( .A(n706), .Y(n697) );
  CLKBUFX2TS U549 ( .A(n2383), .Y(n2380) );
  CLKBUFX2TS U550 ( .A(n2069), .Y(n2067) );
  CLKBUFX2TS U551 ( .A(n2069), .Y(n2065) );
  CLKBUFX2TS U552 ( .A(n2071), .Y(n2061) );
  CLKBUFX2TS U553 ( .A(n2071), .Y(n2063) );
  CLKBUFX2TS U554 ( .A(n680), .Y(n679) );
  CLKBUFX2TS U555 ( .A(n681), .Y(n678) );
  CLKBUFX2TS U556 ( .A(n681), .Y(n677) );
  CLKBUFX2TS U557 ( .A(n338), .Y(n2027) );
  CLKBUFX2TS U558 ( .A(n537), .Y(n535) );
  CLKBUFX2TS U559 ( .A(n537), .Y(n534) );
  CLKBUFX2TS U560 ( .A(n1384), .Y(n533) );
  CLKBUFX2TS U561 ( .A(n538), .Y(n532) );
  CLKBUFX2TS U562 ( .A(n538), .Y(n531) );
  CLKBUFX2TS U563 ( .A(n539), .Y(n530) );
  CLKBUFX2TS U564 ( .A(n539), .Y(n529) );
  CLKBUFX2TS U565 ( .A(n540), .Y(n536) );
  CLKBUFX2TS U566 ( .A(n447), .Y(n440) );
  CLKBUFX2TS U567 ( .A(n449), .Y(n441) );
  CLKBUFX2TS U568 ( .A(n449), .Y(n442) );
  CLKBUFX2TS U569 ( .A(n514), .Y(n505) );
  CLKBUFX2TS U570 ( .A(n511), .Y(n506) );
  CLKBUFX2TS U571 ( .A(n511), .Y(n507) );
  CLKBUFX2TS U572 ( .A(n510), .Y(n508) );
  CLKBUFX2TS U573 ( .A(n510), .Y(n509) );
  INVX2TS U574 ( .A(n2089), .Y(n2075) );
  INVX2TS U575 ( .A(n2089), .Y(n2073) );
  INVX2TS U576 ( .A(n340), .Y(n2085) );
  INVX2TS U577 ( .A(n2091), .Y(n2083) );
  INVX2TS U578 ( .A(n2089), .Y(n2081) );
  INVX2TS U579 ( .A(n340), .Y(n2079) );
  INVX2TS U580 ( .A(n2089), .Y(n2077) );
  CLKBUFX2TS U581 ( .A(n2385), .Y(n2373) );
  CLKBUFX2TS U582 ( .A(n2385), .Y(n2375) );
  CLKBUFX2TS U583 ( .A(n2385), .Y(n2374) );
  CLKBUFX2TS U584 ( .A(n2383), .Y(n2381) );
  CLKBUFX2TS U585 ( .A(n557), .Y(n555) );
  CLKBUFX2TS U586 ( .A(n459), .Y(n452) );
  CLKBUFX2TS U587 ( .A(n461), .Y(n453) );
  CLKBUFX2TS U588 ( .A(n461), .Y(n454) );
  CLKBUFX2TS U589 ( .A(n460), .Y(n455) );
  CLKBUFX2TS U590 ( .A(n460), .Y(n456) );
  CLKBUFX2TS U591 ( .A(n459), .Y(n457) );
  CLKBUFX2TS U592 ( .A(n459), .Y(n458) );
  CLKBUFX2TS U593 ( .A(n1552), .Y(n428) );
  CLKBUFX2TS U594 ( .A(n438), .Y(n429) );
  CLKBUFX2TS U595 ( .A(n438), .Y(n430) );
  CLKBUFX2TS U596 ( .A(n437), .Y(n431) );
  CLKBUFX2TS U597 ( .A(n437), .Y(n432) );
  CLKBUFX2TS U598 ( .A(n439), .Y(n433) );
  CLKBUFX2TS U599 ( .A(n448), .Y(n443) );
  CLKBUFX2TS U600 ( .A(n448), .Y(n444) );
  CLKBUFX2TS U601 ( .A(n447), .Y(n445) );
  CLKBUFX2TS U602 ( .A(n447), .Y(n446) );
  CLKBUFX2TS U603 ( .A(n436), .Y(n434) );
  CLKBUFX2TS U604 ( .A(n436), .Y(n435) );
  CLKBUFX2TS U605 ( .A(n2106), .Y(n2102) );
  CLKBUFX2TS U606 ( .A(n2106), .Y(n2101) );
  CLKBUFX2TS U607 ( .A(n2107), .Y(n2094) );
  CLKBUFX2TS U608 ( .A(n2107), .Y(n2099) );
  INVX2TS U609 ( .A(n474), .Y(n464) );
  INVX2TS U610 ( .A(n476), .Y(n472) );
  INVX2TS U611 ( .A(n476), .Y(n473) );
  INVX2TS U612 ( .A(n475), .Y(n465) );
  INVX2TS U613 ( .A(n474), .Y(n466) );
  INVX2TS U614 ( .A(n474), .Y(n467) );
  INVX2TS U615 ( .A(n474), .Y(n468) );
  INVX2TS U616 ( .A(n475), .Y(n469) );
  INVX2TS U617 ( .A(n475), .Y(n470) );
  INVX2TS U618 ( .A(n475), .Y(n471) );
  CLKBUFX2TS U619 ( .A(n2384), .Y(n2376) );
  CLKBUFX2TS U620 ( .A(n2384), .Y(n2377) );
  CLKBUFX2TS U621 ( .A(n2383), .Y(n2382) );
  CLKBUFX2TS U622 ( .A(n502), .Y(n489) );
  CLKBUFX2TS U623 ( .A(n502), .Y(n490) );
  CLKBUFX2TS U624 ( .A(n501), .Y(n494) );
  CLKBUFX2TS U625 ( .A(n502), .Y(n492) );
  CLKBUFX2TS U626 ( .A(n501), .Y(n493) );
  CLKBUFX2TS U627 ( .A(n501), .Y(n495) );
  CLKBUFX2TS U628 ( .A(n500), .Y(n496) );
  CLKBUFX2TS U629 ( .A(n500), .Y(n497) );
  CLKBUFX2TS U630 ( .A(n502), .Y(n491) );
  CLKBUFX2TS U631 ( .A(n500), .Y(n498) );
  CLKBUFX2TS U632 ( .A(n500), .Y(n499) );
  INVX2TS U633 ( .A(n488), .Y(n487) );
  CLKBUFX2TS U634 ( .A(n2384), .Y(n2378) );
  CLKBUFX2TS U635 ( .A(n2384), .Y(n2379) );
  NOR2BX1TS U636 ( .AN(n1115), .B(n2368), .Y(n1186) );
  NOR2X1TS U637 ( .A(n2363), .B(n1332), .Y(n1364) );
  CLKBUFX2TS U638 ( .A(n1247), .Y(n704) );
  CLKBUFX2TS U639 ( .A(n1247), .Y(n705) );
  CLKBUFX2TS U640 ( .A(n1247), .Y(n706) );
  CLKBUFX2TS U641 ( .A(n1044), .Y(n905) );
  CLKBUFX2TS U642 ( .A(n1043), .Y(n916) );
  CLKBUFX2TS U643 ( .A(n1044), .Y(n906) );
  CLKBUFX2TS U644 ( .A(n1043), .Y(n917) );
  CLKBUFX2TS U645 ( .A(n1044), .Y(n907) );
  CLKBUFX2TS U646 ( .A(n1043), .Y(n918) );
  CLKBUFX2TS U647 ( .A(n695), .Y(n693) );
  CLKBUFX2TS U648 ( .A(n694), .Y(n692) );
  CLKBUFX2TS U649 ( .A(n694), .Y(n691) );
  CLKBUFX2TS U650 ( .A(n695), .Y(n690) );
  CLKBUFX2TS U651 ( .A(n695), .Y(n689) );
  CLKBUFX2TS U652 ( .A(n696), .Y(n688) );
  CLKBUFX2TS U653 ( .A(n696), .Y(n687) );
  CLKBUFX2TS U654 ( .A(n1717), .Y(n1660) );
  CLKBUFX2TS U655 ( .A(n1717), .Y(n1589) );
  CLKBUFX2TS U656 ( .A(n2008), .Y(n1518) );
  CLKBUFX2TS U657 ( .A(n2007), .Y(n1515) );
  CLKBUFX2TS U658 ( .A(n2007), .Y(n1505) );
  CLKBUFX2TS U659 ( .A(n2008), .Y(n1502) );
  CLKBUFX2TS U660 ( .A(n2008), .Y(n1492) );
  CLKBUFX2TS U661 ( .A(n585), .Y(n584) );
  CLKBUFX2TS U662 ( .A(n585), .Y(n583) );
  CLKBUFX2TS U663 ( .A(n586), .Y(n582) );
  CLKBUFX2TS U664 ( .A(n586), .Y(n581) );
  CLKBUFX2TS U665 ( .A(n587), .Y(n580) );
  CLKBUFX2TS U666 ( .A(n585), .Y(n579) );
  CLKBUFX2TS U667 ( .A(n586), .Y(n578) );
  NAND2X1TS U668 ( .A(n1374), .B(n2377), .Y(n1464) );
  CLKBUFX2TS U669 ( .A(n477), .Y(n476) );
  CLKBUFX2TS U670 ( .A(n515), .Y(n514) );
  CLKBUFX2TS U671 ( .A(n515), .Y(n513) );
  CLKBUFX2TS U672 ( .A(n515), .Y(n512) );
  CLKBUFX2TS U673 ( .A(n540), .Y(n538) );
  CLKBUFX2TS U674 ( .A(n1384), .Y(n539) );
  CLKBUFX2TS U675 ( .A(n450), .Y(n449) );
  CLKBUFX2TS U676 ( .A(n685), .Y(n682) );
  CLKBUFX2TS U677 ( .A(n685), .Y(n683) );
  CLKBUFX2TS U678 ( .A(n540), .Y(n537) );
  CLKBUFX2TS U679 ( .A(n516), .Y(n511) );
  CLKBUFX2TS U680 ( .A(n516), .Y(n510) );
  CLKBUFX2TS U681 ( .A(n686), .Y(n680) );
  CLKBUFX2TS U682 ( .A(n686), .Y(n681) );
  CLKBUFX2TS U683 ( .A(n339), .Y(n556) );
  CLKBUFX2TS U684 ( .A(n2047), .Y(n2031) );
  CLKBUFX2TS U685 ( .A(n2047), .Y(n2029) );
  CLKBUFX2TS U686 ( .A(n426), .Y(n416) );
  CLKBUFX2TS U687 ( .A(n425), .Y(n417) );
  CLKBUFX2TS U688 ( .A(n425), .Y(n418) );
  CLKBUFX2TS U689 ( .A(n424), .Y(n419) );
  CLKBUFX2TS U690 ( .A(n424), .Y(n420) );
  CLKBUFX2TS U691 ( .A(n423), .Y(n421) );
  CLKBUFX2TS U692 ( .A(n423), .Y(n422) );
  CLKBUFX2TS U693 ( .A(n2045), .Y(n2041) );
  CLKBUFX2TS U694 ( .A(n2043), .Y(n2039) );
  CLKBUFX2TS U695 ( .A(n2043), .Y(n2037) );
  CLKBUFX2TS U696 ( .A(n2045), .Y(n2035) );
  CLKBUFX2TS U697 ( .A(n2045), .Y(n2033) );
  CLKBUFX2TS U698 ( .A(n564), .Y(n563) );
  CLKBUFX2TS U699 ( .A(n565), .Y(n562) );
  CLKBUFX2TS U700 ( .A(n565), .Y(n561) );
  CLKBUFX2TS U701 ( .A(n565), .Y(n560) );
  CLKBUFX2TS U702 ( .A(n566), .Y(n559) );
  CLKBUFX2TS U703 ( .A(n566), .Y(n558) );
  CLKBUFX2TS U704 ( .A(n1003), .Y(n2071) );
  CLKBUFX2TS U705 ( .A(n2386), .Y(n2383) );
  CLKBUFX2TS U706 ( .A(n340), .Y(n2091) );
  CLKBUFX2TS U707 ( .A(n340), .Y(n2089) );
  CLKBUFX2TS U708 ( .A(n1325), .Y(n1283) );
  CLKBUFX2TS U709 ( .A(n1368), .Y(n1188) );
  CLKBUFX2TS U710 ( .A(n1368), .Y(n1187) );
  CLKBUFX2TS U711 ( .A(n1374), .Y(n1006) );
  CLKBUFX2TS U712 ( .A(n1374), .Y(n1002) );
  CLKBUFX2TS U713 ( .A(n1472), .Y(n995) );
  CLKBUFX2TS U714 ( .A(n1472), .Y(n993) );
  CLKBUFX2TS U715 ( .A(n1385), .Y(n517) );
  CLKBUFX2TS U716 ( .A(n527), .Y(n518) );
  CLKBUFX2TS U717 ( .A(n527), .Y(n519) );
  CLKBUFX2TS U718 ( .A(n526), .Y(n520) );
  CLKBUFX2TS U719 ( .A(n526), .Y(n521) );
  CLKBUFX2TS U720 ( .A(n525), .Y(n522) );
  CLKBUFX2TS U721 ( .A(n525), .Y(n523) );
  CLKBUFX2TS U722 ( .A(n525), .Y(n524) );
  CLKBUFX2TS U723 ( .A(n1325), .Y(n1324) );
  CLKBUFX2TS U724 ( .A(n477), .Y(n474) );
  CLKBUFX2TS U725 ( .A(n1552), .Y(n438) );
  CLKBUFX2TS U726 ( .A(n462), .Y(n461) );
  CLKBUFX2TS U727 ( .A(n1552), .Y(n437) );
  CLKBUFX2TS U728 ( .A(n2110), .Y(n2103) );
  CLKBUFX2TS U729 ( .A(n2110), .Y(n2104) );
  CLKBUFX2TS U730 ( .A(n2109), .Y(n2106) );
  CLKBUFX2TS U731 ( .A(n2109), .Y(n2107) );
  CLKBUFX2TS U732 ( .A(n2110), .Y(n2105) );
  CLKBUFX2TS U733 ( .A(n451), .Y(n448) );
  CLKBUFX2TS U734 ( .A(n463), .Y(n460) );
  CLKBUFX2TS U735 ( .A(n451), .Y(n447) );
  CLKBUFX2TS U736 ( .A(n463), .Y(n459) );
  CLKBUFX2TS U737 ( .A(n439), .Y(n436) );
  CLKBUFX2TS U738 ( .A(n339), .Y(n557) );
  CLKBUFX2TS U739 ( .A(n348), .Y(n344) );
  CLKBUFX2TS U740 ( .A(n348), .Y(n345) );
  CLKBUFX2TS U741 ( .A(n347), .Y(n346) );
  CLKBUFX2TS U742 ( .A(n2386), .Y(n2385) );
  CLKBUFX2TS U743 ( .A(n2108), .Y(n2093) );
  CLKBUFX2TS U744 ( .A(n2109), .Y(n2108) );
  CLKBUFX2TS U745 ( .A(n503), .Y(n488) );
  CLKBUFX2TS U746 ( .A(n504), .Y(n503) );
  CLKBUFX2TS U747 ( .A(n2386), .Y(n2384) );
  CLKBUFX2TS U748 ( .A(n504), .Y(n501) );
  CLKBUFX2TS U749 ( .A(n504), .Y(n500) );
  CLKBUFX2TS U750 ( .A(n504), .Y(n502) );
  NOR2X1TS U751 ( .A(n2363), .B(n641), .Y(n1323) );
  NOR2X1TS U752 ( .A(n2362), .B(n750), .Y(n1234) );
  NAND2X1TS U753 ( .A(n162), .B(n1282), .Y(n1247) );
  CLKBUFX2TS U754 ( .A(n1329), .Y(n585) );
  CLKBUFX2TS U755 ( .A(n1329), .Y(n586) );
  CLKBUFX2TS U756 ( .A(n1329), .Y(n587) );
  CLKBUFX2TS U757 ( .A(n1040), .Y(n1717) );
  CLKBUFX2TS U758 ( .A(n1040), .Y(n2007) );
  CLKBUFX2TS U759 ( .A(n1040), .Y(n2008) );
  CLKBUFX2TS U760 ( .A(n1249), .Y(n694) );
  CLKBUFX2TS U761 ( .A(n1249), .Y(n695) );
  CLKBUFX2TS U762 ( .A(n1249), .Y(n696) );
  CLKBUFX2TS U763 ( .A(n1250), .Y(n685) );
  CLKBUFX2TS U764 ( .A(n576), .Y(n575) );
  CLKBUFX2TS U765 ( .A(n577), .Y(n574) );
  CLKBUFX2TS U766 ( .A(n576), .Y(n573) );
  CLKBUFX2TS U767 ( .A(n576), .Y(n572) );
  CLKBUFX2TS U768 ( .A(n577), .Y(n571) );
  CLKBUFX2TS U769 ( .A(n577), .Y(n570) );
  CLKBUFX2TS U770 ( .A(n576), .Y(n569) );
  CLKBUFX2TS U771 ( .A(n577), .Y(n568) );
  CLKBUFX2TS U772 ( .A(n714), .Y(n713) );
  CLKBUFX2TS U773 ( .A(n714), .Y(n712) );
  CLKBUFX2TS U774 ( .A(n737), .Y(n711) );
  CLKBUFX2TS U775 ( .A(n595), .Y(n593) );
  CLKBUFX2TS U776 ( .A(n737), .Y(n710) );
  CLKBUFX2TS U777 ( .A(n595), .Y(n592) );
  CLKBUFX2TS U778 ( .A(n738), .Y(n709) );
  CLKBUFX2TS U779 ( .A(n598), .Y(n591) );
  CLKBUFX2TS U780 ( .A(n598), .Y(n590) );
  CLKBUFX2TS U781 ( .A(n714), .Y(n708) );
  CLKBUFX2TS U782 ( .A(n631), .Y(n589) );
  CLKBUFX2TS U783 ( .A(n737), .Y(n707) );
  CLKBUFX2TS U784 ( .A(n631), .Y(n588) );
  CLKBUFX2TS U785 ( .A(n676), .Y(n673) );
  CLKBUFX2TS U786 ( .A(n674), .Y(n672) );
  CLKBUFX2TS U787 ( .A(n674), .Y(n671) );
  CLKBUFX2TS U788 ( .A(n675), .Y(n670) );
  CLKBUFX2TS U789 ( .A(n675), .Y(n669) );
  CLKBUFX2TS U790 ( .A(n676), .Y(n668) );
  CLKBUFX2TS U791 ( .A(n676), .Y(n667) );
  CLKBUFX2TS U792 ( .A(n895), .Y(n894) );
  CLKBUFX2TS U793 ( .A(n895), .Y(n893) );
  CLKBUFX2TS U794 ( .A(n896), .Y(n892) );
  CLKBUFX2TS U795 ( .A(n896), .Y(n891) );
  CLKBUFX2TS U796 ( .A(n897), .Y(n890) );
  CLKBUFX2TS U797 ( .A(n895), .Y(n889) );
  CLKBUFX2TS U798 ( .A(n896), .Y(n888) );
  CLKBUFX2TS U799 ( .A(n664), .Y(n663) );
  CLKBUFX2TS U800 ( .A(n664), .Y(n662) );
  CLKBUFX2TS U801 ( .A(n665), .Y(n661) );
  CLKBUFX2TS U802 ( .A(n665), .Y(n660) );
  CLKBUFX2TS U803 ( .A(n665), .Y(n659) );
  CLKBUFX2TS U804 ( .A(n666), .Y(n658) );
  CLKBUFX2TS U805 ( .A(n666), .Y(n657) );
  CLKBUFX2TS U806 ( .A(n884), .Y(n883) );
  CLKBUFX2TS U807 ( .A(n884), .Y(n882) );
  CLKBUFX2TS U808 ( .A(n886), .Y(n881) );
  CLKBUFX2TS U809 ( .A(n886), .Y(n879) );
  CLKBUFX2TS U810 ( .A(n886), .Y(n878) );
  CLKBUFX2TS U811 ( .A(n887), .Y(n877) );
  CLKBUFX2TS U812 ( .A(n887), .Y(n876) );
  INVX2TS U813 ( .A(n1475), .Y(n810) );
  OR2X2TS U814 ( .A(n334), .B(n2365), .Y(n339) );
  AOI21X1TS U815 ( .A0(n806), .A1(n276), .B0(n2091), .Y(n1692) );
  OR2X2TS U816 ( .A(n272), .B(n334), .Y(n1590) );
  NOR2X1TS U817 ( .A(n1573), .B(n316), .Y(n1688) );
  INVX2TS U818 ( .A(n305), .Y(n813) );
  NAND2X1TS U819 ( .A(n1460), .B(n813), .Y(n1003) );
  CLKBUFX2TS U820 ( .A(n1005), .Y(n2047) );
  CLKBUFX2TS U821 ( .A(n1005), .Y(n2043) );
  CLKBUFX2TS U822 ( .A(n1005), .Y(n2045) );
  CLKBUFX2TS U823 ( .A(n1385), .Y(n527) );
  CLKBUFX2TS U824 ( .A(n1385), .Y(n526) );
  CLKBUFX2TS U825 ( .A(n426), .Y(n425) );
  CLKBUFX2TS U826 ( .A(n1332), .Y(n566) );
  CLKBUFX2TS U827 ( .A(n1478), .Y(n1325) );
  CLKBUFX2TS U828 ( .A(n1478), .Y(n1368) );
  CLKBUFX2TS U829 ( .A(n1478), .Y(n1374) );
  CLKBUFX2TS U830 ( .A(n1368), .Y(n1472) );
  CLKBUFX2TS U831 ( .A(n528), .Y(n525) );
  CLKBUFX2TS U832 ( .A(n427), .Y(n424) );
  CLKBUFX2TS U833 ( .A(n427), .Y(n423) );
  CLKBUFX2TS U834 ( .A(n567), .Y(n564) );
  CLKBUFX2TS U835 ( .A(n567), .Y(n565) );
  CLKBUFX2TS U836 ( .A(n1386), .Y(n515) );
  CLKBUFX2TS U837 ( .A(n1551), .Y(n450) );
  INVX2TS U838 ( .A(reset), .Y(n2386) );
  INVX2TS U839 ( .A(n1547), .Y(n477) );
  CLKBUFX2TS U840 ( .A(n746), .Y(n745) );
  CLKBUFX2TS U841 ( .A(n747), .Y(n744) );
  CLKBUFX2TS U842 ( .A(n747), .Y(n743) );
  CLKBUFX2TS U843 ( .A(n748), .Y(n742) );
  CLKBUFX2TS U844 ( .A(n638), .Y(n637) );
  CLKBUFX2TS U845 ( .A(n639), .Y(n636) );
  CLKBUFX2TS U846 ( .A(n639), .Y(n635) );
  CLKBUFX2TS U847 ( .A(n640), .Y(n634) );
  CLKBUFX2TS U848 ( .A(n640), .Y(n633) );
  CLKBUFX2TS U849 ( .A(n640), .Y(n632) );
  CLKBUFX2TS U850 ( .A(n1250), .Y(n686) );
  CLKBUFX2TS U851 ( .A(n1386), .Y(n516) );
  CLKBUFX2TS U852 ( .A(n1384), .Y(n540) );
  CLKBUFX2TS U853 ( .A(n863), .Y(n855) );
  CLKBUFX2TS U854 ( .A(n862), .Y(n856) );
  CLKBUFX2TS U855 ( .A(n862), .Y(n857) );
  CLKBUFX2TS U856 ( .A(n865), .Y(n858) );
  CLKBUFX2TS U857 ( .A(n861), .Y(n859) );
  CLKBUFX2TS U858 ( .A(n861), .Y(n860) );
  CLKBUFX2TS U859 ( .A(n838), .Y(n836) );
  CLKBUFX2TS U860 ( .A(n838), .Y(n834) );
  CLKBUFX2TS U861 ( .A(n840), .Y(n829) );
  CLKBUFX2TS U862 ( .A(n840), .Y(n826) );
  CLKBUFX2TS U863 ( .A(n841), .Y(n823) );
  CLKBUFX2TS U864 ( .A(n841), .Y(n817) );
  NOR2X1TS U865 ( .A(n374), .B(n2364), .Y(n1740) );
  NOR2X1TS U866 ( .A(n395), .B(n2364), .Y(n1728) );
  NAND2X1TS U867 ( .A(n289), .B(n2382), .Y(n1371) );
  CLKBUFX2TS U868 ( .A(n351), .Y(n349) );
  CLKBUFX2TS U869 ( .A(n352), .Y(n348) );
  CLKBUFX2TS U870 ( .A(n352), .Y(n347) );
  CLKBUFX2TS U871 ( .A(n807), .Y(n2110) );
  CLKBUFX2TS U872 ( .A(n807), .Y(n2109) );
  CLKBUFX2TS U873 ( .A(n1550), .Y(n462) );
  CLKBUFX2TS U874 ( .A(n358), .Y(n357) );
  CLKBUFX2TS U875 ( .A(n359), .Y(n356) );
  CLKBUFX2TS U876 ( .A(n359), .Y(n355) );
  CLKBUFX2TS U877 ( .A(n358), .Y(n354) );
  CLKBUFX2TS U878 ( .A(n379), .Y(n377) );
  CLKBUFX2TS U879 ( .A(n380), .Y(n376) );
  CLKBUFX2TS U880 ( .A(n381), .Y(n375) );
  CLKBUFX2TS U881 ( .A(n400), .Y(n398) );
  CLKBUFX2TS U882 ( .A(n401), .Y(n397) );
  CLKBUFX2TS U883 ( .A(n402), .Y(n396) );
  CLKBUFX2TS U884 ( .A(n350), .Y(n343) );
  CLKBUFX2TS U885 ( .A(n351), .Y(n350) );
  CLKBUFX2TS U886 ( .A(n863), .Y(n854) );
  CLKBUFX2TS U887 ( .A(n1551), .Y(n451) );
  CLKBUFX2TS U888 ( .A(n1550), .Y(n463) );
  CLKBUFX2TS U889 ( .A(n1552), .Y(n439) );
  INVX2TS U890 ( .A(n1575), .Y(n814) );
  CLKBUFX2TS U891 ( .A(n379), .Y(n378) );
  CLKBUFX2TS U892 ( .A(n400), .Y(n399) );
  NOR2X1TS U893 ( .A(n353), .B(n2363), .Y(n1752) );
  INVX2TS U894 ( .A(n1446), .Y(n504) );
  CLKBUFX2TS U895 ( .A(n2118), .Y(n2116) );
  CLKBUFX2TS U896 ( .A(n2118), .Y(n2115) );
  CLKBUFX2TS U897 ( .A(n2119), .Y(n2113) );
  CLKBUFX2TS U898 ( .A(n2119), .Y(n2114) );
  CLKBUFX2TS U899 ( .A(n2120), .Y(n2112) );
  CLKBUFX2TS U900 ( .A(n2120), .Y(n2111) );
  NOR2BX1TS U901 ( .AN(n1286), .B(n177), .Y(n1250) );
  CLKBUFX2TS U902 ( .A(n1246), .Y(n714) );
  CLKBUFX2TS U903 ( .A(n1246), .Y(n737) );
  CLKBUFX2TS U904 ( .A(n1246), .Y(n738) );
  CLKBUFX2TS U905 ( .A(n1111), .Y(n895) );
  CLKBUFX2TS U906 ( .A(n1111), .Y(n896) );
  CLKBUFX2TS U907 ( .A(n1111), .Y(n897) );
  CLKBUFX2TS U908 ( .A(n1328), .Y(n594) );
  CLKBUFX2TS U909 ( .A(n1328), .Y(n595) );
  CLKBUFX2TS U910 ( .A(n1328), .Y(n598) );
  CLKBUFX2TS U911 ( .A(n1328), .Y(n631) );
  CLKBUFX2TS U912 ( .A(n1287), .Y(n674) );
  CLKBUFX2TS U913 ( .A(n1287), .Y(n675) );
  CLKBUFX2TS U914 ( .A(n1287), .Y(n676) );
  CLKBUFX2TS U915 ( .A(n1112), .Y(n884) );
  CLKBUFX2TS U916 ( .A(n1112), .Y(n886) );
  CLKBUFX2TS U917 ( .A(n1112), .Y(n887) );
  CLKBUFX2TS U918 ( .A(n1288), .Y(n664) );
  CLKBUFX2TS U919 ( .A(n1288), .Y(n665) );
  CLKBUFX2TS U920 ( .A(n1288), .Y(n666) );
  CLKBUFX2TS U921 ( .A(n1331), .Y(n576) );
  CLKBUFX2TS U922 ( .A(n1331), .Y(n577) );
  CLKBUFX2TS U923 ( .A(n805), .Y(n804) );
  CLKBUFX2TS U924 ( .A(n805), .Y(n803) );
  CLKBUFX2TS U925 ( .A(n809), .Y(n755) );
  CLKBUFX2TS U926 ( .A(n809), .Y(n754) );
  CLKBUFX2TS U927 ( .A(n815), .Y(n753) );
  CLKBUFX2TS U928 ( .A(n815), .Y(n752) );
  CLKBUFX2TS U929 ( .A(n654), .Y(n653) );
  CLKBUFX2TS U930 ( .A(n655), .Y(n652) );
  CLKBUFX2TS U931 ( .A(n656), .Y(n651) );
  CLKBUFX2TS U932 ( .A(n655), .Y(n650) );
  CLKBUFX2TS U933 ( .A(n655), .Y(n644) );
  CLKBUFX2TS U934 ( .A(n656), .Y(n643) );
  CLKBUFX2TS U935 ( .A(n656), .Y(n642) );
  CLKBUFX2TS U936 ( .A(n875), .Y(n872) );
  CLKBUFX2TS U937 ( .A(n873), .Y(n871) );
  CLKBUFX2TS U938 ( .A(n873), .Y(n870) );
  CLKBUFX2TS U939 ( .A(n874), .Y(n869) );
  CLKBUFX2TS U940 ( .A(n874), .Y(n868) );
  CLKBUFX2TS U941 ( .A(n875), .Y(n867) );
  CLKBUFX2TS U942 ( .A(n875), .Y(n866) );
  INVX2TS U943 ( .A(n1285), .Y(n822) );
  NOR2X1TS U944 ( .A(n339), .B(n825), .Y(n1460) );
  NOR2X1TS U945 ( .A(n1590), .B(n113), .Y(n1595) );
  AND2X2TS U946 ( .A(n1709), .B(n832), .Y(n1697) );
  NOR3X1TS U947 ( .A(n1663), .B(n835), .C(n557), .Y(n1675) );
  NAND2X1TS U948 ( .A(n113), .B(n124), .Y(n1661) );
  NAND2X1TS U949 ( .A(n1711), .B(n541), .Y(n1547) );
  NAND2X1TS U950 ( .A(n816), .B(n292), .Y(n1573) );
  INVX2TS U951 ( .A(n1451), .Y(n835) );
  NOR2X1TS U952 ( .A(n113), .B(n555), .Y(n1551) );
  NOR2X1TS U953 ( .A(n1451), .B(n554), .Y(n1384) );
  NAND2BX1TS U954 ( .AN(n124), .B(n1710), .Y(n1694) );
  AND2X2TS U955 ( .A(n1675), .B(n831), .Y(n1386) );
  INVX2TS U956 ( .A(n1576), .Y(n816) );
  CLKBUFX2TS U957 ( .A(n1191), .Y(n838) );
  CLKBUFX2TS U958 ( .A(n1191), .Y(n839) );
  CLKBUFX2TS U959 ( .A(n1191), .Y(n840) );
  CLKBUFX2TS U960 ( .A(n1191), .Y(n841) );
  CLKBUFX2TS U961 ( .A(n750), .Y(n748) );
  CLKBUFX2TS U962 ( .A(n750), .Y(n749) );
  CLKBUFX2TS U963 ( .A(n1291), .Y(n640) );
  CLKBUFX2TS U964 ( .A(n865), .Y(n862) );
  CLKBUFX2TS U965 ( .A(n863), .Y(n861) );
  CLKBUFX2TS U966 ( .A(n865), .Y(n863) );
  CLKBUFX2TS U967 ( .A(n751), .Y(n746) );
  CLKBUFX2TS U968 ( .A(n751), .Y(n747) );
  CLKBUFX2TS U969 ( .A(n641), .Y(n638) );
  CLKBUFX2TS U970 ( .A(n641), .Y(n639) );
  CLKBUFX2TS U971 ( .A(n1553), .Y(n426) );
  CLKBUFX2TS U972 ( .A(n1041), .Y(n1478) );
  CLKBUFX2TS U973 ( .A(n864), .Y(n853) );
  CLKBUFX2TS U974 ( .A(n865), .Y(n864) );
  AND2X2TS U975 ( .A(n1710), .B(n124), .Y(n1709) );
  AND2X2TS U976 ( .A(n1688), .B(n831), .Y(n1682) );
  CLKBUFX2TS U977 ( .A(n1553), .Y(n427) );
  CLKBUFX2TS U978 ( .A(n1332), .Y(n567) );
  CLKBUFX2TS U979 ( .A(n1385), .Y(n528) );
  NAND2X1TS U980 ( .A(n1527), .B(n2386), .Y(n1529) );
  NAND2X1TS U981 ( .A(n2376), .B(n172), .Y(n1376) );
  NOR2X1TS U982 ( .A(n1576), .B(n293), .Y(n1575) );
  NOR2X1TS U983 ( .A(n125), .B(n555), .Y(n1550) );
  NOR2X1TS U984 ( .A(n832), .B(n555), .Y(n1552) );
  INVX2TS U985 ( .A(n1663), .Y(n807) );
  CLKBUFX2TS U986 ( .A(n383), .Y(n381) );
  CLKBUFX2TS U987 ( .A(n1736), .Y(n402) );
  CLKBUFX2TS U988 ( .A(n362), .Y(n359) );
  CLKBUFX2TS U989 ( .A(n383), .Y(n380) );
  CLKBUFX2TS U990 ( .A(n404), .Y(n401) );
  CLKBUFX2TS U991 ( .A(n362), .Y(n358) );
  CLKBUFX2TS U992 ( .A(n383), .Y(n379) );
  CLKBUFX2TS U993 ( .A(n404), .Y(n400) );
  CLKBUFX2TS U994 ( .A(n360), .Y(n353) );
  CLKBUFX2TS U995 ( .A(n361), .Y(n360) );
  CLKBUFX2TS U996 ( .A(n382), .Y(n374) );
  CLKBUFX2TS U997 ( .A(n1748), .Y(n382) );
  CLKBUFX2TS U998 ( .A(n403), .Y(n395) );
  CLKBUFX2TS U999 ( .A(n1736), .Y(n403) );
  CLKBUFX2TS U1000 ( .A(n1762), .Y(n351) );
  CLKBUFX2TS U1001 ( .A(n1762), .Y(n352) );
  NOR2X1TS U1002 ( .A(n392), .B(n2364), .Y(n1741) );
  NOR2X1TS U1003 ( .A(n414), .B(n2365), .Y(n1729) );
  NOR2X1TS U1004 ( .A(n371), .B(n2364), .Y(n1753) );
  CLKBUFX2TS U1005 ( .A(n2121), .Y(n2119) );
  CLKBUFX2TS U1006 ( .A(n2121), .Y(n2120) );
  CLKBUFX2TS U1007 ( .A(n2121), .Y(n2117) );
  CLKBUFX2TS U1008 ( .A(n2121), .Y(n2118) );
  NAND2X1TS U1009 ( .A(n1724), .B(n2117), .Y(n1714) );
  CLKBUFX2TS U1010 ( .A(n367), .Y(n365) );
  CLKBUFX2TS U1011 ( .A(n368), .Y(n364) );
  CLKBUFX2TS U1012 ( .A(n368), .Y(n363) );
  CLKBUFX2TS U1013 ( .A(n388), .Y(n386) );
  CLKBUFX2TS U1014 ( .A(n389), .Y(n385) );
  CLKBUFX2TS U1015 ( .A(n389), .Y(n384) );
  CLKBUFX2TS U1016 ( .A(n411), .Y(n409) );
  CLKBUFX2TS U1017 ( .A(n412), .Y(n408) );
  CLKBUFX2TS U1018 ( .A(n412), .Y(n407) );
  CLKBUFX2TS U1019 ( .A(n413), .Y(n406) );
  CLKBUFX2TS U1020 ( .A(n413), .Y(n405) );
  CLKBUFX2TS U1021 ( .A(n388), .Y(n387) );
  CLKBUFX2TS U1022 ( .A(n411), .Y(n410) );
  CLKBUFX2TS U1023 ( .A(n367), .Y(n366) );
  NOR2X1TS U1024 ( .A(n177), .B(n2366), .Y(n1380) );
  NAND3X1TS U1025 ( .A(n797), .B(n1366), .C(n1364), .Y(n1328) );
  NAND3X1TS U1026 ( .A(n1326), .B(n798), .C(n1323), .Y(n1287) );
  NAND3X1TS U1027 ( .A(n820), .B(n1189), .C(n1186), .Y(n1111) );
  NAND2X1TS U1028 ( .A(n165), .B(n1323), .Y(n1288) );
  NAND2X1TS U1029 ( .A(n169), .B(n1186), .Y(n1112) );
  AOI221X1TS U1030 ( .A0(n171), .A1(n1513), .B0(n1475), .B1(n822), .C0(n2371), 
        .Y(n1286) );
  AOI221X1TS U1031 ( .A0(n170), .A1(n1474), .B0(n1475), .B1(n117), .C0(n2371), 
        .Y(n1473) );
  CLKBUFX2TS U1032 ( .A(n1193), .Y(n805) );
  CLKBUFX2TS U1033 ( .A(n1193), .Y(n808) );
  CLKBUFX2TS U1034 ( .A(n1193), .Y(n809) );
  CLKBUFX2TS U1035 ( .A(n1193), .Y(n815) );
  CLKBUFX2TS U1036 ( .A(n1290), .Y(n654) );
  CLKBUFX2TS U1037 ( .A(n1290), .Y(n655) );
  CLKBUFX2TS U1038 ( .A(n1290), .Y(n656) );
  CLKBUFX2TS U1039 ( .A(n1114), .Y(n873) );
  CLKBUFX2TS U1040 ( .A(n1114), .Y(n874) );
  CLKBUFX2TS U1041 ( .A(n1114), .Y(n875) );
  CLKBUFX2TS U1042 ( .A(n1194), .Y(n750) );
  NAND2X1TS U1043 ( .A(n293), .B(n831), .Y(n1689) );
  NOR3X1TS U1044 ( .A(n833), .B(n1662), .C(n1661), .Y(n1711) );
  AND2X2TS U1045 ( .A(n1709), .B(n281), .Y(n1698) );
  NAND2X1TS U1046 ( .A(n120), .B(n1234), .Y(n1191) );
  NAND2X1TS U1047 ( .A(n334), .B(n885), .Y(n1439) );
  NOR2X1TS U1048 ( .A(n837), .B(n9), .Y(n1539) );
  INVX2TS U1049 ( .A(n1676), .Y(n837) );
  INVX2TS U1050 ( .A(n257), .Y(n831) );
  INVX2TS U1051 ( .A(n1569), .Y(n825) );
  AND2X2TS U1052 ( .A(n1675), .B(n258), .Y(n1385) );
  CLKBUFX2TS U1053 ( .A(n1115), .Y(n865) );
  NOR2X1TS U1054 ( .A(n983), .B(n984), .Y(n3644) );
  NOR2X1TS U1055 ( .A(n986), .B(n984), .Y(n3642) );
  AND2X2TS U1056 ( .A(n1688), .B(n258), .Y(n1681) );
  CLKBUFX2TS U1057 ( .A(n1291), .Y(n641) );
  CLKBUFX2TS U1058 ( .A(n1194), .Y(n751) );
  CLKBUFX2TS U1059 ( .A(n850), .Y(n849) );
  CLKBUFX2TS U1060 ( .A(n850), .Y(n848) );
  CLKBUFX2TS U1061 ( .A(n851), .Y(n847) );
  CLKBUFX2TS U1062 ( .A(n851), .Y(n846) );
  CLKBUFX2TS U1063 ( .A(n852), .Y(n845) );
  CLKBUFX2TS U1064 ( .A(n852), .Y(n843) );
  CLKBUFX2TS U1065 ( .A(n852), .Y(n842) );
  XNOR2X1TS U1066 ( .A(n1448), .B(n885), .Y(n997) );
  NAND3BX1TS U1067 ( .AN(n115), .B(n992), .C(n1001), .Y(n1429) );
  NAND2X1TS U1068 ( .A(n1449), .B(n1450), .Y(n992) );
  NAND2X1TS U1069 ( .A(n1725), .B(n739), .Y(n1762) );
  INVX2TS U1070 ( .A(n1662), .Y(n832) );
  CLKBUFX2TS U1071 ( .A(n372), .Y(n371) );
  CLKBUFX2TS U1072 ( .A(n393), .Y(n392) );
  CLKBUFX2TS U1073 ( .A(n1760), .Y(n361) );
  CLKBUFX2TS U1074 ( .A(n1760), .Y(n362) );
  CLKBUFX2TS U1075 ( .A(n1748), .Y(n383) );
  CLKBUFX2TS U1076 ( .A(n1736), .Y(n404) );
  XNOR2X1TS U1077 ( .A(n997), .B(n998), .Y(n983) );
  NOR2X1TS U1078 ( .A(n138), .B(n2365), .Y(n1724) );
  NOR3X1TS U1079 ( .A(n1435), .B(n2362), .C(n825), .Y(n1434) );
  NOR2X1TS U1080 ( .A(n885), .B(n293), .Y(n1422) );
  CLKBUFX2TS U1081 ( .A(n372), .Y(n369) );
  CLKBUFX2TS U1082 ( .A(n372), .Y(n370) );
  CLKBUFX2TS U1083 ( .A(n393), .Y(n390) );
  CLKBUFX2TS U1084 ( .A(n393), .Y(n391) );
  CLKBUFX2TS U1085 ( .A(n414), .Y(n413) );
  CLKBUFX2TS U1086 ( .A(n394), .Y(n388) );
  CLKBUFX2TS U1087 ( .A(n415), .Y(n411) );
  CLKBUFX2TS U1088 ( .A(n373), .Y(n367) );
  CLKBUFX2TS U1089 ( .A(n373), .Y(n368) );
  CLKBUFX2TS U1090 ( .A(n394), .Y(n389) );
  CLKBUFX2TS U1091 ( .A(n415), .Y(n412) );
  CLKBUFX2TS U1092 ( .A(n739), .Y(n2121) );
  INVX2TS U1093 ( .A(n2243), .Y(n2242) );
  INVX2TS U1094 ( .A(n2246), .Y(n2245) );
  INVX2TS U1095 ( .A(n2249), .Y(n2248) );
  INVX2TS U1096 ( .A(n2252), .Y(n2251) );
  INVX2TS U1097 ( .A(n2256), .Y(n2254) );
  INVX2TS U1098 ( .A(n2258), .Y(n2257) );
  INVX2TS U1099 ( .A(n2261), .Y(n2260) );
  INVX2TS U1100 ( .A(n2265), .Y(n2263) );
  INVX2TS U1101 ( .A(n2267), .Y(n2266) );
  INVX2TS U1102 ( .A(n2270), .Y(n2269) );
  INVX2TS U1103 ( .A(n2273), .Y(n2272) );
  INVX2TS U1104 ( .A(n2276), .Y(n2275) );
  INVX2TS U1105 ( .A(n2279), .Y(n2278) );
  INVX2TS U1106 ( .A(n2282), .Y(n2281) );
  INVX2TS U1107 ( .A(n2286), .Y(n2284) );
  INVX2TS U1108 ( .A(n2289), .Y(n2287) );
  INVX2TS U1109 ( .A(n2291), .Y(n2290) );
  INVX2TS U1110 ( .A(n2294), .Y(n2293) );
  INVX2TS U1111 ( .A(n2297), .Y(n2296) );
  INVX2TS U1112 ( .A(n2301), .Y(n2299) );
  INVX2TS U1113 ( .A(n2303), .Y(n2302) );
  INVX2TS U1114 ( .A(n2307), .Y(n2305) );
  INVX2TS U1115 ( .A(n2310), .Y(n2308) );
  INVX2TS U1116 ( .A(n2312), .Y(n2311) );
  INVX2TS U1117 ( .A(n2315), .Y(n2314) );
  INVX2TS U1118 ( .A(n2318), .Y(n2317) );
  INVX2TS U1119 ( .A(n2321), .Y(n2320) );
  INVX2TS U1120 ( .A(n2325), .Y(n2323) );
  INVX2TS U1121 ( .A(n2327), .Y(n2326) );
  INVX2TS U1122 ( .A(n2331), .Y(n2329) );
  INVX2TS U1123 ( .A(n2333), .Y(n2332) );
  INVX2TS U1124 ( .A(n2336), .Y(n2335) );
  INVX2TS U1125 ( .A(n2124), .Y(n2122) );
  INVX2TS U1126 ( .A(n2126), .Y(n2125) );
  INVX2TS U1127 ( .A(n2130), .Y(n2128) );
  INVX2TS U1128 ( .A(n2132), .Y(n2131) );
  INVX2TS U1129 ( .A(n2135), .Y(n2134) );
  INVX2TS U1130 ( .A(n2139), .Y(n2137) );
  INVX2TS U1131 ( .A(n2141), .Y(n2140) );
  INVX2TS U1132 ( .A(n2144), .Y(n2143) );
  INVX2TS U1133 ( .A(n2148), .Y(n2146) );
  INVX2TS U1134 ( .A(n2150), .Y(n2149) );
  INVX2TS U1135 ( .A(n2153), .Y(n2152) );
  INVX2TS U1136 ( .A(n2156), .Y(n2155) );
  INVX2TS U1137 ( .A(n2159), .Y(n2158) );
  INVX2TS U1138 ( .A(n2163), .Y(n2161) );
  INVX2TS U1139 ( .A(n2165), .Y(n2164) );
  INVX2TS U1140 ( .A(n2168), .Y(n2167) );
  INVX2TS U1141 ( .A(n2172), .Y(n2170) );
  INVX2TS U1142 ( .A(n2174), .Y(n2173) );
  INVX2TS U1143 ( .A(n2178), .Y(n2176) );
  INVX2TS U1144 ( .A(n2180), .Y(n2179) );
  INVX2TS U1145 ( .A(n2183), .Y(n2182) );
  INVX2TS U1146 ( .A(n2186), .Y(n2185) );
  INVX2TS U1147 ( .A(n2189), .Y(n2188) );
  INVX2TS U1148 ( .A(n2192), .Y(n2191) );
  INVX2TS U1149 ( .A(n2196), .Y(n2194) );
  INVX2TS U1150 ( .A(n2198), .Y(n2197) );
  INVX2TS U1151 ( .A(n2201), .Y(n2200) );
  INVX2TS U1152 ( .A(n2204), .Y(n2203) );
  INVX2TS U1153 ( .A(n2207), .Y(n2206) );
  INVX2TS U1154 ( .A(n2211), .Y(n2209) );
  INVX2TS U1155 ( .A(n2213), .Y(n2212) );
  INVX2TS U1156 ( .A(n2216), .Y(n2215) );
  CLKBUFX2TS U1157 ( .A(n2224), .Y(n2225) );
  CLKBUFX2TS U1158 ( .A(n2226), .Y(n2227) );
  CLKBUFX2TS U1159 ( .A(n2228), .Y(n2229) );
  CLKBUFX2TS U1160 ( .A(n2230), .Y(n2231) );
  CLKBUFX2TS U1161 ( .A(n2236), .Y(n2237) );
  CLKBUFX2TS U1162 ( .A(n2239), .Y(n2240) );
  CLKBUFX2TS U1163 ( .A(n2344), .Y(n2345) );
  CLKBUFX2TS U1164 ( .A(n2346), .Y(n2347) );
  CLKBUFX2TS U1165 ( .A(n2350), .Y(n2351) );
  CLKBUFX2TS U1166 ( .A(n2354), .Y(n2355) );
  CLKBUFX2TS U1167 ( .A(n2356), .Y(n2357) );
  CLKBUFX2TS U1168 ( .A(n2359), .Y(n2360) );
  CLKBUFX2TS U1169 ( .A(n2232), .Y(n2233) );
  CLKBUFX2TS U1170 ( .A(n2234), .Y(n2235) );
  CLKBUFX2TS U1171 ( .A(n2236), .Y(n2238) );
  CLKBUFX2TS U1172 ( .A(n2239), .Y(n2241) );
  CLKBUFX2TS U1173 ( .A(n2348), .Y(n2349) );
  CLKBUFX2TS U1174 ( .A(n2352), .Y(n2353) );
  CLKBUFX2TS U1175 ( .A(n2356), .Y(n2358) );
  CLKBUFX2TS U1176 ( .A(n2359), .Y(n2361) );
  NOR2X1TS U1177 ( .A(n332), .B(n2365), .Y(n1382) );
  INVX2TS U1178 ( .A(requesterAddressIn_WEST[0]), .Y(n2218) );
  INVX2TS U1179 ( .A(requesterAddressIn_WEST[1]), .Y(n2219) );
  INVX2TS U1180 ( .A(requesterAddressIn_WEST[2]), .Y(n2220) );
  INVX2TS U1181 ( .A(requesterAddressIn_WEST[3]), .Y(n2221) );
  INVX2TS U1182 ( .A(requesterAddressIn_WEST[4]), .Y(n2222) );
  INVX2TS U1183 ( .A(requesterAddressIn_WEST[5]), .Y(n2223) );
  NOR2X1TS U1184 ( .A(n308), .B(n9), .Y(n1039) );
  INVX2TS U1185 ( .A(n1284), .Y(n801) );
  INVX2TS U1186 ( .A(n330), .Y(n797) );
  XNOR2X1TS U1187 ( .A(n189), .B(n144), .Y(n1543) );
  XNOR2X1TS U1188 ( .A(n833), .B(n175), .Y(n998) );
  OAI22X1TS U1189 ( .A0(n366), .A1(n950), .B0(n360), .B1(n982), .Y(N10083) );
  OAI22X1TS U1190 ( .A0(n366), .A1(n949), .B0(n357), .B1(n981), .Y(N10084) );
  OAI22X1TS U1191 ( .A0(n366), .A1(n948), .B0(n357), .B1(n980), .Y(N10085) );
  OAI22X1TS U1192 ( .A0(n365), .A1(n947), .B0(n357), .B1(n979), .Y(N10086) );
  OAI22X1TS U1193 ( .A0(n365), .A1(n946), .B0(n357), .B1(n978), .Y(N10087) );
  OAI22X1TS U1194 ( .A0(n365), .A1(n945), .B0(n356), .B1(n977), .Y(N10088) );
  OAI22X1TS U1195 ( .A0(n365), .A1(n944), .B0(n356), .B1(n976), .Y(N10089) );
  OAI22X1TS U1196 ( .A0(n364), .A1(n943), .B0(n356), .B1(n975), .Y(N10090) );
  OAI22X1TS U1197 ( .A0(n364), .A1(n942), .B0(n356), .B1(n974), .Y(N10091) );
  OAI22X1TS U1198 ( .A0(n364), .A1(n941), .B0(n355), .B1(n973), .Y(N10092) );
  OAI22X1TS U1199 ( .A0(n364), .A1(n940), .B0(n355), .B1(n972), .Y(N10093) );
  OAI22X1TS U1200 ( .A0(n363), .A1(n939), .B0(n355), .B1(n971), .Y(N10094) );
  OAI22X1TS U1201 ( .A0(n363), .A1(n938), .B0(n355), .B1(n970), .Y(N10095) );
  OAI22X1TS U1202 ( .A0(n363), .A1(n937), .B0(n361), .B1(n969), .Y(N10096) );
  OAI22X1TS U1203 ( .A0(n363), .A1(n936), .B0(n1760), .B1(n968), .Y(N10097) );
  OAI22X1TS U1204 ( .A0(n369), .A1(n935), .B0(n359), .B1(n967), .Y(N10098) );
  OAI22X1TS U1205 ( .A0(n373), .A1(n934), .B0(n359), .B1(n966), .Y(N10099) );
  OAI22X1TS U1206 ( .A0(n373), .A1(n933), .B0(n360), .B1(n965), .Y(N10100) );
  OAI22X1TS U1207 ( .A0(n369), .A1(n932), .B0(n362), .B1(n964), .Y(N10101) );
  OAI22X1TS U1208 ( .A0(n367), .A1(n931), .B0(n1760), .B1(n963), .Y(N10102) );
  OAI22X1TS U1209 ( .A0(n372), .A1(n930), .B0(n358), .B1(n962), .Y(N10103) );
  OAI22X1TS U1210 ( .A0(n1759), .A1(n929), .B0(n360), .B1(n961), .Y(N10104) );
  OAI22X1TS U1211 ( .A0(n370), .A1(n928), .B0(n362), .B1(n960), .Y(N10105) );
  OAI22X1TS U1212 ( .A0(n370), .A1(n927), .B0(n361), .B1(n959), .Y(N10106) );
  OAI22X1TS U1213 ( .A0(n370), .A1(n926), .B0(n361), .B1(n958), .Y(N10107) );
  OAI22X1TS U1214 ( .A0(n367), .A1(n925), .B0(n354), .B1(n957), .Y(N10108) );
  OAI22X1TS U1215 ( .A0(n368), .A1(n924), .B0(n354), .B1(n956), .Y(N10109) );
  OAI22X1TS U1216 ( .A0(n370), .A1(n923), .B0(n354), .B1(n955), .Y(N10110) );
  OAI22X1TS U1217 ( .A0(n369), .A1(n922), .B0(n354), .B1(n954), .Y(N10111) );
  OAI22X1TS U1218 ( .A0(n368), .A1(n921), .B0(n353), .B1(n953), .Y(N10112) );
  OAI22X1TS U1219 ( .A0(n371), .A1(n920), .B0(n353), .B1(n952), .Y(N10113) );
  OAI22X1TS U1220 ( .A0(n369), .A1(n919), .B0(n353), .B1(n951), .Y(N10114) );
  OAI22X1TS U1221 ( .A0(n387), .A1(n950), .B0(n378), .B1(n982), .Y(N10117) );
  OAI22X1TS U1222 ( .A0(n387), .A1(n949), .B0(n377), .B1(n981), .Y(N10118) );
  OAI22X1TS U1223 ( .A0(n387), .A1(n948), .B0(n377), .B1(n980), .Y(N10119) );
  OAI22X1TS U1224 ( .A0(n386), .A1(n947), .B0(n377), .B1(n979), .Y(N10120) );
  OAI22X1TS U1225 ( .A0(n386), .A1(n946), .B0(n377), .B1(n978), .Y(N10121) );
  OAI22X1TS U1226 ( .A0(n386), .A1(n945), .B0(n380), .B1(n977), .Y(N10122) );
  OAI22X1TS U1227 ( .A0(n386), .A1(n944), .B0(n378), .B1(n976), .Y(N10123) );
  OAI22X1TS U1228 ( .A0(n385), .A1(n943), .B0(n379), .B1(n975), .Y(N10124) );
  OAI22X1TS U1229 ( .A0(n385), .A1(n942), .B0(n382), .B1(n974), .Y(N10125) );
  OAI22X1TS U1230 ( .A0(n385), .A1(n941), .B0(n376), .B1(n973), .Y(N10126) );
  OAI22X1TS U1231 ( .A0(n385), .A1(n940), .B0(n376), .B1(n972), .Y(N10127) );
  OAI22X1TS U1232 ( .A0(n384), .A1(n939), .B0(n376), .B1(n971), .Y(N10128) );
  OAI22X1TS U1233 ( .A0(n384), .A1(n938), .B0(n376), .B1(n970), .Y(N10129) );
  OAI22X1TS U1234 ( .A0(n384), .A1(n937), .B0(n375), .B1(n969), .Y(N10130) );
  OAI22X1TS U1235 ( .A0(n384), .A1(n936), .B0(n375), .B1(n968), .Y(N10131) );
  OAI22X1TS U1236 ( .A0(n390), .A1(n935), .B0(n375), .B1(n967), .Y(N10132) );
  OAI22X1TS U1237 ( .A0(n394), .A1(n934), .B0(n375), .B1(n966), .Y(N10133) );
  OAI22X1TS U1238 ( .A0(n394), .A1(n933), .B0(n380), .B1(n965), .Y(N10134) );
  OAI22X1TS U1239 ( .A0(n390), .A1(n932), .B0(n382), .B1(n964), .Y(N10135) );
  OAI22X1TS U1240 ( .A0(n388), .A1(n931), .B0(n1748), .B1(n963), .Y(N10136) );
  OAI22X1TS U1241 ( .A0(n393), .A1(n930), .B0(n1748), .B1(n962), .Y(N10137) );
  OAI22X1TS U1242 ( .A0(n1747), .A1(n929), .B0(n381), .B1(n961), .Y(N10138) );
  OAI22X1TS U1243 ( .A0(n391), .A1(n928), .B0(n380), .B1(n960), .Y(N10139) );
  OAI22X1TS U1244 ( .A0(n391), .A1(n927), .B0(n382), .B1(n959), .Y(N10140) );
  OAI22X1TS U1245 ( .A0(n391), .A1(n926), .B0(n381), .B1(n958), .Y(N10141) );
  OAI22X1TS U1246 ( .A0(n388), .A1(n925), .B0(n381), .B1(n957), .Y(N10142) );
  OAI22X1TS U1247 ( .A0(n389), .A1(n924), .B0(n378), .B1(n956), .Y(N10143) );
  OAI22X1TS U1248 ( .A0(n391), .A1(n923), .B0(n383), .B1(n955), .Y(N10144) );
  OAI22X1TS U1249 ( .A0(n390), .A1(n922), .B0(n379), .B1(n954), .Y(N10145) );
  OAI22X1TS U1250 ( .A0(n389), .A1(n921), .B0(n374), .B1(n953), .Y(N10146) );
  OAI22X1TS U1251 ( .A0(n392), .A1(n920), .B0(n374), .B1(n952), .Y(N10147) );
  OAI22X1TS U1252 ( .A0(n390), .A1(n919), .B0(n374), .B1(n951), .Y(N10148) );
  OAI22X1TS U1253 ( .A0(n410), .A1(n950), .B0(n399), .B1(n982), .Y(N10151) );
  OAI22X1TS U1254 ( .A0(n410), .A1(n949), .B0(n398), .B1(n981), .Y(N10152) );
  OAI22X1TS U1255 ( .A0(n410), .A1(n948), .B0(n398), .B1(n980), .Y(N10153) );
  OAI22X1TS U1256 ( .A0(n409), .A1(n947), .B0(n398), .B1(n979), .Y(N10154) );
  OAI22X1TS U1257 ( .A0(n409), .A1(n946), .B0(n398), .B1(n978), .Y(N10155) );
  OAI22X1TS U1258 ( .A0(n409), .A1(n945), .B0(n397), .B1(n977), .Y(N10156) );
  OAI22X1TS U1259 ( .A0(n409), .A1(n944), .B0(n397), .B1(n976), .Y(N10157) );
  OAI22X1TS U1260 ( .A0(n408), .A1(n943), .B0(n397), .B1(n975), .Y(N10158) );
  OAI22X1TS U1261 ( .A0(n408), .A1(n942), .B0(n397), .B1(n974), .Y(N10159) );
  OAI22X1TS U1262 ( .A0(n408), .A1(n941), .B0(n401), .B1(n973), .Y(N10160) );
  OAI22X1TS U1263 ( .A0(n408), .A1(n940), .B0(n400), .B1(n972), .Y(N10161) );
  OAI22X1TS U1264 ( .A0(n407), .A1(n939), .B0(n403), .B1(n971), .Y(N10162) );
  OAI22X1TS U1265 ( .A0(n407), .A1(n938), .B0(n1736), .B1(n970), .Y(N10163) );
  OAI22X1TS U1266 ( .A0(n407), .A1(n937), .B0(n401), .B1(n969), .Y(N10164) );
  OAI22X1TS U1267 ( .A0(n407), .A1(n936), .B0(n402), .B1(n968), .Y(N10165) );
  OAI22X1TS U1268 ( .A0(n412), .A1(n935), .B0(n399), .B1(n967), .Y(N10166) );
  OAI22X1TS U1269 ( .A0(n411), .A1(n934), .B0(n404), .B1(n966), .Y(N10167) );
  OAI22X1TS U1270 ( .A0(n412), .A1(n933), .B0(n396), .B1(n965), .Y(N10168) );
  OAI22X1TS U1271 ( .A0(n414), .A1(n932), .B0(n396), .B1(n964), .Y(N10169) );
  OAI22X1TS U1272 ( .A0(n415), .A1(n931), .B0(n396), .B1(n963), .Y(N10170) );
  OAI22X1TS U1273 ( .A0(n411), .A1(n930), .B0(n396), .B1(n962), .Y(N10171) );
  OAI22X1TS U1274 ( .A0(n413), .A1(n929), .B0(n402), .B1(n961), .Y(N10172) );
  OAI22X1TS U1275 ( .A0(n406), .A1(n928), .B0(n403), .B1(n960), .Y(N10173) );
  OAI22X1TS U1276 ( .A0(n406), .A1(n927), .B0(n403), .B1(n959), .Y(N10174) );
  OAI22X1TS U1277 ( .A0(n406), .A1(n926), .B0(n400), .B1(n958), .Y(N10175) );
  OAI22X1TS U1278 ( .A0(n413), .A1(n925), .B0(n402), .B1(n957), .Y(N10176) );
  OAI22X1TS U1279 ( .A0(n405), .A1(n924), .B0(n401), .B1(n956), .Y(N10177) );
  OAI22X1TS U1280 ( .A0(n405), .A1(n923), .B0(n399), .B1(n955), .Y(N10178) );
  OAI22X1TS U1281 ( .A0(n406), .A1(n922), .B0(n404), .B1(n954), .Y(N10179) );
  OAI22X1TS U1282 ( .A0(n405), .A1(n921), .B0(n395), .B1(n953), .Y(N10180) );
  OAI22X1TS U1283 ( .A0(n415), .A1(n920), .B0(n395), .B1(n952), .Y(N10181) );
  OAI22X1TS U1284 ( .A0(n405), .A1(n919), .B0(n395), .B1(n951), .Y(N10182) );
  OAI22X1TS U1285 ( .A0(n2120), .A1(n950), .B0(n343), .B1(n982), .Y(N10185) );
  OAI22X1TS U1286 ( .A0(n2117), .A1(n949), .B0(n343), .B1(n981), .Y(N10186) );
  OAI22X1TS U1287 ( .A0(n2119), .A1(n948), .B0(n343), .B1(n980), .Y(N10187) );
  OAI22X1TS U1288 ( .A0(n2117), .A1(n947), .B0(n349), .B1(n979), .Y(N10188) );
  OAI22X1TS U1289 ( .A0(n2117), .A1(n946), .B0(n352), .B1(n978), .Y(N10189) );
  OAI22X1TS U1290 ( .A0(n2120), .A1(n945), .B0(n351), .B1(n977), .Y(N10190) );
  OAI22X1TS U1291 ( .A0(n2118), .A1(n944), .B0(n1762), .B1(n976), .Y(N10191)
         );
  OAI22X1TS U1292 ( .A0(n2116), .A1(n943), .B0(n349), .B1(n975), .Y(N10192) );
  OAI22X1TS U1293 ( .A0(n2116), .A1(n942), .B0(n349), .B1(n974), .Y(N10193) );
  OAI22X1TS U1294 ( .A0(n2116), .A1(n941), .B0(n348), .B1(n973), .Y(N10194) );
  OAI22X1TS U1295 ( .A0(n2116), .A1(n940), .B0(n347), .B1(n972), .Y(N10195) );
  OAI22X1TS U1296 ( .A0(n2115), .A1(n939), .B0(n351), .B1(n971), .Y(N10196) );
  OAI22X1TS U1297 ( .A0(n2115), .A1(n938), .B0(n1762), .B1(n970), .Y(N10197)
         );
  OAI22X1TS U1298 ( .A0(n2115), .A1(n937), .B0(n350), .B1(n969), .Y(N10198) );
  OAI22X1TS U1299 ( .A0(n2115), .A1(n936), .B0(n349), .B1(n968), .Y(N10199) );
  OAI22X1TS U1300 ( .A0(n2114), .A1(n935), .B0(n348), .B1(n967), .Y(N10200) );
  OAI22X1TS U1301 ( .A0(n2114), .A1(n934), .B0(n350), .B1(n966), .Y(N10201) );
  OAI22X1TS U1302 ( .A0(n2114), .A1(n933), .B0(n347), .B1(n965), .Y(N10202) );
  OAI22X1TS U1303 ( .A0(n2113), .A1(n932), .B0(n352), .B1(n964), .Y(N10203) );
  OAI22X1TS U1304 ( .A0(n2113), .A1(n931), .B0(n344), .B1(n963), .Y(N10204) );
  OAI22X1TS U1305 ( .A0(n2113), .A1(n930), .B0(n344), .B1(n962), .Y(N10205) );
  OAI22X1TS U1306 ( .A0(n2113), .A1(n929), .B0(n344), .B1(n961), .Y(N10206) );
  OAI22X1TS U1307 ( .A0(n2112), .A1(n928), .B0(n344), .B1(n960), .Y(N10207) );
  OAI22X1TS U1308 ( .A0(n2112), .A1(n927), .B0(n345), .B1(n959), .Y(N10208) );
  OAI22X1TS U1309 ( .A0(n2114), .A1(n926), .B0(n345), .B1(n958), .Y(N10209) );
  OAI22X1TS U1310 ( .A0(n2112), .A1(n925), .B0(n345), .B1(n957), .Y(N10210) );
  OAI22X1TS U1311 ( .A0(n2112), .A1(n924), .B0(n345), .B1(n956), .Y(N10211) );
  OAI22X1TS U1312 ( .A0(n2111), .A1(n923), .B0(n346), .B1(n955), .Y(N10212) );
  OAI22X1TS U1313 ( .A0(n2111), .A1(n922), .B0(n346), .B1(n954), .Y(N10213) );
  OAI22X1TS U1314 ( .A0(n2111), .A1(n921), .B0(n346), .B1(n953), .Y(N10214) );
  OAI22X1TS U1315 ( .A0(n2111), .A1(n920), .B0(n346), .B1(n952), .Y(N10215) );
  OAI22X1TS U1316 ( .A0(n2118), .A1(n919), .B0(n347), .B1(n951), .Y(N10216) );
  NAND2X1TS U1317 ( .A(n1488), .B(n116), .Y(n1244) );
  NOR2X1TS U1318 ( .A(n1545), .B(n175), .Y(n1541) );
  AOI31X1TS U1319 ( .A0(n1474), .A1(n171), .A2(n1487), .B0(n2372), .Y(n1500)
         );
  AOI31X1TS U1320 ( .A0(n170), .A1(n123), .A2(n1513), .B0(n2372), .Y(n1538) );
  OA21XLTS U1321 ( .A0(n810), .A1(n1326), .B0(n1526), .Y(n1327) );
  AOI31X1TS U1322 ( .A0(n1501), .A1(n171), .A2(n1474), .B0(n2372), .Y(n1526)
         );
  AOI221X1TS U1323 ( .A0(n170), .A1(n1487), .B0(n1475), .B1(n795), .C0(n2370), 
        .Y(n1486) );
  INVX2TS U1324 ( .A(n1447), .Y(n833) );
  AOI21X1TS U1325 ( .A0(n833), .A1(n299), .B0(n1662), .Y(n1691) );
  NAND3BX1TS U1326 ( .AN(n1501), .B(n1539), .C(n170), .Y(n1569) );
  XOR2X1TS U1327 ( .A(n999), .B(n134), .Y(n986) );
  NAND2X1TS U1328 ( .A(n991), .B(n992), .Y(n999) );
  INVX2TS U1329 ( .A(n1690), .Y(n885) );
  NAND3X1TS U1330 ( .A(n987), .B(n2373), .C(n988), .Y(n984) );
  XNOR2X1TS U1331 ( .A(n137), .B(n990), .Y(n988) );
  OR3X1TS U1332 ( .A(n983), .B(n986), .C(n985), .Y(n987) );
  AOI21X1TS U1333 ( .A0(n991), .A1(n992), .B0(n135), .Y(n990) );
  NOR2X1TS U1334 ( .A(n837), .B(n175), .Y(n1474) );
  CLKBUFX2TS U1335 ( .A(n1190), .Y(n850) );
  CLKBUFX2TS U1336 ( .A(n1190), .Y(n851) );
  CLKBUFX2TS U1337 ( .A(n1190), .Y(n852) );
  NOR2X1TS U1338 ( .A(n985), .B(n984), .Y(n3643) );
  OAI221XLTS U1339 ( .A0(n814), .A1(n31), .B0(n816), .B1(n3), .C0(n1680), .Y(
        n3202) );
  AOI222XLTS U1340 ( .A0(n141), .A1(requesterAddressIn_WEST[0]), .B0(
        requesterAddressIn_EAST[0]), .B1(n1681), .C0(
        requesterAddressIn_SOUTH[0]), .C1(n1682), .Y(n1680) );
  OAI221XLTS U1341 ( .A0(n814), .A1(n32), .B0(n816), .B1(n4), .C0(n1683), .Y(
        n3201) );
  AOI222XLTS U1342 ( .A0(n1578), .A1(requesterAddressIn_WEST[1]), .B0(
        requesterAddressIn_EAST[1]), .B1(n1681), .C0(
        requesterAddressIn_SOUTH[1]), .C1(n1682), .Y(n1683) );
  OAI221XLTS U1343 ( .A0(n814), .A1(n33), .B0(n320), .B1(n5), .C0(n1684), .Y(
        n3200) );
  AOI222XLTS U1344 ( .A0(n141), .A1(requesterAddressIn_WEST[2]), .B0(
        requesterAddressIn_EAST[2]), .B1(n1681), .C0(
        requesterAddressIn_SOUTH[2]), .C1(n1682), .Y(n1684) );
  OAI221XLTS U1345 ( .A0(n814), .A1(n34), .B0(n320), .B1(n6), .C0(n1685), .Y(
        n3199) );
  AOI222XLTS U1346 ( .A0(n1578), .A1(requesterAddressIn_WEST[3]), .B0(
        requesterAddressIn_EAST[3]), .B1(n279), .C0(
        requesterAddressIn_SOUTH[3]), .C1(n296), .Y(n1685) );
  OAI221XLTS U1347 ( .A0(n266), .A1(n35), .B0(n320), .B1(n7), .C0(n1686), .Y(
        n3198) );
  AOI222XLTS U1348 ( .A0(n141), .A1(requesterAddressIn_WEST[4]), .B0(
        requesterAddressIn_EAST[4]), .B1(n279), .C0(
        requesterAddressIn_SOUTH[4]), .C1(n296), .Y(n1686) );
  OAI221XLTS U1349 ( .A0(n266), .A1(n36), .B0(n320), .B1(n8), .C0(n1687), .Y(
        n3197) );
  AOI222XLTS U1350 ( .A0(n1578), .A1(requesterAddressIn_WEST[5]), .B0(
        requesterAddressIn_EAST[5]), .B1(n279), .C0(
        requesterAddressIn_SOUTH[5]), .C1(n296), .Y(n1687) );
  AND2X2TS U1351 ( .A(n1539), .B(n1501), .Y(n1513) );
  NOR2X1TS U1352 ( .A(n1244), .B(n328), .Y(n1243) );
  XOR2X1TS U1353 ( .A(n997), .B(n317), .Y(n1001) );
  OAI22X1TS U1354 ( .A0(n392), .A1(n2), .B0(n378), .B1(n27), .Y(N10020) );
  OAI22X1TS U1355 ( .A0(n414), .A1(n2), .B0(n399), .B1(n27), .Y(N10030) );
  OAI22X1TS U1356 ( .A0(n2119), .A1(n2), .B0(n343), .B1(n27), .Y(N10040) );
  OAI22X1TS U1357 ( .A0(n174), .A1(n31), .B0(n1376), .B1(n2218), .Y(n3203) );
  OAI22X1TS U1358 ( .A0(n172), .A1(n32), .B0(n1376), .B1(n2219), .Y(n3204) );
  OAI22X1TS U1359 ( .A0(n173), .A1(n33), .B0(n319), .B1(n2220), .Y(n3205) );
  OAI22X1TS U1360 ( .A0(n174), .A1(n34), .B0(n319), .B1(n2221), .Y(n3206) );
  OAI22X1TS U1361 ( .A0(n172), .A1(n35), .B0(n319), .B1(n2222), .Y(n3207) );
  OAI22X1TS U1362 ( .A0(n173), .A1(n36), .B0(n319), .B1(n2223), .Y(n3208) );
  NOR2X1TS U1363 ( .A(n1001), .B(n175), .Y(n996) );
  OAI32X1TS U1364 ( .A0(n1427), .A1(n553), .A2(n830), .B0(n490), .B1(n30), .Y(
        n3344) );
  INVX2TS U1365 ( .A(n1428), .Y(n830) );
  OAI21X1TS U1366 ( .A0(n1001), .A1(n114), .B0(n1429), .Y(n1427) );
  NAND2X1TS U1367 ( .A(n1761), .B(n1759), .Y(n1760) );
  NAND2X1TS U1368 ( .A(n1749), .B(n1747), .Y(n1748) );
  NAND2X1TS U1369 ( .A(n1737), .B(n1735), .Y(n1736) );
  CLKBUFX2TS U1370 ( .A(n1759), .Y(n372) );
  CLKBUFX2TS U1371 ( .A(n1747), .Y(n393) );
  CLKBUFX2TS U1372 ( .A(n1735), .Y(n414) );
  INVX2TS U1373 ( .A(n1723), .Y(n739) );
  NOR3BX1TS U1374 ( .AN(n366), .B(n2367), .C(n1761), .Y(n1750) );
  NOR3BX1TS U1375 ( .AN(n387), .B(n2368), .C(n1749), .Y(n1738) );
  NOR3BX1TS U1376 ( .AN(n410), .B(n2367), .C(n1737), .Y(n1726) );
  NOR2X1TS U1377 ( .A(n1440), .B(n298), .Y(n1435) );
  AOI211X1TS U1378 ( .A0(n1677), .A1(n1436), .B0(n1424), .C0(n1678), .Y(n1420)
         );
  NAND2X1TS U1379 ( .A(n2375), .B(n1426), .Y(n1678) );
  OAI22X1TS U1380 ( .A0(n371), .A1(n2), .B0(n358), .B1(n27), .Y(N10010) );
  NOR2BX1TS U1381 ( .AN(n135), .B(n317), .Y(n1436) );
  OR2X2TS U1382 ( .A(n1679), .B(n298), .Y(n1426) );
  AND3X2TS U1383 ( .A(n135), .B(n118), .C(n1677), .Y(n1424) );
  NAND2X1TS U1384 ( .A(n1723), .B(n1724), .Y(n1715) );
  AOI31X1TS U1385 ( .A0(n4621), .A1(n318), .A2(n1436), .B0(n1437), .Y(n1433)
         );
  CLKBUFX2TS U1386 ( .A(cacheAddressIn_WEST[0]), .Y(n2224) );
  CLKBUFX2TS U1387 ( .A(cacheAddressIn_EAST[0]), .Y(n2344) );
  CLKBUFX2TS U1388 ( .A(cacheAddressIn_WEST[1]), .Y(n2226) );
  CLKBUFX2TS U1389 ( .A(cacheAddressIn_EAST[1]), .Y(n2346) );
  CLKBUFX2TS U1390 ( .A(cacheAddressIn_WEST[2]), .Y(n2228) );
  CLKBUFX2TS U1391 ( .A(cacheAddressIn_EAST[2]), .Y(n2348) );
  CLKBUFX2TS U1392 ( .A(cacheAddressIn_WEST[3]), .Y(n2230) );
  CLKBUFX2TS U1393 ( .A(cacheAddressIn_EAST[3]), .Y(n2350) );
  CLKBUFX2TS U1394 ( .A(cacheAddressIn_WEST[4]), .Y(n2232) );
  CLKBUFX2TS U1395 ( .A(cacheAddressIn_EAST[4]), .Y(n2352) );
  CLKBUFX2TS U1396 ( .A(cacheAddressIn_WEST[5]), .Y(n2234) );
  CLKBUFX2TS U1397 ( .A(cacheAddressIn_EAST[5]), .Y(n2354) );
  CLKBUFX2TS U1398 ( .A(cacheAddressIn_WEST[6]), .Y(n2236) );
  CLKBUFX2TS U1399 ( .A(cacheAddressIn_EAST[6]), .Y(n2356) );
  CLKBUFX2TS U1400 ( .A(cacheAddressIn_WEST[7]), .Y(n2239) );
  CLKBUFX2TS U1401 ( .A(cacheAddressIn_EAST[7]), .Y(n2359) );
  CLKBUFX2TS U1402 ( .A(n2127), .Y(n2126) );
  CLKBUFX2TS U1403 ( .A(n2133), .Y(n2132) );
  CLKBUFX2TS U1404 ( .A(n2136), .Y(n2135) );
  CLKBUFX2TS U1405 ( .A(n2142), .Y(n2141) );
  CLKBUFX2TS U1406 ( .A(n2145), .Y(n2144) );
  CLKBUFX2TS U1407 ( .A(n2151), .Y(n2150) );
  CLKBUFX2TS U1408 ( .A(n2154), .Y(n2153) );
  CLKBUFX2TS U1409 ( .A(n2157), .Y(n2156) );
  CLKBUFX2TS U1410 ( .A(n2160), .Y(n2159) );
  CLKBUFX2TS U1411 ( .A(n2166), .Y(n2165) );
  CLKBUFX2TS U1412 ( .A(n2169), .Y(n2168) );
  CLKBUFX2TS U1413 ( .A(n2175), .Y(n2174) );
  CLKBUFX2TS U1414 ( .A(n2181), .Y(n2180) );
  CLKBUFX2TS U1415 ( .A(n2184), .Y(n2183) );
  CLKBUFX2TS U1416 ( .A(n2187), .Y(n2186) );
  CLKBUFX2TS U1417 ( .A(n2190), .Y(n2189) );
  CLKBUFX2TS U1418 ( .A(n2193), .Y(n2192) );
  CLKBUFX2TS U1419 ( .A(n2199), .Y(n2198) );
  CLKBUFX2TS U1420 ( .A(n2202), .Y(n2201) );
  CLKBUFX2TS U1421 ( .A(n2205), .Y(n2204) );
  CLKBUFX2TS U1422 ( .A(n2208), .Y(n2207) );
  CLKBUFX2TS U1423 ( .A(n2214), .Y(n2213) );
  CLKBUFX2TS U1424 ( .A(n2217), .Y(n2216) );
  CLKBUFX2TS U1425 ( .A(n2244), .Y(n2243) );
  CLKBUFX2TS U1426 ( .A(n2247), .Y(n2246) );
  CLKBUFX2TS U1427 ( .A(n2250), .Y(n2249) );
  CLKBUFX2TS U1428 ( .A(n2253), .Y(n2252) );
  CLKBUFX2TS U1429 ( .A(n2259), .Y(n2258) );
  CLKBUFX2TS U1430 ( .A(n2262), .Y(n2261) );
  CLKBUFX2TS U1431 ( .A(n2268), .Y(n2267) );
  CLKBUFX2TS U1432 ( .A(n2271), .Y(n2270) );
  CLKBUFX2TS U1433 ( .A(n2274), .Y(n2273) );
  CLKBUFX2TS U1434 ( .A(n2277), .Y(n2276) );
  CLKBUFX2TS U1435 ( .A(n2280), .Y(n2279) );
  CLKBUFX2TS U1436 ( .A(n2283), .Y(n2282) );
  CLKBUFX2TS U1437 ( .A(n2292), .Y(n2291) );
  CLKBUFX2TS U1438 ( .A(n2295), .Y(n2294) );
  CLKBUFX2TS U1439 ( .A(n2298), .Y(n2297) );
  CLKBUFX2TS U1440 ( .A(n2304), .Y(n2303) );
  CLKBUFX2TS U1441 ( .A(n2313), .Y(n2312) );
  CLKBUFX2TS U1442 ( .A(n2316), .Y(n2315) );
  CLKBUFX2TS U1443 ( .A(n2319), .Y(n2318) );
  CLKBUFX2TS U1444 ( .A(n2322), .Y(n2321) );
  CLKBUFX2TS U1445 ( .A(n2328), .Y(n2327) );
  CLKBUFX2TS U1446 ( .A(n2334), .Y(n2333) );
  CLKBUFX2TS U1447 ( .A(n2337), .Y(n2336) );
  CLKBUFX2TS U1448 ( .A(n1747), .Y(n394) );
  CLKBUFX2TS U1449 ( .A(n1735), .Y(n415) );
  CLKBUFX2TS U1450 ( .A(n1759), .Y(n373) );
  NOR2X1TS U1451 ( .A(n185), .B(n2366), .Y(n1381) );
  NOR2X1TS U1452 ( .A(n190), .B(n2366), .Y(n1379) );
  NOR2X1TS U1453 ( .A(n181), .B(n2366), .Y(n1378) );
  CLKBUFX2TS U1454 ( .A(n2124), .Y(n2123) );
  CLKBUFX2TS U1455 ( .A(n2130), .Y(n2129) );
  CLKBUFX2TS U1456 ( .A(n2139), .Y(n2138) );
  CLKBUFX2TS U1457 ( .A(n2148), .Y(n2147) );
  CLKBUFX2TS U1458 ( .A(n2163), .Y(n2162) );
  CLKBUFX2TS U1459 ( .A(n2172), .Y(n2171) );
  CLKBUFX2TS U1460 ( .A(n2178), .Y(n2177) );
  CLKBUFX2TS U1461 ( .A(n2196), .Y(n2195) );
  CLKBUFX2TS U1462 ( .A(n2211), .Y(n2210) );
  CLKBUFX2TS U1463 ( .A(n2256), .Y(n2255) );
  CLKBUFX2TS U1464 ( .A(n2265), .Y(n2264) );
  CLKBUFX2TS U1465 ( .A(n2286), .Y(n2285) );
  CLKBUFX2TS U1466 ( .A(n2289), .Y(n2288) );
  CLKBUFX2TS U1467 ( .A(n2301), .Y(n2300) );
  CLKBUFX2TS U1468 ( .A(n2307), .Y(n2306) );
  CLKBUFX2TS U1469 ( .A(n2310), .Y(n2309) );
  CLKBUFX2TS U1470 ( .A(n2325), .Y(n2324) );
  CLKBUFX2TS U1471 ( .A(n2331), .Y(n2330) );
  INVX2TS U1472 ( .A(requesterAddressIn_EAST[0]), .Y(n2338) );
  INVX2TS U1473 ( .A(requesterAddressIn_EAST[1]), .Y(n2339) );
  INVX2TS U1474 ( .A(requesterAddressIn_EAST[2]), .Y(n2340) );
  INVX2TS U1475 ( .A(requesterAddressIn_EAST[3]), .Y(n2341) );
  INVX2TS U1476 ( .A(requesterAddressIn_EAST[4]), .Y(n2342) );
  INVX2TS U1477 ( .A(requesterAddressIn_EAST[5]), .Y(n2343) );
  NAND3X1TS U1478 ( .A(n134), .B(n123), .C(n342), .Y(n1440) );
  INVX2TS U1479 ( .A(n185), .Y(n798) );
  NAND2X1TS U1480 ( .A(n1677), .B(n134), .Y(n1679) );
  INVX2TS U1481 ( .A(n181), .Y(n820) );
  XNOR2X1TS U1482 ( .A(n1541), .B(n910), .Y(n1540) );
  OAI221XLTS U1483 ( .A0(n2244), .A1(n849), .B0(n2123), .B1(n836), .C0(n1192), 
        .Y(n3545) );
  AOI22X1TS U1484 ( .A0(n1827), .A1(n804), .B0(n746), .B1(n1891), .Y(n1192) );
  OAI221XLTS U1485 ( .A0(n2247), .A1(n849), .B0(n2127), .B1(n836), .C0(n1195), 
        .Y(n3544) );
  AOI22X1TS U1486 ( .A0(n1828), .A1(n804), .B0(n745), .B1(n1892), .Y(n1195) );
  OAI221XLTS U1487 ( .A0(n2250), .A1(n849), .B0(n2129), .B1(n836), .C0(n1196), 
        .Y(n3543) );
  AOI22X1TS U1488 ( .A0(n1829), .A1(n804), .B0(n745), .B1(n1893), .Y(n1196) );
  OAI221XLTS U1489 ( .A0(n2253), .A1(n849), .B0(n2133), .B1(n836), .C0(n1197), 
        .Y(n3542) );
  AOI22X1TS U1490 ( .A0(n1830), .A1(n804), .B0(n745), .B1(n1894), .Y(n1197) );
  OAI221XLTS U1491 ( .A0(n2255), .A1(n848), .B0(n2136), .B1(n834), .C0(n1198), 
        .Y(n3541) );
  AOI22X1TS U1492 ( .A0(n1831), .A1(n803), .B0(n745), .B1(n1895), .Y(n1198) );
  OAI221XLTS U1493 ( .A0(n2259), .A1(n848), .B0(n2138), .B1(n834), .C0(n1199), 
        .Y(n3540) );
  AOI22X1TS U1494 ( .A0(n1832), .A1(n803), .B0(n744), .B1(n1896), .Y(n1199) );
  OAI221XLTS U1495 ( .A0(n2262), .A1(n848), .B0(n2142), .B1(n834), .C0(n1200), 
        .Y(n3539) );
  AOI22X1TS U1496 ( .A0(n1833), .A1(n803), .B0(n744), .B1(n1897), .Y(n1200) );
  OAI221XLTS U1497 ( .A0(n2264), .A1(n848), .B0(n2145), .B1(n834), .C0(n1201), 
        .Y(n3538) );
  AOI22X1TS U1498 ( .A0(n1834), .A1(n803), .B0(n744), .B1(n1898), .Y(n1201) );
  OAI221XLTS U1499 ( .A0(n2268), .A1(n847), .B0(n2147), .B1(n839), .C0(n1202), 
        .Y(n3537) );
  AOI22X1TS U1500 ( .A0(n1835), .A1(n808), .B0(n744), .B1(n1899), .Y(n1202) );
  OAI221XLTS U1501 ( .A0(n2271), .A1(n847), .B0(n2151), .B1(n839), .C0(n1203), 
        .Y(n3536) );
  AOI22X1TS U1502 ( .A0(n1836), .A1(n808), .B0(n743), .B1(n1900), .Y(n1203) );
  OAI221XLTS U1503 ( .A0(n2274), .A1(n847), .B0(n2154), .B1(n841), .C0(n1204), 
        .Y(n3535) );
  AOI22X1TS U1504 ( .A0(n1837), .A1(n808), .B0(n743), .B1(n1901), .Y(n1204) );
  OAI221XLTS U1505 ( .A0(n2277), .A1(n847), .B0(n2157), .B1(n841), .C0(n1205), 
        .Y(n3534) );
  AOI22X1TS U1506 ( .A0(n1838), .A1(n809), .B0(n743), .B1(n1902), .Y(n1205) );
  OAI221XLTS U1507 ( .A0(n2280), .A1(n846), .B0(n2160), .B1(n839), .C0(n1206), 
        .Y(n3533) );
  AOI22X1TS U1508 ( .A0(n1839), .A1(n808), .B0(n743), .B1(n1903), .Y(n1206) );
  OAI221XLTS U1509 ( .A0(n2283), .A1(n846), .B0(n2162), .B1(n839), .C0(n1207), 
        .Y(n3532) );
  AOI22X1TS U1510 ( .A0(n1840), .A1(n809), .B0(n742), .B1(n1904), .Y(n1207) );
  OAI221XLTS U1511 ( .A0(n2285), .A1(n846), .B0(n2166), .B1(n838), .C0(n1208), 
        .Y(n3531) );
  AOI22X1TS U1512 ( .A0(n1841), .A1(n815), .B0(n742), .B1(n1905), .Y(n1208) );
  OAI221XLTS U1513 ( .A0(n2288), .A1(n846), .B0(n2169), .B1(n840), .C0(n1209), 
        .Y(n3530) );
  AOI22X1TS U1514 ( .A0(n1842), .A1(n805), .B0(n742), .B1(n1906), .Y(n1209) );
  OAI221XLTS U1515 ( .A0(n2292), .A1(n852), .B0(n2171), .B1(n829), .C0(n1210), 
        .Y(n3529) );
  AOI22X1TS U1516 ( .A0(n1843), .A1(n755), .B0(n742), .B1(n1907), .Y(n1210) );
  OAI221XLTS U1517 ( .A0(n2295), .A1(n850), .B0(n2175), .B1(n829), .C0(n1211), 
        .Y(n3528) );
  AOI22X1TS U1518 ( .A0(n1844), .A1(n755), .B0(n748), .B1(n1908), .Y(n1211) );
  OAI221XLTS U1519 ( .A0(n2298), .A1(n850), .B0(n2177), .B1(n829), .C0(n1212), 
        .Y(n3527) );
  AOI22X1TS U1520 ( .A0(n1845), .A1(n755), .B0(n748), .B1(n1909), .Y(n1212) );
  OAI221XLTS U1521 ( .A0(n2300), .A1(n851), .B0(n2181), .B1(n829), .C0(n1213), 
        .Y(n3526) );
  AOI22X1TS U1522 ( .A0(n1846), .A1(n755), .B0(n747), .B1(n1910), .Y(n1213) );
  OAI221XLTS U1523 ( .A0(n2304), .A1(n845), .B0(n2184), .B1(n826), .C0(n1214), 
        .Y(n3525) );
  AOI22X1TS U1524 ( .A0(n1847), .A1(n754), .B0(n751), .B1(n1911), .Y(n1214) );
  OAI221XLTS U1525 ( .A0(n2306), .A1(n845), .B0(n2187), .B1(n826), .C0(n1215), 
        .Y(n3524) );
  AOI22X1TS U1526 ( .A0(n1848), .A1(n754), .B0(n749), .B1(n1912), .Y(n1215) );
  OAI221XLTS U1527 ( .A0(n2309), .A1(n845), .B0(n2190), .B1(n826), .C0(n1216), 
        .Y(n3523) );
  AOI22X1TS U1528 ( .A0(n1849), .A1(n754), .B0(n749), .B1(n1913), .Y(n1216) );
  OAI221XLTS U1529 ( .A0(n2313), .A1(n845), .B0(n2193), .B1(n826), .C0(n1217), 
        .Y(n3522) );
  AOI22X1TS U1530 ( .A0(n1850), .A1(n754), .B0(n749), .B1(n1914), .Y(n1217) );
  OAI221XLTS U1531 ( .A0(n2316), .A1(n843), .B0(n2195), .B1(n823), .C0(n1218), 
        .Y(n3521) );
  AOI22X1TS U1532 ( .A0(n1851), .A1(n753), .B0(n748), .B1(n1915), .Y(n1218) );
  OAI221XLTS U1533 ( .A0(n2319), .A1(n843), .B0(n2199), .B1(n823), .C0(n1227), 
        .Y(n3520) );
  AOI22X1TS U1534 ( .A0(n1852), .A1(n753), .B0(n747), .B1(n1916), .Y(n1227) );
  OAI221XLTS U1535 ( .A0(n2322), .A1(n843), .B0(n2202), .B1(n823), .C0(n1228), 
        .Y(n3519) );
  AOI22X1TS U1536 ( .A0(n1853), .A1(n753), .B0(n749), .B1(n1917), .Y(n1228) );
  OAI221XLTS U1537 ( .A0(n2324), .A1(n843), .B0(n2205), .B1(n823), .C0(n1229), 
        .Y(n3518) );
  AOI22X1TS U1538 ( .A0(n1854), .A1(n753), .B0(n746), .B1(n1918), .Y(n1229) );
  OAI221XLTS U1539 ( .A0(n2328), .A1(n842), .B0(n2208), .B1(n817), .C0(n1230), 
        .Y(n3517) );
  AOI22X1TS U1540 ( .A0(n1855), .A1(n752), .B0(n751), .B1(n1919), .Y(n1230) );
  OAI221XLTS U1541 ( .A0(n2330), .A1(n842), .B0(n2210), .B1(n817), .C0(n1231), 
        .Y(n3516) );
  AOI22X1TS U1542 ( .A0(n1856), .A1(n752), .B0(n750), .B1(n1920), .Y(n1231) );
  OAI221XLTS U1543 ( .A0(n2334), .A1(n842), .B0(n2214), .B1(n817), .C0(n1232), 
        .Y(n3515) );
  AOI22X1TS U1544 ( .A0(n1857), .A1(n752), .B0(n746), .B1(n1921), .Y(n1232) );
  OAI221XLTS U1545 ( .A0(n2337), .A1(n842), .B0(n2217), .B1(n817), .C0(n1233), 
        .Y(n3514) );
  AOI22X1TS U1546 ( .A0(n1858), .A1(n752), .B0(n1194), .B1(n1922), .Y(n1233)
         );
  OAI221XLTS U1547 ( .A0(n1660), .A1(n80), .B0(n1324), .B1(n630), .C0(n1042), 
        .Y(n3609) );
  OAI221XLTS U1548 ( .A0(n1660), .A1(n81), .B0(n1324), .B1(n629), .C0(n1045), 
        .Y(n3608) );
  OAI221XLTS U1549 ( .A0(n2244), .A1(n894), .B0(n2123), .B1(n883), .C0(n1113), 
        .Y(n3577) );
  AOI2BB2X1TS U1550 ( .B0(n1763), .B1(n1114), .A0N(n864), .A1N(n1103), .Y(
        n1113) );
  OAI221XLTS U1551 ( .A0(n2247), .A1(n894), .B0(n2127), .B1(n883), .C0(n1116), 
        .Y(n3576) );
  AOI2BB2X1TS U1552 ( .B0(n1765), .B1(n875), .A0N(n855), .A1N(n1102), .Y(n1116) );
  OAI221XLTS U1553 ( .A0(n2250), .A1(n894), .B0(n2129), .B1(n883), .C0(n1117), 
        .Y(n3575) );
  AOI2BB2X1TS U1554 ( .B0(n1767), .B1(n873), .A0N(n855), .A1N(n1101), .Y(n1117) );
  OAI221XLTS U1555 ( .A0(n2253), .A1(n894), .B0(n2133), .B1(n883), .C0(n1118), 
        .Y(n3574) );
  AOI2BB2X1TS U1556 ( .B0(n1769), .B1(n874), .A0N(n855), .A1N(n1100), .Y(n1118) );
  OAI221XLTS U1557 ( .A0(n2255), .A1(n893), .B0(n2136), .B1(n884), .C0(n1119), 
        .Y(n3573) );
  AOI2BB2X1TS U1558 ( .B0(n1771), .B1(n872), .A0N(n856), .A1N(n1099), .Y(n1119) );
  OAI221XLTS U1559 ( .A0(n2259), .A1(n893), .B0(n2138), .B1(n887), .C0(n1120), 
        .Y(n3572) );
  AOI2BB2X1TS U1560 ( .B0(n1773), .B1(n872), .A0N(n856), .A1N(n1098), .Y(n1120) );
  OAI221XLTS U1561 ( .A0(n2262), .A1(n893), .B0(n2142), .B1(n884), .C0(n1121), 
        .Y(n3571) );
  AOI2BB2X1TS U1562 ( .B0(n1775), .B1(n872), .A0N(n856), .A1N(n1097), .Y(n1121) );
  OAI221XLTS U1563 ( .A0(n2264), .A1(n893), .B0(n2145), .B1(n887), .C0(n1122), 
        .Y(n3570) );
  AOI2BB2X1TS U1564 ( .B0(n1777), .B1(n872), .A0N(n856), .A1N(n1096), .Y(n1122) );
  OAI221XLTS U1565 ( .A0(n2268), .A1(n892), .B0(n2147), .B1(n882), .C0(n1123), 
        .Y(n3569) );
  AOI2BB2X1TS U1566 ( .B0(n1779), .B1(n871), .A0N(n857), .A1N(n1095), .Y(n1123) );
  OAI221XLTS U1567 ( .A0(n2271), .A1(n892), .B0(n2151), .B1(n882), .C0(n1124), 
        .Y(n3568) );
  AOI2BB2X1TS U1568 ( .B0(n1781), .B1(n871), .A0N(n857), .A1N(n1094), .Y(n1124) );
  OAI221XLTS U1569 ( .A0(n2274), .A1(n892), .B0(n2154), .B1(n882), .C0(n1125), 
        .Y(n3567) );
  AOI2BB2X1TS U1570 ( .B0(n1783), .B1(n871), .A0N(n857), .A1N(n1093), .Y(n1125) );
  OAI221XLTS U1571 ( .A0(n2277), .A1(n892), .B0(n2157), .B1(n882), .C0(n1126), 
        .Y(n3566) );
  AOI2BB2X1TS U1572 ( .B0(n1785), .B1(n871), .A0N(n857), .A1N(n1092), .Y(n1126) );
  OAI221XLTS U1573 ( .A0(n2280), .A1(n891), .B0(n2160), .B1(n881), .C0(n1127), 
        .Y(n3565) );
  AOI2BB2X1TS U1574 ( .B0(n1787), .B1(n870), .A0N(n858), .A1N(n1091), .Y(n1127) );
  OAI221XLTS U1575 ( .A0(n2283), .A1(n891), .B0(n2162), .B1(n881), .C0(n1128), 
        .Y(n3564) );
  AOI2BB2X1TS U1576 ( .B0(n1789), .B1(n870), .A0N(n858), .A1N(n1090), .Y(n1128) );
  OAI221XLTS U1577 ( .A0(n2285), .A1(n891), .B0(n2166), .B1(n881), .C0(n1129), 
        .Y(n3563) );
  AOI2BB2X1TS U1578 ( .B0(n1791), .B1(n870), .A0N(n858), .A1N(n1089), .Y(n1129) );
  OAI221XLTS U1579 ( .A0(n2288), .A1(n891), .B0(n2169), .B1(n881), .C0(n1130), 
        .Y(n3562) );
  AOI2BB2X1TS U1580 ( .B0(n1793), .B1(n870), .A0N(n858), .A1N(n1088), .Y(n1130) );
  OAI221XLTS U1581 ( .A0(n2292), .A1(n890), .B0(n2171), .B1(n879), .C0(n1131), 
        .Y(n3561) );
  AOI2BB2X1TS U1582 ( .B0(n1795), .B1(n869), .A0N(n864), .A1N(n1087), .Y(n1131) );
  OAI221XLTS U1583 ( .A0(n2295), .A1(n890), .B0(n2175), .B1(n879), .C0(n1132), 
        .Y(n3560) );
  AOI2BB2X1TS U1584 ( .B0(n1797), .B1(n869), .A0N(n864), .A1N(n1086), .Y(n1132) );
  OAI221XLTS U1585 ( .A0(n2298), .A1(n890), .B0(n2177), .B1(n879), .C0(n1133), 
        .Y(n3559) );
  AOI2BB2X1TS U1586 ( .B0(n1799), .B1(n869), .A0N(n1115), .A1N(n1085), .Y(
        n1133) );
  OAI221XLTS U1587 ( .A0(n2300), .A1(n890), .B0(n2181), .B1(n879), .C0(n1134), 
        .Y(n3558) );
  AOI2BB2X1TS U1588 ( .B0(n1801), .B1(n869), .A0N(n859), .A1N(n1084), .Y(n1134) );
  OAI221XLTS U1589 ( .A0(n2304), .A1(n897), .B0(n2184), .B1(n878), .C0(n1135), 
        .Y(n3557) );
  AOI2BB2X1TS U1590 ( .B0(n1803), .B1(n868), .A0N(n859), .A1N(n1083), .Y(n1135) );
  OAI221XLTS U1591 ( .A0(n2306), .A1(n897), .B0(n2187), .B1(n878), .C0(n1168), 
        .Y(n3556) );
  AOI2BB2X1TS U1592 ( .B0(n1805), .B1(n868), .A0N(n859), .A1N(n1082), .Y(n1168) );
  OAI221XLTS U1593 ( .A0(n2309), .A1(n897), .B0(n2190), .B1(n878), .C0(n1176), 
        .Y(n3555) );
  AOI2BB2X1TS U1594 ( .B0(n1807), .B1(n868), .A0N(n859), .A1N(n1081), .Y(n1176) );
  OAI221XLTS U1595 ( .A0(n2313), .A1(n895), .B0(n2193), .B1(n878), .C0(n1177), 
        .Y(n3554) );
  AOI2BB2X1TS U1596 ( .B0(n1809), .B1(n868), .A0N(n860), .A1N(n1080), .Y(n1177) );
  OAI221XLTS U1597 ( .A0(n2316), .A1(n889), .B0(n2195), .B1(n877), .C0(n1178), 
        .Y(n3553) );
  AOI2BB2X1TS U1598 ( .B0(n1811), .B1(n867), .A0N(n860), .A1N(n1079), .Y(n1178) );
  OAI221XLTS U1599 ( .A0(n2319), .A1(n889), .B0(n2199), .B1(n877), .C0(n1179), 
        .Y(n3552) );
  AOI2BB2X1TS U1600 ( .B0(n1813), .B1(n867), .A0N(n860), .A1N(n1078), .Y(n1179) );
  OAI221XLTS U1601 ( .A0(n2322), .A1(n889), .B0(n2202), .B1(n877), .C0(n1180), 
        .Y(n3551) );
  AOI2BB2X1TS U1602 ( .B0(n1815), .B1(n867), .A0N(n860), .A1N(n1077), .Y(n1180) );
  OAI221XLTS U1603 ( .A0(n2324), .A1(n889), .B0(n2205), .B1(n877), .C0(n1181), 
        .Y(n3550) );
  AOI2BB2X1TS U1604 ( .B0(n1817), .B1(n867), .A0N(n863), .A1N(n1076), .Y(n1181) );
  OAI221XLTS U1605 ( .A0(n2328), .A1(n888), .B0(n2208), .B1(n876), .C0(n1182), 
        .Y(n3549) );
  AOI2BB2X1TS U1606 ( .B0(n1819), .B1(n866), .A0N(n861), .A1N(n1075), .Y(n1182) );
  OAI221XLTS U1607 ( .A0(n2330), .A1(n888), .B0(n2210), .B1(n876), .C0(n1183), 
        .Y(n3548) );
  AOI2BB2X1TS U1608 ( .B0(n1821), .B1(n866), .A0N(n862), .A1N(n1074), .Y(n1183) );
  OAI221XLTS U1609 ( .A0(n2334), .A1(n888), .B0(n2214), .B1(n876), .C0(n1184), 
        .Y(n3547) );
  AOI2BB2X1TS U1610 ( .B0(n1823), .B1(n866), .A0N(n862), .A1N(n1073), .Y(n1184) );
  OAI221XLTS U1611 ( .A0(n2337), .A1(n888), .B0(n2217), .B1(n876), .C0(n1185), 
        .Y(n3546) );
  AOI2BB2X1TS U1612 ( .B0(n1825), .B1(n866), .A0N(n861), .A1N(n1072), .Y(n1185) );
  OAI221XLTS U1613 ( .A0(n2243), .A1(n713), .B0(n2124), .B1(n703), .C0(n1248), 
        .Y(n3513) );
  AOI22X1TS U1614 ( .A0(n1764), .A1(n694), .B0(n680), .B1(n1763), .Y(n1248) );
  OAI221XLTS U1615 ( .A0(n2243), .A1(n594), .B0(n2123), .B1(n584), .C0(n1330), 
        .Y(n3449) );
  AOI22X1TS U1616 ( .A0(n575), .A1(n736), .B0(n564), .B1(n1764), .Y(n1330) );
  OAI221XLTS U1617 ( .A0(n2246), .A1(n713), .B0(n2126), .B1(n703), .C0(n1251), 
        .Y(n3512) );
  OAI221XLTS U1618 ( .A0(n2246), .A1(n594), .B0(n2126), .B1(n584), .C0(n1333), 
        .Y(n3448) );
  AOI22X1TS U1619 ( .A0(n575), .A1(n735), .B0(n563), .B1(n1766), .Y(n1333) );
  OAI221XLTS U1620 ( .A0(n2249), .A1(n713), .B0(n2130), .B1(n703), .C0(n1252), 
        .Y(n3511) );
  OAI221XLTS U1621 ( .A0(n2249), .A1(n631), .B0(n2129), .B1(n584), .C0(n1334), 
        .Y(n3447) );
  AOI22X1TS U1622 ( .A0(n575), .A1(n734), .B0(n563), .B1(n1768), .Y(n1334) );
  OAI221XLTS U1623 ( .A0(n2252), .A1(n713), .B0(n2132), .B1(n703), .C0(n1253), 
        .Y(n3510) );
  OAI221XLTS U1624 ( .A0(n2252), .A1(n631), .B0(n2132), .B1(n584), .C0(n1335), 
        .Y(n3446) );
  AOI22X1TS U1625 ( .A0(n575), .A1(n733), .B0(n563), .B1(n1770), .Y(n1335) );
  OAI221XLTS U1626 ( .A0(n2256), .A1(n712), .B0(n2135), .B1(n702), .C0(n1254), 
        .Y(n3509) );
  AOI22X1TS U1627 ( .A0(n1772), .A1(n693), .B0(n679), .B1(n1771), .Y(n1254) );
  OAI221XLTS U1628 ( .A0(n2255), .A1(n594), .B0(n2135), .B1(n583), .C0(n1336), 
        .Y(n3445) );
  AOI22X1TS U1629 ( .A0(n574), .A1(n732), .B0(n563), .B1(n1772), .Y(n1336) );
  OAI221XLTS U1630 ( .A0(n2258), .A1(n712), .B0(n2139), .B1(n702), .C0(n1255), 
        .Y(n3508) );
  OAI221XLTS U1631 ( .A0(n2258), .A1(n594), .B0(n2138), .B1(n583), .C0(n1337), 
        .Y(n3444) );
  AOI22X1TS U1632 ( .A0(n574), .A1(n731), .B0(n562), .B1(n1774), .Y(n1337) );
  OAI221XLTS U1633 ( .A0(n2261), .A1(n712), .B0(n2141), .B1(n702), .C0(n1256), 
        .Y(n3507) );
  OAI221XLTS U1634 ( .A0(n2261), .A1(n595), .B0(n2141), .B1(n583), .C0(n1338), 
        .Y(n3443) );
  AOI22X1TS U1635 ( .A0(n574), .A1(n730), .B0(n562), .B1(n1776), .Y(n1338) );
  OAI221XLTS U1636 ( .A0(n2265), .A1(n712), .B0(n2144), .B1(n702), .C0(n1257), 
        .Y(n3506) );
  OAI221XLTS U1637 ( .A0(n2264), .A1(n598), .B0(n2144), .B1(n583), .C0(n1339), 
        .Y(n3442) );
  AOI22X1TS U1638 ( .A0(n574), .A1(n729), .B0(n562), .B1(n1778), .Y(n1339) );
  OAI221XLTS U1639 ( .A0(n2267), .A1(n711), .B0(n2148), .B1(n701), .C0(n1258), 
        .Y(n3505) );
  AOI22X1TS U1640 ( .A0(n1780), .A1(n692), .B0(n678), .B1(n1779), .Y(n1258) );
  OAI221XLTS U1641 ( .A0(n2267), .A1(n593), .B0(n2147), .B1(n582), .C0(n1340), 
        .Y(n3441) );
  AOI22X1TS U1642 ( .A0(n573), .A1(n728), .B0(n562), .B1(n1780), .Y(n1340) );
  OAI221XLTS U1643 ( .A0(n2270), .A1(n711), .B0(n2150), .B1(n701), .C0(n1259), 
        .Y(n3504) );
  OAI221XLTS U1644 ( .A0(n2270), .A1(n593), .B0(n2150), .B1(n582), .C0(n1341), 
        .Y(n3440) );
  AOI22X1TS U1645 ( .A0(n573), .A1(n727), .B0(n561), .B1(n1782), .Y(n1341) );
  OAI221XLTS U1646 ( .A0(n2273), .A1(n711), .B0(n2153), .B1(n701), .C0(n1260), 
        .Y(n3503) );
  OAI221XLTS U1647 ( .A0(n2273), .A1(n593), .B0(n2153), .B1(n582), .C0(n1342), 
        .Y(n3439) );
  AOI22X1TS U1648 ( .A0(n573), .A1(n726), .B0(n561), .B1(n1784), .Y(n1342) );
  OAI221XLTS U1649 ( .A0(n2276), .A1(n711), .B0(n2156), .B1(n701), .C0(n1261), 
        .Y(n3502) );
  OAI221XLTS U1650 ( .A0(n2276), .A1(n593), .B0(n2156), .B1(n582), .C0(n1343), 
        .Y(n3438) );
  AOI22X1TS U1651 ( .A0(n573), .A1(n725), .B0(n561), .B1(n1786), .Y(n1343) );
  OAI221XLTS U1652 ( .A0(n2279), .A1(n710), .B0(n2159), .B1(n700), .C0(n1262), 
        .Y(n3501) );
  AOI22X1TS U1653 ( .A0(n1788), .A1(n691), .B0(n677), .B1(n1787), .Y(n1262) );
  OAI221XLTS U1654 ( .A0(n2279), .A1(n592), .B0(n2159), .B1(n581), .C0(n1344), 
        .Y(n3437) );
  AOI22X1TS U1655 ( .A0(n572), .A1(n724), .B0(n561), .B1(n1788), .Y(n1344) );
  OAI221XLTS U1656 ( .A0(n2282), .A1(n710), .B0(n2163), .B1(n700), .C0(n1263), 
        .Y(n3500) );
  OAI221XLTS U1657 ( .A0(n2282), .A1(n592), .B0(n2162), .B1(n581), .C0(n1345), 
        .Y(n3436) );
  AOI22X1TS U1658 ( .A0(n572), .A1(n723), .B0(n565), .B1(n1790), .Y(n1345) );
  OAI221XLTS U1659 ( .A0(n2286), .A1(n710), .B0(n2165), .B1(n700), .C0(n1264), 
        .Y(n3499) );
  OAI221XLTS U1660 ( .A0(n2285), .A1(n592), .B0(n2165), .B1(n581), .C0(n1346), 
        .Y(n3435) );
  AOI22X1TS U1661 ( .A0(n572), .A1(n722), .B0(n567), .B1(n1792), .Y(n1346) );
  OAI221XLTS U1662 ( .A0(n2289), .A1(n710), .B0(n2168), .B1(n700), .C0(n1265), 
        .Y(n3498) );
  OAI221XLTS U1663 ( .A0(n2288), .A1(n592), .B0(n2168), .B1(n581), .C0(n1347), 
        .Y(n3434) );
  AOI22X1TS U1664 ( .A0(n572), .A1(n721), .B0(n564), .B1(n1794), .Y(n1347) );
  OAI221XLTS U1665 ( .A0(n2291), .A1(n709), .B0(n2172), .B1(n705), .C0(n1266), 
        .Y(n3497) );
  AOI22X1TS U1666 ( .A0(n1796), .A1(n690), .B0(n684), .B1(n1795), .Y(n1266) );
  OAI221XLTS U1667 ( .A0(n2291), .A1(n591), .B0(n2171), .B1(n580), .C0(n1348), 
        .Y(n3433) );
  AOI22X1TS U1668 ( .A0(n571), .A1(n720), .B0(n567), .B1(n1796), .Y(n1348) );
  OAI221XLTS U1669 ( .A0(n2294), .A1(n709), .B0(n2174), .B1(n706), .C0(n1267), 
        .Y(n3496) );
  OAI221XLTS U1670 ( .A0(n2294), .A1(n591), .B0(n2174), .B1(n580), .C0(n1349), 
        .Y(n3432) );
  AOI22X1TS U1671 ( .A0(n571), .A1(n719), .B0(n560), .B1(n1798), .Y(n1349) );
  OAI221XLTS U1672 ( .A0(n2297), .A1(n709), .B0(n2178), .B1(n704), .C0(n1268), 
        .Y(n3495) );
  OAI221XLTS U1673 ( .A0(n2297), .A1(n591), .B0(n2177), .B1(n580), .C0(n1350), 
        .Y(n3431) );
  AOI22X1TS U1674 ( .A0(n571), .A1(n718), .B0(n560), .B1(n1800), .Y(n1350) );
  OAI221XLTS U1675 ( .A0(n2301), .A1(n709), .B0(n2180), .B1(n704), .C0(n1269), 
        .Y(n3494) );
  OAI221XLTS U1676 ( .A0(n2300), .A1(n591), .B0(n2180), .B1(n580), .C0(n1351), 
        .Y(n3430) );
  AOI22X1TS U1677 ( .A0(n571), .A1(n717), .B0(n560), .B1(n1802), .Y(n1351) );
  OAI221XLTS U1678 ( .A0(n2303), .A1(n714), .B0(n2183), .B1(n699), .C0(n1270), 
        .Y(n3493) );
  AOI22X1TS U1679 ( .A0(n1804), .A1(n689), .B0(n686), .B1(n1803), .Y(n1270) );
  OAI221XLTS U1680 ( .A0(n2303), .A1(n590), .B0(n2183), .B1(n587), .C0(n1352), 
        .Y(n3429) );
  AOI22X1TS U1681 ( .A0(n570), .A1(n716), .B0(n560), .B1(n1804), .Y(n1352) );
  OAI221XLTS U1682 ( .A0(n2307), .A1(n738), .B0(n2186), .B1(n699), .C0(n1271), 
        .Y(n3492) );
  OAI221XLTS U1683 ( .A0(n2306), .A1(n590), .B0(n2186), .B1(n587), .C0(n1353), 
        .Y(n3428) );
  AOI22X1TS U1684 ( .A0(n570), .A1(n793), .B0(n559), .B1(n1806), .Y(n1353) );
  OAI221XLTS U1685 ( .A0(n2310), .A1(n738), .B0(n2189), .B1(n699), .C0(n1272), 
        .Y(n3491) );
  OAI221XLTS U1686 ( .A0(n2309), .A1(n590), .B0(n2189), .B1(n587), .C0(n1354), 
        .Y(n3427) );
  AOI22X1TS U1687 ( .A0(n570), .A1(n792), .B0(n559), .B1(n1808), .Y(n1354) );
  OAI221XLTS U1688 ( .A0(n2312), .A1(n738), .B0(n2192), .B1(n699), .C0(n1273), 
        .Y(n3490) );
  OAI221XLTS U1689 ( .A0(n2312), .A1(n590), .B0(n2192), .B1(n585), .C0(n1355), 
        .Y(n3426) );
  AOI22X1TS U1690 ( .A0(n570), .A1(n791), .B0(n559), .B1(n1810), .Y(n1355) );
  OAI221XLTS U1691 ( .A0(n2315), .A1(n708), .B0(n2196), .B1(n698), .C0(n1274), 
        .Y(n3489) );
  AOI22X1TS U1692 ( .A0(n1812), .A1(n688), .B0(n682), .B1(n1811), .Y(n1274) );
  OAI221XLTS U1693 ( .A0(n2315), .A1(n589), .B0(n2195), .B1(n579), .C0(n1356), 
        .Y(n3425) );
  AOI22X1TS U1694 ( .A0(n569), .A1(n790), .B0(n559), .B1(n1812), .Y(n1356) );
  OAI221XLTS U1695 ( .A0(n2318), .A1(n708), .B0(n2198), .B1(n698), .C0(n1275), 
        .Y(n3488) );
  OAI221XLTS U1696 ( .A0(n2318), .A1(n589), .B0(n2198), .B1(n579), .C0(n1357), 
        .Y(n3424) );
  AOI22X1TS U1697 ( .A0(n569), .A1(n789), .B0(n558), .B1(n1814), .Y(n1357) );
  OAI221XLTS U1698 ( .A0(n2321), .A1(n708), .B0(n2201), .B1(n698), .C0(n1276), 
        .Y(n3487) );
  OAI221XLTS U1699 ( .A0(n2321), .A1(n589), .B0(n2201), .B1(n579), .C0(n1358), 
        .Y(n3423) );
  AOI22X1TS U1700 ( .A0(n569), .A1(n788), .B0(n558), .B1(n1816), .Y(n1358) );
  OAI221XLTS U1701 ( .A0(n2325), .A1(n708), .B0(n2204), .B1(n698), .C0(n1277), 
        .Y(n3486) );
  OAI221XLTS U1702 ( .A0(n2324), .A1(n589), .B0(n2204), .B1(n579), .C0(n1359), 
        .Y(n3422) );
  AOI22X1TS U1703 ( .A0(n569), .A1(n787), .B0(n558), .B1(n1818), .Y(n1359) );
  OAI221XLTS U1704 ( .A0(n2327), .A1(n707), .B0(n2207), .B1(n697), .C0(n1278), 
        .Y(n3485) );
  AOI22X1TS U1705 ( .A0(n1820), .A1(n687), .B0(n686), .B1(n1819), .Y(n1278) );
  OAI221XLTS U1706 ( .A0(n2327), .A1(n588), .B0(n2207), .B1(n578), .C0(n1360), 
        .Y(n3421) );
  AOI22X1TS U1707 ( .A0(n568), .A1(n786), .B0(n558), .B1(n1820), .Y(n1360) );
  OAI221XLTS U1708 ( .A0(n2331), .A1(n707), .B0(n2211), .B1(n697), .C0(n1279), 
        .Y(n3484) );
  OAI221XLTS U1709 ( .A0(n2330), .A1(n588), .B0(n2210), .B1(n578), .C0(n1361), 
        .Y(n3420) );
  AOI22X1TS U1710 ( .A0(n568), .A1(n785), .B0(n566), .B1(n1822), .Y(n1361) );
  OAI221XLTS U1711 ( .A0(n2333), .A1(n707), .B0(n2213), .B1(n697), .C0(n1280), 
        .Y(n3483) );
  OAI221XLTS U1712 ( .A0(n2333), .A1(n588), .B0(n2213), .B1(n578), .C0(n1362), 
        .Y(n3419) );
  AOI22X1TS U1713 ( .A0(n568), .A1(n784), .B0(n1332), .B1(n1824), .Y(n1362) );
  OAI221XLTS U1714 ( .A0(n2336), .A1(n707), .B0(n2216), .B1(n697), .C0(n1281), 
        .Y(n3482) );
  OAI221XLTS U1715 ( .A0(n2336), .A1(n588), .B0(n2216), .B1(n578), .C0(n1363), 
        .Y(n3418) );
  AOI22X1TS U1716 ( .A0(n568), .A1(n783), .B0(n566), .B1(n1826), .Y(n1363) );
  OAI221XLTS U1717 ( .A0(n2243), .A1(n676), .B0(n2123), .B1(n663), .C0(n1289), 
        .Y(n3481) );
  AOI22X1TS U1718 ( .A0(n1931), .A1(n653), .B0(n638), .B1(n1827), .Y(n1289) );
  OAI221XLTS U1719 ( .A0(n2246), .A1(n674), .B0(n2126), .B1(n663), .C0(n1292), 
        .Y(n3480) );
  AOI22X1TS U1720 ( .A0(n1932), .A1(n653), .B0(n637), .B1(n1828), .Y(n1292) );
  OAI221XLTS U1721 ( .A0(n2249), .A1(n674), .B0(n2129), .B1(n663), .C0(n1293), 
        .Y(n3479) );
  AOI22X1TS U1722 ( .A0(n1933), .A1(n653), .B0(n637), .B1(n1829), .Y(n1293) );
  OAI221XLTS U1723 ( .A0(n2252), .A1(n675), .B0(n2132), .B1(n663), .C0(n1294), 
        .Y(n3478) );
  AOI22X1TS U1724 ( .A0(n1934), .A1(n653), .B0(n637), .B1(n1830), .Y(n1294) );
  OAI221XLTS U1725 ( .A0(n2255), .A1(n673), .B0(n2135), .B1(n664), .C0(n1295), 
        .Y(n3477) );
  AOI22X1TS U1726 ( .A0(n1935), .A1(n654), .B0(n637), .B1(n1831), .Y(n1295) );
  OAI221XLTS U1727 ( .A0(n2258), .A1(n673), .B0(n2138), .B1(n666), .C0(n1296), 
        .Y(n3476) );
  AOI22X1TS U1728 ( .A0(n1936), .A1(n654), .B0(n636), .B1(n1832), .Y(n1296) );
  OAI221XLTS U1729 ( .A0(n2261), .A1(n673), .B0(n2141), .B1(n664), .C0(n1297), 
        .Y(n3475) );
  AOI22X1TS U1730 ( .A0(n1937), .A1(n655), .B0(n636), .B1(n1833), .Y(n1297) );
  OAI221XLTS U1731 ( .A0(n2264), .A1(n673), .B0(n2144), .B1(n666), .C0(n1298), 
        .Y(n3474) );
  AOI22X1TS U1732 ( .A0(n1938), .A1(n656), .B0(n636), .B1(n1834), .Y(n1298) );
  OAI221XLTS U1733 ( .A0(n2267), .A1(n672), .B0(n2147), .B1(n662), .C0(n1299), 
        .Y(n3473) );
  AOI22X1TS U1734 ( .A0(n1939), .A1(n652), .B0(n636), .B1(n1835), .Y(n1299) );
  OAI221XLTS U1735 ( .A0(n2270), .A1(n672), .B0(n2150), .B1(n662), .C0(n1300), 
        .Y(n3472) );
  AOI22X1TS U1736 ( .A0(n1940), .A1(n652), .B0(n635), .B1(n1836), .Y(n1300) );
  OAI221XLTS U1737 ( .A0(n2273), .A1(n672), .B0(n2153), .B1(n662), .C0(n1301), 
        .Y(n3471) );
  AOI22X1TS U1738 ( .A0(n1941), .A1(n652), .B0(n635), .B1(n1837), .Y(n1301) );
  OAI221XLTS U1739 ( .A0(n2276), .A1(n672), .B0(n2156), .B1(n662), .C0(n1302), 
        .Y(n3470) );
  AOI22X1TS U1740 ( .A0(n1942), .A1(n652), .B0(n635), .B1(n1838), .Y(n1302) );
  OAI221XLTS U1741 ( .A0(n2279), .A1(n671), .B0(n2159), .B1(n661), .C0(n1303), 
        .Y(n3469) );
  AOI22X1TS U1742 ( .A0(n1943), .A1(n651), .B0(n635), .B1(n1839), .Y(n1303) );
  OAI221XLTS U1743 ( .A0(n2282), .A1(n671), .B0(n2162), .B1(n661), .C0(n1304), 
        .Y(n3468) );
  AOI22X1TS U1744 ( .A0(n1944), .A1(n651), .B0(n639), .B1(n1840), .Y(n1304) );
  OAI221XLTS U1745 ( .A0(n2285), .A1(n671), .B0(n2165), .B1(n661), .C0(n1305), 
        .Y(n3467) );
  AOI22X1TS U1746 ( .A0(n1945), .A1(n651), .B0(n1291), .B1(n1841), .Y(n1305)
         );
  OAI221XLTS U1747 ( .A0(n2288), .A1(n671), .B0(n2168), .B1(n661), .C0(n1306), 
        .Y(n3466) );
  AOI22X1TS U1748 ( .A0(n1946), .A1(n651), .B0(n638), .B1(n1842), .Y(n1306) );
  OAI221XLTS U1749 ( .A0(n2291), .A1(n670), .B0(n2171), .B1(n660), .C0(n1307), 
        .Y(n3465) );
  AOI22X1TS U1750 ( .A0(n1947), .A1(n650), .B0(n641), .B1(n1843), .Y(n1307) );
  OAI221XLTS U1751 ( .A0(n2294), .A1(n670), .B0(n2174), .B1(n660), .C0(n1308), 
        .Y(n3464) );
  AOI22X1TS U1752 ( .A0(n1948), .A1(n650), .B0(n634), .B1(n1844), .Y(n1308) );
  OAI221XLTS U1753 ( .A0(n2297), .A1(n670), .B0(n2177), .B1(n660), .C0(n1309), 
        .Y(n3463) );
  AOI22X1TS U1754 ( .A0(n1949), .A1(n650), .B0(n634), .B1(n1845), .Y(n1309) );
  OAI221XLTS U1755 ( .A0(n2300), .A1(n670), .B0(n2180), .B1(n660), .C0(n1310), 
        .Y(n3462) );
  AOI22X1TS U1756 ( .A0(n1950), .A1(n650), .B0(n634), .B1(n1846), .Y(n1310) );
  OAI221XLTS U1757 ( .A0(n2303), .A1(n669), .B0(n2183), .B1(n659), .C0(n1311), 
        .Y(n3461) );
  AOI22X1TS U1758 ( .A0(n1951), .A1(n644), .B0(n634), .B1(n1847), .Y(n1311) );
  OAI221XLTS U1759 ( .A0(n2306), .A1(n669), .B0(n2186), .B1(n659), .C0(n1312), 
        .Y(n3460) );
  AOI22X1TS U1760 ( .A0(n1952), .A1(n644), .B0(n633), .B1(n1848), .Y(n1312) );
  OAI221XLTS U1761 ( .A0(n2309), .A1(n669), .B0(n2189), .B1(n659), .C0(n1313), 
        .Y(n3459) );
  AOI22X1TS U1762 ( .A0(n1953), .A1(n644), .B0(n633), .B1(n1849), .Y(n1313) );
  OAI221XLTS U1763 ( .A0(n2312), .A1(n669), .B0(n2192), .B1(n659), .C0(n1314), 
        .Y(n3458) );
  AOI22X1TS U1764 ( .A0(n1954), .A1(n644), .B0(n633), .B1(n1850), .Y(n1314) );
  OAI221XLTS U1765 ( .A0(n2315), .A1(n668), .B0(n2195), .B1(n658), .C0(n1315), 
        .Y(n3457) );
  AOI22X1TS U1766 ( .A0(n1955), .A1(n643), .B0(n633), .B1(n1851), .Y(n1315) );
  OAI221XLTS U1767 ( .A0(n2318), .A1(n668), .B0(n2198), .B1(n658), .C0(n1316), 
        .Y(n3456) );
  AOI22X1TS U1768 ( .A0(n1956), .A1(n643), .B0(n632), .B1(n1852), .Y(n1316) );
  OAI221XLTS U1769 ( .A0(n2321), .A1(n668), .B0(n2201), .B1(n658), .C0(n1317), 
        .Y(n3455) );
  AOI22X1TS U1770 ( .A0(n1957), .A1(n643), .B0(n632), .B1(n1853), .Y(n1317) );
  OAI221XLTS U1771 ( .A0(n2324), .A1(n668), .B0(n2204), .B1(n658), .C0(n1318), 
        .Y(n3454) );
  AOI22X1TS U1772 ( .A0(n1958), .A1(n643), .B0(n632), .B1(n1854), .Y(n1318) );
  OAI221XLTS U1773 ( .A0(n2327), .A1(n667), .B0(n2207), .B1(n657), .C0(n1319), 
        .Y(n3453) );
  AOI22X1TS U1774 ( .A0(n1959), .A1(n642), .B0(n632), .B1(n1855), .Y(n1319) );
  OAI221XLTS U1775 ( .A0(n2330), .A1(n667), .B0(n2210), .B1(n657), .C0(n1320), 
        .Y(n3452) );
  AOI22X1TS U1776 ( .A0(n1960), .A1(n642), .B0(n640), .B1(n1856), .Y(n1320) );
  OAI221XLTS U1777 ( .A0(n2333), .A1(n667), .B0(n2213), .B1(n657), .C0(n1321), 
        .Y(n3451) );
  AOI22X1TS U1778 ( .A0(n1961), .A1(n642), .B0(n1291), .B1(n1857), .Y(n1321)
         );
  OAI221XLTS U1779 ( .A0(n2336), .A1(n667), .B0(n2216), .B1(n657), .C0(n1322), 
        .Y(n3450) );
  AOI22X1TS U1780 ( .A0(n1962), .A1(n642), .B0(n639), .B1(n1858), .Y(n1322) );
  OAI221XLTS U1781 ( .A0(n1660), .A1(n82), .B0(n1283), .B1(n628), .C0(n1046), 
        .Y(n3607) );
  OAI221XLTS U1782 ( .A0(n1660), .A1(n83), .B0(n1283), .B1(n627), .C0(n1047), 
        .Y(n3606) );
  AOI22X1TS U1783 ( .A0(n915), .A1(n2251), .B0(n904), .B1(n2131), .Y(n1047) );
  OAI221XLTS U1784 ( .A0(n1589), .A1(n84), .B0(n1283), .B1(n626), .C0(n1048), 
        .Y(n3605) );
  AOI22X1TS U1785 ( .A0(n914), .A1(n2254), .B0(n903), .B1(n2134), .Y(n1048) );
  OAI221XLTS U1786 ( .A0(n1589), .A1(n85), .B0(n1283), .B1(n625), .C0(n1049), 
        .Y(n3604) );
  OAI221XLTS U1787 ( .A0(n1589), .A1(n86), .B0(n1188), .B1(n624), .C0(n1050), 
        .Y(n3603) );
  OAI221XLTS U1788 ( .A0(n1589), .A1(n87), .B0(n1188), .B1(n623), .C0(n1051), 
        .Y(n3602) );
  OAI221XLTS U1789 ( .A0(n2007), .A1(n88), .B0(n1188), .B1(n622), .C0(n1052), 
        .Y(n3601) );
  AOI22X1TS U1790 ( .A0(n913), .A1(n2266), .B0(n902), .B1(n2146), .Y(n1052) );
  OAI221XLTS U1791 ( .A0(n2008), .A1(n89), .B0(n1188), .B1(n621), .C0(n1053), 
        .Y(n3600) );
  OAI221XLTS U1792 ( .A0(n2007), .A1(n90), .B0(n1187), .B1(n620), .C0(n1054), 
        .Y(n3599) );
  OAI221XLTS U1793 ( .A0(n1717), .A1(n91), .B0(n1187), .B1(n619), .C0(n1055), 
        .Y(n3598) );
  OAI221XLTS U1794 ( .A0(n1518), .A1(n92), .B0(n1187), .B1(n618), .C0(n1056), 
        .Y(n3597) );
  AOI22X1TS U1795 ( .A0(n917), .A1(n2278), .B0(n901), .B1(n2158), .Y(n1056) );
  OAI221XLTS U1796 ( .A0(n1518), .A1(n93), .B0(n1187), .B1(n617), .C0(n1057), 
        .Y(n3596) );
  OAI221XLTS U1797 ( .A0(n1518), .A1(n94), .B0(n1006), .B1(n616), .C0(n1058), 
        .Y(n3595) );
  OAI221XLTS U1798 ( .A0(n1518), .A1(n95), .B0(n1006), .B1(n615), .C0(n1059), 
        .Y(n3594) );
  OAI221XLTS U1799 ( .A0(n1515), .A1(n96), .B0(n1006), .B1(n614), .C0(n1060), 
        .Y(n3593) );
  AOI22X1TS U1800 ( .A0(n912), .A1(n2290), .B0(n900), .B1(n2170), .Y(n1060) );
  OAI221XLTS U1801 ( .A0(n1515), .A1(n97), .B0(n1006), .B1(n613), .C0(n1061), 
        .Y(n3592) );
  OAI221XLTS U1802 ( .A0(n1515), .A1(n98), .B0(n1002), .B1(n612), .C0(n1062), 
        .Y(n3591) );
  OAI221XLTS U1803 ( .A0(n1515), .A1(n99), .B0(n1002), .B1(n611), .C0(n1063), 
        .Y(n3590) );
  OAI221XLTS U1804 ( .A0(n1505), .A1(n100), .B0(n1002), .B1(n610), .C0(n1064), 
        .Y(n3589) );
  AOI22X1TS U1805 ( .A0(n911), .A1(n2302), .B0(n907), .B1(n2182), .Y(n1064) );
  OAI221XLTS U1806 ( .A0(n1505), .A1(n101), .B0(n1002), .B1(n609), .C0(n1065), 
        .Y(n3588) );
  OAI221XLTS U1807 ( .A0(n1505), .A1(n102), .B0(n995), .B1(n608), .C0(n1066), 
        .Y(n3587) );
  OAI221XLTS U1808 ( .A0(n1505), .A1(n103), .B0(n995), .B1(n607), .C0(n1067), 
        .Y(n3586) );
  OAI221XLTS U1809 ( .A0(n1502), .A1(n104), .B0(n995), .B1(n606), .C0(n1068), 
        .Y(n3585) );
  AOI22X1TS U1810 ( .A0(n909), .A1(n2314), .B0(n899), .B1(n2194), .Y(n1068) );
  OAI221XLTS U1811 ( .A0(n1502), .A1(n105), .B0(n995), .B1(n605), .C0(n1069), 
        .Y(n3584) );
  OAI221XLTS U1812 ( .A0(n1502), .A1(n106), .B0(n993), .B1(n604), .C0(n1070), 
        .Y(n3583) );
  OAI221XLTS U1813 ( .A0(n1502), .A1(n107), .B0(n993), .B1(n603), .C0(n1071), 
        .Y(n3582) );
  OAI221XLTS U1814 ( .A0(n1492), .A1(n108), .B0(n993), .B1(n602), .C0(n1104), 
        .Y(n3581) );
  OAI221XLTS U1815 ( .A0(n1492), .A1(n109), .B0(n993), .B1(n601), .C0(n1105), 
        .Y(n3580) );
  OAI221XLTS U1816 ( .A0(n1492), .A1(n110), .B0(n1472), .B1(n600), .C0(n1106), 
        .Y(n3579) );
  OAI221XLTS U1817 ( .A0(n1492), .A1(n111), .B0(n1325), .B1(n599), .C0(n1107), 
        .Y(n3578) );
  AOI22X1TS U1818 ( .A0(n908), .A1(n2335), .B0(n898), .B1(n2215), .Y(n1107) );
  AOI21X1TS U1819 ( .A0(n115), .A1(n996), .B0(n1000), .Y(n991) );
  OA21XLTS U1820 ( .A0(n996), .A1(n114), .B0(n910), .Y(n1000) );
  OAI22X1TS U1821 ( .A0(n1226), .A1(n855), .B0(n1476), .B1(n326), .Y(n3325) );
  AOI222XLTS U1822 ( .A0(n1859), .A1(n182), .B0(n152), .B1(n2345), .C0(n2224), 
        .C1(n167), .Y(n1476) );
  OAI22X1TS U1823 ( .A0(n1225), .A1(n854), .B0(n1479), .B1(n326), .Y(n3324) );
  AOI222XLTS U1824 ( .A0(n1861), .A1(n183), .B0(n153), .B1(n2347), .C0(n2226), 
        .C1(n168), .Y(n1479) );
  OAI22X1TS U1825 ( .A0(n1224), .A1(n854), .B0(n1480), .B1(n326), .Y(n3323) );
  AOI222XLTS U1826 ( .A0(n1863), .A1(n10), .B0(n152), .B1(n2348), .C0(n2228), 
        .C1(n169), .Y(n1480) );
  OAI22X1TS U1827 ( .A0(n1223), .A1(n854), .B0(n1481), .B1(n326), .Y(n3322) );
  AOI222XLTS U1828 ( .A0(n1865), .A1(n181), .B0(n153), .B1(n2351), .C0(n2230), 
        .C1(n167), .Y(n1481) );
  OAI22X1TS U1829 ( .A0(n1222), .A1(n854), .B0(n1482), .B1(n327), .Y(n3321) );
  AOI222XLTS U1830 ( .A0(n1867), .A1(n182), .B0(n152), .B1(n2352), .C0(n2233), 
        .C1(n168), .Y(n1482) );
  OAI22X1TS U1831 ( .A0(n1221), .A1(n853), .B0(n1483), .B1(n327), .Y(n3320) );
  AOI222XLTS U1832 ( .A0(n1869), .A1(n183), .B0(n153), .B1(n2355), .C0(n2235), 
        .C1(n169), .Y(n1483) );
  OAI22X1TS U1833 ( .A0(n1220), .A1(n853), .B0(n1484), .B1(n327), .Y(n3319) );
  AOI222XLTS U1834 ( .A0(n1871), .A1(n10), .B0(n152), .B1(n2357), .C0(n2238), 
        .C1(n167), .Y(n1484) );
  OAI22X1TS U1835 ( .A0(n1219), .A1(n853), .B0(n1485), .B1(n327), .Y(n3318) );
  AOI222XLTS U1836 ( .A0(n1873), .A1(n181), .B0(n153), .B1(n2360), .C0(n2241), 
        .C1(n168), .Y(n1485) );
  OAI22X1TS U1837 ( .A0(n48), .A1(n158), .B0(n1503), .B1(n324), .Y(n3309) );
  AOI222XLTS U1838 ( .A0(n1860), .A1(n178), .B0(n150), .B1(n2345), .C0(
        cacheAddressIn_WEST[0]), .C1(n160), .Y(n1503) );
  OAI22X1TS U1839 ( .A0(n49), .A1(n288), .B0(n1528), .B1(n1529), .Y(n3293) );
  AOI222XLTS U1840 ( .A0(n332), .A1(n782), .B0(n268), .B1(
        cacheAddressIn_EAST[0]), .C0(n2225), .C1(n794), .Y(n1528) );
  OAI22X1TS U1841 ( .A0(n50), .A1(n159), .B0(n1506), .B1(n324), .Y(n3308) );
  AOI222XLTS U1842 ( .A0(n1862), .A1(n179), .B0(n151), .B1(n2347), .C0(
        cacheAddressIn_WEST[1]), .C1(n161), .Y(n1506) );
  OAI22X1TS U1843 ( .A0(n51), .A1(n287), .B0(n1531), .B1(n260), .Y(n3292) );
  AOI222XLTS U1844 ( .A0(n332), .A1(n781), .B0(n267), .B1(
        cacheAddressIn_EAST[1]), .C0(n2227), .C1(n303), .Y(n1531) );
  OAI22X1TS U1845 ( .A0(n52), .A1(n157), .B0(n1507), .B1(n324), .Y(n3307) );
  AOI222XLTS U1846 ( .A0(n1864), .A1(n801), .B0(n150), .B1(
        cacheAddressIn_EAST[2]), .C0(cacheAddressIn_WEST[2]), .C1(n162), .Y(
        n1507) );
  OAI22X1TS U1847 ( .A0(n53), .A1(n288), .B0(n1532), .B1(n1529), .Y(n3291) );
  AOI222XLTS U1848 ( .A0(n333), .A1(n780), .B0(n267), .B1(n2349), .C0(n2229), 
        .C1(n303), .Y(n1532) );
  OAI22X1TS U1849 ( .A0(n54), .A1(n158), .B0(n1508), .B1(n324), .Y(n3306) );
  AOI222XLTS U1850 ( .A0(n1866), .A1(n177), .B0(n150), .B1(n2351), .C0(
        cacheAddressIn_WEST[3]), .C1(n160), .Y(n1508) );
  OAI22X1TS U1851 ( .A0(n55), .A1(n287), .B0(n1533), .B1(n260), .Y(n3290) );
  AOI222XLTS U1852 ( .A0(n331), .A1(n779), .B0(n267), .B1(
        cacheAddressIn_EAST[3]), .C0(n2231), .C1(n303), .Y(n1533) );
  OAI22X1TS U1853 ( .A0(n56), .A1(n159), .B0(n1509), .B1(n325), .Y(n3305) );
  AOI222XLTS U1854 ( .A0(n1868), .A1(n178), .B0(n151), .B1(
        cacheAddressIn_EAST[4]), .C0(n2233), .C1(n161), .Y(n1509) );
  OAI22X1TS U1855 ( .A0(n57), .A1(n288), .B0(n1534), .B1(n1529), .Y(n3289) );
  AOI222XLTS U1856 ( .A0(n333), .A1(n778), .B0(n267), .B1(n2353), .C0(
        cacheAddressIn_WEST[4]), .C1(n304), .Y(n1534) );
  OAI22X1TS U1857 ( .A0(n58), .A1(n157), .B0(n1510), .B1(n325), .Y(n3304) );
  AOI222XLTS U1858 ( .A0(n1870), .A1(n179), .B0(n151), .B1(n2355), .C0(n2235), 
        .C1(n162), .Y(n1510) );
  OAI22X1TS U1859 ( .A0(n59), .A1(n287), .B0(n1535), .B1(n260), .Y(n3288) );
  AOI222XLTS U1860 ( .A0(n331), .A1(n777), .B0(n268), .B1(
        cacheAddressIn_EAST[5]), .C0(cacheAddressIn_WEST[5]), .C1(n304), .Y(
        n1535) );
  OAI22X1TS U1861 ( .A0(n60), .A1(n158), .B0(n1511), .B1(n325), .Y(n3303) );
  AOI222XLTS U1862 ( .A0(n1872), .A1(n801), .B0(n150), .B1(n2357), .C0(n2238), 
        .C1(n160), .Y(n1511) );
  OAI22X1TS U1863 ( .A0(n61), .A1(n288), .B0(n1536), .B1(n1529), .Y(n3287) );
  AOI222XLTS U1864 ( .A0(n333), .A1(n776), .B0(n268), .B1(n2358), .C0(n2237), 
        .C1(n304), .Y(n1536) );
  OAI22X1TS U1865 ( .A0(n62), .A1(n159), .B0(n1512), .B1(n325), .Y(n3302) );
  AOI222XLTS U1866 ( .A0(n1874), .A1(n177), .B0(n151), .B1(n2360), .C0(n2241), 
        .C1(n161), .Y(n1512) );
  OAI22X1TS U1867 ( .A0(n63), .A1(n287), .B0(n1537), .B1(n260), .Y(n3286) );
  AOI222XLTS U1868 ( .A0(n331), .A1(n775), .B0(n268), .B1(n2361), .C0(n2240), 
        .C1(n304), .Y(n1537) );
  OAI22X1TS U1869 ( .A0(n64), .A1(n155), .B0(n1516), .B1(n322), .Y(n3301) );
  AOI222XLTS U1870 ( .A0(n1923), .A1(n186), .B0(n148), .B1(n2344), .C0(n2225), 
        .C1(n163), .Y(n1516) );
  OAI22X1TS U1871 ( .A0(n65), .A1(n156), .B0(n1519), .B1(n322), .Y(n3300) );
  AOI222XLTS U1872 ( .A0(n1924), .A1(n187), .B0(n149), .B1(n2346), .C0(n2227), 
        .C1(n164), .Y(n1519) );
  OAI22X1TS U1873 ( .A0(n66), .A1(n154), .B0(n1520), .B1(n322), .Y(n3299) );
  AOI222XLTS U1874 ( .A0(n1925), .A1(n184), .B0(n148), .B1(n2349), .C0(n2229), 
        .C1(n165), .Y(n1520) );
  OAI22X1TS U1875 ( .A0(n67), .A1(n155), .B0(n1521), .B1(n322), .Y(n3298) );
  AOI222XLTS U1876 ( .A0(n1926), .A1(n185), .B0(n148), .B1(n2350), .C0(n2231), 
        .C1(n163), .Y(n1521) );
  OAI22X1TS U1877 ( .A0(n68), .A1(n156), .B0(n1522), .B1(n323), .Y(n3297) );
  AOI222XLTS U1878 ( .A0(n1927), .A1(n186), .B0(n149), .B1(n2353), .C0(n2232), 
        .C1(n164), .Y(n1522) );
  OAI22X1TS U1879 ( .A0(n69), .A1(n154), .B0(n1523), .B1(n323), .Y(n3296) );
  AOI222XLTS U1880 ( .A0(n1928), .A1(n187), .B0(n149), .B1(n2354), .C0(n2234), 
        .C1(n165), .Y(n1523) );
  OAI22X1TS U1881 ( .A0(n70), .A1(n155), .B0(n1524), .B1(n323), .Y(n3295) );
  AOI222XLTS U1882 ( .A0(n1929), .A1(n184), .B0(n148), .B1(n2358), .C0(n2237), 
        .C1(n163), .Y(n1524) );
  OAI22X1TS U1883 ( .A0(n71), .A1(n156), .B0(n1525), .B1(n323), .Y(n3294) );
  AOI222XLTS U1884 ( .A0(n1930), .A1(n185), .B0(n149), .B1(n2361), .C0(n2240), 
        .C1(n164), .Y(n1525) );
  AOI222XLTS U1885 ( .A0(n1875), .A1(n136), .B0(n2344), .B1(n285), .C0(n2224), 
        .C1(n270), .Y(n1463) );
  OAI22X1TS U1886 ( .A0(n1324), .A1(n37), .B0(n1465), .B1(n1464), .Y(n3332) );
  AOI222XLTS U1887 ( .A0(n1876), .A1(n136), .B0(n2346), .B1(n285), .C0(n2226), 
        .C1(n270), .Y(n1465) );
  OAI22X1TS U1888 ( .A0(n1324), .A1(n38), .B0(n1466), .B1(n1464), .Y(n3331) );
  AOI222XLTS U1889 ( .A0(n1877), .A1(n310), .B0(n2349), .B1(n286), .C0(n2228), 
        .C1(n271), .Y(n1466) );
  OAI22X1TS U1890 ( .A0(n1478), .A1(n39), .B0(n1467), .B1(n1464), .Y(n3330) );
  AOI222XLTS U1891 ( .A0(n1878), .A1(n309), .B0(n2350), .B1(n285), .C0(n2230), 
        .C1(n270), .Y(n1467) );
  OAI22X1TS U1892 ( .A0(n1472), .A1(n40), .B0(n1468), .B1(n1464), .Y(n3329) );
  AOI222XLTS U1893 ( .A0(n1879), .A1(n308), .B0(n2353), .B1(n286), .C0(n2233), 
        .C1(n271), .Y(n1468) );
  OAI22X1TS U1894 ( .A0(n1325), .A1(n41), .B0(n1469), .B1(n321), .Y(n3328) );
  AOI222XLTS U1895 ( .A0(n1880), .A1(n308), .B0(n2354), .B1(n286), .C0(n2235), 
        .C1(n271), .Y(n1469) );
  OAI22X1TS U1896 ( .A0(n1374), .A1(n42), .B0(n1470), .B1(n321), .Y(n3327) );
  AOI222XLTS U1897 ( .A0(n1881), .A1(n310), .B0(n2358), .B1(n285), .C0(n2238), 
        .C1(n270), .Y(n1470) );
  OAI22X1TS U1898 ( .A0(n1041), .A1(n43), .B0(n1471), .B1(n321), .Y(n3326) );
  AOI222XLTS U1899 ( .A0(n1882), .A1(n309), .B0(n2361), .B1(n286), .C0(n2241), 
        .C1(n271), .Y(n1471) );
  NAND2X1TS U1900 ( .A(n1676), .B(n880), .Y(n1501) );
  NOR2X1TS U1901 ( .A(n1501), .B(n910), .Y(n1487) );
  OAI32X1TS U1902 ( .A0(n1430), .A1(n2369), .A2(n811), .B0(n1431), .B1(n45), 
        .Y(n3343) );
  INVX2TS U1903 ( .A(n1431), .Y(n811) );
  NAND3BX1TS U1904 ( .AN(n1432), .B(n1433), .C(n1434), .Y(n1431) );
  OAI21X1TS U1905 ( .A0(n1437), .A1(n1441), .B0(n844), .Y(n1438) );
  INVX2TS U1906 ( .A(n1435), .Y(n821) );
  OAI221XLTS U1907 ( .A0(n1082), .A1(n2077), .B0(n1146), .B1(n2071), .C0(n1027), .Y(n3620) );
  AOI22X1TS U1908 ( .A0(n2305), .A1(n2033), .B0(n2185), .B1(n2011), .Y(n1027)
         );
  OAI221XLTS U1909 ( .A0(n1081), .A1(n2077), .B0(n1145), .B1(n2059), .C0(n1028), .Y(n3619) );
  OAI221XLTS U1910 ( .A0(n1080), .A1(n2077), .B0(n1144), .B1(n2051), .C0(n1029), .Y(n3618) );
  OAI221XLTS U1911 ( .A0(n1079), .A1(n2075), .B0(n1143), .B1(n2051), .C0(n1030), .Y(n3617) );
  AOI22X1TS U1912 ( .A0(n2314), .A1(n2031), .B0(n2194), .B1(n2010), .Y(n1030)
         );
  OAI221XLTS U1913 ( .A0(n1078), .A1(n2075), .B0(n1142), .B1(n2051), .C0(n1031), .Y(n3616) );
  OAI221XLTS U1914 ( .A0(n1077), .A1(n2075), .B0(n1141), .B1(n2051), .C0(n1032), .Y(n3615) );
  OAI221XLTS U1915 ( .A0(n1076), .A1(n2075), .B0(n1140), .B1(n2049), .C0(n1033), .Y(n3614) );
  OAI221XLTS U1916 ( .A0(n1075), .A1(n2073), .B0(n1139), .B1(n2049), .C0(n1034), .Y(n3613) );
  OAI221XLTS U1917 ( .A0(n1074), .A1(n2073), .B0(n1138), .B1(n2049), .C0(n1035), .Y(n3612) );
  OAI221XLTS U1918 ( .A0(n1073), .A1(n2073), .B0(n1137), .B1(n2049), .C0(n1036), .Y(n3611) );
  OAI221XLTS U1919 ( .A0(n1072), .A1(n2073), .B0(n1136), .B1(n2061), .C0(n1037), .Y(n3610) );
  AOI22X1TS U1920 ( .A0(n2335), .A1(n2029), .B0(n2215), .B1(n2009), .Y(n1037)
         );
  OAI221XLTS U1921 ( .A0(n1103), .A1(n2087), .B0(n1167), .B1(n2059), .C0(n1004), .Y(n3641) );
  AOI22X1TS U1922 ( .A0(n2242), .A1(n2043), .B0(n2122), .B1(n2019), .Y(n1004)
         );
  OAI221XLTS U1923 ( .A0(n1102), .A1(n2087), .B0(n1166), .B1(n2059), .C0(n1007), .Y(n3640) );
  OAI221XLTS U1924 ( .A0(n1101), .A1(n2087), .B0(n1165), .B1(n2059), .C0(n1008), .Y(n3639) );
  OAI221XLTS U1925 ( .A0(n1100), .A1(n2087), .B0(n1164), .B1(n2057), .C0(n1009), .Y(n3638) );
  OAI221XLTS U1926 ( .A0(n1099), .A1(n2085), .B0(n1163), .B1(n2057), .C0(n1010), .Y(n3637) );
  AOI22X1TS U1927 ( .A0(n2254), .A1(n2041), .B0(n2134), .B1(n2017), .Y(n1010)
         );
  OAI221XLTS U1928 ( .A0(n1098), .A1(n2085), .B0(n1162), .B1(n2057), .C0(n1011), .Y(n3636) );
  OAI221XLTS U1929 ( .A0(n1097), .A1(n2085), .B0(n1161), .B1(n2057), .C0(n1012), .Y(n3635) );
  OAI221XLTS U1930 ( .A0(n1096), .A1(n2085), .B0(n1160), .B1(n2055), .C0(n1013), .Y(n3634) );
  OAI221XLTS U1931 ( .A0(n1095), .A1(n2083), .B0(n1159), .B1(n2055), .C0(n1014), .Y(n3633) );
  AOI22X1TS U1932 ( .A0(n2266), .A1(n2039), .B0(n2146), .B1(n2015), .Y(n1014)
         );
  OAI221XLTS U1933 ( .A0(n1094), .A1(n2083), .B0(n1158), .B1(n2055), .C0(n1015), .Y(n3632) );
  OAI221XLTS U1934 ( .A0(n1093), .A1(n2083), .B0(n1157), .B1(n2055), .C0(n1016), .Y(n3631) );
  OAI221XLTS U1935 ( .A0(n1092), .A1(n2083), .B0(n1156), .B1(n2053), .C0(n1017), .Y(n3630) );
  OAI221XLTS U1936 ( .A0(n1091), .A1(n2081), .B0(n1155), .B1(n2053), .C0(n1018), .Y(n3629) );
  AOI22X1TS U1937 ( .A0(n2278), .A1(n2037), .B0(n2158), .B1(n2013), .Y(n1018)
         );
  OAI221XLTS U1938 ( .A0(n1090), .A1(n2081), .B0(n1154), .B1(n2053), .C0(n1019), .Y(n3628) );
  OAI221XLTS U1939 ( .A0(n1089), .A1(n2081), .B0(n1153), .B1(n2053), .C0(n1020), .Y(n3627) );
  OAI221XLTS U1940 ( .A0(n1088), .A1(n2081), .B0(n1152), .B1(n2065), .C0(n1021), .Y(n3626) );
  OAI221XLTS U1941 ( .A0(n1087), .A1(n2079), .B0(n1151), .B1(n2067), .C0(n1022), .Y(n3625) );
  AOI22X1TS U1942 ( .A0(n2290), .A1(n2035), .B0(n2170), .B1(n2012), .Y(n1022)
         );
  OAI221XLTS U1943 ( .A0(n1086), .A1(n2079), .B0(n1150), .B1(n2065), .C0(n1023), .Y(n3624) );
  OAI221XLTS U1944 ( .A0(n1085), .A1(n2079), .B0(n1149), .B1(n2065), .C0(n1024), .Y(n3623) );
  OAI221XLTS U1945 ( .A0(n1084), .A1(n2079), .B0(n1148), .B1(n2063), .C0(n1025), .Y(n3622) );
  OAI221XLTS U1946 ( .A0(n1083), .A1(n2077), .B0(n1147), .B1(n2065), .C0(n1026), .Y(n3621) );
  OAI221XLTS U1947 ( .A0(n2014), .A1(n2094), .B0(n490), .B1(n44), .C0(n1674), 
        .Y(n3209) );
  AOI222XLTS U1948 ( .A0(n2225), .A1(n539), .B0(cacheAddressIn_EAST[0]), .B1(
        n528), .C0(cacheAddressIn_SOUTH[0]), .C1(n505), .Y(n1674) );
  OAI221XLTS U1949 ( .A0(n2016), .A1(n2103), .B0(n488), .B1(n37), .C0(n1673), 
        .Y(n3210) );
  AOI222XLTS U1950 ( .A0(n2227), .A1(n539), .B0(cacheAddressIn_EAST[1]), .B1(
        n525), .C0(cacheAddressIn_SOUTH[1]), .C1(n505), .Y(n1673) );
  OAI221XLTS U1951 ( .A0(n2018), .A1(n2103), .B0(n488), .B1(n38), .C0(n1672), 
        .Y(n3211) );
  AOI222XLTS U1952 ( .A0(n2229), .A1(n538), .B0(cacheAddressIn_EAST[2]), .B1(
        n528), .C0(cacheAddressIn_SOUTH[2]), .C1(n505), .Y(n1672) );
  OAI221XLTS U1953 ( .A0(n2020), .A1(n2103), .B0(n488), .B1(n39), .C0(n1671), 
        .Y(n3212) );
  AOI222XLTS U1954 ( .A0(n2231), .A1(n538), .B0(cacheAddressIn_EAST[3]), .B1(
        n528), .C0(cacheAddressIn_SOUTH[3]), .C1(n505), .Y(n1671) );
  OAI221XLTS U1955 ( .A0(n2022), .A1(n2106), .B0(n489), .B1(n40), .C0(n1670), 
        .Y(n3213) );
  AOI222XLTS U1956 ( .A0(n2232), .A1(n536), .B0(cacheAddressIn_EAST[4]), .B1(
        n517), .C0(cacheAddressIn_SOUTH[4]), .C1(n510), .Y(n1670) );
  OAI221XLTS U1957 ( .A0(n2024), .A1(n2108), .B0(n489), .B1(n41), .C0(n1669), 
        .Y(n3214) );
  AOI222XLTS U1958 ( .A0(n2234), .A1(n536), .B0(cacheAddressIn_EAST[5]), .B1(
        n517), .C0(cacheAddressIn_SOUTH[5]), .C1(n514), .Y(n1669) );
  OAI221XLTS U1959 ( .A0(n2026), .A1(n2104), .B0(n490), .B1(n42), .C0(n1668), 
        .Y(n3215) );
  AOI222XLTS U1960 ( .A0(n2237), .A1(n536), .B0(cacheAddressIn_EAST[6]), .B1(
        n517), .C0(cacheAddressIn_SOUTH[6]), .C1(n514), .Y(n1668) );
  OAI221XLTS U1961 ( .A0(n2028), .A1(n2104), .B0(n489), .B1(n43), .C0(n1667), 
        .Y(n3216) );
  AOI222XLTS U1962 ( .A0(n2240), .A1(n536), .B0(cacheAddressIn_EAST[7]), .B1(
        n517), .C0(cacheAddressIn_SOUTH[7]), .C1(n516), .Y(n1667) );
  OAI221XLTS U1963 ( .A0(n2030), .A1(n2108), .B0(n630), .B1(n491), .C0(n1417), 
        .Y(n3346) );
  AOI222XLTS U1964 ( .A0(n535), .A1(n2122), .B0(n518), .B1(n2242), .C0(
        dataIn_SOUTH[0]), .C1(n513), .Y(n1417) );
  OAI221XLTS U1965 ( .A0(n2032), .A1(n2107), .B0(n629), .B1(n491), .C0(n1416), 
        .Y(n3347) );
  AOI222XLTS U1966 ( .A0(n535), .A1(n2125), .B0(n518), .B1(n2245), .C0(
        dataIn_SOUTH[1]), .C1(n513), .Y(n1416) );
  OAI221XLTS U1967 ( .A0(n2034), .A1(n2107), .B0(n628), .B1(n492), .C0(n1415), 
        .Y(n3348) );
  AOI222XLTS U1968 ( .A0(n535), .A1(n2128), .B0(n518), .B1(n2248), .C0(
        dataIn_SOUTH[2]), .C1(n514), .Y(n1415) );
  OAI221XLTS U1969 ( .A0(n2036), .A1(n2106), .B0(n627), .B1(n493), .C0(n1414), 
        .Y(n3349) );
  AOI222XLTS U1970 ( .A0(n535), .A1(n2131), .B0(n518), .B1(n2251), .C0(
        dataIn_SOUTH[3]), .C1(n511), .Y(n1414) );
  OAI221XLTS U1971 ( .A0(n2038), .A1(n2104), .B0(n626), .B1(n493), .C0(n1413), 
        .Y(n3350) );
  AOI222XLTS U1972 ( .A0(n534), .A1(n2134), .B0(n519), .B1(n2254), .C0(
        dataIn_SOUTH[4]), .C1(n513), .Y(n1413) );
  OAI221XLTS U1973 ( .A0(n2040), .A1(n2103), .B0(n625), .B1(n494), .C0(n1412), 
        .Y(n3351) );
  AOI222XLTS U1974 ( .A0(n534), .A1(n2137), .B0(n519), .B1(n2257), .C0(
        dataIn_SOUTH[5]), .C1(n513), .Y(n1412) );
  OAI221XLTS U1975 ( .A0(n2042), .A1(n2105), .B0(n624), .B1(n494), .C0(n1411), 
        .Y(n3352) );
  AOI222XLTS U1976 ( .A0(n534), .A1(n2140), .B0(n519), .B1(n2260), .C0(
        dataIn_SOUTH[6]), .C1(n1386), .Y(n1411) );
  OAI221XLTS U1977 ( .A0(n2044), .A1(n2105), .B0(n623), .B1(n494), .C0(n1410), 
        .Y(n3353) );
  AOI222XLTS U1978 ( .A0(n534), .A1(n2143), .B0(n519), .B1(n2263), .C0(
        dataIn_SOUTH[7]), .C1(n1386), .Y(n1410) );
  OAI221XLTS U1979 ( .A0(n2046), .A1(n2104), .B0(n622), .B1(n492), .C0(n1409), 
        .Y(n3354) );
  AOI222XLTS U1980 ( .A0(n537), .A1(n2146), .B0(n520), .B1(n2266), .C0(
        dataIn_SOUTH[8]), .C1(n512), .Y(n1409) );
  OAI221XLTS U1981 ( .A0(n2048), .A1(n2110), .B0(n621), .B1(n492), .C0(n1408), 
        .Y(n3355) );
  AOI222XLTS U1982 ( .A0(n1384), .A1(n2149), .B0(n520), .B1(n2269), .C0(
        dataIn_SOUTH[9]), .C1(n512), .Y(n1408) );
  OAI221XLTS U1983 ( .A0(n2050), .A1(n2105), .B0(n620), .B1(n493), .C0(n1407), 
        .Y(n3356) );
  AOI222XLTS U1984 ( .A0(n540), .A1(n2152), .B0(n520), .B1(n2272), .C0(
        dataIn_SOUTH[10]), .C1(n512), .Y(n1407) );
  OAI221XLTS U1985 ( .A0(n2052), .A1(n2108), .B0(n619), .B1(n501), .C0(n1406), 
        .Y(n3357) );
  AOI222XLTS U1986 ( .A0(n537), .A1(n2155), .B0(n520), .B1(n2275), .C0(
        dataIn_SOUTH[11]), .C1(n515), .Y(n1406) );
  OAI221XLTS U1987 ( .A0(n2054), .A1(n2105), .B0(n618), .B1(n503), .C0(n1405), 
        .Y(n3358) );
  AOI222XLTS U1988 ( .A0(n533), .A1(n2158), .B0(n521), .B1(n2278), .C0(
        dataIn_SOUTH[12]), .C1(n511), .Y(n1405) );
  OAI221XLTS U1989 ( .A0(n2056), .A1(n2102), .B0(n617), .B1(n496), .C0(n1404), 
        .Y(n3359) );
  AOI222XLTS U1990 ( .A0(n533), .A1(n2161), .B0(n521), .B1(n2281), .C0(
        dataIn_SOUTH[13]), .C1(n510), .Y(n1404) );
  OAI221XLTS U1991 ( .A0(n2058), .A1(n2102), .B0(n616), .B1(n496), .C0(n1403), 
        .Y(n3360) );
  AOI222XLTS U1992 ( .A0(n533), .A1(n2164), .B0(n521), .B1(n2284), .C0(
        dataIn_SOUTH[14]), .C1(n516), .Y(n1403) );
  OAI221XLTS U1993 ( .A0(n2060), .A1(n2102), .B0(n615), .B1(n495), .C0(n1402), 
        .Y(n3361) );
  AOI222XLTS U1994 ( .A0(n533), .A1(n2167), .B0(n521), .B1(n2287), .C0(
        dataIn_SOUTH[15]), .C1(n512), .Y(n1402) );
  OAI221XLTS U1995 ( .A0(n2062), .A1(n2102), .B0(n614), .B1(n495), .C0(n1401), 
        .Y(n3362) );
  AOI222XLTS U1996 ( .A0(n532), .A1(n2170), .B0(n527), .B1(n2290), .C0(
        dataIn_SOUTH[16]), .C1(n506), .Y(n1401) );
  OAI221XLTS U1997 ( .A0(n2064), .A1(n2101), .B0(n613), .B1(n495), .C0(n1400), 
        .Y(n3363) );
  AOI222XLTS U1998 ( .A0(n532), .A1(n2173), .B0(n526), .B1(n2293), .C0(
        dataIn_SOUTH[17]), .C1(n506), .Y(n1400) );
  OAI221XLTS U1999 ( .A0(n2066), .A1(n2101), .B0(n612), .B1(n503), .C0(n1399), 
        .Y(n3364) );
  AOI222XLTS U2000 ( .A0(n532), .A1(n2176), .B0(n527), .B1(n2296), .C0(
        dataIn_SOUTH[18]), .C1(n506), .Y(n1399) );
  OAI221XLTS U2001 ( .A0(n2068), .A1(n2101), .B0(n611), .B1(n498), .C0(n1398), 
        .Y(n3365) );
  AOI222XLTS U2002 ( .A0(n532), .A1(n2179), .B0(n526), .B1(n2299), .C0(
        dataIn_SOUTH[19]), .C1(n506), .Y(n1398) );
  OAI221XLTS U2003 ( .A0(n2070), .A1(n2101), .B0(n610), .B1(n498), .C0(n1397), 
        .Y(n3366) );
  AOI222XLTS U2004 ( .A0(n531), .A1(n2182), .B0(n522), .B1(n2302), .C0(
        dataIn_SOUTH[20]), .C1(n507), .Y(n1397) );
  OAI221XLTS U2005 ( .A0(n2072), .A1(n2099), .B0(n609), .B1(n498), .C0(n1396), 
        .Y(n3367) );
  AOI222XLTS U2006 ( .A0(n531), .A1(n2185), .B0(n522), .B1(n2305), .C0(
        dataIn_SOUTH[21]), .C1(n507), .Y(n1396) );
  OAI221XLTS U2007 ( .A0(n2074), .A1(n2099), .B0(n608), .B1(n498), .C0(n1395), 
        .Y(n3368) );
  AOI222XLTS U2008 ( .A0(n531), .A1(n2188), .B0(n522), .B1(n2308), .C0(
        dataIn_SOUTH[22]), .C1(n507), .Y(n1395) );
  OAI221XLTS U2009 ( .A0(n2076), .A1(n2099), .B0(n607), .B1(n496), .C0(n1394), 
        .Y(n3369) );
  AOI222XLTS U2010 ( .A0(n531), .A1(n2191), .B0(n522), .B1(n2311), .C0(
        dataIn_SOUTH[23]), .C1(n507), .Y(n1394) );
  OAI221XLTS U2011 ( .A0(n2078), .A1(n2094), .B0(n606), .B1(n497), .C0(n1393), 
        .Y(n3370) );
  AOI222XLTS U2012 ( .A0(n530), .A1(n2194), .B0(n523), .B1(n2314), .C0(
        dataIn_SOUTH[24]), .C1(n508), .Y(n1393) );
  OAI221XLTS U2013 ( .A0(n2080), .A1(n2094), .B0(n605), .B1(n497), .C0(n1392), 
        .Y(n3371) );
  AOI222XLTS U2014 ( .A0(n530), .A1(n2197), .B0(n523), .B1(n2317), .C0(
        dataIn_SOUTH[25]), .C1(n508), .Y(n1392) );
  OAI221XLTS U2015 ( .A0(n2082), .A1(n2094), .B0(n604), .B1(n497), .C0(n1391), 
        .Y(n3372) );
  AOI222XLTS U2016 ( .A0(n530), .A1(n2200), .B0(n523), .B1(n2320), .C0(
        dataIn_SOUTH[26]), .C1(n508), .Y(n1391) );
  OAI221XLTS U2017 ( .A0(n2084), .A1(n2099), .B0(n603), .B1(n499), .C0(n1390), 
        .Y(n3373) );
  AOI222XLTS U2018 ( .A0(n530), .A1(n2203), .B0(n523), .B1(n2323), .C0(
        dataIn_SOUTH[27]), .C1(n508), .Y(n1390) );
  OAI221XLTS U2019 ( .A0(n2086), .A1(n2093), .B0(n602), .B1(n499), .C0(n1389), 
        .Y(n3374) );
  AOI222XLTS U2020 ( .A0(n529), .A1(n2206), .B0(n524), .B1(n2326), .C0(
        dataIn_SOUTH[28]), .C1(n509), .Y(n1389) );
  OAI221XLTS U2021 ( .A0(n2088), .A1(n2093), .B0(n601), .B1(n499), .C0(n1388), 
        .Y(n3375) );
  AOI222XLTS U2022 ( .A0(n529), .A1(n2209), .B0(n524), .B1(n2329), .C0(
        dataIn_SOUTH[29]), .C1(n509), .Y(n1388) );
  OAI221XLTS U2023 ( .A0(n2090), .A1(n2093), .B0(n600), .B1(n491), .C0(n1387), 
        .Y(n3376) );
  AOI222XLTS U2024 ( .A0(n529), .A1(n2212), .B0(n524), .B1(n2332), .C0(
        dataIn_SOUTH[30]), .C1(n509), .Y(n1387) );
  OAI221XLTS U2025 ( .A0(n2092), .A1(n2109), .B0(n599), .B1(n499), .C0(n1383), 
        .Y(n3377) );
  AOI222XLTS U2026 ( .A0(n529), .A1(n2215), .B0(n524), .B1(n2335), .C0(
        dataIn_SOUTH[31]), .C1(n509), .Y(n1383) );
  OAI211X1TS U2027 ( .A0(n2338), .A1(n1694), .B0(n1695), .C0(n1696), .Y(n3190)
         );
  AOI22X1TS U2028 ( .A0(requesterAddressIn_NORTH[0]), .A1(n1697), .B0(n1698), 
        .B1(requesterAddressIn_SOUTH[0]), .Y(n1695) );
  AOI222XLTS U2029 ( .A0(prevRequesterAddress_A[0]), .A1(n273), .B0(
        \requesterAddressBuffer[0][0] ), .B1(n261), .C0(n143), .C1(
        requesterAddressIn_WEST[0]), .Y(n1696) );
  OAI211X1TS U2030 ( .A0(n2339), .A1(n1694), .B0(n1699), .C0(n1700), .Y(n3189)
         );
  AOI22X1TS U2031 ( .A0(requesterAddressIn_NORTH[1]), .A1(n1697), .B0(n1698), 
        .B1(requesterAddressIn_SOUTH[1]), .Y(n1699) );
  AOI222XLTS U2032 ( .A0(prevRequesterAddress_A[1]), .A1(n274), .B0(
        \requesterAddressBuffer[0][1] ), .B1(n261), .C0(n1595), .C1(
        requesterAddressIn_WEST[1]), .Y(n1700) );
  OAI211X1TS U2033 ( .A0(n2340), .A1(n1694), .B0(n1701), .C0(n1702), .Y(n3188)
         );
  AOI22X1TS U2034 ( .A0(requesterAddressIn_NORTH[2]), .A1(n1697), .B0(n1698), 
        .B1(requesterAddressIn_SOUTH[2]), .Y(n1701) );
  AOI222XLTS U2035 ( .A0(prevRequesterAddress_A[2]), .A1(n273), .B0(
        \requesterAddressBuffer[0][2] ), .B1(n261), .C0(n143), .C1(
        requesterAddressIn_WEST[2]), .Y(n1702) );
  OAI211X1TS U2036 ( .A0(n2341), .A1(n280), .B0(n1703), .C0(n1704), .Y(n3187)
         );
  AOI22X1TS U2037 ( .A0(requesterAddressIn_NORTH[3]), .A1(n297), .B0(n315), 
        .B1(requesterAddressIn_SOUTH[3]), .Y(n1703) );
  AOI222XLTS U2038 ( .A0(prevRequesterAddress_A[3]), .A1(n274), .B0(
        \requesterAddressBuffer[0][3] ), .B1(n261), .C0(n1595), .C1(
        requesterAddressIn_WEST[3]), .Y(n1704) );
  OAI211X1TS U2039 ( .A0(n2342), .A1(n280), .B0(n1705), .C0(n1706), .Y(n3186)
         );
  AOI22X1TS U2040 ( .A0(requesterAddressIn_NORTH[4]), .A1(n297), .B0(n315), 
        .B1(requesterAddressIn_SOUTH[4]), .Y(n1705) );
  AOI222XLTS U2041 ( .A0(prevRequesterAddress_A[4]), .A1(n273), .B0(
        \requesterAddressBuffer[0][4] ), .B1(n262), .C0(n143), .C1(
        requesterAddressIn_WEST[4]), .Y(n1706) );
  OAI211X1TS U2042 ( .A0(n2343), .A1(n280), .B0(n1707), .C0(n1708), .Y(n3185)
         );
  AOI22X1TS U2043 ( .A0(requesterAddressIn_NORTH[5]), .A1(n297), .B0(n315), 
        .B1(requesterAddressIn_SOUTH[5]), .Y(n1707) );
  AOI222XLTS U2044 ( .A0(prevRequesterAddress_A[5]), .A1(n274), .B0(
        \requesterAddressBuffer[0][5] ), .B1(n262), .C0(n1595), .C1(
        requesterAddressIn_WEST[5]), .Y(n1708) );
  OAI211X1TS U2045 ( .A0(n1974), .A1(n1547), .B0(n1548), .C0(n1549), .Y(n3277)
         );
  AOI222XLTS U2046 ( .A0(n458), .A1(n2360), .B0(n446), .B1(n2240), .C0(
        cacheAddressIn_SOUTH[7]), .C1(n435), .Y(n1549) );
  AOI22X1TS U2047 ( .A0(cacheAddressIn_NORTH[7]), .A1(n422), .B0(n487), .B1(
        n775), .Y(n1548) );
  OAI211X1TS U2048 ( .A0(n1975), .A1(n464), .B0(n1658), .C0(n1659), .Y(n3218)
         );
  AOI222XLTS U2049 ( .A0(n460), .A1(n2242), .B0(n449), .B1(n2122), .C0(n436), 
        .C1(dataIn_SOUTH[0]), .Y(n1659) );
  AOI22X1TS U2050 ( .A0(dataIn_NORTH[0]), .A1(n426), .B0(n482), .B1(n736), .Y(
        n1658) );
  OAI211X1TS U2051 ( .A0(n1976), .A1(n464), .B0(n1656), .C0(n1657), .Y(n3219)
         );
  AOI222XLTS U2052 ( .A0(n461), .A1(n2245), .B0(n450), .B1(n2125), .C0(n439), 
        .C1(dataIn_SOUTH[1]), .Y(n1657) );
  AOI22X1TS U2053 ( .A0(dataIn_NORTH[1]), .A1(n424), .B0(n486), .B1(n735), .Y(
        n1656) );
  OAI211X1TS U2054 ( .A0(n1977), .A1(n464), .B0(n1654), .C0(n1655), .Y(n3220)
         );
  AOI222XLTS U2055 ( .A0(n462), .A1(n2248), .B0(n448), .B1(n2128), .C0(n439), 
        .C1(dataIn_SOUTH[2]), .Y(n1655) );
  AOI22X1TS U2056 ( .A0(dataIn_NORTH[2]), .A1(n423), .B0(n486), .B1(n734), .Y(
        n1654) );
  OAI211X1TS U2057 ( .A0(n1978), .A1(n465), .B0(n1652), .C0(n1653), .Y(n3221)
         );
  AOI222XLTS U2058 ( .A0(n460), .A1(n2251), .B0(n448), .B1(n2131), .C0(n436), 
        .C1(dataIn_SOUTH[3]), .Y(n1653) );
  AOI22X1TS U2059 ( .A0(dataIn_NORTH[3]), .A1(n424), .B0(n486), .B1(n733), .Y(
        n1652) );
  OAI211X1TS U2060 ( .A0(n1979), .A1(n465), .B0(n1650), .C0(n1651), .Y(n3222)
         );
  AOI222XLTS U2061 ( .A0(n462), .A1(n2254), .B0(n450), .B1(n2134), .C0(n428), 
        .C1(dataIn_SOUTH[4]), .Y(n1651) );
  AOI22X1TS U2062 ( .A0(dataIn_NORTH[4]), .A1(n1553), .B0(n486), .B1(n732), 
        .Y(n1650) );
  OAI211X1TS U2063 ( .A0(n1980), .A1(n465), .B0(n1648), .C0(n1649), .Y(n3223)
         );
  AOI222XLTS U2064 ( .A0(n1550), .A1(n2257), .B0(n1551), .B1(n2137), .C0(n428), 
        .C1(dataIn_SOUTH[5]), .Y(n1649) );
  AOI22X1TS U2065 ( .A0(dataIn_NORTH[5]), .A1(n425), .B0(n485), .B1(n731), .Y(
        n1648) );
  OAI211X1TS U2066 ( .A0(n1981), .A1(n465), .B0(n1646), .C0(n1647), .Y(n3224)
         );
  AOI222XLTS U2067 ( .A0(n461), .A1(n2260), .B0(n449), .B1(n2140), .C0(n428), 
        .C1(dataIn_SOUTH[6]), .Y(n1647) );
  AOI22X1TS U2068 ( .A0(dataIn_NORTH[6]), .A1(n1553), .B0(n485), .B1(n730), 
        .Y(n1646) );
  OAI211X1TS U2069 ( .A0(n1982), .A1(n466), .B0(n1644), .C0(n1645), .Y(n3225)
         );
  AOI222XLTS U2070 ( .A0(n1550), .A1(n2263), .B0(n1551), .B1(n2143), .C0(n428), 
        .C1(dataIn_SOUTH[7]), .Y(n1645) );
  AOI22X1TS U2071 ( .A0(dataIn_NORTH[7]), .A1(n425), .B0(n485), .B1(n729), .Y(
        n1644) );
  OAI211X1TS U2072 ( .A0(n1983), .A1(n466), .B0(n1642), .C0(n1643), .Y(n3226)
         );
  AOI222XLTS U2073 ( .A0(n463), .A1(n2266), .B0(n451), .B1(n2146), .C0(n429), 
        .C1(dataIn_SOUTH[8]), .Y(n1643) );
  AOI22X1TS U2074 ( .A0(dataIn_NORTH[8]), .A1(n427), .B0(n485), .B1(n728), .Y(
        n1642) );
  OAI211X1TS U2075 ( .A0(n1984), .A1(n466), .B0(n1640), .C0(n1641), .Y(n3227)
         );
  AOI222XLTS U2076 ( .A0(n459), .A1(n2269), .B0(n447), .B1(n2149), .C0(n429), 
        .C1(dataIn_SOUTH[9]), .Y(n1641) );
  AOI22X1TS U2077 ( .A0(dataIn_NORTH[9]), .A1(n423), .B0(n484), .B1(n727), .Y(
        n1640) );
  OAI211X1TS U2078 ( .A0(n1985), .A1(n466), .B0(n1638), .C0(n1639), .Y(n3228)
         );
  AOI222XLTS U2079 ( .A0(n463), .A1(n2272), .B0(n451), .B1(n2152), .C0(n429), 
        .C1(dataIn_SOUTH[10]), .Y(n1639) );
  AOI22X1TS U2080 ( .A0(dataIn_NORTH[10]), .A1(n426), .B0(n484), .B1(n726), 
        .Y(n1638) );
  OAI211X1TS U2081 ( .A0(n1986), .A1(n467), .B0(n1636), .C0(n1637), .Y(n3229)
         );
  AOI222XLTS U2082 ( .A0(n462), .A1(n2275), .B0(n450), .B1(n2155), .C0(n429), 
        .C1(dataIn_SOUTH[11]), .Y(n1637) );
  AOI22X1TS U2083 ( .A0(dataIn_NORTH[11]), .A1(n427), .B0(n484), .B1(n725), 
        .Y(n1636) );
  OAI211X1TS U2084 ( .A0(n1987), .A1(n467), .B0(n1634), .C0(n1635), .Y(n3230)
         );
  AOI222XLTS U2085 ( .A0(n452), .A1(n2278), .B0(n440), .B1(n2158), .C0(n430), 
        .C1(dataIn_SOUTH[12]), .Y(n1635) );
  AOI22X1TS U2086 ( .A0(dataIn_NORTH[12]), .A1(n416), .B0(n484), .B1(n724), 
        .Y(n1634) );
  OAI211X1TS U2087 ( .A0(n1988), .A1(n467), .B0(n1632), .C0(n1633), .Y(n3231)
         );
  AOI222XLTS U2088 ( .A0(n452), .A1(n2281), .B0(n440), .B1(n2161), .C0(n430), 
        .C1(dataIn_SOUTH[13]), .Y(n1633) );
  AOI22X1TS U2089 ( .A0(dataIn_NORTH[13]), .A1(n416), .B0(n483), .B1(n723), 
        .Y(n1632) );
  OAI211X1TS U2090 ( .A0(n1989), .A1(n467), .B0(n1630), .C0(n1631), .Y(n3232)
         );
  AOI222XLTS U2091 ( .A0(n452), .A1(n2284), .B0(n440), .B1(n2164), .C0(n430), 
        .C1(dataIn_SOUTH[14]), .Y(n1631) );
  AOI22X1TS U2092 ( .A0(dataIn_NORTH[14]), .A1(n416), .B0(n483), .B1(n722), 
        .Y(n1630) );
  OAI211X1TS U2093 ( .A0(n1990), .A1(n468), .B0(n1628), .C0(n1629), .Y(n3233)
         );
  AOI222XLTS U2094 ( .A0(n452), .A1(n2287), .B0(n440), .B1(n2167), .C0(n430), 
        .C1(dataIn_SOUTH[15]), .Y(n1629) );
  AOI22X1TS U2095 ( .A0(dataIn_NORTH[15]), .A1(n416), .B0(n483), .B1(n721), 
        .Y(n1628) );
  OAI211X1TS U2096 ( .A0(n1991), .A1(n468), .B0(n1626), .C0(n1627), .Y(n3234)
         );
  AOI222XLTS U2097 ( .A0(n453), .A1(n2290), .B0(n441), .B1(n2170), .C0(n431), 
        .C1(dataIn_SOUTH[16]), .Y(n1627) );
  AOI22X1TS U2098 ( .A0(dataIn_NORTH[16]), .A1(n417), .B0(n483), .B1(n720), 
        .Y(n1626) );
  OAI211X1TS U2099 ( .A0(n1992), .A1(n468), .B0(n1624), .C0(n1625), .Y(n3235)
         );
  AOI222XLTS U2100 ( .A0(n453), .A1(n2293), .B0(n441), .B1(n2173), .C0(n431), 
        .C1(dataIn_SOUTH[17]), .Y(n1625) );
  AOI22X1TS U2101 ( .A0(dataIn_NORTH[17]), .A1(n417), .B0(n482), .B1(n719), 
        .Y(n1624) );
  OAI211X1TS U2102 ( .A0(n1993), .A1(n468), .B0(n1622), .C0(n1623), .Y(n3236)
         );
  AOI222XLTS U2103 ( .A0(n453), .A1(n2296), .B0(n441), .B1(n2176), .C0(n431), 
        .C1(dataIn_SOUTH[18]), .Y(n1623) );
  AOI22X1TS U2104 ( .A0(dataIn_NORTH[18]), .A1(n417), .B0(n482), .B1(n718), 
        .Y(n1622) );
  OAI211X1TS U2105 ( .A0(n1994), .A1(n469), .B0(n1620), .C0(n1621), .Y(n3237)
         );
  AOI222XLTS U2106 ( .A0(n453), .A1(n2299), .B0(n441), .B1(n2179), .C0(n431), 
        .C1(dataIn_SOUTH[19]), .Y(n1621) );
  AOI22X1TS U2107 ( .A0(dataIn_NORTH[19]), .A1(n417), .B0(n482), .B1(n717), 
        .Y(n1620) );
  OAI211X1TS U2108 ( .A0(n1995), .A1(n469), .B0(n1618), .C0(n1619), .Y(n3238)
         );
  AOI222XLTS U2109 ( .A0(n454), .A1(n2302), .B0(n442), .B1(n2182), .C0(n432), 
        .C1(dataIn_SOUTH[20]), .Y(n1619) );
  AOI22X1TS U2110 ( .A0(dataIn_NORTH[20]), .A1(n418), .B0(n481), .B1(n716), 
        .Y(n1618) );
  OAI211X1TS U2111 ( .A0(n1996), .A1(n469), .B0(n1616), .C0(n1617), .Y(n3239)
         );
  AOI222XLTS U2112 ( .A0(n454), .A1(n2305), .B0(n442), .B1(n2185), .C0(n432), 
        .C1(dataIn_SOUTH[21]), .Y(n1617) );
  AOI22X1TS U2113 ( .A0(dataIn_NORTH[21]), .A1(n418), .B0(n481), .B1(n793), 
        .Y(n1616) );
  OAI211X1TS U2114 ( .A0(n1997), .A1(n469), .B0(n1614), .C0(n1615), .Y(n3240)
         );
  AOI222XLTS U2115 ( .A0(n454), .A1(n2308), .B0(n442), .B1(n2188), .C0(n432), 
        .C1(dataIn_SOUTH[22]), .Y(n1615) );
  AOI22X1TS U2116 ( .A0(dataIn_NORTH[22]), .A1(n418), .B0(n481), .B1(n792), 
        .Y(n1614) );
  OAI211X1TS U2117 ( .A0(n1998), .A1(n470), .B0(n1612), .C0(n1613), .Y(n3241)
         );
  AOI222XLTS U2118 ( .A0(n454), .A1(n2311), .B0(n442), .B1(n2191), .C0(n432), 
        .C1(dataIn_SOUTH[23]), .Y(n1613) );
  AOI22X1TS U2119 ( .A0(dataIn_NORTH[23]), .A1(n418), .B0(n481), .B1(n791), 
        .Y(n1612) );
  OAI211X1TS U2120 ( .A0(n1999), .A1(n470), .B0(n1610), .C0(n1611), .Y(n3242)
         );
  AOI222XLTS U2121 ( .A0(n455), .A1(n2314), .B0(n443), .B1(n2194), .C0(n438), 
        .C1(dataIn_SOUTH[24]), .Y(n1611) );
  AOI22X1TS U2122 ( .A0(dataIn_NORTH[24]), .A1(n419), .B0(n480), .B1(n790), 
        .Y(n1610) );
  OAI211X1TS U2123 ( .A0(n2000), .A1(n470), .B0(n1608), .C0(n1609), .Y(n3243)
         );
  AOI222XLTS U2124 ( .A0(n455), .A1(n2317), .B0(n443), .B1(n2197), .C0(n437), 
        .C1(dataIn_SOUTH[25]), .Y(n1609) );
  AOI22X1TS U2125 ( .A0(dataIn_NORTH[25]), .A1(n419), .B0(n480), .B1(n789), 
        .Y(n1608) );
  OAI211X1TS U2126 ( .A0(n2001), .A1(n470), .B0(n1606), .C0(n1607), .Y(n3244)
         );
  AOI222XLTS U2127 ( .A0(n455), .A1(n2320), .B0(n443), .B1(n2200), .C0(n438), 
        .C1(dataIn_SOUTH[26]), .Y(n1607) );
  AOI22X1TS U2128 ( .A0(dataIn_NORTH[26]), .A1(n419), .B0(n480), .B1(n788), 
        .Y(n1606) );
  OAI211X1TS U2129 ( .A0(n2002), .A1(n471), .B0(n1604), .C0(n1605), .Y(n3245)
         );
  AOI222XLTS U2130 ( .A0(n455), .A1(n2323), .B0(n443), .B1(n2203), .C0(n437), 
        .C1(dataIn_SOUTH[27]), .Y(n1605) );
  AOI22X1TS U2131 ( .A0(dataIn_NORTH[27]), .A1(n419), .B0(n480), .B1(n787), 
        .Y(n1604) );
  OAI211X1TS U2132 ( .A0(n2003), .A1(n471), .B0(n1602), .C0(n1603), .Y(n3246)
         );
  AOI222XLTS U2133 ( .A0(n456), .A1(n2326), .B0(n444), .B1(n2206), .C0(n433), 
        .C1(dataIn_SOUTH[28]), .Y(n1603) );
  AOI22X1TS U2134 ( .A0(dataIn_NORTH[28]), .A1(n420), .B0(n479), .B1(n786), 
        .Y(n1602) );
  OAI211X1TS U2135 ( .A0(n2004), .A1(n471), .B0(n1600), .C0(n1601), .Y(n3247)
         );
  AOI222XLTS U2136 ( .A0(n456), .A1(n2329), .B0(n444), .B1(n2209), .C0(n433), 
        .C1(dataIn_SOUTH[29]), .Y(n1601) );
  AOI22X1TS U2137 ( .A0(dataIn_NORTH[29]), .A1(n420), .B0(n479), .B1(n785), 
        .Y(n1600) );
  OAI211X1TS U2138 ( .A0(n2005), .A1(n471), .B0(n1598), .C0(n1599), .Y(n3248)
         );
  AOI222XLTS U2139 ( .A0(n456), .A1(n2332), .B0(n444), .B1(n2212), .C0(n433), 
        .C1(dataIn_SOUTH[30]), .Y(n1599) );
  AOI22X1TS U2140 ( .A0(dataIn_NORTH[30]), .A1(n420), .B0(n479), .B1(n784), 
        .Y(n1598) );
  OAI211X1TS U2141 ( .A0(n2006), .A1(n472), .B0(n1596), .C0(n1597), .Y(n3249)
         );
  AOI222XLTS U2142 ( .A0(n456), .A1(n2335), .B0(n444), .B1(n2215), .C0(n433), 
        .C1(dataIn_SOUTH[31]), .Y(n1597) );
  AOI22X1TS U2143 ( .A0(dataIn_NORTH[31]), .A1(n420), .B0(n479), .B1(n783), 
        .Y(n1596) );
  OAI211X1TS U2144 ( .A0(n1967), .A1(n472), .B0(n1566), .C0(n1567), .Y(n3270)
         );
  AOI222XLTS U2145 ( .A0(n457), .A1(n2345), .B0(n445), .B1(n2225), .C0(
        cacheAddressIn_SOUTH[0]), .C1(n434), .Y(n1567) );
  AOI22X1TS U2146 ( .A0(cacheAddressIn_NORTH[0]), .A1(n421), .B0(n478), .B1(
        n782), .Y(n1566) );
  OAI211X1TS U2147 ( .A0(n1968), .A1(n472), .B0(n1564), .C0(n1565), .Y(n3271)
         );
  AOI222XLTS U2148 ( .A0(n457), .A1(n2347), .B0(n445), .B1(n2227), .C0(
        cacheAddressIn_SOUTH[1]), .C1(n434), .Y(n1565) );
  AOI22X1TS U2149 ( .A0(cacheAddressIn_NORTH[1]), .A1(n421), .B0(n478), .B1(
        n781), .Y(n1564) );
  OAI211X1TS U2150 ( .A0(n1969), .A1(n472), .B0(n1562), .C0(n1563), .Y(n3272)
         );
  AOI222XLTS U2151 ( .A0(n457), .A1(n2348), .B0(n445), .B1(n2229), .C0(
        cacheAddressIn_SOUTH[2]), .C1(n434), .Y(n1563) );
  AOI22X1TS U2152 ( .A0(cacheAddressIn_NORTH[2]), .A1(n421), .B0(n478), .B1(
        n780), .Y(n1562) );
  OAI211X1TS U2153 ( .A0(n1970), .A1(n473), .B0(n1560), .C0(n1561), .Y(n3273)
         );
  AOI222XLTS U2154 ( .A0(n457), .A1(n2351), .B0(n445), .B1(n2231), .C0(
        cacheAddressIn_SOUTH[3]), .C1(n434), .Y(n1561) );
  AOI22X1TS U2155 ( .A0(cacheAddressIn_NORTH[3]), .A1(n421), .B0(n478), .B1(
        n779), .Y(n1560) );
  OAI211X1TS U2156 ( .A0(n1971), .A1(n473), .B0(n1558), .C0(n1559), .Y(n3274)
         );
  AOI222XLTS U2157 ( .A0(n458), .A1(n2352), .B0(n446), .B1(n2232), .C0(
        cacheAddressIn_SOUTH[4]), .C1(n435), .Y(n1559) );
  AOI22X1TS U2158 ( .A0(cacheAddressIn_NORTH[4]), .A1(n422), .B0(n1446), .B1(
        n778), .Y(n1558) );
  OAI211X1TS U2159 ( .A0(n1972), .A1(n473), .B0(n1556), .C0(n1557), .Y(n3275)
         );
  AOI222XLTS U2160 ( .A0(n458), .A1(n2355), .B0(n446), .B1(n2234), .C0(
        cacheAddressIn_SOUTH[5]), .C1(n435), .Y(n1557) );
  AOI22X1TS U2161 ( .A0(cacheAddressIn_NORTH[5]), .A1(n422), .B0(n1446), .B1(
        n777), .Y(n1556) );
  OAI211X1TS U2162 ( .A0(n1973), .A1(n473), .B0(n1554), .C0(n1555), .Y(n3276)
         );
  AOI222XLTS U2163 ( .A0(n458), .A1(n2357), .B0(n446), .B1(n2237), .C0(
        cacheAddressIn_SOUTH[6]), .C1(n435), .Y(n1555) );
  AOI22X1TS U2164 ( .A0(cacheAddressIn_NORTH[6]), .A1(n422), .B0(n1446), .B1(
        n776), .Y(n1554) );
  XOR2X1TS U2165 ( .A(n994), .B(n114), .Y(n985) );
  XNOR2X1TS U2166 ( .A(n996), .B(n122), .Y(n994) );
  AOI2BB2X1TS U2167 ( .B0(n112), .B1(n316), .A0N(n316), .A1N(n1665), .Y(n1428)
         );
  OAI22X1TS U2168 ( .A0(n2095), .A1(n464), .B0(n476), .B1(n1712), .Y(n3184) );
  AOI221X1TS U2169 ( .A0(n1175), .A1(n336), .B0(n292), .B1(n1445), .C0(n2371), 
        .Y(n1712) );
  OAI22X1TS U2170 ( .A0(n72), .A1(n302), .B0(n1490), .B1(n282), .Y(n3317) );
  AOI222XLTS U2171 ( .A0(n1883), .A1(n191), .B0(n146), .B1(n2345), .C0(n2224), 
        .C1(n120), .Y(n1490) );
  OAI22X1TS U2172 ( .A0(n73), .A1(n301), .B0(n1493), .B1(n282), .Y(n3316) );
  AOI222XLTS U2173 ( .A0(n1884), .A1(n828), .B0(n147), .B1(n2347), .C0(n2226), 
        .C1(n1243), .Y(n1493) );
  OAI22X1TS U2174 ( .A0(n74), .A1(n302), .B0(n1494), .B1(n282), .Y(n3315) );
  AOI222XLTS U2175 ( .A0(n1885), .A1(n189), .B0(n146), .B1(n2348), .C0(n2228), 
        .C1(n121), .Y(n1494) );
  OAI22X1TS U2176 ( .A0(n75), .A1(n301), .B0(n1495), .B1(n282), .Y(n3314) );
  AOI222XLTS U2177 ( .A0(n1886), .A1(n190), .B0(n147), .B1(n2351), .C0(n2230), 
        .C1(n1243), .Y(n1495) );
  OAI22X1TS U2178 ( .A0(n76), .A1(n302), .B0(n1496), .B1(n283), .Y(n3313) );
  AOI222XLTS U2179 ( .A0(n1887), .A1(n191), .B0(n146), .B1(n2352), .C0(n2233), 
        .C1(n120), .Y(n1496) );
  OAI22X1TS U2180 ( .A0(n77), .A1(n301), .B0(n1497), .B1(n283), .Y(n3312) );
  AOI222XLTS U2181 ( .A0(n1888), .A1(n328), .B0(n147), .B1(n2355), .C0(n2235), 
        .C1(n1243), .Y(n1497) );
  OAI22X1TS U2182 ( .A0(n78), .A1(n302), .B0(n1498), .B1(n283), .Y(n3311) );
  AOI222XLTS U2183 ( .A0(n1889), .A1(n189), .B0(n146), .B1(n2357), .C0(n2238), 
        .C1(n121), .Y(n1498) );
  OAI22X1TS U2184 ( .A0(n79), .A1(n301), .B0(n1499), .B1(n283), .Y(n3310) );
  AOI222XLTS U2185 ( .A0(n1890), .A1(n190), .B0(n147), .B1(n2360), .C0(n2241), 
        .C1(n121), .Y(n1499) );
  OAI22X1TS U2186 ( .A0(n174), .A1(n46), .B0(n2367), .B1(n1571), .Y(n3267) );
  AOI21X1TS U2187 ( .A0(n1963), .A1(n310), .B0(n1377), .Y(n1571) );
  OAI22X1TS U2188 ( .A0(n172), .A1(n47), .B0(n2367), .B1(n1572), .Y(n3266) );
  AOI21X1TS U2189 ( .A0(n1964), .A1(n309), .B0(n1377), .Y(n1572) );
  OAI22X1TS U2190 ( .A0(n1174), .A1(n173), .B0(n1375), .B1(n1376), .Y(n3384)
         );
  AOI2BB2X1TS U2191 ( .B0(n1377), .B1(n112), .A0N(n989), .A1N(n1172), .Y(n1375) );
  OAI22X1TS U2192 ( .A0(n2097), .A1(n2093), .B0(n1663), .B1(n1664), .Y(n3217)
         );
  AOI221X1TS U2193 ( .A0(n1174), .A1(n337), .B0(n1428), .B1(n341), .C0(n2371), 
        .Y(n1664) );
  NAND2X1TS U2194 ( .A(n3677), .B(n741), .Y(n1735) );
  NAND2X1TS U2195 ( .A(n3678), .B(n740), .Y(n1747) );
  NAND2X1TS U2196 ( .A(n3678), .B(n3677), .Y(n1759) );
  OAI22X1TS U2197 ( .A0(n1175), .A1(n289), .B0(n1370), .B1(n1371), .Y(n3385)
         );
  AOI222XLTS U2198 ( .A0(n336), .A1(n768), .B0(memWrite_EAST), .B1(n277), .C0(
        memWrite_WEST), .C1(n305), .Y(n1370) );
  OAI22X1TS U2199 ( .A0(n1242), .A1(n291), .B0(n1452), .B1(n263), .Y(n3341) );
  AOI222XLTS U2200 ( .A0(n335), .A1(n767), .B0(n2344), .B1(n277), .C0(
        cacheAddressIn_WEST[0]), .C1(n305), .Y(n1452) );
  OAI22X1TS U2201 ( .A0(n1241), .A1(n290), .B0(n1453), .B1(n264), .Y(n3340) );
  AOI222XLTS U2202 ( .A0(n337), .A1(n766), .B0(n2346), .B1(n275), .C0(
        cacheAddressIn_WEST[1]), .C1(n307), .Y(n1453) );
  OAI22X1TS U2203 ( .A0(n1240), .A1(n291), .B0(n1454), .B1(n1371), .Y(n3339)
         );
  AOI222XLTS U2204 ( .A0(n336), .A1(n765), .B0(n2349), .B1(n275), .C0(
        cacheAddressIn_WEST[2]), .C1(n306), .Y(n1454) );
  OAI22X1TS U2205 ( .A0(n1239), .A1(n290), .B0(n1455), .B1(n263), .Y(n3338) );
  AOI222XLTS U2206 ( .A0(n335), .A1(n764), .B0(n2350), .B1(n276), .C0(
        cacheAddressIn_WEST[3]), .C1(n307), .Y(n1455) );
  OAI22X1TS U2207 ( .A0(n1238), .A1(n291), .B0(n1456), .B1(n264), .Y(n3337) );
  AOI222XLTS U2208 ( .A0(n337), .A1(n763), .B0(n2353), .B1(n277), .C0(
        cacheAddressIn_WEST[4]), .C1(n306), .Y(n1456) );
  OAI22X1TS U2209 ( .A0(n1237), .A1(n290), .B0(n1457), .B1(n1371), .Y(n3336)
         );
  AOI222XLTS U2210 ( .A0(n336), .A1(n762), .B0(n2354), .B1(n276), .C0(
        cacheAddressIn_WEST[5]), .C1(n307), .Y(n1457) );
  OAI22X1TS U2211 ( .A0(n1236), .A1(n291), .B0(n1458), .B1(n263), .Y(n3335) );
  AOI222XLTS U2212 ( .A0(n335), .A1(n761), .B0(n2358), .B1(n277), .C0(
        cacheAddressIn_WEST[6]), .C1(n306), .Y(n1458) );
  OAI22X1TS U2213 ( .A0(n1235), .A1(n290), .B0(n1459), .B1(n264), .Y(n3334) );
  AOI222XLTS U2214 ( .A0(n335), .A1(n760), .B0(n2361), .B1(n276), .C0(
        cacheAddressIn_WEST[7]), .C1(n307), .Y(n1459) );
  OAI222X1TS U2215 ( .A0(n1713), .A1(n1661), .B0(memWrite_EAST), .B1(n125), 
        .C0(memWrite_WEST), .C1(n113), .Y(n1445) );
  OAI2BB1X1TS U2216 ( .A0N(requesterAddressOut_SOUTH[0]), .A1N(n131), .B0(
        n1746), .Y(n3166) );
  AOI22X1TS U2217 ( .A0(n314), .A1(prevRequesterAddress_B[0]), .B0(n295), .B1(
        prevRequesterAddress_A[0]), .Y(n1746) );
  OAI2BB1X1TS U2218 ( .A0N(requesterAddressOut_SOUTH[1]), .A1N(n1738), .B0(
        n1745), .Y(n3167) );
  AOI22X1TS U2219 ( .A0(n1740), .A1(prevRequesterAddress_B[1]), .B0(n1741), 
        .B1(prevRequesterAddress_A[1]), .Y(n1745) );
  OAI2BB1X1TS U2220 ( .A0N(requesterAddressOut_SOUTH[2]), .A1N(n131), .B0(
        n1744), .Y(n3168) );
  AOI22X1TS U2221 ( .A0(n1740), .A1(prevRequesterAddress_B[2]), .B0(n1741), 
        .B1(prevRequesterAddress_A[2]), .Y(n1744) );
  OAI2BB1X1TS U2222 ( .A0N(requesterAddressOut_SOUTH[3]), .A1N(n1738), .B0(
        n1743), .Y(n3169) );
  AOI22X1TS U2223 ( .A0(n1740), .A1(prevRequesterAddress_B[3]), .B0(n1741), 
        .B1(prevRequesterAddress_A[3]), .Y(n1743) );
  OAI2BB1X1TS U2224 ( .A0N(requesterAddressOut_SOUTH[4]), .A1N(n131), .B0(
        n1742), .Y(n3170) );
  AOI22X1TS U2225 ( .A0(n314), .A1(prevRequesterAddress_B[4]), .B0(n295), .B1(
        prevRequesterAddress_A[4]), .Y(n1742) );
  OAI2BB1X1TS U2226 ( .A0N(requesterAddressOut_SOUTH[5]), .A1N(n1738), .B0(
        n1739), .Y(n3171) );
  AOI22X1TS U2227 ( .A0(n314), .A1(prevRequesterAddress_B[5]), .B0(n295), .B1(
        prevRequesterAddress_A[5]), .Y(n1739) );
  OAI2BB1X1TS U2228 ( .A0N(requesterAddressOut_EAST[0]), .A1N(n133), .B0(n1734), .Y(n3172) );
  AOI22X1TS U2229 ( .A0(n278), .A1(prevRequesterAddress_B[0]), .B0(n313), .B1(
        prevRequesterAddress_A[0]), .Y(n1734) );
  OAI2BB1X1TS U2230 ( .A0N(requesterAddressOut_EAST[1]), .A1N(n1726), .B0(
        n1733), .Y(n3173) );
  AOI22X1TS U2231 ( .A0(n1728), .A1(prevRequesterAddress_B[1]), .B0(n1729), 
        .B1(prevRequesterAddress_A[1]), .Y(n1733) );
  OAI2BB1X1TS U2232 ( .A0N(requesterAddressOut_EAST[2]), .A1N(n133), .B0(n1732), .Y(n3174) );
  AOI22X1TS U2233 ( .A0(n1728), .A1(prevRequesterAddress_B[2]), .B0(n1729), 
        .B1(prevRequesterAddress_A[2]), .Y(n1732) );
  OAI2BB1X1TS U2234 ( .A0N(requesterAddressOut_EAST[3]), .A1N(n1726), .B0(
        n1731), .Y(n3175) );
  AOI22X1TS U2235 ( .A0(n1728), .A1(prevRequesterAddress_B[3]), .B0(n1729), 
        .B1(prevRequesterAddress_A[3]), .Y(n1731) );
  OAI2BB1X1TS U2236 ( .A0N(requesterAddressOut_EAST[4]), .A1N(n133), .B0(n1730), .Y(n3176) );
  AOI22X1TS U2237 ( .A0(n278), .A1(prevRequesterAddress_B[4]), .B0(n313), .B1(
        prevRequesterAddress_A[4]), .Y(n1730) );
  OAI2BB1X1TS U2238 ( .A0N(requesterAddressOut_EAST[5]), .A1N(n1726), .B0(
        n1727), .Y(n3177) );
  AOI22X1TS U2239 ( .A0(n278), .A1(prevRequesterAddress_B[5]), .B0(n313), .B1(
        prevRequesterAddress_A[5]), .Y(n1727) );
  OAI32X1TS U2240 ( .A0(n1418), .A1(n2369), .A2(n802), .B0(n1419), .B1(n30), 
        .Y(n3345) );
  AOI21X1TS U2241 ( .A0(n1422), .A1(n1423), .B0(memRead_WEST), .Y(n1418) );
  INVX2TS U2242 ( .A(n1419), .Y(n802) );
  NAND2X1TS U2243 ( .A(n1420), .B(n1421), .Y(n1419) );
  OAI221XLTS U2244 ( .A0(n552), .A1(n1569), .B0(n2368), .B1(n813), .C0(n1570), 
        .Y(n3268) );
  AOI22X1TS U2245 ( .A0(\requesterPortBuffer[0][1] ), .A1(n1460), .B0(n1966), 
        .B1(n487), .Y(n1570) );
  OAI211X1TS U2246 ( .A0(n837), .A1(n1573), .B0(n140), .C0(n1574), .Y(n3265)
         );
  AOI22X1TS U2247 ( .A0(n1575), .A1(n2096), .B0(prevRequesterPort_B[0]), .B1(
        n1576), .Y(n1574) );
  OAI211X1TS U2248 ( .A0(n1666), .A1(n1573), .B0(n140), .C0(n1577), .Y(n3264)
         );
  AOI22X1TS U2249 ( .A0(n1575), .A1(n2100), .B0(prevRequesterPort_B[1]), .B1(
        n1576), .Y(n1577) );
  OAI211X1TS U2250 ( .A0(n832), .A1(n1590), .B0(n142), .C0(n1594), .Y(n3250)
         );
  AOI22X1TS U2251 ( .A0(n262), .A1(\requesterPortBuffer[0][0] ), .B0(n274), 
        .B1(n740), .Y(n1594) );
  OAI211X1TS U2252 ( .A0(n125), .A1(n1590), .B0(n142), .C0(n1591), .Y(n3251)
         );
  AOI22X1TS U2253 ( .A0(n262), .A1(\requesterPortBuffer[0][1] ), .B0(n273), 
        .B1(n741), .Y(n1591) );
  INVX2TS U2254 ( .A(n1568), .Y(n645) );
  AOI222XLTS U2255 ( .A0(n487), .A1(\requesterPortBuffer[2][0] ), .B0(n1460), 
        .B1(\requesterPortBuffer[0][0] ), .C0(n2376), .C1(n306), .Y(n1568) );
  INVX2TS U2256 ( .A(n1444), .Y(n596) );
  AOI32X1TS U2257 ( .A0(n551), .A1(n1429), .A2(n1445), .B0(n487), .B1(n2098), 
        .Y(n1444) );
  NOR2X1TS U2258 ( .A(prevRequesterPort_B[1]), .B(prevRequesterPort_B[0]), .Y(
        n1761) );
  NOR2X1TS U2259 ( .A(n26), .B(prevRequesterPort_B[1]), .Y(n1749) );
  NOR2X1TS U2260 ( .A(n1), .B(prevRequesterPort_B[0]), .Y(n1737) );
  OAI21X1TS U2261 ( .A0(n1424), .A1(n1425), .B0(n844), .Y(n1423) );
  OAI2BB1X1TS U2262 ( .A0N(requesterAddressOut_NORTH[0]), .A1N(n129), .B0(
        n1758), .Y(n3160) );
  AOI22X1TS U2263 ( .A0(n312), .A1(prevRequesterAddress_B[0]), .B0(n265), .B1(
        prevRequesterAddress_A[0]), .Y(n1758) );
  OAI2BB1X1TS U2264 ( .A0N(requesterAddressOut_NORTH[1]), .A1N(n1750), .B0(
        n1757), .Y(n3161) );
  AOI22X1TS U2265 ( .A0(n1752), .A1(prevRequesterAddress_B[1]), .B0(n1753), 
        .B1(prevRequesterAddress_A[1]), .Y(n1757) );
  OAI2BB1X1TS U2266 ( .A0N(requesterAddressOut_NORTH[2]), .A1N(n129), .B0(
        n1756), .Y(n3162) );
  AOI22X1TS U2267 ( .A0(n1752), .A1(prevRequesterAddress_B[2]), .B0(n1753), 
        .B1(prevRequesterAddress_A[2]), .Y(n1756) );
  OAI2BB1X1TS U2268 ( .A0N(requesterAddressOut_NORTH[3]), .A1N(n1750), .B0(
        n1755), .Y(n3163) );
  AOI22X1TS U2269 ( .A0(n1752), .A1(prevRequesterAddress_B[3]), .B0(n1753), 
        .B1(prevRequesterAddress_A[3]), .Y(n1755) );
  OAI2BB1X1TS U2270 ( .A0N(requesterAddressOut_NORTH[4]), .A1N(n129), .B0(
        n1754), .Y(n3164) );
  AOI22X1TS U2271 ( .A0(n312), .A1(prevRequesterAddress_B[4]), .B0(n265), .B1(
        prevRequesterAddress_A[4]), .Y(n1754) );
  OAI2BB1X1TS U2272 ( .A0N(requesterAddressOut_NORTH[5]), .A1N(n1750), .B0(
        n1751), .Y(n3165) );
  AOI22X1TS U2273 ( .A0(n312), .A1(prevRequesterAddress_B[5]), .B0(n265), .B1(
        prevRequesterAddress_A[5]), .Y(n1751) );
  OAI221XLTS U2274 ( .A0(n3), .A1(n1714), .B0(n256), .B1(n1715), .C0(n1722), 
        .Y(n3178) );
  NAND2X1TS U2275 ( .A(requesterAddressOut_WEST[0]), .B(n139), .Y(n1722) );
  OAI221XLTS U2276 ( .A0(n4), .A1(n1714), .B0(n255), .B1(n1715), .C0(n1721), 
        .Y(n3179) );
  NAND2X1TS U2277 ( .A(requesterAddressOut_WEST[1]), .B(n138), .Y(n1721) );
  OAI221XLTS U2278 ( .A0(n5), .A1(n1714), .B0(n254), .B1(n1715), .C0(n1720), 
        .Y(n3180) );
  NAND2X1TS U2279 ( .A(requesterAddressOut_WEST[2]), .B(n139), .Y(n1720) );
  OAI221XLTS U2280 ( .A0(n6), .A1(n311), .B0(n253), .B1(n294), .C0(n1719), .Y(
        n3181) );
  NAND2X1TS U2281 ( .A(requesterAddressOut_WEST[3]), .B(n138), .Y(n1719) );
  OAI221XLTS U2282 ( .A0(n7), .A1(n311), .B0(n252), .B1(n294), .C0(n1718), .Y(
        n3182) );
  NAND2X1TS U2283 ( .A(requesterAddressOut_WEST[4]), .B(n139), .Y(n1718) );
  OAI221XLTS U2284 ( .A0(n8), .A1(n311), .B0(n251), .B1(n294), .C0(n1716), .Y(
        n3183) );
  NAND2X1TS U2285 ( .A(requesterAddressOut_WEST[5]), .B(n138), .Y(n1716) );
  INVX2TS U2286 ( .A(dataIn_WEST[0]), .Y(n2124) );
  INVX2TS U2287 ( .A(dataIn_EAST[0]), .Y(n2244) );
  INVX2TS U2288 ( .A(dataIn_WEST[1]), .Y(n2127) );
  INVX2TS U2289 ( .A(dataIn_EAST[1]), .Y(n2247) );
  INVX2TS U2290 ( .A(dataIn_WEST[2]), .Y(n2130) );
  INVX2TS U2291 ( .A(dataIn_EAST[2]), .Y(n2250) );
  INVX2TS U2292 ( .A(dataIn_WEST[3]), .Y(n2133) );
  INVX2TS U2293 ( .A(dataIn_EAST[3]), .Y(n2253) );
  INVX2TS U2294 ( .A(dataIn_WEST[4]), .Y(n2136) );
  INVX2TS U2295 ( .A(dataIn_EAST[4]), .Y(n2256) );
  INVX2TS U2296 ( .A(dataIn_WEST[5]), .Y(n2139) );
  INVX2TS U2297 ( .A(dataIn_EAST[5]), .Y(n2259) );
  INVX2TS U2298 ( .A(dataIn_WEST[6]), .Y(n2142) );
  INVX2TS U2299 ( .A(dataIn_EAST[6]), .Y(n2262) );
  INVX2TS U2300 ( .A(dataIn_WEST[7]), .Y(n2145) );
  INVX2TS U2301 ( .A(dataIn_EAST[7]), .Y(n2265) );
  INVX2TS U2302 ( .A(dataIn_WEST[8]), .Y(n2148) );
  INVX2TS U2303 ( .A(dataIn_EAST[8]), .Y(n2268) );
  INVX2TS U2304 ( .A(dataIn_WEST[9]), .Y(n2151) );
  INVX2TS U2305 ( .A(dataIn_EAST[9]), .Y(n2271) );
  INVX2TS U2306 ( .A(dataIn_WEST[10]), .Y(n2154) );
  INVX2TS U2307 ( .A(dataIn_EAST[10]), .Y(n2274) );
  INVX2TS U2308 ( .A(dataIn_WEST[11]), .Y(n2157) );
  INVX2TS U2309 ( .A(dataIn_EAST[11]), .Y(n2277) );
  INVX2TS U2310 ( .A(dataIn_WEST[12]), .Y(n2160) );
  INVX2TS U2311 ( .A(dataIn_EAST[12]), .Y(n2280) );
  INVX2TS U2312 ( .A(dataIn_WEST[13]), .Y(n2163) );
  INVX2TS U2313 ( .A(dataIn_EAST[13]), .Y(n2283) );
  INVX2TS U2314 ( .A(dataIn_WEST[14]), .Y(n2166) );
  INVX2TS U2315 ( .A(dataIn_EAST[14]), .Y(n2286) );
  INVX2TS U2316 ( .A(dataIn_WEST[15]), .Y(n2169) );
  INVX2TS U2317 ( .A(dataIn_EAST[15]), .Y(n2289) );
  INVX2TS U2318 ( .A(dataIn_WEST[16]), .Y(n2172) );
  INVX2TS U2319 ( .A(dataIn_EAST[16]), .Y(n2292) );
  INVX2TS U2320 ( .A(dataIn_WEST[17]), .Y(n2175) );
  INVX2TS U2321 ( .A(dataIn_EAST[17]), .Y(n2295) );
  INVX2TS U2322 ( .A(dataIn_WEST[18]), .Y(n2178) );
  INVX2TS U2323 ( .A(dataIn_EAST[18]), .Y(n2298) );
  INVX2TS U2324 ( .A(dataIn_WEST[19]), .Y(n2181) );
  INVX2TS U2325 ( .A(dataIn_EAST[19]), .Y(n2301) );
  INVX2TS U2326 ( .A(dataIn_WEST[20]), .Y(n2184) );
  INVX2TS U2327 ( .A(dataIn_EAST[20]), .Y(n2304) );
  INVX2TS U2328 ( .A(dataIn_WEST[21]), .Y(n2187) );
  INVX2TS U2329 ( .A(dataIn_EAST[21]), .Y(n2307) );
  INVX2TS U2330 ( .A(dataIn_WEST[22]), .Y(n2190) );
  INVX2TS U2331 ( .A(dataIn_EAST[22]), .Y(n2310) );
  INVX2TS U2332 ( .A(dataIn_WEST[23]), .Y(n2193) );
  INVX2TS U2333 ( .A(dataIn_EAST[23]), .Y(n2313) );
  INVX2TS U2334 ( .A(dataIn_WEST[24]), .Y(n2196) );
  INVX2TS U2335 ( .A(dataIn_EAST[24]), .Y(n2316) );
  INVX2TS U2336 ( .A(dataIn_WEST[25]), .Y(n2199) );
  INVX2TS U2337 ( .A(dataIn_EAST[25]), .Y(n2319) );
  INVX2TS U2338 ( .A(dataIn_WEST[26]), .Y(n2202) );
  INVX2TS U2339 ( .A(dataIn_EAST[26]), .Y(n2322) );
  INVX2TS U2340 ( .A(dataIn_WEST[27]), .Y(n2205) );
  INVX2TS U2341 ( .A(dataIn_EAST[27]), .Y(n2325) );
  INVX2TS U2342 ( .A(dataIn_WEST[28]), .Y(n2208) );
  INVX2TS U2343 ( .A(dataIn_EAST[28]), .Y(n2328) );
  INVX2TS U2344 ( .A(dataIn_WEST[29]), .Y(n2211) );
  INVX2TS U2345 ( .A(dataIn_EAST[29]), .Y(n2331) );
  INVX2TS U2346 ( .A(dataIn_WEST[30]), .Y(n2214) );
  INVX2TS U2347 ( .A(dataIn_EAST[30]), .Y(n2334) );
  INVX2TS U2348 ( .A(dataIn_WEST[31]), .Y(n2217) );
  INVX2TS U2349 ( .A(dataIn_EAST[31]), .Y(n2337) );
  AND2X2TS U2350 ( .A(n1931), .B(n546), .Y(n3417) );
  AND2X2TS U2351 ( .A(n1932), .B(n541), .Y(n3416) );
  AND2X2TS U2352 ( .A(n1933), .B(n541), .Y(n3415) );
  AND2X2TS U2353 ( .A(n1934), .B(n542), .Y(n3414) );
  AND2X2TS U2354 ( .A(n1935), .B(n542), .Y(n3413) );
  AND2X2TS U2355 ( .A(n1936), .B(n542), .Y(n3412) );
  AND2X2TS U2356 ( .A(n1937), .B(n542), .Y(n3411) );
  AND2X2TS U2357 ( .A(n1938), .B(n543), .Y(n3410) );
  AND2X2TS U2358 ( .A(n1939), .B(n543), .Y(n3409) );
  AND2X2TS U2359 ( .A(n1940), .B(n543), .Y(n3408) );
  AND2X2TS U2360 ( .A(n1941), .B(n543), .Y(n3407) );
  AND2X2TS U2361 ( .A(n1942), .B(n544), .Y(n3406) );
  AND2X2TS U2362 ( .A(n1943), .B(n544), .Y(n3405) );
  AND2X2TS U2363 ( .A(n1944), .B(n544), .Y(n3404) );
  AND2X2TS U2364 ( .A(n1945), .B(n544), .Y(n3403) );
  AND2X2TS U2365 ( .A(n1946), .B(n545), .Y(n3402) );
  AND2X2TS U2366 ( .A(n1947), .B(n545), .Y(n3401) );
  AND2X2TS U2367 ( .A(n1948), .B(n545), .Y(n3400) );
  AND2X2TS U2368 ( .A(n1949), .B(n545), .Y(n3399) );
  AND2X2TS U2369 ( .A(n1950), .B(n546), .Y(n3398) );
  AND2X2TS U2370 ( .A(n1951), .B(n546), .Y(n3397) );
  AND2X2TS U2371 ( .A(n1952), .B(n546), .Y(n3396) );
  AND2X2TS U2372 ( .A(n1953), .B(n547), .Y(n3395) );
  AND2X2TS U2373 ( .A(n1954), .B(n547), .Y(n3394) );
  AND2X2TS U2374 ( .A(n1955), .B(n547), .Y(n3393) );
  AND2X2TS U2375 ( .A(n1956), .B(n547), .Y(n3392) );
  AND2X2TS U2376 ( .A(n1957), .B(n548), .Y(n3391) );
  AND2X2TS U2377 ( .A(n1958), .B(n548), .Y(n3390) );
  AND2X2TS U2378 ( .A(n1959), .B(n548), .Y(n3389) );
  AND2X2TS U2379 ( .A(n1960), .B(n548), .Y(n3388) );
  AND2X2TS U2380 ( .A(n1961), .B(n549), .Y(n3387) );
  AND2X2TS U2381 ( .A(n1962), .B(n549), .Y(n3386) );
  AND2X2TS U2382 ( .A(\requesterPortBuffer[7][1] ), .B(n541), .Y(n3252) );
  AND2X2TS U2383 ( .A(n1923), .B(n549), .Y(n3285) );
  AND2X2TS U2384 ( .A(n1924), .B(n550), .Y(n3284) );
  AND2X2TS U2385 ( .A(n1925), .B(n550), .Y(n3283) );
  AND2X2TS U2386 ( .A(n1926), .B(n550), .Y(n3282) );
  AND2X2TS U2387 ( .A(n1927), .B(n550), .Y(n3281) );
  AND2X2TS U2388 ( .A(n1928), .B(n551), .Y(n3280) );
  AND2X2TS U2389 ( .A(n1929), .B(n551), .Y(n3279) );
  AND2X2TS U2390 ( .A(n1930), .B(n551), .Y(n3278) );
  AND2X2TS U2391 ( .A(\requesterPortBuffer[7][0] ), .B(n549), .Y(n3253) );
  INVX2TS U2392 ( .A(n1582), .Y(n715) );
  AOI32X1TS U2393 ( .A0(\requesterPortBuffer[5][1] ), .A1(n2377), .A2(n191), 
        .B0(n1379), .B1(n1964), .Y(n1582) );
  INVX2TS U2394 ( .A(n1581), .Y(n648) );
  AOI32X1TS U2395 ( .A0(\requesterPortBuffer[5][0] ), .A1(n2380), .A2(n828), 
        .B0(n1379), .B1(n1963), .Y(n1581) );
  OAI32X1TS U2396 ( .A0(n1378), .A1(n2370), .A2(n1171), .B0(n1173), .B1(n819), 
        .Y(n3383) );
  INVX2TS U2397 ( .A(n1378), .Y(n819) );
  OAI32X1TS U2398 ( .A0(n1381), .A1(n2369), .A2(n1965), .B0(n1170), .B1(n799), 
        .Y(n3380) );
  INVX2TS U2399 ( .A(n1381), .Y(n799) );
  OAI32X1TS U2400 ( .A0(n1380), .A1(n2370), .A2(n1169), .B0(n1171), .B1(n800), 
        .Y(n3381) );
  INVX2TS U2401 ( .A(n1380), .Y(n800) );
  OAI32X1TS U2402 ( .A0(n1382), .A1(n2369), .A2(n1175), .B0(n1169), .B1(n796), 
        .Y(n3379) );
  INVX2TS U2403 ( .A(n1382), .Y(n796) );
  OAI32X1TS U2404 ( .A0(n1379), .A1(n2370), .A2(n1170), .B0(n1172), .B1(n827), 
        .Y(n3382) );
  INVX2TS U2405 ( .A(n1379), .Y(n827) );
  NOR2X1TS U2406 ( .A(n1965), .B(n555), .Y(n3378) );
  INVX2TS U2407 ( .A(n1587), .Y(n646) );
  AOI32X1TS U2408 ( .A0(\requesterPortBuffer[0][0] ), .A1(n2381), .A2(n333), 
        .B0(n1382), .B1(\requesterPortBuffer[6][0] ), .Y(n1587) );
  INVX2TS U2409 ( .A(n1588), .Y(n647) );
  AOI32X1TS U2410 ( .A0(\requesterPortBuffer[0][1] ), .A1(n2380), .A2(n331), 
        .B0(n1382), .B1(\requesterPortBuffer[6][1] ), .Y(n1588) );
  INVX2TS U2411 ( .A(n1585), .Y(n597) );
  AOI32X1TS U2412 ( .A0(\requesterPortBuffer[7][0] ), .A1(n2376), .A2(n186), 
        .B0(n1381), .B1(\requesterPortBuffer[5][0] ), .Y(n1585) );
  INVX2TS U2413 ( .A(n1586), .Y(n759) );
  AOI32X1TS U2414 ( .A0(\requesterPortBuffer[7][1] ), .A1(n2379), .A2(n187), 
        .B0(n1381), .B1(\requesterPortBuffer[5][1] ), .Y(n1586) );
  INVX2TS U2415 ( .A(n1579), .Y(n757) );
  AOI32X1TS U2416 ( .A0(\requesterPortBuffer[4][0] ), .A1(n2378), .A2(n182), 
        .B0(n1378), .B1(\requesterPortBuffer[2][0] ), .Y(n1579) );
  INVX2TS U2417 ( .A(n1583), .Y(n758) );
  AOI32X1TS U2418 ( .A0(\requesterPortBuffer[6][0] ), .A1(n2379), .A2(n178), 
        .B0(n1380), .B1(\requesterPortBuffer[4][0] ), .Y(n1583) );
  INVX2TS U2419 ( .A(n1584), .Y(n756) );
  AOI32X1TS U2420 ( .A0(\requesterPortBuffer[6][1] ), .A1(n2378), .A2(n179), 
        .B0(n1380), .B1(\requesterPortBuffer[4][1] ), .Y(n1584) );
  INVX2TS U2421 ( .A(n1580), .Y(n649) );
  AOI32X1TS U2422 ( .A0(\requesterPortBuffer[4][1] ), .A1(n2377), .A2(n183), 
        .B0(n1378), .B1(n1966), .Y(n1580) );
  INVX2TS U2423 ( .A(n880), .Y(n828) );
  NOR2X1TS U2424 ( .A(n122), .B(n4621), .Y(n1677) );
endmodule


module outputPortArbiter_0 ( clk, reset, selectBit_NORTH, 
        destinationAddressIn_NORTH, requesterAddressIn_NORTH, readIn_NORTH, 
        writeIn_NORTH, dataIn_NORTH, selectBit_SOUTH, 
        destinationAddressIn_SOUTH, requesterAddressIn_SOUTH, readIn_SOUTH, 
        writeIn_SOUTH, dataIn_SOUTH, selectBit_EAST, destinationAddressIn_EAST, 
        requesterAddressIn_EAST, readIn_EAST, writeIn_EAST, dataIn_EAST, 
        selectBit_WEST, destinationAddressIn_WEST, requesterAddressIn_WEST, 
        readIn_WEST, writeIn_WEST, dataIn_WEST, readReady, 
        readRequesterAddress, cacheDataOut, destinationAddressOut, 
        requesterAddressOut, readOut, writeOut, dataOut );
  input [13:0] destinationAddressIn_NORTH;
  input [5:0] requesterAddressIn_NORTH;
  input [31:0] dataIn_NORTH;
  input [13:0] destinationAddressIn_SOUTH;
  input [5:0] requesterAddressIn_SOUTH;
  input [31:0] dataIn_SOUTH;
  input [13:0] destinationAddressIn_EAST;
  input [5:0] requesterAddressIn_EAST;
  input [31:0] dataIn_EAST;
  input [13:0] destinationAddressIn_WEST;
  input [5:0] requesterAddressIn_WEST;
  input [31:0] dataIn_WEST;
  input [5:0] readRequesterAddress;
  input [31:0] cacheDataOut;
  output [13:0] destinationAddressOut;
  output [5:0] requesterAddressOut;
  output [31:0] dataOut;
  input clk, reset, selectBit_NORTH, readIn_NORTH, writeIn_NORTH,
         selectBit_SOUTH, readIn_SOUTH, writeIn_SOUTH, selectBit_EAST,
         readIn_EAST, writeIn_EAST, selectBit_WEST, readIn_WEST, writeIn_WEST,
         readReady;
  output readOut, writeOut;
  wire   N4718, n2888, n5327, n2886, n5326, n2889, n2883, n2887, n5323, n2569,
         n2567, n2566, n2578, n2638, n2624, n2617, n2577, n2544, n2541, n2540,
         n2537, n2535, n2703, n2692, n2691, n2689, n2511, n2507, n2731, n2574,
         n2499, n2496, n2493, n2770, n2768, n2764, n2754, n2748, n2746, n2739,
         n2486, n2484, n2482, n2480, n2802, n2834, n2833, n2832, n2829, n2825,
         n2814, n2811, n2807, n2806, n2457, n2455, n2453, n2570, n2565, n2573,
         n2568, n2564, n2563, n2575, n2882, n2881, n2879, n2610, n2609, n2608,
         n2607, n2606, n2605, n2604, n2603, n2602, n2601, n2600, n2599, n2598,
         n2597, n2596, n2595, n2594, n2593, n2592, n2591, n2590, n2589, n2588,
         n2587, n2586, n2585, n2584, n2583, n2582, n2581, n2580, n2579, n2561,
         n2560, n2559, n2557, n2556, n2555, n2554, n2552, n2551, n2550, n2549,
         n2642, n2640, n2639, n2637, n2635, n2634, n2633, n2631, n2628, n2627,
         n2626, n2625, n2623, n2620, n2618, n2616, n2615, n2614, n2612, n2611,
         n2870, n2869, n2868, n2867, n2866, n2865, n2674, n2672, n2671, n2670,
         n2669, n2668, n2667, n2666, n2665, n2664, n2662, n2661, n2660, n2657,
         n2656, n2655, n2654, n2653, n2652, n2651, n2650, n2649, n2648, n2647,
         n2646, n2645, n2644, n2576, n2534, n2533, n2532, n2531, n2530, n2529,
         n2528, n2527, n2526, n2525, n2524, n2523, n2522, n2521, n2860, n2859,
         n2706, n2705, n2700, n2698, n2696, n2695, n2694, n2690, n2687, n2686,
         n2685, n2684, n2677, n2675, n2736, n2734, n2733, n2725, n2723, n2720,
         n2718, n2715, n2713, n2504, n2498, n2497, n2494, n2850,
         \requesterAddressbuffer[2][2] , n2849, \requesterAddressbuffer[2][3] ,
         n2847, \requesterAddressbuffer[2][5] , n2769, n2760, n2743, n2492,
         n2491, n2489, n2488, n2487, n2485, n2483, n2481, n2846, n2845, n2844,
         n2843, n2842, n2841, n2801, n2799, n2798, n2796, n2795, n2793, n2791,
         n2790, n2789, n2788, n2787, n2786, n2785, n2784, n2781, n2779, n2778,
         n2777, n2776, n2774, n2773, n2772, n2771, n2572, n2478, n2477, n2476,
         n2475, n2474, n2473, n2472, n2471, n2470, n2469, n2468, n2467, n2466,
         n2465, n2840, \requesterAddressbuffer[0][0] , n2839,
         \requesterAddressbuffer[0][1] , n2838, \requesterAddressbuffer[0][2] ,
         n2836, \requesterAddressbuffer[0][4] , n2571, n2464, n2460, n2458,
         n2454, n2451, n2880, n2878, n2877, n2562, n2558, n2553, n2876,
         \requesterAddressbuffer[6][0] , n2875, \requesterAddressbuffer[6][1] ,
         n2874, \requesterAddressbuffer[6][2] , n2873,
         \requesterAddressbuffer[6][3] , n2872, \requesterAddressbuffer[6][4] ,
         n2871, \requesterAddressbuffer[6][5] , n2641, n2636, n2632, n2630,
         n2629, n2622, n2621, n2619, n2613, n2548, n2547, n2546, n2545, n2543,
         n2542, n2539, n2538, n2536, n2673, n2663, n2659, n2658, n2643, n2864,
         n2863, n2862, n2861, n2704, n2702, n2701, n2699, n2697, n2693, n2688,
         n2683, n2682, n2681, n2680, n2679, n2678, n2676, n2520, n2519, n2518,
         n2517, n2516, n2515, n2514, n2513, n2512, n2510, n2509, n2508, n2858,
         \requesterAddressbuffer[3][0] , n2857, \requesterAddressbuffer[3][1] ,
         n2856, \requesterAddressbuffer[3][2] , n2855,
         \requesterAddressbuffer[3][3] , n2854, \requesterAddressbuffer[3][4] ,
         n2853, \requesterAddressbuffer[3][5] , n2738, n2737, n2735, n2732,
         n2730, n2729, n2728, n2727, n2726, n2724, n2722, n2721, n2719, n2717,
         n2716, n2714, n2712, n2711, n2710, n2709, n2708, n2707, n2506, n2505,
         n2503, n2502, n2501, n2500, n2495, n2852,
         \requesterAddressbuffer[2][0] , n2851, \requesterAddressbuffer[2][1] ,
         n2848, \requesterAddressbuffer[2][4] , n2767, n2766, n2765, n2763,
         n2762, n2761, n2759, n2758, n2757, n2756, n2755, n2753, n2752, n2751,
         n2750, n2749, n2747, n2745, n2744, n2742, n2741, n2740, n2490, n2479,
         n2800, n2797, n2794, n2792, n2783, n2782, n2780, n2775, n2837,
         \requesterAddressbuffer[0][3] , n2835, \requesterAddressbuffer[0][5] ,
         n2831, n2830, n2828, n2827, n2826, n2824, n2823, n2822, n2821, n2820,
         n2819, n2818, n2817, n2816, n2815, n2813, n2812, n2810, n2809, n2808,
         n2805, n2804, n2803, n2463, n2462, n2461, n2459, n2456, n2452, n2885,
         n2449, n2434, n2431, n2450, n2448, n2447, n2446, n2445, n2444, n2443,
         n2442, n2441, n2440, n2439, n2438, n2437, n2436, n2435, n2433, n2432,
         n2430, n2429, n2428, n2427, n2426, n2425, n2424, n2423, n2422, n2421,
         n2420, n2419, n2418, n2417, n2416, n2415, n2414, n2413, n2412, n2411,
         n2410, n2409, n2408, n2407, n2406, n2405, n2404, n2403, n2402, n2401,
         n2400, n2399, n2398, n2397, n2884, n496, n497, n498, n499, n500, n502,
         n504, n506, n510, n513, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n538, n539, n540, n542, n547, n549, n550, n552, n553, n558,
         n583, n585, n586, n587, n615, n616, n617, n618, n619, n620, n621,
         n625, n626, n627, n709, n710, n713, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n728, n730, n731, n744, n778, n825, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n956, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1545, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1818, n1819, n1820,
         n1821, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n501, n503, n505, n507, n508, n509, n511, n512, n514, n515, n516,
         n536, n537, n541, n543, n544, n545, n546, n548, n551, n554, n555,
         n556, n557, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n584, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n622,
         n623, n624, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n711, n712, n714, n715, n716,
         n717, n727, n729, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n886, n919, n936,
         n955, n957, n970, n986, n1402, n1531, n1544, n1546, n1585, n1653,
         n1654, n1669, n1728, n1817, n1822, n1894, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392;
  wire   [0:7] readOutbuffer;
  wire   [0:7] writeOutbuffer;

  DFFNSRX2TS \destinationAddressbuffer_reg[2][6]  ( .D(n2486), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2290) );
  DFFNSRX2TS \destinationAddressbuffer_reg[2][8]  ( .D(n2484), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2310) );
  DFFNSRX2TS \destinationAddressbuffer_reg[2][10]  ( .D(n2482), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n2324) );
  DFFNSRX2TS \destinationAddressbuffer_reg[2][12]  ( .D(n2480), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n2338) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][7]  ( .D(n2457), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2302) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][9]  ( .D(n2455), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2318) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][11]  ( .D(n2453), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n2332) );
  DFFNSRX2TS \destinationAddressbuffer_reg[2][7]  ( .D(n2485), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2297) );
  DFFNSRX2TS \destinationAddressbuffer_reg[2][9]  ( .D(n2483), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2313) );
  DFFNSRX2TS \destinationAddressbuffer_reg[2][11]  ( .D(n2481), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n2329) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][6]  ( .D(n2458), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2289) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][10]  ( .D(n2454), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n2323) );
  DFFNSRX2TS \destinationAddressbuffer_reg[2][13]  ( .D(n2479), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n2352) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][8]  ( .D(n2456), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2312) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][12]  ( .D(n2452), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n2344) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][7]  ( .D(n2499), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2298) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][10]  ( .D(n2496), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n2322) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][13]  ( .D(n2493), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n2348) );
  DFFNSRX2TS \destinationAddressbuffer_reg[5][6]  ( .D(n2528), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2295) );
  DFFNSRX2TS \destinationAddressbuffer_reg[5][7]  ( .D(n2527), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2301) );
  DFFNSRX2TS \destinationAddressbuffer_reg[5][8]  ( .D(n2526), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2307) );
  DFFNSRX2TS \destinationAddressbuffer_reg[5][9]  ( .D(n2525), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2317) );
  DFFNSRX2TS \destinationAddressbuffer_reg[5][10]  ( .D(n2524), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n2321) );
  DFFNSRX2TS \destinationAddressbuffer_reg[5][11]  ( .D(n2523), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n2331) );
  DFFNSRX2TS \destinationAddressbuffer_reg[5][12]  ( .D(n2522), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n2337) );
  DFFNSRX2TS \destinationAddressbuffer_reg[5][13]  ( .D(n2521), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n2347) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][8]  ( .D(n2498), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2305) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][9]  ( .D(n2497), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2319) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][12]  ( .D(n2494), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n2341) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][6]  ( .D(n2500), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2294) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][11]  ( .D(n2495), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n2334) );
  DFFNSRX2TS \destinationAddressbuffer_reg[6][7]  ( .D(n2541), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2300) );
  DFFNSRX2TS \destinationAddressbuffer_reg[6][8]  ( .D(n2540), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2306) );
  DFFNSRX2TS \destinationAddressbuffer_reg[6][11]  ( .D(n2537), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n2330) );
  DFFNSRX2TS \destinationAddressbuffer_reg[6][13]  ( .D(n2535), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n2350) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][9]  ( .D(n2511), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2314) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][13]  ( .D(n2507), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n2346) );
  DFFNSRX2TS \destinationAddressbuffer_reg[6][6]  ( .D(n2542), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2296) );
  DFFNSRX2TS \destinationAddressbuffer_reg[6][9]  ( .D(n2539), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2320) );
  DFFNSRX2TS \destinationAddressbuffer_reg[6][10]  ( .D(n2538), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n2328) );
  DFFNSRX2TS \destinationAddressbuffer_reg[6][12]  ( .D(n2536), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n2340) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][6]  ( .D(n2514), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2292) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][7]  ( .D(n2513), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2304) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][8]  ( .D(n2512), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2308) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][10]  ( .D(n2510), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n2326) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][11]  ( .D(n2509), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n2336) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][12]  ( .D(n2508), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n2342) );
  DFFNSRX2TS \dataoutbuffer_reg[4][3]  ( .D(n2703), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2932) );
  DFFNSRX2TS \dataoutbuffer_reg[4][14]  ( .D(n2692), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3031) );
  DFFNSRX2TS \dataoutbuffer_reg[4][15]  ( .D(n2691), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3040) );
  DFFNSRX2TS \dataoutbuffer_reg[4][17]  ( .D(n2689), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3058) );
  DFFNSRX2TS \dataoutbuffer_reg[4][0]  ( .D(n2706), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2908) );
  DFFNSRX2TS \dataoutbuffer_reg[4][1]  ( .D(n2705), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2919) );
  DFFNSRX2TS \dataoutbuffer_reg[4][6]  ( .D(n2700), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2960) );
  DFFNSRX2TS \dataoutbuffer_reg[4][8]  ( .D(n2698), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2982) );
  DFFNSRX2TS \dataoutbuffer_reg[4][10]  ( .D(n2696), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n2998) );
  DFFNSRX2TS \dataoutbuffer_reg[4][11]  ( .D(n2695), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3005) );
  DFFNSRX2TS \dataoutbuffer_reg[4][12]  ( .D(n2694), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3016) );
  DFFNSRX2TS \dataoutbuffer_reg[4][16]  ( .D(n2690), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3054) );
  DFFNSRX2TS \dataoutbuffer_reg[4][19]  ( .D(n2687), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3081) );
  DFFNSRX2TS \dataoutbuffer_reg[4][20]  ( .D(n2686), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3086) );
  DFFNSRX2TS \dataoutbuffer_reg[4][21]  ( .D(n2685), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3095) );
  DFFNSRX2TS \dataoutbuffer_reg[4][22]  ( .D(n2684), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3106) );
  DFFNSRX2TS \dataoutbuffer_reg[4][29]  ( .D(n2677), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3165) );
  DFFNSRX2TS \dataoutbuffer_reg[4][31]  ( .D(n2675), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3189) );
  DFFNSRX2TS \dataoutbuffer_reg[4][2]  ( .D(n2704), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2927) );
  DFFNSRX2TS \dataoutbuffer_reg[4][4]  ( .D(n2702), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2943) );
  DFFNSRX2TS \dataoutbuffer_reg[4][5]  ( .D(n2701), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2954) );
  DFFNSRX2TS \dataoutbuffer_reg[4][7]  ( .D(n2699), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2970) );
  DFFNSRX2TS \dataoutbuffer_reg[4][9]  ( .D(n2697), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2988) );
  DFFNSRX2TS \dataoutbuffer_reg[4][13]  ( .D(n2693), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3028) );
  DFFNSRX2TS \dataoutbuffer_reg[4][18]  ( .D(n2688), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3073) );
  DFFNSRX2TS \dataoutbuffer_reg[4][23]  ( .D(n2683), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3116) );
  DFFNSRX2TS \dataoutbuffer_reg[4][24]  ( .D(n2682), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3127) );
  DFFNSRX2TS \dataoutbuffer_reg[4][25]  ( .D(n2681), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3132) );
  DFFNSRX2TS \dataoutbuffer_reg[4][26]  ( .D(n2680), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3145) );
  DFFNSRX2TS \dataoutbuffer_reg[4][27]  ( .D(n2679), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3152) );
  DFFNSRX2TS \dataoutbuffer_reg[4][28]  ( .D(n2678), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3163) );
  DFFNSRX2TS \dataoutbuffer_reg[4][30]  ( .D(n2676), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3181) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][0]  ( .D(n2520), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2360) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][1]  ( .D(n2519), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2365) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][2]  ( .D(n2518), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2378) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][3]  ( .D(n2517), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2383) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][4]  ( .D(n2516), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2392) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][5]  ( .D(n2515), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2896) );
  DFFNSRX2TS \dataoutbuffer_reg[5][2]  ( .D(n2672), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2926) );
  DFFNSRX2TS \dataoutbuffer_reg[5][3]  ( .D(n2671), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2931) );
  DFFNSRX2TS \dataoutbuffer_reg[5][4]  ( .D(n2670), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2942) );
  DFFNSRX2TS \dataoutbuffer_reg[5][5]  ( .D(n2669), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2949) );
  DFFNSRX2TS \dataoutbuffer_reg[5][6]  ( .D(n2668), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2962) );
  DFFNSRX2TS \dataoutbuffer_reg[5][7]  ( .D(n2667), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2969) );
  DFFNSRX2TS \dataoutbuffer_reg[5][8]  ( .D(n2666), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2978) );
  DFFNSRX2TS \dataoutbuffer_reg[5][9]  ( .D(n2665), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2989) );
  DFFNSRX2TS \dataoutbuffer_reg[5][10]  ( .D(n2664), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3000) );
  DFFNSRX2TS \dataoutbuffer_reg[5][12]  ( .D(n2662), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3014) );
  DFFNSRX2TS \dataoutbuffer_reg[5][13]  ( .D(n2661), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3023) );
  DFFNSRX2TS \dataoutbuffer_reg[5][14]  ( .D(n2660), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3036) );
  DFFNSRX2TS \dataoutbuffer_reg[5][17]  ( .D(n2657), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3059) );
  DFFNSRX2TS \dataoutbuffer_reg[5][18]  ( .D(n2656), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3070) );
  DFFNSRX2TS \dataoutbuffer_reg[5][19]  ( .D(n2655), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3077) );
  DFFNSRX2TS \dataoutbuffer_reg[5][20]  ( .D(n2654), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3090) );
  DFFNSRX2TS \dataoutbuffer_reg[5][21]  ( .D(n2653), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3097) );
  DFFNSRX2TS \dataoutbuffer_reg[5][22]  ( .D(n2652), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3104) );
  DFFNSRX2TS \dataoutbuffer_reg[5][23]  ( .D(n2651), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3115) );
  DFFNSRX2TS \dataoutbuffer_reg[5][24]  ( .D(n2650), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3122) );
  DFFNSRX2TS \dataoutbuffer_reg[5][25]  ( .D(n2649), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3129) );
  DFFNSRX2TS \dataoutbuffer_reg[5][26]  ( .D(n2648), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3144) );
  DFFNSRX2TS \dataoutbuffer_reg[5][27]  ( .D(n2647), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3153) );
  DFFNSRX2TS \dataoutbuffer_reg[5][28]  ( .D(n2646), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3156) );
  DFFNSRX2TS \dataoutbuffer_reg[5][29]  ( .D(n2645), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3167) );
  DFFNSRX2TS \dataoutbuffer_reg[5][30]  ( .D(n2644), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3178) );
  DFFNSRX2TS \destinationAddressbuffer_reg[5][0]  ( .D(n2534), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2357) );
  DFFNSRX2TS \destinationAddressbuffer_reg[5][1]  ( .D(n2533), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2364) );
  DFFNSRX2TS \destinationAddressbuffer_reg[5][2]  ( .D(n2532), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2373) );
  DFFNSRX2TS \destinationAddressbuffer_reg[5][3]  ( .D(n2531), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2382) );
  DFFNSRX2TS \destinationAddressbuffer_reg[5][4]  ( .D(n2530), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2391) );
  DFFNSRX2TS \destinationAddressbuffer_reg[5][5]  ( .D(n2529), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2893) );
  DFFNSRX2TS \dataoutbuffer_reg[5][1]  ( .D(n2673), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2916) );
  DFFNSRX2TS \dataoutbuffer_reg[5][11]  ( .D(n2663), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3008) );
  DFFNSRX2TS \dataoutbuffer_reg[5][15]  ( .D(n2659), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3046) );
  DFFNSRX2TS \dataoutbuffer_reg[5][16]  ( .D(n2658), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3051) );
  DFFNSRX2TS \dataoutbuffer_reg[5][31]  ( .D(n2643), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3186) );
  DFFNSRX2TS \requesterAddressbuffer_reg[2][2]  ( .D(n2850), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][2] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[2][3]  ( .D(n2849), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][3] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[2][5]  ( .D(n2847), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][5] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[0][0]  ( .D(n2840), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][0] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[0][1]  ( .D(n2839), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][1] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[0][2]  ( .D(n2838), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][2] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[0][4]  ( .D(n2836), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][4] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[2][0]  ( .D(n2852), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][0] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[2][1]  ( .D(n2851), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][1] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[2][4]  ( .D(n2848), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][4] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[0][3]  ( .D(n2837), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][3] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[0][5]  ( .D(n2835), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][5] ) );
  DFFNSRX2TS \readOutbuffer_reg[3]  ( .D(n2566), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[3]) );
  DFFNSRX2TS \readOutbuffer_reg[6]  ( .D(n2569), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n28) );
  DFFNSRX2TS \readOutbuffer_reg[5]  ( .D(n2568), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n29) );
  DFFNSRX2TS \readOutbuffer_reg[1]  ( .D(n2564), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n20) );
  DFFNSRX2TS \requesterAddressbuffer_reg[5][0]  ( .D(n2870), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n27) );
  DFFNSRX2TS \requesterAddressbuffer_reg[5][1]  ( .D(n2869), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n25) );
  DFFNSRX2TS \requesterAddressbuffer_reg[5][2]  ( .D(n2868), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n24) );
  DFFNSRX2TS \requesterAddressbuffer_reg[5][3]  ( .D(n2867), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n26) );
  DFFNSRX2TS \requesterAddressbuffer_reg[5][4]  ( .D(n2866), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n23) );
  DFFNSRX2TS \requesterAddressbuffer_reg[5][5]  ( .D(n2865), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n22) );
  DFFNSRX2TS \writeOutbuffer_reg[5]  ( .D(n2576), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n21) );
  DFFNSRX2TS \requesterAddressbuffer_reg[4][4]  ( .D(n2860), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n31) );
  DFFNSRX2TS \requesterAddressbuffer_reg[4][5]  ( .D(n2859), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n30) );
  DFFNSRX2TS \requesterAddressbuffer_reg[4][0]  ( .D(n2864), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n35) );
  DFFNSRX2TS \requesterAddressbuffer_reg[4][1]  ( .D(n2863), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n33) );
  DFFNSRX2TS \requesterAddressbuffer_reg[4][2]  ( .D(n2862), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n32) );
  DFFNSRX2TS \requesterAddressbuffer_reg[4][3]  ( .D(n2861), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n34) );
  DFFNSRX2TS \writeOutbuffer_reg[2]  ( .D(n2573), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[2]), .QN(n156) );
  DFFNSRX2TS \dataoutbuffer_reg[3][7]  ( .D(n2731), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n111), .QN(n2968) );
  DFFNSRX2TS \dataoutbuffer_reg[2][0]  ( .D(n2770), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n149), .QN(n2909) );
  DFFNSRX2TS \dataoutbuffer_reg[2][2]  ( .D(n2768), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n148), .QN(n2925) );
  DFFNSRX2TS \dataoutbuffer_reg[2][6]  ( .D(n2764), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n147), .QN(n2959) );
  DFFNSRX2TS \dataoutbuffer_reg[2][16]  ( .D(n2754), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n146), .QN(n3049) );
  DFFNSRX2TS \dataoutbuffer_reg[2][22]  ( .D(n2748), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n145), .QN(n3103) );
  DFFNSRX2TS \dataoutbuffer_reg[2][24]  ( .D(n2746), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n144), .QN(n3121) );
  DFFNSRX2TS \dataoutbuffer_reg[2][31]  ( .D(n2739), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n143), .QN(n3184) );
  DFFNSRX2TS \dataoutbuffer_reg[0][0]  ( .D(n2834), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n110), .QN(n2907) );
  DFFNSRX2TS \dataoutbuffer_reg[0][1]  ( .D(n2833), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n109), .QN(n2914) );
  DFFNSRX2TS \dataoutbuffer_reg[0][2]  ( .D(n2832), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n108), .QN(n2923) );
  DFFNSRX2TS \dataoutbuffer_reg[0][5]  ( .D(n2829), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n107), .QN(n2950) );
  DFFNSRX2TS \dataoutbuffer_reg[0][9]  ( .D(n2825), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n106), .QN(n2986) );
  DFFNSRX2TS \dataoutbuffer_reg[0][20]  ( .D(n2814), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n105), .QN(n3085) );
  DFFNSRX2TS \dataoutbuffer_reg[0][23]  ( .D(n2811), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n104), .QN(n3112) );
  DFFNSRX2TS \dataoutbuffer_reg[0][27]  ( .D(n2807), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n103), .QN(n3148) );
  DFFNSRX2TS \dataoutbuffer_reg[0][28]  ( .D(n2806), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n102), .QN(n3157) );
  DFFNSRX2TS \dataoutbuffer_reg[3][2]  ( .D(n2736), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n101), .QN(n2924) );
  DFFNSRX2TS \dataoutbuffer_reg[3][4]  ( .D(n2734), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n100), .QN(n2944) );
  DFFNSRX2TS \dataoutbuffer_reg[3][5]  ( .D(n2733), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n99), .QN(n2951) );
  DFFNSRX2TS \dataoutbuffer_reg[3][13]  ( .D(n2725), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n98), .QN(n3025) );
  DFFNSRX2TS \dataoutbuffer_reg[3][15]  ( .D(n2723), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n97), .QN(n3043) );
  DFFNSRX2TS \dataoutbuffer_reg[3][18]  ( .D(n2720), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n96), .QN(n3068) );
  DFFNSRX2TS \dataoutbuffer_reg[3][20]  ( .D(n2718), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n95), .QN(n3084) );
  DFFNSRX2TS \dataoutbuffer_reg[3][23]  ( .D(n2715), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n94), .QN(n3111) );
  DFFNSRX2TS \dataoutbuffer_reg[3][25]  ( .D(n2713), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n93), .QN(n3135) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][2]  ( .D(n2504), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n92), .QN(n2377) );
  DFFNSRX2TS \dataoutbuffer_reg[2][1]  ( .D(n2769), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n142), .QN(n2913) );
  DFFNSRX2TS \dataoutbuffer_reg[2][10]  ( .D(n2760), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n141), .QN(n2996) );
  DFFNSRX2TS \dataoutbuffer_reg[2][27]  ( .D(n2743), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n140), .QN(n3147) );
  DFFNSRX2TS \destinationAddressbuffer_reg[2][0]  ( .D(n2492), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n139), .QN(n2359) );
  DFFNSRX2TS \destinationAddressbuffer_reg[2][1]  ( .D(n2491), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n138), .QN(n2366) );
  DFFNSRX2TS \destinationAddressbuffer_reg[2][3]  ( .D(n2489), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n137), .QN(n2380) );
  DFFNSRX2TS \destinationAddressbuffer_reg[2][4]  ( .D(n2488), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n136), .QN(n2389) );
  DFFNSRX2TS \destinationAddressbuffer_reg[2][5]  ( .D(n2487), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n135), .QN(n2895) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][0]  ( .D(n2464), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n91), .QN(n2355) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][4]  ( .D(n2460), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n90), .QN(n2393) );
  DFFNSRX2TS \dataoutbuffer_reg[3][0]  ( .D(n2738), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n89), .QN(n2911) );
  DFFNSRX2TS \dataoutbuffer_reg[3][1]  ( .D(n2737), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n88), .QN(n2920) );
  DFFNSRX2TS \dataoutbuffer_reg[3][3]  ( .D(n2735), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n87), .QN(n2934) );
  DFFNSRX2TS \dataoutbuffer_reg[3][6]  ( .D(n2732), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n86), .QN(n2961) );
  DFFNSRX2TS \dataoutbuffer_reg[3][8]  ( .D(n2730), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n85), .QN(n2983) );
  DFFNSRX2TS \dataoutbuffer_reg[3][9]  ( .D(n2729), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n84), .QN(n2990) );
  DFFNSRX2TS \dataoutbuffer_reg[3][10]  ( .D(n2728), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n83), .QN(n2999) );
  DFFNSRX2TS \dataoutbuffer_reg[3][11]  ( .D(n2727), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n82), .QN(n3006) );
  DFFNSRX2TS \dataoutbuffer_reg[3][12]  ( .D(n2726), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n81), .QN(n3017) );
  DFFNSRX2TS \dataoutbuffer_reg[3][14]  ( .D(n2724), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n80), .QN(n3033) );
  DFFNSRX2TS \dataoutbuffer_reg[3][16]  ( .D(n2722), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n79), .QN(n3055) );
  DFFNSRX2TS \dataoutbuffer_reg[3][17]  ( .D(n2721), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n78), .QN(n3064) );
  DFFNSRX2TS \dataoutbuffer_reg[3][19]  ( .D(n2719), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n77), .QN(n3076) );
  DFFNSRX2TS \dataoutbuffer_reg[3][21]  ( .D(n2717), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n76), .QN(n3096) );
  DFFNSRX2TS \dataoutbuffer_reg[3][22]  ( .D(n2716), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n75), .QN(n3107) );
  DFFNSRX2TS \dataoutbuffer_reg[3][24]  ( .D(n2714), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n74), .QN(n3123) );
  DFFNSRX2TS \dataoutbuffer_reg[3][26]  ( .D(n2712), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n73), .QN(n3139) );
  DFFNSRX2TS \dataoutbuffer_reg[3][27]  ( .D(n2711), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n72), .QN(n3150) );
  DFFNSRX2TS \dataoutbuffer_reg[3][28]  ( .D(n2710), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n71), .QN(n3159) );
  DFFNSRX2TS \dataoutbuffer_reg[3][29]  ( .D(n2709), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n70), .QN(n3170) );
  DFFNSRX2TS \dataoutbuffer_reg[3][30]  ( .D(n2708), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n69), .QN(n3175) );
  DFFNSRX2TS \dataoutbuffer_reg[3][31]  ( .D(n2707), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n68), .QN(n3188) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][0]  ( .D(n2506), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n67), .QN(n2356) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][1]  ( .D(n2505), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n66), .QN(n2363) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][3]  ( .D(n2503), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n65), .QN(n2381) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][4]  ( .D(n2502), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n64), .QN(n2394) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][5]  ( .D(n2501), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n63), .QN(n2892) );
  DFFNSRX2TS \dataoutbuffer_reg[2][3]  ( .D(n2767), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n134), .QN(n2938) );
  DFFNSRX2TS \dataoutbuffer_reg[2][4]  ( .D(n2766), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n133), .QN(n2945) );
  DFFNSRX2TS \dataoutbuffer_reg[2][5]  ( .D(n2765), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n132), .QN(n2952) );
  DFFNSRX2TS \dataoutbuffer_reg[2][7]  ( .D(n2763), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n131), .QN(n2974) );
  DFFNSRX2TS \dataoutbuffer_reg[2][8]  ( .D(n2762), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n130), .QN(n2979) );
  DFFNSRX2TS \dataoutbuffer_reg[2][9]  ( .D(n2761), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n129), .QN(n2992) );
  DFFNSRX2TS \dataoutbuffer_reg[2][11]  ( .D(n2759), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n128), .QN(n3004) );
  DFFNSRX2TS \dataoutbuffer_reg[2][12]  ( .D(n2758), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n127), .QN(n3019) );
  DFFNSRX2TS \dataoutbuffer_reg[2][13]  ( .D(n2757), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n126), .QN(n3026) );
  DFFNSRX2TS \dataoutbuffer_reg[2][14]  ( .D(n2756), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n125), .QN(n3037) );
  DFFNSRX2TS \dataoutbuffer_reg[2][15]  ( .D(n2755), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n124), .QN(n3044) );
  DFFNSRX2TS \dataoutbuffer_reg[2][17]  ( .D(n2753), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n123), .QN(n3060) );
  DFFNSRX2TS \dataoutbuffer_reg[2][18]  ( .D(n2752), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n122), .QN(n3069) );
  DFFNSRX2TS \dataoutbuffer_reg[2][19]  ( .D(n2751), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n121), .QN(n3082) );
  DFFNSRX2TS \dataoutbuffer_reg[2][20]  ( .D(n2750), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n120), .QN(n3087) );
  DFFNSRX2TS \dataoutbuffer_reg[2][21]  ( .D(n2749), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n119), .QN(n3100) );
  DFFNSRX2TS \dataoutbuffer_reg[2][23]  ( .D(n2747), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n118), .QN(n3114) );
  DFFNSRX2TS \dataoutbuffer_reg[2][25]  ( .D(n2745), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n117), .QN(n3136) );
  DFFNSRX2TS \dataoutbuffer_reg[2][26]  ( .D(n2744), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n116), .QN(n3143) );
  DFFNSRX2TS \dataoutbuffer_reg[2][28]  ( .D(n2742), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n115), .QN(n3161) );
  DFFNSRX2TS \dataoutbuffer_reg[2][29]  ( .D(n2741), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n114), .QN(n3172) );
  DFFNSRX2TS \dataoutbuffer_reg[2][30]  ( .D(n2740), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n113), .QN(n3179) );
  DFFNSRX2TS \destinationAddressbuffer_reg[2][2]  ( .D(n2490), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n112), .QN(n2372) );
  DFFNSRX2TS \dataoutbuffer_reg[0][3]  ( .D(n2831), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n62), .QN(n2936) );
  DFFNSRX2TS \dataoutbuffer_reg[0][4]  ( .D(n2830), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n61), .QN(n2947) );
  DFFNSRX2TS \dataoutbuffer_reg[0][6]  ( .D(n2828), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n60), .QN(n2963) );
  DFFNSRX2TS \dataoutbuffer_reg[0][7]  ( .D(n2827), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n59), .QN(n2972) );
  DFFNSRX2TS \dataoutbuffer_reg[0][8]  ( .D(n2826), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n58), .QN(n2977) );
  DFFNSRX2TS \dataoutbuffer_reg[0][10]  ( .D(n2824), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n57), .QN(n2997) );
  DFFNSRX2TS \dataoutbuffer_reg[0][11]  ( .D(n2823), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n56), .QN(n3010) );
  DFFNSRX2TS \dataoutbuffer_reg[0][12]  ( .D(n2822), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n55), .QN(n3015) );
  DFFNSRX2TS \dataoutbuffer_reg[0][13]  ( .D(n2821), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n54), .QN(n3022) );
  DFFNSRX2TS \dataoutbuffer_reg[0][14]  ( .D(n2820), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n53), .QN(n3035) );
  DFFNSRX2TS \dataoutbuffer_reg[0][15]  ( .D(n2819), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n52), .QN(n3042) );
  DFFNSRX2TS \dataoutbuffer_reg[0][16]  ( .D(n2818), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n51), .QN(n3053) );
  DFFNSRX2TS \dataoutbuffer_reg[0][17]  ( .D(n2817), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n50), .QN(n3062) );
  DFFNSRX2TS \dataoutbuffer_reg[0][18]  ( .D(n2816), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n49), .QN(n3071) );
  DFFNSRX2TS \dataoutbuffer_reg[0][19]  ( .D(n2815), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n48), .QN(n3080) );
  DFFNSRX2TS \dataoutbuffer_reg[0][21]  ( .D(n2813), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n47), .QN(n3094) );
  DFFNSRX2TS \dataoutbuffer_reg[0][22]  ( .D(n2812), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n46), .QN(n3109) );
  DFFNSRX2TS \dataoutbuffer_reg[0][24]  ( .D(n2810), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n45), .QN(n3125) );
  DFFNSRX2TS \dataoutbuffer_reg[0][25]  ( .D(n2809), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n44), .QN(n3134) );
  DFFNSRX2TS \dataoutbuffer_reg[0][26]  ( .D(n2808), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n43), .QN(n3141) );
  DFFNSRX2TS \dataoutbuffer_reg[0][29]  ( .D(n2805), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n42), .QN(n3166) );
  DFFNSRX2TS \dataoutbuffer_reg[0][30]  ( .D(n2804), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n41), .QN(n3177) );
  DFFNSRX2TS \dataoutbuffer_reg[0][31]  ( .D(n2803), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n40), .QN(n3190) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][1]  ( .D(n2463), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n39), .QN(n2369) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][2]  ( .D(n2462), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n38), .QN(n2374) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][3]  ( .D(n2461), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n37), .QN(n2385) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][5]  ( .D(n2459), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n36), .QN(n2898) );
  DFFNSRX2TS \writeOutbuffer_reg[0]  ( .D(n2571), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[0]), .QN(n158) );
  DFFNSRX2TS \writeOutbuffer_reg[3]  ( .D(n2574), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[3]), .QN(n157) );
  DFFNSRX2TS \writeOutbuffer_reg[6]  ( .D(n2577), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[6]), .QN(n154) );
  DFFNSRX2TS \writeOutbuffer_reg[4]  ( .D(n2575), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[4]), .QN(n155) );
  DFFNSRX2TS \readOutbuffer_reg[7]  ( .D(n2570), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[7]), .QN(n152) );
  DFFNSRX2TS \readOutbuffer_reg[2]  ( .D(n2565), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[2]), .QN(n153) );
  DFFNSRX2TS \readOutbuffer_reg[4]  ( .D(n2567), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[4]), .QN(n151) );
  DFFNSRX2TS \read_reg_reg[0]  ( .D(n2889), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n9), .QN(n14) );
  DFFNSRX2TS full_reg_reg ( .D(N4718), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        n2285), .QN(n150) );
  DFFNSRX2TS writeOut_reg ( .D(n2449), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        writeOut), .QN(n2288) );
  DFFNSRX2TS \requesterAddressOut_reg[0]  ( .D(n2434), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[0]), .QN(n2284) );
  DFFNSRX2TS \requesterAddressOut_reg[3]  ( .D(n2431), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[3]), .QN(n2283) );
  DFFNSRX2TS readOut_reg ( .D(n2450), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        readOut), .QN(n2286) );
  DFFNSRX2TS \destinationAddressOut_reg[0]  ( .D(n2440), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[0]), .QN(n2361) );
  DFFNSRX2TS \destinationAddressOut_reg[1]  ( .D(n2439), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[1]), .QN(n2370) );
  DFFNSRX2TS \destinationAddressOut_reg[2]  ( .D(n2438), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[2]), .QN(n2379) );
  DFFNSRX2TS \destinationAddressOut_reg[3]  ( .D(n2437), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[3]), .QN(n2388) );
  DFFNSRX2TS \destinationAddressOut_reg[4]  ( .D(n2436), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[4]), .QN(n2890) );
  DFFNSRX2TS \destinationAddressOut_reg[5]  ( .D(n2435), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[5]), .QN(n2899) );
  DFFNSRX2TS \requesterAddressOut_reg[1]  ( .D(n2433), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[1]), .QN(n2900) );
  DFFNSRX2TS \requesterAddressOut_reg[2]  ( .D(n2432), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[2]), .QN(n2901) );
  DFFNSRX2TS \requesterAddressOut_reg[4]  ( .D(n2430), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[4]), .QN(n2902) );
  DFFNSRX2TS \requesterAddressOut_reg[5]  ( .D(n2429), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[5]), .QN(n2903) );
  DFFNSRX2TS \dataOut_reg[0]  ( .D(n2428), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[0]), .QN(n2912) );
  DFFNSRX2TS \dataOut_reg[1]  ( .D(n2427), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[1]), .QN(n2921) );
  DFFNSRX2TS \dataOut_reg[2]  ( .D(n2426), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[2]), .QN(n2930) );
  DFFNSRX2TS \dataOut_reg[3]  ( .D(n2425), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[3]), .QN(n2939) );
  DFFNSRX2TS \dataOut_reg[4]  ( .D(n2424), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[4]), .QN(n2948) );
  DFFNSRX2TS \dataOut_reg[5]  ( .D(n2423), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[5]), .QN(n2957) );
  DFFNSRX2TS \dataOut_reg[6]  ( .D(n2422), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[6]), .QN(n2966) );
  DFFNSRX2TS \dataOut_reg[7]  ( .D(n2421), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[7]), .QN(n2975) );
  DFFNSRX2TS \dataOut_reg[8]  ( .D(n2420), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[8]), .QN(n2984) );
  DFFNSRX2TS \dataOut_reg[9]  ( .D(n2419), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[9]), .QN(n2993) );
  DFFNSRX2TS \dataOut_reg[10]  ( .D(n2418), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[10]), .QN(n3002) );
  DFFNSRX2TS \dataOut_reg[11]  ( .D(n2417), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[11]), .QN(n3011) );
  DFFNSRX2TS \dataOut_reg[12]  ( .D(n2416), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[12]), .QN(n3020) );
  DFFNSRX2TS \dataOut_reg[13]  ( .D(n2415), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[13]), .QN(n3029) );
  DFFNSRX2TS \dataOut_reg[14]  ( .D(n2414), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[14]), .QN(n3038) );
  DFFNSRX2TS \dataOut_reg[15]  ( .D(n2413), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[15]), .QN(n3047) );
  DFFNSRX2TS \dataOut_reg[16]  ( .D(n2412), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[16]), .QN(n3056) );
  DFFNSRX2TS \dataOut_reg[17]  ( .D(n2411), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[17]), .QN(n3065) );
  DFFNSRX2TS \dataOut_reg[18]  ( .D(n2410), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[18]), .QN(n3074) );
  DFFNSRX2TS \dataOut_reg[19]  ( .D(n2409), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[19]), .QN(n3083) );
  DFFNSRX2TS \dataOut_reg[20]  ( .D(n2408), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[20]), .QN(n3092) );
  DFFNSRX2TS \dataOut_reg[21]  ( .D(n2407), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[21]), .QN(n3101) );
  DFFNSRX2TS \dataOut_reg[22]  ( .D(n2406), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[22]), .QN(n3110) );
  DFFNSRX2TS \dataOut_reg[23]  ( .D(n2405), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[23]), .QN(n3119) );
  DFFNSRX2TS \dataOut_reg[24]  ( .D(n2404), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[24]), .QN(n3128) );
  DFFNSRX2TS \dataOut_reg[25]  ( .D(n2403), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[25]), .QN(n3137) );
  DFFNSRX2TS \dataOut_reg[26]  ( .D(n2402), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[26]), .QN(n3146) );
  DFFNSRX2TS \dataOut_reg[27]  ( .D(n2401), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[27]), .QN(n3155) );
  DFFNSRX2TS \dataOut_reg[28]  ( .D(n2400), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[28]), .QN(n3164) );
  DFFNSRX2TS \dataOut_reg[29]  ( .D(n2399), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[29]), .QN(n3173) );
  DFFNSRX2TS \dataOut_reg[30]  ( .D(n2398), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[30]), .QN(n3182) );
  DFFNSRX2TS \dataOut_reg[31]  ( .D(n2397), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[31]), .QN(n3191) );
  DFFNSRX2TS \destinationAddressOut_reg[6]  ( .D(n2448), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[6]) );
  DFFNSRX2TS \destinationAddressOut_reg[7]  ( .D(n2447), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[7]) );
  DFFNSRX2TS \destinationAddressOut_reg[8]  ( .D(n2446), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[8]) );
  DFFNSRX2TS \destinationAddressOut_reg[9]  ( .D(n2445), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[9]) );
  DFFNSRX2TS \destinationAddressOut_reg[10]  ( .D(n2444), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[10]) );
  DFFNSRX2TS \destinationAddressOut_reg[11]  ( .D(n2443), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[11]) );
  DFFNSRX2TS \destinationAddressOut_reg[12]  ( .D(n2442), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[12]) );
  DFFNSRX2TS \destinationAddressOut_reg[13]  ( .D(n2441), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[13]) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][13]  ( .D(n2549), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n2349) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][6]  ( .D(n2472), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2291) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][7]  ( .D(n2471), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2303) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][8]  ( .D(n2470), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2311) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][9]  ( .D(n2469), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2315) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][10]  ( .D(n2468), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n2327) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][11]  ( .D(n2467), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n2333) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][12]  ( .D(n2466), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n2343) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][4]  ( .D(n2558), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2396) );
  DFFNSRXLTS \dataoutbuffer_reg[1][0]  ( .D(n2802), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2905) );
  DFFNSRXLTS \dataoutbuffer_reg[7][0]  ( .D(n2610), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2910) );
  DFFNSRXLTS \dataoutbuffer_reg[7][1]  ( .D(n2609), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2915) );
  DFFNSRXLTS \dataoutbuffer_reg[7][2]  ( .D(n2608), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2928) );
  DFFNSRXLTS \dataoutbuffer_reg[7][3]  ( .D(n2607), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2933) );
  DFFNSRXLTS \dataoutbuffer_reg[7][4]  ( .D(n2606), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2946) );
  DFFNSRXLTS \dataoutbuffer_reg[7][5]  ( .D(n2605), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2955) );
  DFFNSRXLTS \dataoutbuffer_reg[7][6]  ( .D(n2604), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2958) );
  DFFNSRXLTS \dataoutbuffer_reg[7][7]  ( .D(n2603), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2973) );
  DFFNSRXLTS \dataoutbuffer_reg[7][8]  ( .D(n2602), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2980) );
  DFFNSRXLTS \dataoutbuffer_reg[7][9]  ( .D(n2601), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2985) );
  DFFNSRXLTS \dataoutbuffer_reg[7][10]  ( .D(n2600), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n2994) );
  DFFNSRXLTS \dataoutbuffer_reg[7][11]  ( .D(n2599), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3007) );
  DFFNSRXLTS \dataoutbuffer_reg[7][12]  ( .D(n2598), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3018) );
  DFFNSRXLTS \dataoutbuffer_reg[7][13]  ( .D(n2597), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3027) );
  DFFNSRXLTS \dataoutbuffer_reg[7][14]  ( .D(n2596), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3030) );
  DFFNSRXLTS \dataoutbuffer_reg[7][15]  ( .D(n2595), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3045) );
  DFFNSRXLTS \dataoutbuffer_reg[7][16]  ( .D(n2594), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3050) );
  DFFNSRXLTS \dataoutbuffer_reg[7][17]  ( .D(n2593), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3061) );
  DFFNSRXLTS \dataoutbuffer_reg[7][18]  ( .D(n2592), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3072) );
  DFFNSRXLTS \dataoutbuffer_reg[7][19]  ( .D(n2591), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3075) );
  DFFNSRXLTS \dataoutbuffer_reg[7][20]  ( .D(n2590), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3088) );
  DFFNSRXLTS \dataoutbuffer_reg[7][21]  ( .D(n2589), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3093) );
  DFFNSRXLTS \dataoutbuffer_reg[7][22]  ( .D(n2588), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3108) );
  DFFNSRXLTS \dataoutbuffer_reg[7][23]  ( .D(n2587), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3113) );
  DFFNSRXLTS \dataoutbuffer_reg[7][24]  ( .D(n2586), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3124) );
  DFFNSRXLTS \dataoutbuffer_reg[7][25]  ( .D(n2585), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3133) );
  DFFNSRXLTS \dataoutbuffer_reg[7][26]  ( .D(n2584), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3142) );
  DFFNSRXLTS \dataoutbuffer_reg[7][27]  ( .D(n2583), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3149) );
  DFFNSRXLTS \dataoutbuffer_reg[7][28]  ( .D(n2582), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3158) );
  DFFNSRXLTS \dataoutbuffer_reg[7][29]  ( .D(n2581), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3171) );
  DFFNSRXLTS \dataoutbuffer_reg[7][30]  ( .D(n2580), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3180) );
  DFFNSRXLTS \dataoutbuffer_reg[7][31]  ( .D(n2579), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3185) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][1]  ( .D(n2561), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2368) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][2]  ( .D(n2560), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2375) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][3]  ( .D(n2559), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2386) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][5]  ( .D(n2557), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2891) );
  DFFNSRXLTS \dataoutbuffer_reg[1][1]  ( .D(n2801), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2917) );
  DFFNSRXLTS \dataoutbuffer_reg[1][3]  ( .D(n2799), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2935) );
  DFFNSRXLTS \dataoutbuffer_reg[1][4]  ( .D(n2798), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2940) );
  DFFNSRXLTS \dataoutbuffer_reg[1][6]  ( .D(n2796), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2964) );
  DFFNSRXLTS \dataoutbuffer_reg[1][7]  ( .D(n2795), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2967) );
  DFFNSRXLTS \dataoutbuffer_reg[1][9]  ( .D(n2793), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2991) );
  DFFNSRXLTS \dataoutbuffer_reg[1][11]  ( .D(n2791), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3009) );
  DFFNSRXLTS \dataoutbuffer_reg[1][12]  ( .D(n2790), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3012) );
  DFFNSRXLTS \dataoutbuffer_reg[1][13]  ( .D(n2789), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3021) );
  DFFNSRXLTS \dataoutbuffer_reg[1][14]  ( .D(n2788), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3034) );
  DFFNSRXLTS \dataoutbuffer_reg[1][15]  ( .D(n2787), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3041) );
  DFFNSRXLTS \dataoutbuffer_reg[1][16]  ( .D(n2786), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3048) );
  DFFNSRXLTS \dataoutbuffer_reg[1][17]  ( .D(n2785), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3063) );
  DFFNSRXLTS \dataoutbuffer_reg[1][18]  ( .D(n2784), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3066) );
  DFFNSRXLTS \dataoutbuffer_reg[1][21]  ( .D(n2781), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3099) );
  DFFNSRXLTS \dataoutbuffer_reg[1][23]  ( .D(n2779), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3117) );
  DFFNSRXLTS \dataoutbuffer_reg[1][24]  ( .D(n2778), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3126) );
  DFFNSRXLTS \dataoutbuffer_reg[1][25]  ( .D(n2777), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3131) );
  DFFNSRXLTS \dataoutbuffer_reg[1][26]  ( .D(n2776), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3138) );
  DFFNSRXLTS \dataoutbuffer_reg[1][28]  ( .D(n2774), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3162) );
  DFFNSRXLTS \dataoutbuffer_reg[1][29]  ( .D(n2773), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3169) );
  DFFNSRXLTS \dataoutbuffer_reg[1][30]  ( .D(n2772), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3174) );
  DFFNSRXLTS \dataoutbuffer_reg[1][31]  ( .D(n2771), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3183) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][0]  ( .D(n2478), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2353) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][1]  ( .D(n2477), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2362) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][2]  ( .D(n2476), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2371) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][3]  ( .D(n2475), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2384) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][5]  ( .D(n2473), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2897) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][0]  ( .D(n2562), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2354) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][0]  ( .D(n2548), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2358) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][1]  ( .D(n2547), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2367) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][2]  ( .D(n2546), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2376) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][3]  ( .D(n2545), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2387) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][5]  ( .D(n2543), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2894) );
  DFFNSRXLTS \dataoutbuffer_reg[1][2]  ( .D(n2800), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2929) );
  DFFNSRXLTS \dataoutbuffer_reg[1][5]  ( .D(n2797), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2956) );
  DFFNSRXLTS \dataoutbuffer_reg[1][8]  ( .D(n2794), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2981) );
  DFFNSRXLTS \dataoutbuffer_reg[1][10]  ( .D(n2792), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n2995) );
  DFFNSRXLTS \dataoutbuffer_reg[1][19]  ( .D(n2783), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3078) );
  DFFNSRXLTS \dataoutbuffer_reg[1][20]  ( .D(n2782), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3089) );
  DFFNSRXLTS \dataoutbuffer_reg[1][22]  ( .D(n2780), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3105) );
  DFFNSRXLTS \dataoutbuffer_reg[1][27]  ( .D(n2775), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3154) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][4]  ( .D(n2544), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2390) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][10]  ( .D(n2552), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n593), .QN(n2325) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][4]  ( .D(n2474), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2395) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][0]  ( .D(n2858), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][0] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][1]  ( .D(n2857), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][1] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][2]  ( .D(n2856), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][2] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][3]  ( .D(n2855), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][3] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][5]  ( .D(n2853), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][5] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][4]  ( .D(n2854), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][4] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[6][1]  ( .D(n2875), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][1] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[6][2]  ( .D(n2874), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][2] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[6][3]  ( .D(n2873), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][3] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[6][4]  ( .D(n2872), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][4] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[6][5]  ( .D(n2871), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][5] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[6][0]  ( .D(n2876), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][0] ) );
  DFFNSRXLTS \writeOutbuffer_reg[7]  ( .D(n2578), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n558) );
  DFFNSRXLTS \requesterAddressbuffer_reg[7][0]  ( .D(n2882), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n585) );
  DFFNSRXLTS \requesterAddressbuffer_reg[7][1]  ( .D(n2881), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n586) );
  DFFNSRXLTS \requesterAddressbuffer_reg[7][3]  ( .D(n2879), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n587) );
  DFFNSRXLTS \requesterAddressbuffer_reg[7][2]  ( .D(n2880), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n625) );
  DFFNSRXLTS \requesterAddressbuffer_reg[7][4]  ( .D(n2878), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n626) );
  DFFNSRXLTS \requesterAddressbuffer_reg[7][5]  ( .D(n2877), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n627) );
  DFFNSRXLTS \readOutbuffer_reg[0]  ( .D(n2563), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n583) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][0]  ( .D(n2846), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n615) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][1]  ( .D(n2845), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n616) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][2]  ( .D(n2844), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n617) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][3]  ( .D(n2843), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n618) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][4]  ( .D(n2842), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n619) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][5]  ( .D(n2841), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n620) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][6]  ( .D(n2556), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2293) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][7]  ( .D(n2555), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2299) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][8]  ( .D(n2554), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2309) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][11]  ( .D(n2551), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n2335) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][9]  ( .D(n2553), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n2316) );
  DFFNSRXLTS \writeOutbuffer_reg[1]  ( .D(n2572), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[1]), .QN(n621) );
  DFFNSRX2TS \read_reg_reg[1]  ( .D(n2883), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n10), .QN(n459) );
  DFFNSRX2TS \read_reg_reg[2]  ( .D(n2884), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n8), .QN(n455) );
  DFFNSRXLTS \dataoutbuffer_reg[6][31]  ( .D(n2611), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3187) );
  DFFNSRXLTS \dataoutbuffer_reg[6][30]  ( .D(n2612), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3176) );
  DFFNSRXLTS \dataoutbuffer_reg[6][29]  ( .D(n2613), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3168) );
  DFFNSRXLTS \dataoutbuffer_reg[6][28]  ( .D(n2614), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3160) );
  DFFNSRXLTS \dataoutbuffer_reg[6][27]  ( .D(n2615), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3151) );
  DFFNSRXLTS \dataoutbuffer_reg[6][26]  ( .D(n2616), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3140) );
  DFFNSRXLTS \dataoutbuffer_reg[6][25]  ( .D(n2617), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3130) );
  DFFNSRXLTS \dataoutbuffer_reg[6][24]  ( .D(n2618), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3120) );
  DFFNSRXLTS \dataoutbuffer_reg[6][23]  ( .D(n2619), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3118) );
  DFFNSRXLTS \dataoutbuffer_reg[6][22]  ( .D(n2620), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3102) );
  DFFNSRXLTS \dataoutbuffer_reg[6][21]  ( .D(n2621), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3098) );
  DFFNSRXLTS \dataoutbuffer_reg[6][20]  ( .D(n2622), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3091) );
  DFFNSRXLTS \dataoutbuffer_reg[6][19]  ( .D(n2623), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3079) );
  DFFNSRXLTS \dataoutbuffer_reg[6][18]  ( .D(n2624), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3067) );
  DFFNSRXLTS \dataoutbuffer_reg[6][17]  ( .D(n2625), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3057) );
  DFFNSRXLTS \dataoutbuffer_reg[6][16]  ( .D(n2626), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3052) );
  DFFNSRXLTS \dataoutbuffer_reg[6][15]  ( .D(n2627), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3039) );
  DFFNSRXLTS \dataoutbuffer_reg[6][14]  ( .D(n2628), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3032) );
  DFFNSRXLTS \dataoutbuffer_reg[6][13]  ( .D(n2629), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3024) );
  DFFNSRXLTS \dataoutbuffer_reg[6][12]  ( .D(n2630), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3013) );
  DFFNSRXLTS \dataoutbuffer_reg[6][11]  ( .D(n2631), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3003) );
  DFFNSRXLTS \dataoutbuffer_reg[6][10]  ( .D(n2632), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n3001) );
  DFFNSRXLTS \dataoutbuffer_reg[6][9]  ( .D(n2633), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2987) );
  DFFNSRXLTS \dataoutbuffer_reg[6][8]  ( .D(n2634), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2976) );
  DFFNSRXLTS \dataoutbuffer_reg[6][7]  ( .D(n2635), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2971) );
  DFFNSRXLTS \dataoutbuffer_reg[6][6]  ( .D(n2636), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2965) );
  DFFNSRXLTS \dataoutbuffer_reg[6][5]  ( .D(n2637), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2953) );
  DFFNSRXLTS \dataoutbuffer_reg[6][4]  ( .D(n2638), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2941) );
  DFFNSRXLTS \dataoutbuffer_reg[6][3]  ( .D(n2639), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2937) );
  DFFNSRXLTS \dataoutbuffer_reg[6][2]  ( .D(n2640), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2922) );
  DFFNSRXLTS \dataoutbuffer_reg[6][1]  ( .D(n2641), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2918) );
  DFFNSRXLTS \dataoutbuffer_reg[6][0]  ( .D(n2642), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2906) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][12]  ( .D(n2550), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n2339) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][13]  ( .D(n2465), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n2351) );
  DFFNSRXLTS empty_reg_reg ( .D(n2885), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        n710), .QN(n2287) );
  DFFNSRXLTS \write_reg_reg[0]  ( .D(n2888), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n13), .QN(n5327) );
  DFFNSRXLTS \write_reg_reg[1]  ( .D(n2887), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n6), .QN(n5323) );
  DFFNSRXLTS \write_reg_reg[2]  ( .D(n2886), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n12), .QN(n5326) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][13]  ( .D(n2451), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n2345) );
  DFFNSRX1TS \dataoutbuffer_reg[5][0]  ( .D(n2674), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n2904) );
  NOR2X1TS U2 ( .A(n528), .B(n1630), .Y(n1553) );
  BUFX3TS U3 ( .A(n3525), .Y(n3520) );
  CLKAND2X2TS U4 ( .A(n435), .B(n1723), .Y(n18) );
  OAI22X2TS U5 ( .A0(n1589), .A1(n578), .B0(n243), .B1(n222), .Y(n1542) );
  AND3X2TS U6 ( .A(n1655), .B(n1727), .C(n525), .Y(n1591) );
  INVX1TS U7 ( .A(n1680), .Y(n456) );
  INVX1TS U8 ( .A(n1680), .Y(n525) );
  NAND3X1TS U9 ( .A(n1631), .B(n1680), .C(n460), .Y(n1568) );
  XOR2X4TS U10 ( .A(n1796), .B(n12), .Y(n1680) );
  AOI2BB1X2TS U11 ( .A0N(n534), .A1N(n1702), .B0(n1576), .Y(n1574) );
  OAI21X2TS U12 ( .A0(n1630), .A1(n1577), .B0(n1701), .Y(n1576) );
  XNOR2X2TS U13 ( .A(selectBit_NORTH), .B(selectBit_EAST), .Y(n2282) );
  NOR2BX1TS U14 ( .AN(n1774), .B(n825), .Y(n1631) );
  INVX1TS U15 ( .A(n1727), .Y(n460) );
  INVX3TS U16 ( .A(n1727), .Y(n524) );
  XOR2X4TS U17 ( .A(n1800), .B(n208), .Y(n1727) );
  INVX1TS U18 ( .A(n1535), .Y(n1) );
  CLKINVX2TS U19 ( .A(n1), .Y(n2) );
  AND3XLTS U20 ( .A(n1567), .B(n1596), .C(n1593), .Y(n992) );
  INVXLTS U21 ( .A(n1596), .Y(n520) );
  BUFX4TS U22 ( .A(n3423), .Y(n3421) );
  AOI21X1TS U23 ( .A0(n718), .A1(n595), .B0(n1773), .Y(n1803) );
  XOR2XLTS U24 ( .A(n1773), .B(n6), .Y(n16) );
  NOR2X2TS U25 ( .A(n718), .B(n595), .Y(n1773) );
  BUFX8TS U26 ( .A(n3310), .Y(n3309) );
  NAND3XLTS U27 ( .A(n524), .B(n1631), .C(n525), .Y(n1596) );
  OAI22X2TS U28 ( .A0(n1605), .A1(n577), .B0(n242), .B1(n542), .Y(n1547) );
  OA21X4TS U29 ( .A0(n160), .A1(n1702), .B0(n1601), .Y(n1605) );
  BUFX4TS U30 ( .A(n747), .Y(n746) );
  AO21X1TS U31 ( .A0(n463), .A1(n241), .B0(n591), .Y(n1550) );
  AOI21X1TS U32 ( .A0(n1628), .A1(n224), .B0(n588), .Y(n1564) );
  CLKBUFX2TS U33 ( .A(n3527), .Y(n3516) );
  CLKBUFX2TS U34 ( .A(n3556), .Y(n3550) );
  CLKBUFX2TS U35 ( .A(n3558), .Y(n3546) );
  CLKBUFX2TS U36 ( .A(n3555), .Y(n3551) );
  NOR2X1TS U37 ( .A(n1554), .B(n1553), .Y(n1556) );
  CLKBUFX2TS U38 ( .A(n3362), .Y(n3348) );
  CLKBUFX2TS U39 ( .A(n3357), .Y(n3355) );
  NOR2X1TS U40 ( .A(n720), .B(n318), .Y(n1798) );
  NAND2X1TS U41 ( .A(n531), .B(n5323), .Y(n1598) );
  XNOR2X1TS U42 ( .A(n317), .B(n1798), .Y(n1800) );
  AOI21X1TS U43 ( .A0(n220), .A1(n224), .B0(n584), .Y(n1571) );
  CLKBUFX2TS U44 ( .A(n3528), .Y(n3515) );
  CLKBUFX2TS U45 ( .A(n3555), .Y(n3552) );
  CLKBUFX2TS U46 ( .A(n3554), .Y(n3553) );
  CLKBUFX2TS U47 ( .A(n3527), .Y(n3517) );
  CLKBUFX2TS U48 ( .A(n829), .Y(n828) );
  CLKBUFX2TS U49 ( .A(n3528), .Y(n3514) );
  NAND2BX1TS U50 ( .AN(n1750), .B(n1729), .Y(n1577) );
  CLKBUFX2TS U51 ( .A(n3330), .Y(n3319) );
  CLKBUFX2TS U52 ( .A(n1564), .Y(n161) );
  NOR3X1TS U53 ( .A(n1561), .B(n1560), .C(n1563), .Y(n1562) );
  AOI21X1TS U54 ( .A0(n1580), .A1(n1726), .B0(n522), .Y(n1582) );
  CLKBUFX2TS U55 ( .A(n3329), .Y(n3325) );
  CLKBUFX2TS U56 ( .A(n748), .Y(n745) );
  AOI222XLTS U57 ( .A0(n4122), .A1(n3551), .B0(n198), .B1(n3531), .C0(n4278), 
        .C1(n3516), .Y(n1617) );
  AOI222XLTS U58 ( .A0(n4086), .A1(n3550), .B0(n468), .B1(n3539), .C0(n4242), 
        .C1(n3522), .Y(n1530) );
  AOI222XLTS U59 ( .A0(n4083), .A1(n3550), .B0(n470), .B1(n3543), .C0(n4239), 
        .C1(n3522), .Y(n1528) );
  AOI222XLTS U60 ( .A0(n4080), .A1(n3549), .B0(n472), .B1(n3542), .C0(n4236), 
        .C1(n3522), .Y(n1526) );
  AOI222XLTS U61 ( .A0(n4077), .A1(n3549), .B0(n474), .B1(n3540), .C0(n4233), 
        .C1(n3522), .Y(n1524) );
  AOI222XLTS U62 ( .A0(n4074), .A1(n3549), .B0(n476), .B1(n3542), .C0(n4230), 
        .C1(n3521), .Y(n1522) );
  AOI222XLTS U63 ( .A0(n4071), .A1(n3549), .B0(n478), .B1(n3540), .C0(n4227), 
        .C1(n3521), .Y(n1520) );
  AOI222XLTS U64 ( .A0(n4068), .A1(n3548), .B0(n479), .B1(n3532), .C0(n4224), 
        .C1(n3521), .Y(n1518) );
  AOI222XLTS U65 ( .A0(n4065), .A1(n3548), .B0(n482), .B1(n3532), .C0(n4221), 
        .C1(n3521), .Y(n1516) );
  AOI222XLTS U66 ( .A0(n4062), .A1(n3548), .B0(n484), .B1(n3532), .C0(n4218), 
        .C1(n3524), .Y(n1514) );
  AOI222XLTS U67 ( .A0(n4059), .A1(n3548), .B0(n486), .B1(n3532), .C0(n4215), 
        .C1(n3530), .Y(n1512) );
  AOI222XLTS U68 ( .A0(n4056), .A1(n3547), .B0(n488), .B1(n3533), .C0(n4212), 
        .C1(n3527), .Y(n1510) );
  AOI222XLTS U69 ( .A0(n4053), .A1(n3547), .B0(n490), .B1(n3533), .C0(n4209), 
        .C1(n891), .Y(n1508) );
  AOI222XLTS U70 ( .A0(n4050), .A1(n3547), .B0(n492), .B1(n3533), .C0(n4206), 
        .C1(n3523), .Y(n1506) );
  AOI222XLTS U71 ( .A0(n4047), .A1(n3557), .B0(n493), .B1(n3533), .C0(n4203), 
        .C1(n3526), .Y(n1504) );
  AOI222XLTS U72 ( .A0(n4044), .A1(n3554), .B0(n501), .B1(n3534), .C0(n4200), 
        .C1(n3528), .Y(n1502) );
  AOI222XLTS U73 ( .A0(n4041), .A1(n3561), .B0(n505), .B1(n3534), .C0(n4197), 
        .C1(n3524), .Y(n1500) );
  AOI222XLTS U74 ( .A0(n4029), .A1(n3557), .B0(n516), .B1(n3543), .C0(n4185), 
        .C1(n3520), .Y(n1492) );
  AOI222XLTS U75 ( .A0(n4026), .A1(n889), .B0(n537), .B1(n3541), .C0(n4182), 
        .C1(n3520), .Y(n1490) );
  AOI222XLTS U76 ( .A0(n4023), .A1(n3559), .B0(n543), .B1(n3541), .C0(n4179), 
        .C1(n3520), .Y(n1488) );
  AOI222XLTS U77 ( .A0(n4020), .A1(n3556), .B0(n545), .B1(n3535), .C0(n4176), 
        .C1(n3520), .Y(n1486) );
  AOI222XLTS U78 ( .A0(n4017), .A1(n3558), .B0(n548), .B1(n3535), .C0(n4173), 
        .C1(n3519), .Y(n1484) );
  AOI222XLTS U79 ( .A0(n4014), .A1(n3558), .B0(n554), .B1(n3535), .C0(n4170), 
        .C1(n3519), .Y(n1482) );
  AOI222XLTS U80 ( .A0(n4011), .A1(n3559), .B0(n556), .B1(n3535), .C0(n4167), 
        .C1(n3519), .Y(n1480) );
  AOI222XLTS U81 ( .A0(n4008), .A1(n3560), .B0(n559), .B1(n3536), .C0(n4164), 
        .C1(n3519), .Y(n1478) );
  AOI222XLTS U82 ( .A0(n4005), .A1(n3554), .B0(n560), .B1(n3536), .C0(n4161), 
        .C1(n3518), .Y(n1476) );
  AOI222XLTS U83 ( .A0(n4002), .A1(n3556), .B0(n563), .B1(n3536), .C0(n4158), 
        .C1(n3518), .Y(n1474) );
  AOI222XLTS U84 ( .A0(n3999), .A1(n3546), .B0(n565), .B1(n3536), .C0(n4155), 
        .C1(n3518), .Y(n1472) );
  AOI222XLTS U85 ( .A0(n3996), .A1(n3546), .B0(n567), .B1(n3537), .C0(n4152), 
        .C1(n3518), .Y(n1470) );
  OAI221XLTS U86 ( .A0(readIn_SOUTH), .A1(n533), .B0(n3834), .B1(n1555), .C0(
        n1556), .Y(n1551) );
  AOI222XLTS U87 ( .A0(n3348), .A1(n4101), .B0(n3341), .B1(n196), .C0(n3320), 
        .C1(n3945), .Y(n950) );
  AOI222XLTS U88 ( .A0(n4085), .A1(n922), .B0(n467), .B1(n923), .C0(n4242), 
        .C1(n250), .Y(n1401) );
  AOI222XLTS U89 ( .A0(n4040), .A1(n3419), .B0(n503), .B1(n3400), .C0(n4197), 
        .C1(n263), .Y(n1371) );
  AOI222XLTS U90 ( .A0(n4082), .A1(n922), .B0(n470), .B1(n3400), .C0(n4239), 
        .C1(n250), .Y(n1399) );
  AOI222XLTS U91 ( .A0(n4079), .A1(n3426), .B0(n472), .B1(n3409), .C0(n4236), 
        .C1(n277), .Y(n1397) );
  AOI222XLTS U92 ( .A0(n4073), .A1(n3427), .B0(n476), .B1(n3400), .C0(n4230), 
        .C1(n249), .Y(n1393) );
  AOI222XLTS U93 ( .A0(n4067), .A1(n3430), .B0(n480), .B1(n923), .C0(n4224), 
        .C1(n277), .Y(n1389) );
  AOI222XLTS U94 ( .A0(n4064), .A1(n3427), .B0(n482), .B1(n3413), .C0(n4221), 
        .C1(n263), .Y(n1387) );
  AOI222XLTS U95 ( .A0(n4055), .A1(n3425), .B0(n488), .B1(n3412), .C0(n4212), 
        .C1(n277), .Y(n1381) );
  AOI222XLTS U96 ( .A0(n4052), .A1(n3424), .B0(n490), .B1(n3412), .C0(n4209), 
        .C1(n263), .Y(n1379) );
  AOI222XLTS U97 ( .A0(n4046), .A1(n3419), .B0(n494), .B1(n3411), .C0(n4203), 
        .C1(n250), .Y(n1375) );
  AOI222XLTS U98 ( .A0(n4043), .A1(n3419), .B0(n495), .B1(n3401), .C0(n4200), 
        .C1(n277), .Y(n1373) );
  AOI222XLTS U99 ( .A0(n4028), .A1(n3418), .B0(n516), .B1(n3401), .C0(n4185), 
        .C1(n249), .Y(n1363) );
  AOI222XLTS U100 ( .A0(n4019), .A1(n3425), .B0(n545), .B1(n3402), .C0(n4176), 
        .C1(n263), .Y(n1357) );
  AOI222XLTS U101 ( .A0(n4016), .A1(n3417), .B0(n548), .B1(n3403), .C0(n4173), 
        .C1(n249), .Y(n1355) );
  AOI222XLTS U102 ( .A0(n4013), .A1(n3417), .B0(n554), .B1(n3402), .C0(n4170), 
        .C1(n250), .Y(n1353) );
  AOI222XLTS U103 ( .A0(n4001), .A1(n3416), .B0(n562), .B1(n3403), .C0(n4158), 
        .C1(n249), .Y(n1345) );
  AOI222XLTS U104 ( .A0(n4121), .A1(n3355), .B0(n3340), .B1(n198), .C0(n3966), 
        .C1(n3320), .Y(n1692) );
  AOI222XLTS U105 ( .A0(n4082), .A1(n3362), .B0(n469), .B1(n3334), .C0(n3927), 
        .C1(n3329), .Y(n1335) );
  AOI222XLTS U106 ( .A0(n4076), .A1(n3358), .B0(n473), .B1(n3334), .C0(n3921), 
        .C1(n3332), .Y(n1331) );
  AOI222XLTS U107 ( .A0(n4073), .A1(n3358), .B0(n475), .B1(n3334), .C0(n3918), 
        .C1(n3326), .Y(n1329) );
  AOI222XLTS U108 ( .A0(n4070), .A1(n3358), .B0(n477), .B1(n3346), .C0(n3915), 
        .C1(n3331), .Y(n1327) );
  AOI222XLTS U109 ( .A0(n4067), .A1(n3359), .B0(n479), .B1(n3345), .C0(n3912), 
        .C1(n3331), .Y(n1325) );
  AOI222XLTS U110 ( .A0(n4064), .A1(n3359), .B0(n481), .B1(n3344), .C0(n3909), 
        .C1(n3330), .Y(n1323) );
  AOI222XLTS U111 ( .A0(n4061), .A1(n3361), .B0(n483), .B1(n3335), .C0(n3906), 
        .C1(n3327), .Y(n1321) );
  AOI222XLTS U112 ( .A0(n4046), .A1(n3353), .B0(n493), .B1(n3346), .C0(n3891), 
        .C1(n3328), .Y(n1311) );
  AOI222XLTS U113 ( .A0(n4031), .A1(n3352), .B0(n512), .B1(n3337), .C0(n3876), 
        .C1(n3324), .Y(n1301) );
  AOI222XLTS U114 ( .A0(n4019), .A1(n3354), .B0(n544), .B1(n3337), .C0(n3864), 
        .C1(n3323), .Y(n1293) );
  AOI222XLTS U115 ( .A0(n4013), .A1(n3351), .B0(n551), .B1(n3337), .C0(n3858), 
        .C1(n3322), .Y(n1289) );
  AOI222XLTS U116 ( .A0(n4007), .A1(n3350), .B0(n557), .B1(n3339), .C0(n3852), 
        .C1(n3322), .Y(n1285) );
  AOI222XLTS U117 ( .A0(n4004), .A1(n3350), .B0(n560), .B1(n3339), .C0(n3849), 
        .C1(n3322), .Y(n1283) );
  AOI222XLTS U118 ( .A0(n3998), .A1(n3350), .B0(n564), .B1(n3339), .C0(n3843), 
        .C1(n3321), .Y(n1279) );
  AOI222XLTS U119 ( .A0(n4085), .A1(n3362), .B0(n468), .B1(n3346), .C0(n3930), 
        .C1(n3326), .Y(n1337) );
  AOI222XLTS U120 ( .A0(n4079), .A1(n3361), .B0(n471), .B1(n3344), .C0(n3924), 
        .C1(n3330), .Y(n1333) );
  AOI222XLTS U121 ( .A0(n4058), .A1(n3359), .B0(n485), .B1(n3335), .C0(n3903), 
        .C1(n3327), .Y(n1319) );
  AOI222XLTS U122 ( .A0(n4055), .A1(n3354), .B0(n487), .B1(n940), .C0(n3900), 
        .C1(n3328), .Y(n1317) );
  AOI222XLTS U123 ( .A0(n4052), .A1(n3354), .B0(n489), .B1(n3335), .C0(n3897), 
        .C1(n3326), .Y(n1315) );
  AOI222XLTS U124 ( .A0(n4049), .A1(n3354), .B0(n491), .B1(n3336), .C0(n3894), 
        .C1(n3327), .Y(n1313) );
  AOI222XLTS U125 ( .A0(n4040), .A1(n3353), .B0(n505), .B1(n3334), .C0(n3885), 
        .C1(n3327), .Y(n1307) );
  AOI222XLTS U126 ( .A0(n4028), .A1(n3352), .B0(n515), .B1(n3336), .C0(n3873), 
        .C1(n3323), .Y(n1299) );
  AOI222XLTS U127 ( .A0(n4025), .A1(n3352), .B0(n537), .B1(n3338), .C0(n3870), 
        .C1(n3323), .Y(n1297) );
  AOI222XLTS U128 ( .A0(n4022), .A1(n3351), .B0(n541), .B1(n3338), .C0(n3867), 
        .C1(n3323), .Y(n1295) );
  AOI222XLTS U129 ( .A0(n4016), .A1(n3351), .B0(n546), .B1(n3338), .C0(n3861), 
        .C1(n3322), .Y(n1291) );
  AOI222XLTS U130 ( .A0(n4010), .A1(n3351), .B0(n555), .B1(n3337), .C0(n3855), 
        .C1(n3324), .Y(n1287) );
  AOI222XLTS U131 ( .A0(n3995), .A1(n3349), .B0(n567), .B1(n3339), .C0(n3840), 
        .C1(n3321), .Y(n1277) );
  AOI222XLTS U132 ( .A0(n3992), .A1(n3349), .B0(n568), .B1(n3336), .C0(n3837), 
        .C1(n3321), .Y(n1275) );
  AOI222XLTS U133 ( .A0(n4043), .A1(n3353), .B0(n501), .B1(n3336), .C0(n3888), 
        .C1(n3326), .Y(n1309) );
  AOI222XLTS U134 ( .A0(n4037), .A1(n3353), .B0(n508), .B1(n3335), .C0(n3882), 
        .C1(n3324), .Y(n1305) );
  AOI222XLTS U135 ( .A0(n4034), .A1(n3352), .B0(n511), .B1(n3345), .C0(n3879), 
        .C1(n3324), .Y(n1303) );
  AOI222XLTS U136 ( .A0(n4001), .A1(n3350), .B0(n563), .B1(n3338), .C0(n3846), 
        .C1(n3321), .Y(n1281) );
  CLKBUFX2TS U137 ( .A(n922), .Y(n3430) );
  CLKBUFX2TS U138 ( .A(n989), .Y(n835) );
  NAND2X1TS U139 ( .A(n447), .B(selectBit_SOUTH), .Y(n1802) );
  INVX2TS U140 ( .A(n454), .Y(n203) );
  OA22X1TS U141 ( .A0(n1562), .A1(n576), .B0(n240), .B1(n243), .Y(n589) );
  CLKBUFX2TS U142 ( .A(n589), .Y(n734) );
  AND2X2TS U143 ( .A(n162), .B(n1555), .Y(n891) );
  INVX2TS U144 ( .A(n903), .Y(n513) );
  OA22X1TS U145 ( .A0(n1574), .A1(n577), .B0(n242), .B1(n7), .Y(n584) );
  OR2X2TS U146 ( .A(n881), .B(n236), .Y(n3) );
  OA22X1TS U147 ( .A0(n1569), .A1(n576), .B0(n1629), .B1(n7), .Y(n588) );
  OA22X1TS U148 ( .A0(n1556), .A1(n577), .B0(n240), .B1(n1629), .Y(n591) );
  INVX2TS U149 ( .A(n1550), .Y(n163) );
  OAI211X1TS U150 ( .A0(n3138), .A1(n847), .B0(n1134), .C0(n1135), .Y(n2776)
         );
  NAND3X1TS U151 ( .A(n1631), .B(n1727), .C(n456), .Y(n1581) );
  NOR3X2TS U152 ( .A(n534), .B(n317), .C(n1802), .Y(n1555) );
  NAND2X2TS U153 ( .A(n532), .B(n254), .Y(n1630) );
  BUFX2TS U154 ( .A(n3330), .Y(n3320) );
  CLKBUFX2TS U155 ( .A(n992), .Y(n804) );
  CLKBUFX2TS U156 ( .A(n925), .Y(n3399) );
  AOI21X1TS U157 ( .A0(n221), .A1(n239), .B0(n499), .Y(n1795) );
  AOI21X1TS U158 ( .A0(n526), .A1(n1726), .B0(n518), .Y(n1601) );
  CLKBUFX2TS U159 ( .A(n3811), .Y(n3809) );
  CLKBUFX2TS U160 ( .A(n865), .Y(n864) );
  CLKBUFX2TS U161 ( .A(n513), .Y(n3733) );
  AND3X2TS U162 ( .A(n219), .B(n1568), .C(n1564), .Y(n922) );
  NAND3X1TS U163 ( .A(n524), .B(n1655), .C(n525), .Y(n1604) );
  OA22X1TS U164 ( .A0(n1597), .A1(n578), .B0(n1629), .B1(n542), .Y(n590) );
  OAI21X1TS U165 ( .A0(n1801), .A1(n160), .B0(n533), .Y(n1678) );
  NOR2X1TS U166 ( .A(n255), .B(n532), .Y(n1726) );
  CLKBUFX2TS U167 ( .A(n3364), .Y(n3357) );
  CLKBUFX2TS U168 ( .A(n3237), .Y(n3230) );
  CLKBUFX2TS U169 ( .A(n1007), .Y(n748) );
  AOI21X1TS U170 ( .A0(n220), .A1(n1725), .B0(n504), .Y(n1586) );
  CLKBUFX2TS U171 ( .A(n3201), .Y(n1817) );
  INVX2TS U172 ( .A(n1584), .Y(n534) );
  INVX2TS U173 ( .A(n18), .Y(n217) );
  CLKBUFX2TS U174 ( .A(n3811), .Y(n3810) );
  CLKBUFX2TS U175 ( .A(n3363), .Y(n3356) );
  CLKBUFX2TS U176 ( .A(n1540), .Y(n572) );
  CLKBUFX2TS U177 ( .A(n3429), .Y(n3422) );
  CLKBUFX2TS U178 ( .A(n1540), .Y(n573) );
  NAND2X1TS U179 ( .A(n1589), .B(n1586), .Y(n1541) );
  AOI222XLTS U180 ( .A0(n3990), .A1(n770), .B0(n4303), .B1(n749), .C0(n4146), 
        .C1(n574), .Y(n1794) );
  AOI222XLTS U181 ( .A0(n4146), .A1(n798), .B0(destinationAddressIn_SOUTH[13]), 
        .B1(n380), .C0(n3991), .C1(n835), .Y(n1772) );
  AOI222XLTS U182 ( .A0(n3987), .A1(n3507), .B0(n4300), .B1(n3514), .C0(n4144), 
        .C1(n3553), .Y(n1626) );
  AOI222XLTS U183 ( .A0(n3837), .A1(n3724), .B0(n568), .B1(n3467), .C0(n3993), 
        .C1(n3450), .Y(n1404) );
  AOI222XLTS U184 ( .A0(n3840), .A1(n3719), .B0(n566), .B1(n3467), .C0(n3996), 
        .C1(n3450), .Y(n1406) );
  AOI222XLTS U185 ( .A0(n3843), .A1(n3719), .B0(n564), .B1(n3468), .C0(n3999), 
        .C1(n3450), .Y(n1408) );
  AOI222XLTS U186 ( .A0(n3846), .A1(n3719), .B0(n562), .B1(n3468), .C0(n4002), 
        .C1(n3450), .Y(n1410) );
  AOI222XLTS U187 ( .A0(n3849), .A1(n3719), .B0(n561), .B1(n3468), .C0(n4005), 
        .C1(n3451), .Y(n1412) );
  AOI222XLTS U188 ( .A0(n3852), .A1(n3720), .B0(n557), .B1(n3468), .C0(n4008), 
        .C1(n3451), .Y(n1414) );
  AOI222XLTS U189 ( .A0(n3855), .A1(n3720), .B0(n555), .B1(n3469), .C0(n4011), 
        .C1(n3453), .Y(n1416) );
  AOI222XLTS U190 ( .A0(n3858), .A1(n3720), .B0(n551), .B1(n3469), .C0(n4014), 
        .C1(n3451), .Y(n1418) );
  AOI222XLTS U191 ( .A0(n3861), .A1(n3720), .B0(n546), .B1(n3469), .C0(n4017), 
        .C1(n3451), .Y(n1420) );
  AOI222XLTS U192 ( .A0(n3864), .A1(n3721), .B0(n544), .B1(n3469), .C0(n4020), 
        .C1(n3452), .Y(n1422) );
  AOI222XLTS U193 ( .A0(n3867), .A1(n3721), .B0(n541), .B1(n3470), .C0(n4023), 
        .C1(n3452), .Y(n1424) );
  AOI222XLTS U194 ( .A0(n3870), .A1(n3721), .B0(n536), .B1(n3470), .C0(n4026), 
        .C1(n3452), .Y(n1426) );
  AOI222XLTS U195 ( .A0(n3873), .A1(n3721), .B0(n515), .B1(n3470), .C0(n4029), 
        .C1(n3452), .Y(n1428) );
  AOI222XLTS U196 ( .A0(n3876), .A1(n3722), .B0(n512), .B1(n3470), .C0(n4032), 
        .C1(n3453), .Y(n1430) );
  AOI222XLTS U197 ( .A0(n3879), .A1(n3722), .B0(n509), .B1(n3471), .C0(n4035), 
        .C1(n3453), .Y(n1432) );
  AOI222XLTS U198 ( .A0(n3882), .A1(n3722), .B0(n507), .B1(n3471), .C0(n4038), 
        .C1(n3453), .Y(n1434) );
  AOI222XLTS U199 ( .A0(n3885), .A1(n3722), .B0(n503), .B1(n3471), .C0(n4041), 
        .C1(n3454), .Y(n1436) );
  AOI222XLTS U200 ( .A0(n3888), .A1(n3723), .B0(n495), .B1(n3471), .C0(n4044), 
        .C1(n3454), .Y(n1438) );
  AOI222XLTS U201 ( .A0(n3891), .A1(n3723), .B0(n494), .B1(n3472), .C0(n4047), 
        .C1(n3454), .Y(n1440) );
  AOI222XLTS U202 ( .A0(n3894), .A1(n3723), .B0(n491), .B1(n3472), .C0(n4050), 
        .C1(n3454), .Y(n1442) );
  AOI222XLTS U203 ( .A0(n3897), .A1(n3723), .B0(n489), .B1(n3472), .C0(n4053), 
        .C1(n3455), .Y(n1444) );
  AOI222XLTS U204 ( .A0(n3900), .A1(n3724), .B0(n487), .B1(n3472), .C0(n4056), 
        .C1(n3455), .Y(n1446) );
  AOI222XLTS U205 ( .A0(n3903), .A1(n3724), .B0(n485), .B1(n3473), .C0(n4059), 
        .C1(n3455), .Y(n1448) );
  AOI222XLTS U206 ( .A0(n3906), .A1(n3724), .B0(n483), .B1(n3473), .C0(n4062), 
        .C1(n3455), .Y(n1450) );
  AOI222XLTS U207 ( .A0(n3909), .A1(n3725), .B0(n481), .B1(n3473), .C0(n4065), 
        .C1(n3456), .Y(n1452) );
  AOI222XLTS U208 ( .A0(n3912), .A1(n3725), .B0(n480), .B1(n3473), .C0(n4068), 
        .C1(n3456), .Y(n1454) );
  AOI222XLTS U209 ( .A0(n3915), .A1(n3725), .B0(n477), .B1(n3474), .C0(n4071), 
        .C1(n3456), .Y(n1456) );
  AOI222XLTS U210 ( .A0(n3918), .A1(n3725), .B0(n475), .B1(n3474), .C0(n4074), 
        .C1(n3456), .Y(n1458) );
  AOI222XLTS U211 ( .A0(n3921), .A1(n3726), .B0(n473), .B1(n3474), .C0(n4077), 
        .C1(n3457), .Y(n1460) );
  AOI222XLTS U212 ( .A0(n3924), .A1(n3726), .B0(n471), .B1(n3474), .C0(n4080), 
        .C1(n3457), .Y(n1462) );
  AOI222XLTS U213 ( .A0(n3927), .A1(n3726), .B0(n469), .B1(n3477), .C0(n4083), 
        .C1(n3457), .Y(n1464) );
  AOI222XLTS U214 ( .A0(n3930), .A1(n3726), .B0(n467), .B1(n3477), .C0(n4086), 
        .C1(n3457), .Y(n1466) );
  AOI222XLTS U215 ( .A0(n3981), .A1(n3507), .B0(n4294), .B1(n3514), .C0(n4138), 
        .C1(n3553), .Y(n1624) );
  AOI222XLTS U216 ( .A0(n4038), .A1(n3559), .B0(n508), .B1(n3534), .C0(n4194), 
        .C1(n3525), .Y(n1498) );
  AOI222XLTS U217 ( .A0(n4035), .A1(n3555), .B0(n511), .B1(n3534), .C0(n4191), 
        .C1(n3525), .Y(n1496) );
  AOI222XLTS U218 ( .A0(n4032), .A1(n3561), .B0(n514), .B1(n3543), .C0(n4188), 
        .C1(n3526), .Y(n1494) );
  AOI222XLTS U219 ( .A0(n3993), .A1(n3546), .B0(n569), .B1(n3537), .C0(n4149), 
        .C1(n3517), .Y(n1468) );
  AOI222XLTS U220 ( .A0(\requesterAddressbuffer[0][5] ), .A1(n238), .B0(n780), 
        .B1(n3948), .C0(n347), .C1(n4379), .Y(n1017) );
  AOI222XLTS U221 ( .A0(n4037), .A1(n3419), .B0(n507), .B1(n3408), .C0(n4194), 
        .C1(n377), .Y(n1369) );
  AOI222XLTS U222 ( .A0(n4025), .A1(n3418), .B0(n536), .B1(n3403), .C0(n4182), 
        .C1(n376), .Y(n1361) );
  AOI222XLTS U223 ( .A0(n3995), .A1(n3415), .B0(n566), .B1(n3404), .C0(n4152), 
        .C1(n278), .Y(n1341) );
  AOI222XLTS U224 ( .A0(n4076), .A1(n3426), .B0(n474), .B1(n3400), .C0(n4233), 
        .C1(n360), .Y(n1395) );
  AOI222XLTS U225 ( .A0(n4070), .A1(n3428), .B0(n478), .B1(n3410), .C0(n4227), 
        .C1(n377), .Y(n1391) );
  AOI222XLTS U226 ( .A0(n4061), .A1(n3425), .B0(n484), .B1(n3408), .C0(n4218), 
        .C1(n376), .Y(n1385) );
  AOI222XLTS U227 ( .A0(n4058), .A1(n3428), .B0(n486), .B1(n3409), .C0(n4215), 
        .C1(n377), .Y(n1383) );
  AOI222XLTS U228 ( .A0(n4049), .A1(n3424), .B0(n492), .B1(n3401), .C0(n4206), 
        .C1(n284), .Y(n1377) );
  AOI222XLTS U229 ( .A0(n4034), .A1(n3418), .B0(n509), .B1(n3410), .C0(n4191), 
        .C1(n376), .Y(n1367) );
  AOI222XLTS U230 ( .A0(n4031), .A1(n3418), .B0(n514), .B1(n3402), .C0(n4188), 
        .C1(n278), .Y(n1365) );
  AOI222XLTS U231 ( .A0(n4022), .A1(n3417), .B0(n543), .B1(n3403), .C0(n4179), 
        .C1(n278), .Y(n1359) );
  AOI222XLTS U232 ( .A0(n4010), .A1(n3417), .B0(n556), .B1(n3402), .C0(n4167), 
        .C1(n359), .Y(n1351) );
  AOI222XLTS U233 ( .A0(n4007), .A1(n3416), .B0(n559), .B1(n3404), .C0(n4164), 
        .C1(n278), .Y(n1349) );
  AOI222XLTS U234 ( .A0(n4004), .A1(n3416), .B0(n561), .B1(n3404), .C0(n4161), 
        .C1(n358), .Y(n1347) );
  AOI222XLTS U235 ( .A0(n3998), .A1(n3416), .B0(n565), .B1(n3404), .C0(n4155), 
        .C1(n375), .Y(n1343) );
  AOI222XLTS U236 ( .A0(n3992), .A1(n3415), .B0(n569), .B1(n3401), .C0(n4149), 
        .C1(n376), .Y(n1339) );
  AOI222XLTS U237 ( .A0(n3990), .A1(n3394), .B0(n4303), .B1(n377), .C0(n4146), 
        .C1(n3425), .Y(n1677) );
  AOI222XLTS U238 ( .A0(n4296), .A1(n1669), .B0(destinationAddressIn_EAST[11]), 
        .B1(n864), .C0(n3985), .C1(n3215), .Y(n1747) );
  AND3X2TS U239 ( .A(n162), .B(n533), .C(n1556), .Y(n4) );
  INVX2TS U240 ( .A(n924), .Y(n374) );
  INVX2TS U241 ( .A(n375), .Y(n247) );
  NAND2X1TS U242 ( .A(n1562), .B(n212), .Y(n1533) );
  INVX2TS U243 ( .A(n1584), .Y(n159) );
  AOI221X1TS U244 ( .A0(n241), .A1(n1773), .B0(n535), .B1(n279), .C0(n239), 
        .Y(n1584) );
  NOR2BX1TS U245 ( .AN(n1593), .B(n257), .Y(n991) );
  NAND2X1TS U246 ( .A(n1605), .B(n1795), .Y(n5) );
  INVX2TS U247 ( .A(n5), .Y(n496) );
  CLKINVX2TS U248 ( .A(n991), .Y(n443) );
  CLKINVX2TS U249 ( .A(n991), .Y(n267) );
  CLKINVX2TS U250 ( .A(n924), .Y(n437) );
  OR2X2TS U251 ( .A(n316), .B(n279), .Y(n7) );
  AND3X2TS U252 ( .A(n211), .B(n1598), .C(n1597), .Y(n11) );
  CLKBUFX2TS U253 ( .A(n871), .Y(n865) );
  NOR3X1TS U254 ( .A(n521), .B(n160), .C(n217), .Y(n959) );
  CLKBUFX2TS U255 ( .A(n959), .Y(n3237) );
  INVX2TS U256 ( .A(n390), .Y(n244) );
  OR3X1TS U257 ( .A(n320), .B(n236), .C(n459), .Y(n15) );
  AND2X2TS U258 ( .A(n5327), .B(n1764), .Y(n17) );
  CLKBUFX2TS U259 ( .A(n755), .Y(n747) );
  CLKINVX2TS U260 ( .A(n1550), .Y(n162) );
  NOR2BX1TS U261 ( .AN(n225), .B(n1729), .Y(n1567) );
  INVX2TS U262 ( .A(n1598), .Y(n256) );
  INVX2TS U263 ( .A(n256), .Y(n257) );
  OR2X2TS U264 ( .A(n872), .B(n13), .Y(n19) );
  CLKINVX1TS U265 ( .A(n159), .Y(n160) );
  INVXLTS U266 ( .A(n181), .Y(n164) );
  INVXLTS U267 ( .A(n185), .Y(n165) );
  INVXLTS U268 ( .A(n189), .Y(n166) );
  INVXLTS U269 ( .A(n193), .Y(n167) );
  CLKBUFX2TS U270 ( .A(readReady), .Y(n168) );
  CLKBUFX2TS U271 ( .A(selectBit_WEST), .Y(n169) );
  INVXLTS U272 ( .A(n579), .Y(n170) );
  CLKBUFX2TS U273 ( .A(selectBit_NORTH), .Y(n171) );
  INVX2TS U274 ( .A(n204), .Y(n172) );
  INVXLTS U275 ( .A(n454), .Y(n204) );
  INVXLTS U276 ( .A(n204), .Y(n173) );
  INVXLTS U277 ( .A(n203), .Y(n174) );
  INVXLTS U278 ( .A(n203), .Y(n175) );
  INVXLTS U279 ( .A(readRequesterAddress[0]), .Y(n176) );
  INVXLTS U280 ( .A(n176), .Y(n177) );
  INVXLTS U281 ( .A(n176), .Y(n178) );
  INVXLTS U282 ( .A(n176), .Y(n179) );
  INVXLTS U283 ( .A(n176), .Y(n180) );
  INVXLTS U284 ( .A(readRequesterAddress[1]), .Y(n181) );
  INVXLTS U285 ( .A(n181), .Y(n182) );
  INVXLTS U286 ( .A(n181), .Y(n183) );
  INVXLTS U287 ( .A(n181), .Y(n184) );
  INVXLTS U288 ( .A(readRequesterAddress[2]), .Y(n185) );
  INVXLTS U289 ( .A(n185), .Y(n186) );
  INVXLTS U290 ( .A(n185), .Y(n187) );
  INVXLTS U291 ( .A(n185), .Y(n188) );
  INVXLTS U292 ( .A(readRequesterAddress[3]), .Y(n189) );
  INVXLTS U293 ( .A(n189), .Y(n190) );
  INVXLTS U294 ( .A(n189), .Y(n191) );
  INVXLTS U295 ( .A(n189), .Y(n192) );
  INVXLTS U296 ( .A(readRequesterAddress[4]), .Y(n193) );
  INVXLTS U297 ( .A(n193), .Y(n194) );
  INVXLTS U298 ( .A(n193), .Y(n195) );
  INVXLTS U299 ( .A(n193), .Y(n196) );
  INVXLTS U300 ( .A(readRequesterAddress[5]), .Y(n197) );
  INVXLTS U301 ( .A(n197), .Y(n198) );
  INVXLTS U302 ( .A(n197), .Y(n199) );
  INVXLTS U303 ( .A(n197), .Y(n200) );
  INVXLTS U304 ( .A(n197), .Y(n201) );
  CLKBUFX2TS U305 ( .A(n454), .Y(n202) );
  INVX2TS U306 ( .A(n1533), .Y(n454) );
  INVXLTS U307 ( .A(n8), .Y(n205) );
  INVXLTS U308 ( .A(n10), .Y(n206) );
  OAI21X1TS U309 ( .A0(n1724), .A1(n253), .B0(n580), .Y(n435) );
  INVXLTS U310 ( .A(n1797), .Y(n207) );
  INVXLTS U311 ( .A(n207), .Y(n208) );
  CLKINVX2TS U312 ( .A(n1586), .Y(n209) );
  INVX1TS U313 ( .A(n209), .Y(n210) );
  AND2X2TS U314 ( .A(n1586), .B(n1656), .Y(n973) );
  CLKBUFX2TS U315 ( .A(n1593), .Y(n211) );
  AOI21X1TS U316 ( .A0(n463), .A1(n1763), .B0(n590), .Y(n1593) );
  CLKBUFX2TS U317 ( .A(n1557), .Y(n212) );
  AND2X2TS U318 ( .A(n1560), .B(n1557), .Y(n908) );
  NAND2X1TS U319 ( .A(n1563), .B(n1557), .Y(n903) );
  AOI21X1TS U320 ( .A0(n1619), .A1(n221), .B0(n589), .Y(n1557) );
  CLKBUFX2TS U321 ( .A(n1571), .Y(n213) );
  INVXLTS U322 ( .A(n535), .Y(n214) );
  INVXLTS U323 ( .A(n530), .Y(n215) );
  CLKBUFX2TS U324 ( .A(n1803), .Y(n447) );
  CLKINVX1TS U325 ( .A(n18), .Y(n216) );
  INVXLTS U326 ( .A(n1567), .Y(n218) );
  INVXLTS U327 ( .A(n218), .Y(n219) );
  INVXLTS U328 ( .A(n19), .Y(n220) );
  INVXLTS U329 ( .A(n19), .Y(n221) );
  INVXLTS U330 ( .A(n1725), .Y(n222) );
  INVXLTS U331 ( .A(n222), .Y(n223) );
  INVXLTS U332 ( .A(n7), .Y(n224) );
  INVXLTS U333 ( .A(n16), .Y(n225) );
  INVXLTS U334 ( .A(n16), .Y(n226) );
  INVXLTS U335 ( .A(n526), .Y(n227) );
  INVX2TS U336 ( .A(n1541), .Y(n502) );
  INVXLTS U337 ( .A(n15), .Y(n228) );
  INVXLTS U338 ( .A(n15), .Y(n229) );
  INVXLTS U339 ( .A(n3), .Y(n230) );
  INVXLTS U340 ( .A(n3786), .Y(n231) );
  INVXLTS U341 ( .A(n3786), .Y(n232) );
  INVX2TS U342 ( .A(n441), .Y(n442) );
  INVXLTS U343 ( .A(n2278), .Y(n233) );
  OAI2BB1X1TS U344 ( .A0N(n2249), .A1N(selectBit_EAST), .B0(n2281), .Y(n2278)
         );
  INVXLTS U345 ( .A(n744), .Y(n234) );
  INVXLTS U346 ( .A(n234), .Y(n235) );
  INVXLTS U347 ( .A(n455), .Y(n236) );
  INVXLTS U348 ( .A(n459), .Y(n237) );
  INVXLTS U349 ( .A(n434), .Y(n238) );
  INVXLTS U350 ( .A(n542), .Y(n239) );
  INVXLTS U351 ( .A(n1619), .Y(n240) );
  INVXLTS U352 ( .A(n240), .Y(n241) );
  INVXLTS U353 ( .A(n17), .Y(n242) );
  INVXLTS U354 ( .A(n17), .Y(n243) );
  INVXLTS U355 ( .A(n244), .Y(n245) );
  INVXLTS U356 ( .A(n244), .Y(n246) );
  INVX1TS U357 ( .A(n375), .Y(n248) );
  CLKINVX1TS U358 ( .A(n248), .Y(n249) );
  CLKINVX1TS U359 ( .A(n248), .Y(n250) );
  CLKBUFX2TS U360 ( .A(n2249), .Y(n251) );
  INVX2TS U361 ( .A(n578), .Y(n252) );
  INVXLTS U362 ( .A(n252), .Y(n253) );
  INVX2TS U363 ( .A(n778), .Y(n254) );
  INVXLTS U364 ( .A(n254), .Y(n255) );
  INVX1TS U365 ( .A(n443), .Y(n258) );
  INVXLTS U366 ( .A(n261), .Y(n259) );
  INVXLTS U367 ( .A(n261), .Y(n260) );
  CLKINVX2TS U368 ( .A(n258), .Y(n261) );
  INVX1TS U369 ( .A(n261), .Y(n262) );
  CLKINVX1TS U370 ( .A(n248), .Y(n263) );
  INVXLTS U371 ( .A(n264), .Y(n383) );
  INVXLTS U372 ( .A(n264), .Y(n382) );
  INVXLTS U373 ( .A(n267), .Y(n381) );
  INVX1TS U374 ( .A(n991), .Y(n264) );
  INVX1TS U375 ( .A(n264), .Y(n265) );
  CLKINVX1TS U376 ( .A(n264), .Y(n266) );
  INVX1TS U377 ( .A(n267), .Y(n268) );
  CLKINVX1TS U378 ( .A(n267), .Y(n269) );
  INVXLTS U379 ( .A(n389), .Y(n390) );
  INVXLTS U380 ( .A(n496), .Y(n270) );
  INVXLTS U381 ( .A(n270), .Y(n271) );
  INVXLTS U382 ( .A(n3773), .Y(n272) );
  INVXLTS U383 ( .A(n272), .Y(n273) );
  INVXLTS U384 ( .A(n272), .Y(n274) );
  INVXLTS U385 ( .A(n1833), .Y(n275) );
  INVXLTS U386 ( .A(n275), .Y(n276) );
  CLKINVX1TS U387 ( .A(n248), .Y(n277) );
  CLKINVX1TS U388 ( .A(n437), .Y(n278) );
  INVXLTS U389 ( .A(n12), .Y(n279) );
  INVXLTS U390 ( .A(n3298), .Y(n280) );
  INVXLTS U391 ( .A(n3298), .Y(n281) );
  INVXLTS U392 ( .A(n3687), .Y(n282) );
  INVXLTS U393 ( .A(n247), .Y(n283) );
  INVXLTS U394 ( .A(n247), .Y(n284) );
  INVXLTS U395 ( .A(n3802), .Y(n285) );
  INVXLTS U396 ( .A(n285), .Y(n286) );
  INVXLTS U397 ( .A(n285), .Y(n287) );
  INVXLTS U398 ( .A(n285), .Y(n288) );
  INVXLTS U399 ( .A(n730), .Y(n289) );
  INVXLTS U400 ( .A(n289), .Y(n290) );
  INVXLTS U401 ( .A(n289), .Y(n291) );
  INVXLTS U402 ( .A(n728), .Y(n292) );
  INVXLTS U403 ( .A(n292), .Y(n293) );
  INVXLTS U404 ( .A(n292), .Y(n294) );
  INVXLTS U405 ( .A(destinationAddressIn_NORTH[7]), .Y(n295) );
  INVXLTS U406 ( .A(destinationAddressIn_NORTH[7]), .Y(n296) );
  INVXLTS U407 ( .A(destinationAddressIn_NORTH[7]), .Y(n297) );
  INVXLTS U408 ( .A(n722), .Y(n298) );
  INVXLTS U409 ( .A(n298), .Y(n299) );
  INVXLTS U410 ( .A(n298), .Y(n300) );
  INVXLTS U411 ( .A(n724), .Y(n301) );
  INVXLTS U412 ( .A(n301), .Y(n302) );
  INVXLTS U413 ( .A(n301), .Y(n303) );
  INVXLTS U414 ( .A(n725), .Y(n304) );
  INVXLTS U415 ( .A(n304), .Y(n305) );
  INVXLTS U416 ( .A(n304), .Y(n306) );
  INVXLTS U417 ( .A(n721), .Y(n307) );
  INVXLTS U418 ( .A(n307), .Y(n308) );
  INVXLTS U419 ( .A(n307), .Y(n309) );
  INVXLTS U420 ( .A(n723), .Y(n310) );
  INVXLTS U421 ( .A(n310), .Y(n311) );
  INVXLTS U422 ( .A(n310), .Y(n312) );
  INVXLTS U423 ( .A(n726), .Y(n313) );
  INVXLTS U424 ( .A(n313), .Y(n314) );
  INVXLTS U425 ( .A(n313), .Y(n315) );
  INVXLTS U426 ( .A(n594), .Y(n316) );
  INVXLTS U427 ( .A(n316), .Y(n317) );
  INVXLTS U428 ( .A(n13), .Y(n318) );
  INVXLTS U429 ( .A(n14), .Y(n319) );
  INVXLTS U430 ( .A(n14), .Y(n320) );
  INVXLTS U431 ( .A(n3802), .Y(n321) );
  INVXLTS U432 ( .A(n321), .Y(n322) );
  INVXLTS U433 ( .A(n321), .Y(n323) );
  INVXLTS U434 ( .A(n321), .Y(n324) );
  INVXLTS U435 ( .A(n238), .Y(n325) );
  INVXLTS U436 ( .A(n325), .Y(n326) );
  INVXLTS U437 ( .A(n325), .Y(n327) );
  INVXLTS U438 ( .A(n325), .Y(n328) );
  INVXLTS U439 ( .A(n452), .Y(n329) );
  INVXLTS U440 ( .A(n329), .Y(n330) );
  INVXLTS U441 ( .A(n329), .Y(n331) );
  INVXLTS U442 ( .A(n329), .Y(n332) );
  INVXLTS U443 ( .A(n452), .Y(n333) );
  INVXLTS U444 ( .A(n333), .Y(n334) );
  INVXLTS U445 ( .A(n333), .Y(n335) );
  INVXLTS U446 ( .A(n333), .Y(n336) );
  INVXLTS U447 ( .A(n452), .Y(n337) );
  INVXLTS U448 ( .A(n337), .Y(n338) );
  INVXLTS U449 ( .A(n337), .Y(n339) );
  INVXLTS U450 ( .A(n337), .Y(n340) );
  INVXLTS U451 ( .A(n496), .Y(n341) );
  INVXLTS U452 ( .A(n341), .Y(n342) );
  INVXLTS U453 ( .A(n341), .Y(n343) );
  INVXLTS U454 ( .A(n341), .Y(n344) );
  INVXLTS U455 ( .A(n496), .Y(n345) );
  INVXLTS U456 ( .A(n345), .Y(n346) );
  INVXLTS U457 ( .A(n345), .Y(n347) );
  INVXLTS U458 ( .A(n345), .Y(n348) );
  INVXLTS U459 ( .A(n432), .Y(n349) );
  INVXLTS U460 ( .A(n349), .Y(n350) );
  INVXLTS U461 ( .A(n349), .Y(n351) );
  INVXLTS U462 ( .A(n349), .Y(n352) );
  INVXLTS U463 ( .A(n433), .Y(n353) );
  INVXLTS U464 ( .A(n353), .Y(n354) );
  INVXLTS U465 ( .A(n353), .Y(n355) );
  INVXLTS U466 ( .A(n353), .Y(n356) );
  INVXLTS U467 ( .A(n437), .Y(n357) );
  INVXLTS U468 ( .A(n437), .Y(n358) );
  INVXLTS U469 ( .A(n437), .Y(n359) );
  INVXLTS U470 ( .A(n374), .Y(n360) );
  INVXLTS U471 ( .A(n4), .Y(n361) );
  INVXLTS U472 ( .A(n361), .Y(n362) );
  INVXLTS U473 ( .A(n361), .Y(n363) );
  INVXLTS U474 ( .A(n361), .Y(n364) );
  INVXLTS U475 ( .A(n361), .Y(n365) );
  INVXLTS U476 ( .A(n449), .Y(n366) );
  INVXLTS U477 ( .A(n449), .Y(n367) );
  INVXLTS U478 ( .A(n449), .Y(n368) );
  INVXLTS U479 ( .A(n4), .Y(n369) );
  INVXLTS U480 ( .A(n369), .Y(n370) );
  INVXLTS U481 ( .A(n369), .Y(n371) );
  INVXLTS U482 ( .A(n369), .Y(n372) );
  INVXLTS U483 ( .A(n369), .Y(n373) );
  AOI222XLTS U484 ( .A0(n4088), .A1(n3547), .B0(n177), .B1(n3538), .C0(n4245), 
        .C1(n3525), .Y(n888) );
  AOI222XLTS U485 ( .A0(n4094), .A1(n3545), .B0(n188), .B1(n3538), .C0(n4251), 
        .C1(n3517), .Y(n896) );
  AOI222XLTS U486 ( .A0(n4097), .A1(n3545), .B0(n192), .B1(n3538), .C0(n4254), 
        .C1(n3516), .Y(n898) );
  AOI222XLTS U487 ( .A0(n4100), .A1(n3545), .B0(n196), .B1(n3537), .C0(n4257), 
        .C1(n3517), .Y(n900) );
  AOI222XLTS U488 ( .A0(n4103), .A1(n3546), .B0(n201), .B1(n3537), .C0(n4260), 
        .C1(n3517), .Y(n902) );
  AOI222XLTS U489 ( .A0(n3966), .A1(n835), .B0(n811), .B1(n198), .C0(n4278), 
        .C1(n381), .Y(n1762) );
  INVX1TS U490 ( .A(n374), .Y(n375) );
  CLKINVX1TS U491 ( .A(n374), .Y(n376) );
  CLKINVX1TS U492 ( .A(n374), .Y(n377) );
  CLKINVX1TS U493 ( .A(n443), .Y(n378) );
  CLKINVX1TS U494 ( .A(n267), .Y(n379) );
  CLKINVX1TS U495 ( .A(n443), .Y(n380) );
  CLKINVX1TS U496 ( .A(n3802), .Y(n384) );
  INVXLTS U497 ( .A(n384), .Y(n385) );
  INVXLTS U498 ( .A(n452), .Y(n386) );
  CLKINVX1TS U499 ( .A(n386), .Y(n387) );
  CLKINVX1TS U500 ( .A(n386), .Y(n388) );
  INVX2TS U501 ( .A(n496), .Y(n389) );
  INVXLTS U502 ( .A(n389), .Y(n391) );
  INVXLTS U503 ( .A(n389), .Y(n392) );
  CLKINVX2TS U543 ( .A(n1542), .Y(n504) );
  CLKINVX2TS U544 ( .A(n1701), .Y(n519) );
  NAND3X1TS U545 ( .A(n2251), .B(n579), .C(n171), .Y(n1814) );
  INVX1TS U546 ( .A(selectBit_NORTH), .Y(n718) );
  CLKBUFX2TS U547 ( .A(n504), .Y(n432) );
  CLKBUFX2TS U548 ( .A(n504), .Y(n433) );
  NOR2X1TS U549 ( .A(n1592), .B(n1630), .Y(n1560) );
  CLKAND2X2TS U550 ( .A(n1553), .B(n163), .Y(n889) );
  OA21XLTS U551 ( .A0(n1678), .A1(n1679), .B0(n1568), .Y(n1569) );
  INVXLTS U552 ( .A(n1568), .Y(n523) );
  OAI22X1TS U553 ( .A0(n1605), .A1(n577), .B0(n242), .B1(n542), .Y(n434) );
  NOR3X1TS U554 ( .A(n1577), .B(n518), .C(n498), .Y(n1549) );
  OAI211X1TS U555 ( .A0(n4102), .A1(n3809), .B0(n1014), .C0(n1015), .Y(n2836)
         );
  OAI211X1TS U556 ( .A0(n4099), .A1(n3810), .B0(n1012), .C0(n1013), .Y(n2837)
         );
  OAI211X1TS U557 ( .A0(n4105), .A1(n3809), .B0(n1016), .C0(n1017), .Y(n2835)
         );
  OAI21XLTS U558 ( .A0(n1724), .A1(n253), .B0(n580), .Y(n436) );
  OAI22X1TS U559 ( .A0(n1589), .A1(n576), .B0(n243), .B1(n222), .Y(n438) );
  CLKBUFX2TS U560 ( .A(n3773), .Y(n3772) );
  CLKBUFX2TS U561 ( .A(n2), .Y(n439) );
  CLKBUFX2TS U562 ( .A(n2), .Y(n440) );
  CLKINVX2TS U563 ( .A(n1591), .Y(n441) );
  OAI211X1TS U564 ( .A0(n2897), .A1(n840), .B0(n1761), .C0(n1762), .Y(n2473)
         );
  INVX2TS U565 ( .A(n1795), .Y(n498) );
  CLKINVX2TS U566 ( .A(n11), .Y(n444) );
  INVXLTS U567 ( .A(n11), .Y(n445) );
  INVXLTS U568 ( .A(n11), .Y(n446) );
  NAND3X1TS U569 ( .A(n1655), .B(n1680), .C(n524), .Y(n1701) );
  AND2XLTS U570 ( .A(n442), .B(n210), .Y(n582) );
  AOI221X2TS U571 ( .A0(n527), .A1(n1726), .B0(n279), .B1(n1656), .C0(n1591), 
        .Y(n1589) );
  NOR3BX1TS U572 ( .AN(n1586), .B(n1592), .C(n442), .Y(n975) );
  CLKINVX2TS U573 ( .A(n373), .Y(n448) );
  CLKINVX2TS U574 ( .A(n3718), .Y(n449) );
  CLKINVX2TS U575 ( .A(n3718), .Y(n450) );
  CLKINVX2TS U576 ( .A(n3756), .Y(n451) );
  INVX2TS U577 ( .A(n1537), .Y(n452) );
  AOI32X1TS U578 ( .A0(n778), .A1(n731), .A2(n171), .B0(n2282), .B1(
        selectBit_SOUTH), .Y(n2281) );
  AND3XLTS U579 ( .A(n1601), .B(n1602), .C(n1795), .Y(n1007) );
  INVXLTS U580 ( .A(n1602), .Y(n530) );
  AOI21X1TS U581 ( .A0(n579), .A1(n447), .B0(n1602), .Y(n1729) );
  NOR2X1TS U582 ( .A(n731), .B(n447), .Y(n1602) );
  CLKINVX2TS U583 ( .A(n174), .Y(n453) );
  CLKBUFX2TS U584 ( .A(n172), .Y(n3741) );
  AND2XLTS U585 ( .A(n252), .B(n4392), .Y(n874) );
  INVX2TS U586 ( .A(n874), .Y(n457) );
  INVX2TS U587 ( .A(n874), .Y(n458) );
  OR2X2TS U588 ( .A(n1813), .B(n713), .Y(n1837) );
  INVX2TS U589 ( .A(n1837), .Y(n461) );
  INVX2TS U590 ( .A(n1837), .Y(n462) );
  CLKBUFX2TS U591 ( .A(n1628), .Y(n463) );
  OAI31XLTS U592 ( .A0(n1628), .A1(n531), .A2(n214), .B0(n1764), .Y(n1629) );
  INVX2TS U593 ( .A(n3729), .Y(n464) );
  INVX2TS U594 ( .A(n1825), .Y(n465) );
  INVX2TS U595 ( .A(n3702), .Y(n466) );
  CLKBUFX2TS U596 ( .A(cacheDataOut[31]), .Y(n467) );
  CLKBUFX2TS U597 ( .A(cacheDataOut[31]), .Y(n468) );
  CLKBUFX2TS U598 ( .A(cacheDataOut[30]), .Y(n469) );
  CLKBUFX2TS U599 ( .A(cacheDataOut[30]), .Y(n470) );
  CLKBUFX2TS U600 ( .A(cacheDataOut[29]), .Y(n471) );
  CLKBUFX2TS U601 ( .A(cacheDataOut[29]), .Y(n472) );
  CLKBUFX2TS U602 ( .A(cacheDataOut[28]), .Y(n473) );
  CLKBUFX2TS U603 ( .A(cacheDataOut[28]), .Y(n474) );
  CLKBUFX2TS U604 ( .A(cacheDataOut[27]), .Y(n475) );
  CLKBUFX2TS U605 ( .A(cacheDataOut[27]), .Y(n476) );
  CLKBUFX2TS U606 ( .A(cacheDataOut[26]), .Y(n477) );
  CLKBUFX2TS U607 ( .A(cacheDataOut[26]), .Y(n478) );
  CLKBUFX2TS U608 ( .A(cacheDataOut[25]), .Y(n479) );
  CLKBUFX2TS U609 ( .A(cacheDataOut[25]), .Y(n480) );
  CLKBUFX2TS U610 ( .A(cacheDataOut[24]), .Y(n481) );
  CLKBUFX2TS U611 ( .A(cacheDataOut[24]), .Y(n482) );
  CLKBUFX2TS U612 ( .A(cacheDataOut[23]), .Y(n483) );
  CLKBUFX2TS U613 ( .A(cacheDataOut[23]), .Y(n484) );
  CLKBUFX2TS U614 ( .A(cacheDataOut[22]), .Y(n485) );
  CLKBUFX2TS U615 ( .A(cacheDataOut[22]), .Y(n486) );
  CLKBUFX2TS U616 ( .A(cacheDataOut[21]), .Y(n487) );
  CLKBUFX2TS U617 ( .A(cacheDataOut[21]), .Y(n488) );
  CLKBUFX2TS U618 ( .A(cacheDataOut[20]), .Y(n489) );
  CLKBUFX2TS U619 ( .A(cacheDataOut[20]), .Y(n490) );
  CLKBUFX2TS U620 ( .A(cacheDataOut[19]), .Y(n491) );
  CLKBUFX2TS U621 ( .A(cacheDataOut[19]), .Y(n492) );
  CLKBUFX2TS U622 ( .A(cacheDataOut[18]), .Y(n493) );
  CLKBUFX2TS U623 ( .A(cacheDataOut[18]), .Y(n494) );
  CLKBUFX2TS U624 ( .A(cacheDataOut[17]), .Y(n495) );
  CLKBUFX2TS U625 ( .A(cacheDataOut[17]), .Y(n501) );
  CLKBUFX2TS U626 ( .A(cacheDataOut[16]), .Y(n503) );
  CLKBUFX2TS U627 ( .A(cacheDataOut[16]), .Y(n505) );
  CLKBUFX2TS U628 ( .A(cacheDataOut[15]), .Y(n507) );
  CLKBUFX2TS U629 ( .A(cacheDataOut[15]), .Y(n508) );
  CLKBUFX2TS U630 ( .A(cacheDataOut[14]), .Y(n509) );
  CLKBUFX2TS U631 ( .A(cacheDataOut[14]), .Y(n511) );
  CLKBUFX2TS U632 ( .A(cacheDataOut[13]), .Y(n512) );
  CLKBUFX2TS U633 ( .A(cacheDataOut[13]), .Y(n514) );
  CLKBUFX2TS U634 ( .A(cacheDataOut[12]), .Y(n515) );
  CLKBUFX2TS U635 ( .A(cacheDataOut[12]), .Y(n516) );
  CLKBUFX2TS U636 ( .A(cacheDataOut[11]), .Y(n536) );
  CLKBUFX2TS U637 ( .A(cacheDataOut[11]), .Y(n537) );
  CLKBUFX2TS U638 ( .A(cacheDataOut[10]), .Y(n541) );
  CLKBUFX2TS U639 ( .A(cacheDataOut[10]), .Y(n543) );
  CLKBUFX2TS U640 ( .A(cacheDataOut[9]), .Y(n544) );
  CLKBUFX2TS U641 ( .A(cacheDataOut[9]), .Y(n545) );
  CLKBUFX2TS U642 ( .A(cacheDataOut[8]), .Y(n546) );
  CLKBUFX2TS U643 ( .A(cacheDataOut[8]), .Y(n548) );
  CLKBUFX2TS U644 ( .A(cacheDataOut[7]), .Y(n551) );
  CLKBUFX2TS U645 ( .A(cacheDataOut[7]), .Y(n554) );
  CLKBUFX2TS U646 ( .A(cacheDataOut[6]), .Y(n555) );
  CLKBUFX2TS U647 ( .A(cacheDataOut[6]), .Y(n556) );
  CLKBUFX2TS U648 ( .A(cacheDataOut[5]), .Y(n557) );
  CLKBUFX2TS U649 ( .A(cacheDataOut[5]), .Y(n559) );
  CLKBUFX2TS U650 ( .A(cacheDataOut[4]), .Y(n560) );
  CLKBUFX2TS U651 ( .A(cacheDataOut[4]), .Y(n561) );
  CLKBUFX2TS U652 ( .A(cacheDataOut[3]), .Y(n562) );
  CLKBUFX2TS U653 ( .A(cacheDataOut[3]), .Y(n563) );
  CLKBUFX2TS U654 ( .A(cacheDataOut[2]), .Y(n564) );
  CLKBUFX2TS U655 ( .A(cacheDataOut[2]), .Y(n565) );
  CLKBUFX2TS U656 ( .A(cacheDataOut[1]), .Y(n566) );
  CLKBUFX2TS U657 ( .A(cacheDataOut[1]), .Y(n567) );
  CLKBUFX2TS U658 ( .A(cacheDataOut[0]), .Y(n568) );
  CLKBUFX2TS U659 ( .A(cacheDataOut[0]), .Y(n569) );
  CLKBUFX2TS U660 ( .A(n885), .Y(n570) );
  CLKBUFX2TS U661 ( .A(n885), .Y(n571) );
  NOR3X1TS U662 ( .A(n528), .B(n522), .C(n217), .Y(n1540) );
  CLKBUFX2TS U663 ( .A(n1549), .Y(n574) );
  CLKBUFX2TS U664 ( .A(n1549), .Y(n575) );
  INVXLTS U665 ( .A(n1549), .Y(n497) );
  CLKBUFX2TS U666 ( .A(n1764), .Y(n517) );
  INVX2TS U667 ( .A(n517), .Y(n576) );
  INVX2TS U668 ( .A(n517), .Y(n577) );
  INVX2TS U669 ( .A(n517), .Y(n578) );
  INVXLTS U670 ( .A(selectBit_SOUTH), .Y(n731) );
  CLKBUFX2TS U671 ( .A(n731), .Y(n579) );
  INVX1TS U672 ( .A(n1540), .Y(n506) );
  INVX1TS U673 ( .A(n1656), .Y(n529) );
  AND3XLTS U674 ( .A(n1571), .B(n526), .C(n1701), .Y(n939) );
  AND2XLTS U675 ( .A(n1571), .B(n519), .Y(n941) );
  CLKBUFX2TS U676 ( .A(n497), .Y(n3816) );
  NAND2XLTS U677 ( .A(n1574), .B(n1571), .Y(n1537) );
  CLKINVX2TS U678 ( .A(n1580), .Y(n528) );
  INVX2TS U679 ( .A(n958), .Y(n580) );
  OA21XLTS U680 ( .A0(n532), .A1(n1679), .B0(n1596), .Y(n1597) );
  AND2XLTS U681 ( .A(n463), .B(n1764), .Y(n1618) );
  INVXLTS U682 ( .A(selectBit_WEST), .Y(n825) );
  OAI31XLTS U683 ( .A0(n2286), .A1(n1804), .A2(n1805), .B0(n1806), .Y(n2450)
         );
  OAI31XLTS U684 ( .A0(n2288), .A1(n1804), .A2(n1805), .B0(n1823), .Y(n2449)
         );
  INVXLTS U685 ( .A(n3217), .Y(n3212) );
  INVXLTS U686 ( .A(n3216), .Y(n3213) );
  INVXLTS U687 ( .A(n3215), .Y(n3214) );
  INVXLTS U688 ( .A(n3382), .Y(n3377) );
  INVXLTS U689 ( .A(n3382), .Y(n3376) );
  CLKBUFX2TS U690 ( .A(n854), .Y(n851) );
  CLKBUFX2TS U691 ( .A(n3382), .Y(n3379) );
  CLKBUFX2TS U692 ( .A(n733), .Y(n727) );
  CLKBUFX2TS U693 ( .A(n733), .Y(n717) );
  CLKBUFX2TS U694 ( .A(n854), .Y(n852) );
  CLKBUFX2TS U695 ( .A(n588), .Y(n3445) );
  CLKBUFX2TS U696 ( .A(n3448), .Y(n3446) );
  CLKBUFX2TS U697 ( .A(n3578), .Y(n3576) );
  BUFX3TS U698 ( .A(n3316), .Y(n3310) );
  NOR2XLTS U699 ( .A(n530), .B(n225), .Y(n1656) );
  OR2XLTS U700 ( .A(n216), .B(n534), .Y(n581) );
  CLKBUFX2TS U701 ( .A(n701), .Y(n696) );
  NAND3XLTS U702 ( .A(n161), .B(n257), .C(n1569), .Y(n1535) );
  NOR3BXLTS U703 ( .AN(n1655), .B(n525), .C(n524), .Y(n1563) );
  NOR3BXLTS U704 ( .AN(n1631), .B(n456), .C(n460), .Y(n1554) );
  NAND2XLTS U705 ( .A(n1729), .B(n1750), .Y(n1592) );
  NOR3BX1TS U706 ( .AN(n213), .B(n1576), .C(n530), .Y(n942) );
  NOR2BXLTS U707 ( .AN(n1564), .B(n257), .Y(n924) );
  NAND2XLTS U708 ( .A(n1602), .B(n225), .Y(n1702) );
  AND2XLTS U709 ( .A(n1561), .B(n1557), .Y(n906) );
  NOR2X1TS U710 ( .A(n6), .B(n12), .Y(n1763) );
  XOR2XLTS U711 ( .A(n318), .B(n720), .Y(n1774) );
  OAI22X1TS U712 ( .A0(n718), .A1(n731), .B0(n2249), .B1(n778), .Y(n1797) );
  NOR2X1TS U713 ( .A(n1774), .B(n825), .Y(n1655) );
  AOI32XLTS U714 ( .A0(n161), .A1(n1565), .A2(n1566), .B0(n3448), .B1(n29), 
        .Y(n2568) );
  AOI32XLTS U715 ( .A0(n1567), .A1(n1568), .A2(n3826), .B0(n1569), .B1(n1570), 
        .Y(n1566) );
  AOI32XLTS U716 ( .A0(n211), .A1(n1594), .A2(n1595), .B0(n851), .B1(n20), .Y(
        n2564) );
  AOI32XLTS U717 ( .A0(n1567), .A1(n1596), .A2(n3827), .B0(n1597), .B1(n1570), 
        .Y(n1595) );
  AND2XLTS U718 ( .A(n2249), .B(n2251), .Y(n1804) );
  INVXLTS U719 ( .A(n1773), .Y(n535) );
  AND2XLTS U720 ( .A(n2250), .B(n255), .Y(n2251) );
  INVXLTS U721 ( .A(n1592), .Y(n527) );
  NOR2X1TS U722 ( .A(n872), .B(n318), .Y(n1628) );
  OAI32XLTS U723 ( .A0(n3829), .A1(n442), .A2(n1592), .B0(n529), .B1(n235), 
        .Y(n1590) );
  NOR2X1TS U724 ( .A(n5326), .B(n317), .Y(n1619) );
  NOR2X1TS U725 ( .A(n12), .B(n5323), .Y(n1725) );
  NOR2X1TS U726 ( .A(n319), .B(n5327), .Y(n2276) );
  NOR3X1TS U727 ( .A(n455), .B(n9), .C(n206), .Y(n1834) );
  OAI211XLTS U728 ( .A0(n4096), .A1(n3810), .B0(n1010), .C0(n1011), .Y(n2838)
         );
  OAI211XLTS U729 ( .A0(n4093), .A1(n3810), .B0(n1008), .C0(n1009), .Y(n2839)
         );
  OAI211XLTS U730 ( .A0(n4090), .A1(n3810), .B0(n1003), .C0(n1004), .Y(n2840)
         );
  OAI211XLTS U731 ( .A0(n3809), .A1(n3997), .B0(n1020), .C0(n1021), .Y(n2833)
         );
  OAI211XLTS U732 ( .A0(n3809), .A1(n3994), .B0(n1018), .C0(n1019), .Y(n2834)
         );
  OAI211XLTS U733 ( .A0(n3803), .A1(n4123), .B0(n1785), .C0(n1786), .Y(n2459)
         );
  OAI211XLTS U734 ( .A0(n3803), .A1(n4117), .B0(n1781), .C0(n1782), .Y(n2461)
         );
  OAI211XLTS U735 ( .A0(n3803), .A1(n4114), .B0(n1779), .C0(n1780), .Y(n2462)
         );
  OAI211XLTS U736 ( .A0(n3804), .A1(n4111), .B0(n1777), .C0(n1778), .Y(n2463)
         );
  OAI211XLTS U737 ( .A0(n3804), .A1(n4087), .B0(n1080), .C0(n1081), .Y(n2803)
         );
  OAI211XLTS U738 ( .A0(n3804), .A1(n4084), .B0(n1078), .C0(n1079), .Y(n2804)
         );
  OAI211XLTS U739 ( .A0(n3805), .A1(n4081), .B0(n1076), .C0(n1077), .Y(n2805)
         );
  OAI211XLTS U740 ( .A0(n3805), .A1(n4072), .B0(n1070), .C0(n1071), .Y(n2808)
         );
  OAI211XLTS U741 ( .A0(n3806), .A1(n4069), .B0(n1068), .C0(n1069), .Y(n2809)
         );
  OAI211XLTS U742 ( .A0(n3806), .A1(n4066), .B0(n1066), .C0(n1067), .Y(n2810)
         );
  OAI211XLTS U743 ( .A0(n3806), .A1(n4060), .B0(n1062), .C0(n1063), .Y(n2812)
         );
  OAI211XLTS U744 ( .A0(n3807), .A1(n4057), .B0(n1060), .C0(n1061), .Y(n2813)
         );
  OAI211XLTS U745 ( .A0(n3807), .A1(n4051), .B0(n1056), .C0(n1057), .Y(n2815)
         );
  OAI211XLTS U746 ( .A0(n3807), .A1(n4048), .B0(n1054), .C0(n1055), .Y(n2816)
         );
  OAI211XLTS U747 ( .A0(n3813), .A1(n4045), .B0(n1052), .C0(n1053), .Y(n2817)
         );
  OAI211XLTS U748 ( .A0(n3812), .A1(n4042), .B0(n1050), .C0(n1051), .Y(n2818)
         );
  OAI211XLTS U749 ( .A0(n3814), .A1(n4039), .B0(n1048), .C0(n1049), .Y(n2819)
         );
  OAI211XLTS U750 ( .A0(n3815), .A1(n4036), .B0(n1046), .C0(n1047), .Y(n2820)
         );
  OAI211XLTS U751 ( .A0(n3811), .A1(n4033), .B0(n1044), .C0(n1045), .Y(n2821)
         );
  OAI211XLTS U752 ( .A0(n3811), .A1(n4030), .B0(n1042), .C0(n1043), .Y(n2822)
         );
  OAI211XLTS U753 ( .A0(n3816), .A1(n4027), .B0(n1040), .C0(n1041), .Y(n2823)
         );
  OAI211XLTS U754 ( .A0(n3816), .A1(n4024), .B0(n1038), .C0(n1039), .Y(n2824)
         );
  OAI211XLTS U755 ( .A0(n3813), .A1(n4018), .B0(n1034), .C0(n1035), .Y(n2826)
         );
  OAI211XLTS U756 ( .A0(n3814), .A1(n4015), .B0(n1032), .C0(n1033), .Y(n2827)
         );
  OAI211XLTS U757 ( .A0(n3812), .A1(n4012), .B0(n1030), .C0(n1031), .Y(n2828)
         );
  OAI211XLTS U758 ( .A0(n3808), .A1(n4006), .B0(n1026), .C0(n1027), .Y(n2830)
         );
  OAI211XLTS U759 ( .A0(n3808), .A1(n4003), .B0(n1024), .C0(n1025), .Y(n2831)
         );
  OAI211XLTS U760 ( .A0(n3803), .A1(n4120), .B0(n1783), .C0(n1784), .Y(n2460)
         );
  OAI211XLTS U761 ( .A0(n3804), .A1(n4108), .B0(n1775), .C0(n1776), .Y(n2464)
         );
  OAI211XLTS U762 ( .A0(n3805), .A1(n4078), .B0(n1074), .C0(n1075), .Y(n2806)
         );
  OAI211XLTS U763 ( .A0(n3805), .A1(n4075), .B0(n1072), .C0(n1073), .Y(n2807)
         );
  OAI211XLTS U764 ( .A0(n3806), .A1(n4063), .B0(n1064), .C0(n1065), .Y(n2811)
         );
  OAI211XLTS U765 ( .A0(n3807), .A1(n4054), .B0(n1058), .C0(n1059), .Y(n2814)
         );
  OAI211XLTS U766 ( .A0(n3814), .A1(n4021), .B0(n1036), .C0(n1037), .Y(n2825)
         );
  OAI211XLTS U767 ( .A0(n3808), .A1(n4009), .B0(n1028), .C0(n1029), .Y(n2829)
         );
  OAI211XLTS U768 ( .A0(n3808), .A1(n4000), .B0(n1022), .C0(n1023), .Y(n2832)
         );
  OAI22XLTS U769 ( .A0(n160), .A1(n235), .B0(n534), .B1(n3835), .Y(n1583) );
  AOI32XLTS U770 ( .A0(n1580), .A1(n1581), .A2(n3826), .B0(n1582), .B1(n1583), 
        .Y(n1579) );
  NOR2X1TS U771 ( .A(n2285), .B(n1804), .Y(n1764) );
  NAND2XLTS U772 ( .A(n3821), .B(n442), .Y(n1587) );
  AOI2BB2XLTS U773 ( .B0(readReady), .B1(selectBit_WEST), .A0N(n2250), .A1N(
        n720), .Y(n2256) );
  OAI211XLTS U774 ( .A0(n3949), .A1(n903), .B0(n917), .C0(n918), .Y(n2871) );
  AOI22XLTS U775 ( .A0(n3467), .A1(n199), .B0(n3461), .B1(n4103), .Y(n917) );
  OAI211XLTS U776 ( .A0(n3946), .A1(n903), .B0(n915), .C0(n916), .Y(n2872) );
  OAI211XLTS U777 ( .A0(n3943), .A1(n464), .B0(n913), .C0(n914), .Y(n2873) );
  OAI211XLTS U778 ( .A0(n3940), .A1(n464), .B0(n911), .C0(n912), .Y(n2874) );
  OAI211XLTS U779 ( .A0(n3937), .A1(n464), .B0(n909), .C0(n910), .Y(n2875) );
  OAI211XLTS U780 ( .A0(n3934), .A1(n464), .B0(n904), .C0(n905), .Y(n2876) );
  AOI22XLTS U781 ( .A0(n3466), .A1(n178), .B0(n3462), .B1(n4088), .Y(n904) );
  OAI211XLTS U782 ( .A0(n3366), .A1(n34), .B0(n947), .C0(n948), .Y(n2861) );
  OAI211XLTS U783 ( .A0(n3365), .A1(n32), .B0(n945), .C0(n946), .Y(n2862) );
  OAI211XLTS U784 ( .A0(n3365), .A1(n33), .B0(n943), .C0(n944), .Y(n2863) );
  OAI211XLTS U785 ( .A0(n3366), .A1(n35), .B0(n937), .C0(n938), .Y(n2864) );
  OAI211XLTS U786 ( .A0(n3366), .A1(n30), .B0(n951), .C0(n952), .Y(n2859) );
  OAI211XLTS U787 ( .A0(n3365), .A1(n31), .B0(n949), .C0(n950), .Y(n2860) );
  OAI211XLTS U788 ( .A0(n3432), .A1(n26), .B0(n930), .C0(n931), .Y(n2867) );
  OAI211XLTS U789 ( .A0(n3431), .A1(n24), .B0(n928), .C0(n929), .Y(n2868) );
  OAI211XLTS U790 ( .A0(n3431), .A1(n25), .B0(n926), .C0(n927), .Y(n2869) );
  OAI211XLTS U791 ( .A0(n3432), .A1(n22), .B0(n934), .C0(n935), .Y(n2865) );
  OAI211XLTS U792 ( .A0(n3431), .A1(n23), .B0(n932), .C0(n933), .Y(n2866) );
  OAI211XLTS U793 ( .A0(n3432), .A1(n27), .B0(n920), .C0(n921), .Y(n2870) );
  OAI211XLTS U794 ( .A0(n838), .A1(n618), .B0(n997), .C0(n998), .Y(n2843) );
  OAI211XLTS U795 ( .A0(n837), .A1(n617), .B0(n995), .C0(n996), .Y(n2844) );
  OAI211XLTS U796 ( .A0(n837), .A1(n616), .B0(n993), .C0(n994), .Y(n2845) );
  OAI211XLTS U797 ( .A0(n838), .A1(n620), .B0(n1001), .C0(n1002), .Y(n2841) );
  OAI211XLTS U798 ( .A0(n837), .A1(n619), .B0(n999), .C0(n1000), .Y(n2842) );
  OAI211XLTS U799 ( .A0(n838), .A1(n615), .B0(n987), .C0(n988), .Y(n2846) );
  OAI211XLTS U800 ( .A0(n3563), .A1(n587), .B0(n897), .C0(n898), .Y(n2879) );
  OAI211XLTS U801 ( .A0(n3562), .A1(n586), .B0(n893), .C0(n894), .Y(n2881) );
  OAI211XLTS U802 ( .A0(n3563), .A1(n627), .B0(n901), .C0(n902), .Y(n2877) );
  OAI211XLTS U803 ( .A0(n3562), .A1(n626), .B0(n899), .C0(n900), .Y(n2878) );
  OAI211XLTS U804 ( .A0(n3562), .A1(n625), .B0(n895), .C0(n896), .Y(n2880) );
  OAI211XLTS U805 ( .A0(n3563), .A1(n585), .B0(n887), .C0(n888), .Y(n2882) );
  OAI211XLTS U806 ( .A0(n3213), .A1(n3841), .B0(n1148), .C0(n1149), .Y(n2769)
         );
  OAI211XLTS U807 ( .A0(n3213), .A1(n3838), .B0(n1146), .C0(n1147), .Y(n2770)
         );
  OAI211XLTS U808 ( .A0(n3204), .A1(n3958), .B0(n1734), .C0(n1735), .Y(n2490)
         );
  OAI211XLTS U809 ( .A0(n3204), .A1(n3964), .B0(n1738), .C0(n1739), .Y(n2488)
         );
  OAI211XLTS U810 ( .A0(n3204), .A1(n3961), .B0(n1736), .C0(n1737), .Y(n2489)
         );
  OAI211XLTS U811 ( .A0(n3204), .A1(n3967), .B0(n1740), .C0(n1741), .Y(n2487)
         );
  OAI211XLTS U812 ( .A0(n3205), .A1(n3928), .B0(n1206), .C0(n1207), .Y(n2740)
         );
  OAI211XLTS U813 ( .A0(n3206), .A1(n3925), .B0(n1204), .C0(n1205), .Y(n2741)
         );
  OAI211XLTS U814 ( .A0(n3206), .A1(n3922), .B0(n1202), .C0(n1203), .Y(n2742)
         );
  OAI211XLTS U815 ( .A0(n3206), .A1(n3916), .B0(n1198), .C0(n1199), .Y(n2744)
         );
  OAI211XLTS U816 ( .A0(n3207), .A1(n3913), .B0(n1196), .C0(n1197), .Y(n2745)
         );
  OAI211XLTS U817 ( .A0(n3207), .A1(n3907), .B0(n1192), .C0(n1193), .Y(n2747)
         );
  OAI211XLTS U818 ( .A0(n3208), .A1(n3901), .B0(n1188), .C0(n1189), .Y(n2749)
         );
  OAI211XLTS U819 ( .A0(n3208), .A1(n3898), .B0(n1186), .C0(n1187), .Y(n2750)
         );
  OAI211XLTS U820 ( .A0(n3208), .A1(n3895), .B0(n1184), .C0(n1185), .Y(n2751)
         );
  OAI211XLTS U821 ( .A0(n3208), .A1(n3892), .B0(n1182), .C0(n1183), .Y(n2752)
         );
  OAI211XLTS U822 ( .A0(n3209), .A1(n3889), .B0(n1180), .C0(n1181), .Y(n2753)
         );
  OAI211XLTS U823 ( .A0(n3209), .A1(n3883), .B0(n1176), .C0(n1177), .Y(n2755)
         );
  OAI211XLTS U824 ( .A0(n3209), .A1(n3880), .B0(n1174), .C0(n1175), .Y(n2756)
         );
  OAI211XLTS U825 ( .A0(n3210), .A1(n3877), .B0(n1172), .C0(n1173), .Y(n2757)
         );
  OAI211XLTS U826 ( .A0(n3210), .A1(n3874), .B0(n1170), .C0(n1171), .Y(n2758)
         );
  OAI211XLTS U827 ( .A0(n3210), .A1(n3871), .B0(n1168), .C0(n1169), .Y(n2759)
         );
  OAI211XLTS U828 ( .A0(n3211), .A1(n3865), .B0(n1164), .C0(n1165), .Y(n2761)
         );
  OAI211XLTS U829 ( .A0(n3211), .A1(n3862), .B0(n1162), .C0(n1163), .Y(n2762)
         );
  OAI211XLTS U830 ( .A0(n3211), .A1(n3859), .B0(n1160), .C0(n1161), .Y(n2763)
         );
  OAI211XLTS U831 ( .A0(n3212), .A1(n3853), .B0(n1156), .C0(n1157), .Y(n2765)
         );
  OAI211XLTS U832 ( .A0(n3212), .A1(n3850), .B0(n1154), .C0(n1155), .Y(n2766)
         );
  OAI211XLTS U833 ( .A0(n3212), .A1(n3847), .B0(n1152), .C0(n1153), .Y(n2767)
         );
  OAI211XLTS U834 ( .A0(n3205), .A1(n3955), .B0(n1732), .C0(n1733), .Y(n2491)
         );
  OAI211XLTS U835 ( .A0(n3205), .A1(n3952), .B0(n1730), .C0(n1731), .Y(n2492)
         );
  OAI211XLTS U836 ( .A0(n3206), .A1(n3919), .B0(n1200), .C0(n1201), .Y(n2743)
         );
  OAI211XLTS U837 ( .A0(n3210), .A1(n3868), .B0(n1166), .C0(n1167), .Y(n2760)
         );
  OAI211XLTS U838 ( .A0(n3205), .A1(n3931), .B0(n1208), .C0(n1209), .Y(n2739)
         );
  OAI211XLTS U839 ( .A0(n3207), .A1(n3910), .B0(n1194), .C0(n1195), .Y(n2746)
         );
  OAI211XLTS U840 ( .A0(n3207), .A1(n3904), .B0(n1190), .C0(n1191), .Y(n2748)
         );
  OAI211XLTS U841 ( .A0(n3209), .A1(n3886), .B0(n1178), .C0(n1179), .Y(n2754)
         );
  OAI211XLTS U842 ( .A0(n3211), .A1(n3856), .B0(n1158), .C0(n1159), .Y(n2764)
         );
  OAI211XLTS U843 ( .A0(n3212), .A1(n3844), .B0(n1150), .C0(n1151), .Y(n2768)
         );
  OAI211XLTS U844 ( .A0(n3946), .A1(n3213), .B0(n982), .C0(n983), .Y(n2848) );
  OAI211XLTS U845 ( .A0(n3949), .A1(n3213), .B0(n984), .C0(n985), .Y(n2847) );
  OAI211XLTS U846 ( .A0(n3937), .A1(n3214), .B0(n976), .C0(n977), .Y(n2851) );
  OAI211XLTS U847 ( .A0(n3934), .A1(n3214), .B0(n971), .C0(n972), .Y(n2852) );
  OAI211XLTS U848 ( .A0(n3943), .A1(n3214), .B0(n980), .C0(n981), .Y(n2849) );
  OAI211XLTS U849 ( .A0(n3940), .A1(n3214), .B0(n978), .C0(n979), .Y(n2850) );
  OAI211XLTS U850 ( .A0(n4105), .A1(n3763), .B0(n968), .C0(n969), .Y(n2853) );
  OAI211XLTS U851 ( .A0(n4099), .A1(n3764), .B0(n964), .C0(n965), .Y(n2855) );
  OAI211XLTS U852 ( .A0(n4096), .A1(n3764), .B0(n962), .C0(n963), .Y(n2856) );
  OAI211XLTS U853 ( .A0(n4093), .A1(n3764), .B0(n960), .C0(n961), .Y(n2857) );
  OAI211XLTS U854 ( .A0(n4090), .A1(n3764), .B0(n953), .C0(n954), .Y(n2858) );
  OAI211XLTS U855 ( .A0(n4102), .A1(n3763), .B0(n966), .C0(n967), .Y(n2854) );
  OAI211XLTS U856 ( .A0(n2392), .A1(n3378), .B0(n1689), .C0(n1690), .Y(n2516)
         );
  INVXLTS U857 ( .A(n3380), .Y(n3378) );
  OAI211XLTS U858 ( .A0(n2896), .A1(n3368), .B0(n1691), .C0(n1692), .Y(n2515)
         );
  OAI211XLTS U859 ( .A0(n3181), .A1(n3376), .B0(n1334), .C0(n1335), .Y(n2676)
         );
  OAI211XLTS U860 ( .A0(n3163), .A1(n3376), .B0(n1330), .C0(n1331), .Y(n2678)
         );
  OAI211XLTS U861 ( .A0(n3152), .A1(n3375), .B0(n1328), .C0(n1329), .Y(n2679)
         );
  OAI211XLTS U862 ( .A0(n3145), .A1(n3375), .B0(n1326), .C0(n1327), .Y(n2680)
         );
  OAI211XLTS U863 ( .A0(n3132), .A1(n3375), .B0(n1324), .C0(n1325), .Y(n2681)
         );
  OAI211XLTS U864 ( .A0(n3127), .A1(n3375), .B0(n1322), .C0(n1323), .Y(n2682)
         );
  OAI211XLTS U865 ( .A0(n3116), .A1(n3374), .B0(n1320), .C0(n1321), .Y(n2683)
         );
  OAI211XLTS U866 ( .A0(n3073), .A1(n3373), .B0(n1310), .C0(n1311), .Y(n2688)
         );
  OAI211XLTS U867 ( .A0(n3028), .A1(n3372), .B0(n1300), .C0(n1301), .Y(n2693)
         );
  OAI211XLTS U868 ( .A0(n2988), .A1(n3371), .B0(n1292), .C0(n1293), .Y(n2697)
         );
  OAI211XLTS U869 ( .A0(n2970), .A1(n3370), .B0(n1288), .C0(n1289), .Y(n2699)
         );
  OAI211XLTS U870 ( .A0(n2954), .A1(n3370), .B0(n1284), .C0(n1285), .Y(n2701)
         );
  OAI211XLTS U871 ( .A0(n2943), .A1(n3370), .B0(n1282), .C0(n1283), .Y(n2702)
         );
  OAI211XLTS U872 ( .A0(n2927), .A1(n3369), .B0(n1278), .C0(n1279), .Y(n2704)
         );
  OAI211XLTS U873 ( .A0(n3189), .A1(n3376), .B0(n1336), .C0(n1337), .Y(n2675)
         );
  OAI211XLTS U874 ( .A0(n3165), .A1(n3376), .B0(n1332), .C0(n1333), .Y(n2677)
         );
  OAI211XLTS U875 ( .A0(n3106), .A1(n3374), .B0(n1318), .C0(n1319), .Y(n2684)
         );
  OAI211XLTS U876 ( .A0(n3095), .A1(n3374), .B0(n1316), .C0(n1317), .Y(n2685)
         );
  OAI211XLTS U877 ( .A0(n3086), .A1(n3374), .B0(n1314), .C0(n1315), .Y(n2686)
         );
  OAI211XLTS U878 ( .A0(n3081), .A1(n3373), .B0(n1312), .C0(n1313), .Y(n2687)
         );
  OAI211XLTS U879 ( .A0(n3054), .A1(n3373), .B0(n1306), .C0(n1307), .Y(n2690)
         );
  OAI211XLTS U880 ( .A0(n3016), .A1(n3371), .B0(n1298), .C0(n1299), .Y(n2694)
         );
  OAI211XLTS U881 ( .A0(n3005), .A1(n3371), .B0(n1296), .C0(n1297), .Y(n2695)
         );
  OAI211XLTS U882 ( .A0(n2998), .A1(n3371), .B0(n1294), .C0(n1295), .Y(n2696)
         );
  OAI211XLTS U883 ( .A0(n2982), .A1(n3370), .B0(n1290), .C0(n1291), .Y(n2698)
         );
  OAI211XLTS U884 ( .A0(n2960), .A1(n3372), .B0(n1286), .C0(n1287), .Y(n2700)
         );
  OAI211XLTS U885 ( .A0(n2919), .A1(n3369), .B0(n1276), .C0(n1277), .Y(n2705)
         );
  OAI211XLTS U886 ( .A0(n2908), .A1(n3369), .B0(n1274), .C0(n1275), .Y(n2706)
         );
  OAI211XLTS U887 ( .A0(n3058), .A1(n3373), .B0(n1308), .C0(n1309), .Y(n2689)
         );
  OAI211XLTS U888 ( .A0(n3040), .A1(n3372), .B0(n1304), .C0(n1305), .Y(n2691)
         );
  OAI211XLTS U889 ( .A0(n3031), .A1(n3372), .B0(n1302), .C0(n1303), .Y(n2692)
         );
  OAI211XLTS U890 ( .A0(n2932), .A1(n3369), .B0(n1280), .C0(n1281), .Y(n2703)
         );
  OAI211XLTS U891 ( .A0(n2383), .A1(n3377), .B0(n1687), .C0(n1688), .Y(n2517)
         );
  OAI211XLTS U892 ( .A0(n2378), .A1(n3377), .B0(n1685), .C0(n1686), .Y(n2518)
         );
  OAI211XLTS U893 ( .A0(n2365), .A1(n3377), .B0(n1683), .C0(n1684), .Y(n2519)
         );
  OAI211XLTS U894 ( .A0(n2360), .A1(n3377), .B0(n1681), .C0(n1682), .Y(n2520)
         );
  OAI211XLTS U895 ( .A0(n2893), .A1(n3434), .B0(n1667), .C0(n1668), .Y(n2529)
         );
  OAI211XLTS U896 ( .A0(n3186), .A1(n3442), .B0(n1400), .C0(n1401), .Y(n2643)
         );
  OAI211XLTS U897 ( .A0(n3051), .A1(n3439), .B0(n1370), .C0(n1371), .Y(n2658)
         );
  OAI211XLTS U898 ( .A0(n3046), .A1(n3438), .B0(n1368), .C0(n1369), .Y(n2659)
         );
  OAI211XLTS U899 ( .A0(n3008), .A1(n3437), .B0(n1360), .C0(n1361), .Y(n2663)
         );
  OAI211XLTS U900 ( .A0(n2916), .A1(n3435), .B0(n1340), .C0(n1341), .Y(n2673)
         );
  OAI211XLTS U901 ( .A0(n3178), .A1(n3442), .B0(n1398), .C0(n1399), .Y(n2644)
         );
  OAI211XLTS U902 ( .A0(n3167), .A1(n3442), .B0(n1396), .C0(n1397), .Y(n2645)
         );
  OAI211XLTS U903 ( .A0(n3156), .A1(n3442), .B0(n1394), .C0(n1395), .Y(n2646)
         );
  OAI211XLTS U904 ( .A0(n3153), .A1(n3441), .B0(n1392), .C0(n1393), .Y(n2647)
         );
  OAI211XLTS U905 ( .A0(n3144), .A1(n3441), .B0(n1390), .C0(n1391), .Y(n2648)
         );
  OAI211XLTS U906 ( .A0(n3129), .A1(n3441), .B0(n1388), .C0(n1389), .Y(n2649)
         );
  OAI211XLTS U907 ( .A0(n3122), .A1(n3441), .B0(n1386), .C0(n1387), .Y(n2650)
         );
  OAI211XLTS U908 ( .A0(n3115), .A1(n3440), .B0(n1384), .C0(n1385), .Y(n2651)
         );
  OAI211XLTS U909 ( .A0(n3104), .A1(n3440), .B0(n1382), .C0(n1383), .Y(n2652)
         );
  OAI211XLTS U910 ( .A0(n3097), .A1(n3440), .B0(n1380), .C0(n1381), .Y(n2653)
         );
  OAI211XLTS U911 ( .A0(n3090), .A1(n3440), .B0(n1378), .C0(n1379), .Y(n2654)
         );
  OAI211XLTS U912 ( .A0(n3077), .A1(n3439), .B0(n1376), .C0(n1377), .Y(n2655)
         );
  OAI211XLTS U913 ( .A0(n3070), .A1(n3439), .B0(n1374), .C0(n1375), .Y(n2656)
         );
  OAI211XLTS U914 ( .A0(n3059), .A1(n3439), .B0(n1372), .C0(n1373), .Y(n2657)
         );
  OAI211XLTS U915 ( .A0(n3036), .A1(n3438), .B0(n1366), .C0(n1367), .Y(n2660)
         );
  OAI211XLTS U916 ( .A0(n3023), .A1(n3438), .B0(n1364), .C0(n1365), .Y(n2661)
         );
  OAI211XLTS U917 ( .A0(n3014), .A1(n3437), .B0(n1362), .C0(n1363), .Y(n2662)
         );
  OAI211XLTS U918 ( .A0(n3000), .A1(n3437), .B0(n1358), .C0(n1359), .Y(n2664)
         );
  OAI211XLTS U919 ( .A0(n2989), .A1(n3437), .B0(n1356), .C0(n1357), .Y(n2665)
         );
  OAI211XLTS U920 ( .A0(n2978), .A1(n3436), .B0(n1354), .C0(n1355), .Y(n2666)
         );
  OAI211XLTS U921 ( .A0(n2969), .A1(n3436), .B0(n1352), .C0(n1353), .Y(n2667)
         );
  OAI211XLTS U922 ( .A0(n2962), .A1(n3438), .B0(n1350), .C0(n1351), .Y(n2668)
         );
  OAI211XLTS U923 ( .A0(n2949), .A1(n3436), .B0(n1348), .C0(n1349), .Y(n2669)
         );
  OAI211XLTS U924 ( .A0(n2942), .A1(n3436), .B0(n1346), .C0(n1347), .Y(n2670)
         );
  OAI211XLTS U925 ( .A0(n2931), .A1(n3435), .B0(n1344), .C0(n1345), .Y(n2671)
         );
  OAI211XLTS U926 ( .A0(n2926), .A1(n3435), .B0(n1342), .C0(n1343), .Y(n2672)
         );
  OAI211XLTS U927 ( .A0(n2904), .A1(n3435), .B0(n1338), .C0(n1339), .Y(n2674)
         );
  OAI211XLTS U928 ( .A0(n2382), .A1(n3443), .B0(n1663), .C0(n1664), .Y(n2531)
         );
  OAI211XLTS U929 ( .A0(n2373), .A1(n3443), .B0(n1661), .C0(n1662), .Y(n2532)
         );
  OAI211XLTS U930 ( .A0(n2364), .A1(n3443), .B0(n1659), .C0(n1660), .Y(n2533)
         );
  OAI211XLTS U931 ( .A0(n2357), .A1(n3443), .B0(n1657), .C0(n1658), .Y(n2534)
         );
  OAI211XLTS U932 ( .A0(n2391), .A1(n3444), .B0(n1665), .C0(n1666), .Y(n2530)
         );
  INVXLTS U933 ( .A(n3445), .Y(n3444) );
  OAI211XLTS U934 ( .A0(n3154), .A1(n847), .B0(n1136), .C0(n1137), .Y(n2775)
         );
  OAI211XLTS U935 ( .A0(n3105), .A1(n846), .B0(n1126), .C0(n1127), .Y(n2780)
         );
  OAI211XLTS U936 ( .A0(n3089), .A1(n846), .B0(n1122), .C0(n1123), .Y(n2782)
         );
  OAI211XLTS U937 ( .A0(n3078), .A1(n845), .B0(n1120), .C0(n1121), .Y(n2783)
         );
  OAI211XLTS U938 ( .A0(n2995), .A1(n843), .B0(n1102), .C0(n1103), .Y(n2792)
         );
  OAI211XLTS U939 ( .A0(n2981), .A1(n842), .B0(n1098), .C0(n1099), .Y(n2794)
         );
  OAI211XLTS U940 ( .A0(n2956), .A1(n842), .B0(n1092), .C0(n1093), .Y(n2797)
         );
  OAI211XLTS U941 ( .A0(n2929), .A1(n841), .B0(n1086), .C0(n1087), .Y(n2800)
         );
  OAI211XLTS U942 ( .A0(n3183), .A1(n848), .B0(n1144), .C0(n1145), .Y(n2771)
         );
  OAI211XLTS U943 ( .A0(n3174), .A1(n848), .B0(n1142), .C0(n1143), .Y(n2772)
         );
  OAI211XLTS U944 ( .A0(n3169), .A1(n848), .B0(n1140), .C0(n1141), .Y(n2773)
         );
  OAI211XLTS U945 ( .A0(n3162), .A1(n848), .B0(n1138), .C0(n1139), .Y(n2774)
         );
  OAI211XLTS U946 ( .A0(n3131), .A1(n847), .B0(n1132), .C0(n1133), .Y(n2777)
         );
  OAI211XLTS U947 ( .A0(n3126), .A1(n847), .B0(n1130), .C0(n1131), .Y(n2778)
         );
  OAI211XLTS U948 ( .A0(n3117), .A1(n846), .B0(n1128), .C0(n1129), .Y(n2779)
         );
  OAI211XLTS U949 ( .A0(n3099), .A1(n846), .B0(n1124), .C0(n1125), .Y(n2781)
         );
  OAI211XLTS U950 ( .A0(n3066), .A1(n845), .B0(n1118), .C0(n1119), .Y(n2784)
         );
  OAI211XLTS U951 ( .A0(n3063), .A1(n845), .B0(n1116), .C0(n1117), .Y(n2785)
         );
  OAI211XLTS U952 ( .A0(n3048), .A1(n845), .B0(n1114), .C0(n1115), .Y(n2786)
         );
  OAI211XLTS U953 ( .A0(n3041), .A1(n844), .B0(n1112), .C0(n1113), .Y(n2787)
         );
  OAI211XLTS U954 ( .A0(n3034), .A1(n844), .B0(n1110), .C0(n1111), .Y(n2788)
         );
  OAI211XLTS U955 ( .A0(n3021), .A1(n844), .B0(n1108), .C0(n1109), .Y(n2789)
         );
  OAI211XLTS U956 ( .A0(n3012), .A1(n843), .B0(n1106), .C0(n1107), .Y(n2790)
         );
  OAI211XLTS U957 ( .A0(n3009), .A1(n843), .B0(n1104), .C0(n1105), .Y(n2791)
         );
  OAI211XLTS U958 ( .A0(n2991), .A1(n843), .B0(n1100), .C0(n1101), .Y(n2793)
         );
  OAI211XLTS U959 ( .A0(n2967), .A1(n842), .B0(n1096), .C0(n1097), .Y(n2795)
         );
  OAI211XLTS U960 ( .A0(n2964), .A1(n844), .B0(n1094), .C0(n1095), .Y(n2796)
         );
  OAI211XLTS U961 ( .A0(n2940), .A1(n842), .B0(n1090), .C0(n1091), .Y(n2798)
         );
  OAI211XLTS U962 ( .A0(n2935), .A1(n841), .B0(n1088), .C0(n1089), .Y(n2799)
         );
  OAI211XLTS U963 ( .A0(n2917), .A1(n841), .B0(n1084), .C0(n1085), .Y(n2801)
         );
  OAI211XLTS U964 ( .A0(n2905), .A1(n841), .B0(n1082), .C0(n1083), .Y(n2802)
         );
  OAI211XLTS U965 ( .A0(n2384), .A1(n849), .B0(n1757), .C0(n1758), .Y(n2475)
         );
  OAI211XLTS U966 ( .A0(n2371), .A1(n849), .B0(n1755), .C0(n1756), .Y(n2476)
         );
  OAI211XLTS U967 ( .A0(n2362), .A1(n849), .B0(n1753), .C0(n1754), .Y(n2477)
         );
  OAI211XLTS U968 ( .A0(n2353), .A1(n849), .B0(n1751), .C0(n1752), .Y(n2478)
         );
  OAI211XLTS U969 ( .A0(n2387), .A1(n716), .B0(n1638), .C0(n1639), .Y(n2545)
         );
  OAI211XLTS U970 ( .A0(n2376), .A1(n716), .B0(n1636), .C0(n1637), .Y(n2546)
         );
  OAI211XLTS U971 ( .A0(n2367), .A1(n715), .B0(n1634), .C0(n1635), .Y(n2547)
         );
  OAI211XLTS U972 ( .A0(n2358), .A1(n715), .B0(n1632), .C0(n1633), .Y(n2548)
         );
  OAI211XLTS U973 ( .A0(n3168), .A1(n714), .B0(n1461), .C0(n1462), .Y(n2613)
         );
  OAI211XLTS U974 ( .A0(n3118), .A1(n712), .B0(n1449), .C0(n1450), .Y(n2619)
         );
  OAI211XLTS U975 ( .A0(n3098), .A1(n711), .B0(n1445), .C0(n1446), .Y(n2621)
         );
  OAI211XLTS U976 ( .A0(n3091), .A1(n711), .B0(n1443), .C0(n1444), .Y(n2622)
         );
  OAI211XLTS U977 ( .A0(n3024), .A1(n707), .B0(n1429), .C0(n1430), .Y(n2629)
         );
  OAI211XLTS U978 ( .A0(n3013), .A1(n707), .B0(n1427), .C0(n1428), .Y(n2630)
         );
  OAI211XLTS U979 ( .A0(n3001), .A1(n706), .B0(n1423), .C0(n1424), .Y(n2632)
         );
  OAI211XLTS U980 ( .A0(n2965), .A1(n705), .B0(n1415), .C0(n1416), .Y(n2636)
         );
  OAI211XLTS U981 ( .A0(n2918), .A1(n704), .B0(n1405), .C0(n1406), .Y(n2641)
         );
  AOI22XLTS U982 ( .A0(n4151), .A1(n3480), .B0(n4307), .B1(n3739), .Y(n1405)
         );
  OAI211XLTS U983 ( .A0(n3187), .A1(n715), .B0(n1465), .C0(n1466), .Y(n2611)
         );
  OAI211XLTS U984 ( .A0(n3176), .A1(n715), .B0(n1463), .C0(n1464), .Y(n2612)
         );
  OAI211XLTS U985 ( .A0(n3160), .A1(n714), .B0(n1459), .C0(n1460), .Y(n2614)
         );
  OAI211XLTS U986 ( .A0(n3151), .A1(n714), .B0(n1457), .C0(n1458), .Y(n2615)
         );
  OAI211XLTS U987 ( .A0(n3140), .A1(n714), .B0(n1455), .C0(n1456), .Y(n2616)
         );
  OAI211XLTS U988 ( .A0(n3120), .A1(n712), .B0(n1451), .C0(n1452), .Y(n2618)
         );
  OAI211XLTS U989 ( .A0(n3102), .A1(n712), .B0(n1447), .C0(n1448), .Y(n2620)
         );
  OAI211XLTS U990 ( .A0(n3079), .A1(n711), .B0(n1441), .C0(n1442), .Y(n2623)
         );
  OAI211XLTS U991 ( .A0(n3057), .A1(n708), .B0(n1437), .C0(n1438), .Y(n2625)
         );
  OAI211XLTS U992 ( .A0(n3052), .A1(n708), .B0(n1435), .C0(n1436), .Y(n2626)
         );
  OAI211XLTS U993 ( .A0(n3039), .A1(n708), .B0(n1433), .C0(n1434), .Y(n2627)
         );
  OAI211XLTS U994 ( .A0(n3032), .A1(n707), .B0(n1431), .C0(n1432), .Y(n2628)
         );
  OAI211XLTS U995 ( .A0(n3003), .A1(n707), .B0(n1425), .C0(n1426), .Y(n2631)
         );
  OAI211XLTS U996 ( .A0(n2987), .A1(n706), .B0(n1421), .C0(n1422), .Y(n2633)
         );
  OAI211XLTS U997 ( .A0(n2976), .A1(n706), .B0(n1419), .C0(n1420), .Y(n2634)
         );
  OAI211XLTS U998 ( .A0(n2971), .A1(n706), .B0(n1417), .C0(n1418), .Y(n2635)
         );
  OAI211XLTS U999 ( .A0(n2953), .A1(n705), .B0(n1413), .C0(n1414), .Y(n2637)
         );
  OAI211XLTS U1000 ( .A0(n2937), .A1(n705), .B0(n1409), .C0(n1410), .Y(n2639)
         );
  OAI211XLTS U1001 ( .A0(n2922), .A1(n704), .B0(n1407), .C0(n1408), .Y(n2640)
         );
  OAI211XLTS U1002 ( .A0(n2906), .A1(n711), .B0(n1403), .C0(n1404), .Y(n2642)
         );
  AOI22XLTS U1003 ( .A0(n4148), .A1(n3480), .B0(n4304), .B1(n454), .Y(n1403)
         );
  OAI211XLTS U1004 ( .A0(n3130), .A1(n712), .B0(n1453), .C0(n1454), .Y(n2617)
         );
  OAI211XLTS U1005 ( .A0(n3067), .A1(n708), .B0(n1439), .C0(n1440), .Y(n2624)
         );
  OAI211XLTS U1006 ( .A0(n2941), .A1(n705), .B0(n1411), .C0(n1412), .Y(n2638)
         );
  OAI211XLTS U1007 ( .A0(n2894), .A1(n704), .B0(n1642), .C0(n1643), .Y(n2543)
         );
  OAI211XLTS U1008 ( .A0(n2390), .A1(n716), .B0(n1640), .C0(n1641), .Y(n2544)
         );
  OAI211XLTS U1009 ( .A0(n2891), .A1(n3565), .B0(n1616), .C0(n1617), .Y(n2557)
         );
  OAI211XLTS U1010 ( .A0(n3185), .A1(n3573), .B0(n1529), .C0(n1530), .Y(n2579)
         );
  OAI211XLTS U1011 ( .A0(n3180), .A1(n3573), .B0(n1527), .C0(n1528), .Y(n2580)
         );
  OAI211XLTS U1012 ( .A0(n3171), .A1(n3573), .B0(n1525), .C0(n1526), .Y(n2581)
         );
  OAI211XLTS U1013 ( .A0(n3158), .A1(n3573), .B0(n1523), .C0(n1524), .Y(n2582)
         );
  OAI211XLTS U1014 ( .A0(n3149), .A1(n3572), .B0(n1521), .C0(n1522), .Y(n2583)
         );
  OAI211XLTS U1015 ( .A0(n3142), .A1(n3572), .B0(n1519), .C0(n1520), .Y(n2584)
         );
  OAI211XLTS U1016 ( .A0(n3133), .A1(n3572), .B0(n1517), .C0(n1518), .Y(n2585)
         );
  OAI211XLTS U1017 ( .A0(n3124), .A1(n3572), .B0(n1515), .C0(n1516), .Y(n2586)
         );
  OAI211XLTS U1018 ( .A0(n3113), .A1(n3571), .B0(n1513), .C0(n1514), .Y(n2587)
         );
  OAI211XLTS U1019 ( .A0(n3108), .A1(n3571), .B0(n1511), .C0(n1512), .Y(n2588)
         );
  OAI211XLTS U1020 ( .A0(n3093), .A1(n3571), .B0(n1509), .C0(n1510), .Y(n2589)
         );
  OAI211XLTS U1021 ( .A0(n3088), .A1(n3571), .B0(n1507), .C0(n1508), .Y(n2590)
         );
  OAI211XLTS U1022 ( .A0(n3075), .A1(n3570), .B0(n1505), .C0(n1506), .Y(n2591)
         );
  OAI211XLTS U1023 ( .A0(n3072), .A1(n3570), .B0(n1503), .C0(n1504), .Y(n2592)
         );
  OAI211XLTS U1024 ( .A0(n3061), .A1(n3570), .B0(n1501), .C0(n1502), .Y(n2593)
         );
  OAI211XLTS U1025 ( .A0(n3050), .A1(n3570), .B0(n1499), .C0(n1500), .Y(n2594)
         );
  OAI211XLTS U1026 ( .A0(n3045), .A1(n3569), .B0(n1497), .C0(n1498), .Y(n2595)
         );
  OAI211XLTS U1027 ( .A0(n3030), .A1(n3569), .B0(n1495), .C0(n1496), .Y(n2596)
         );
  OAI211XLTS U1028 ( .A0(n3027), .A1(n3569), .B0(n1493), .C0(n1494), .Y(n2597)
         );
  OAI211XLTS U1029 ( .A0(n3018), .A1(n3568), .B0(n1491), .C0(n1492), .Y(n2598)
         );
  OAI211XLTS U1030 ( .A0(n3007), .A1(n3568), .B0(n1489), .C0(n1490), .Y(n2599)
         );
  OAI211XLTS U1031 ( .A0(n2994), .A1(n3568), .B0(n1487), .C0(n1488), .Y(n2600)
         );
  OAI211XLTS U1032 ( .A0(n2985), .A1(n3568), .B0(n1485), .C0(n1486), .Y(n2601)
         );
  OAI211XLTS U1033 ( .A0(n2980), .A1(n3567), .B0(n1483), .C0(n1484), .Y(n2602)
         );
  OAI211XLTS U1034 ( .A0(n2973), .A1(n3567), .B0(n1481), .C0(n1482), .Y(n2603)
         );
  OAI211XLTS U1035 ( .A0(n2958), .A1(n3569), .B0(n1479), .C0(n1480), .Y(n2604)
         );
  OAI211XLTS U1036 ( .A0(n2955), .A1(n3567), .B0(n1477), .C0(n1478), .Y(n2605)
         );
  OAI211XLTS U1037 ( .A0(n2946), .A1(n3567), .B0(n1475), .C0(n1476), .Y(n2606)
         );
  OAI211XLTS U1038 ( .A0(n2933), .A1(n3566), .B0(n1473), .C0(n1474), .Y(n2607)
         );
  OAI211XLTS U1039 ( .A0(n2928), .A1(n3566), .B0(n1471), .C0(n1472), .Y(n2608)
         );
  OAI211XLTS U1040 ( .A0(n2915), .A1(n3566), .B0(n1469), .C0(n1470), .Y(n2609)
         );
  OAI211XLTS U1041 ( .A0(n2910), .A1(n3566), .B0(n1467), .C0(n1468), .Y(n2610)
         );
  OAI211XLTS U1042 ( .A0(n2354), .A1(n3574), .B0(n1606), .C0(n1607), .Y(n2562)
         );
  OAI211XLTS U1043 ( .A0(n2386), .A1(n3574), .B0(n1612), .C0(n1613), .Y(n2559)
         );
  OAI211XLTS U1044 ( .A0(n2375), .A1(n3574), .B0(n1610), .C0(n1611), .Y(n2560)
         );
  OAI211XLTS U1045 ( .A0(n2368), .A1(n3574), .B0(n1608), .C0(n1609), .Y(n2561)
         );
  OAI211XLTS U1046 ( .A0(n2396), .A1(n3575), .B0(n1614), .C0(n1615), .Y(n2558)
         );
  INVXLTS U1047 ( .A(n3577), .Y(n3575) );
  OAI211XLTS U1048 ( .A0(n3757), .A1(n4120), .B0(n1711), .C0(n1712), .Y(n2502)
         );
  OAI211XLTS U1049 ( .A0(n3757), .A1(n4117), .B0(n1709), .C0(n1710), .Y(n2503)
         );
  OAI211XLTS U1050 ( .A0(n3757), .A1(n4114), .B0(n1707), .C0(n1708), .Y(n2504)
         );
  OAI211XLTS U1051 ( .A0(n3757), .A1(n4123), .B0(n1713), .C0(n1714), .Y(n2501)
         );
  OAI211XLTS U1052 ( .A0(n3763), .A1(n3997), .B0(n1212), .C0(n1213), .Y(n2737)
         );
  OAI211XLTS U1053 ( .A0(n3763), .A1(n3994), .B0(n1210), .C0(n1211), .Y(n2738)
         );
  OAI211XLTS U1054 ( .A0(n3765), .A1(n4111), .B0(n1705), .C0(n1706), .Y(n2505)
         );
  OAI211XLTS U1055 ( .A0(n3767), .A1(n4108), .B0(n1703), .C0(n1704), .Y(n2506)
         );
  OAI211XLTS U1056 ( .A0(n3766), .A1(n4087), .B0(n1272), .C0(n1273), .Y(n2707)
         );
  OAI211XLTS U1057 ( .A0(n3770), .A1(n4084), .B0(n1270), .C0(n1271), .Y(n2708)
         );
  OAI211XLTS U1058 ( .A0(n3769), .A1(n4081), .B0(n1268), .C0(n1269), .Y(n2709)
         );
  OAI211XLTS U1059 ( .A0(n3765), .A1(n4078), .B0(n1266), .C0(n1267), .Y(n2710)
         );
  OAI211XLTS U1060 ( .A0(n3768), .A1(n4075), .B0(n1264), .C0(n1265), .Y(n2711)
         );
  OAI211XLTS U1061 ( .A0(n3769), .A1(n4072), .B0(n1262), .C0(n1263), .Y(n2712)
         );
  OAI211XLTS U1062 ( .A0(n3767), .A1(n4066), .B0(n1258), .C0(n1259), .Y(n2714)
         );
  OAI211XLTS U1063 ( .A0(n3768), .A1(n4060), .B0(n1254), .C0(n1255), .Y(n2716)
         );
  OAI211XLTS U1064 ( .A0(n3758), .A1(n4057), .B0(n1252), .C0(n1253), .Y(n2717)
         );
  OAI211XLTS U1065 ( .A0(n3758), .A1(n4051), .B0(n1248), .C0(n1249), .Y(n2719)
         );
  OAI211XLTS U1066 ( .A0(n3759), .A1(n4045), .B0(n1244), .C0(n1245), .Y(n2721)
         );
  OAI211XLTS U1067 ( .A0(n3759), .A1(n4042), .B0(n1242), .C0(n1243), .Y(n2722)
         );
  OAI211XLTS U1068 ( .A0(n3759), .A1(n4036), .B0(n1238), .C0(n1239), .Y(n2724)
         );
  OAI211XLTS U1069 ( .A0(n3760), .A1(n4030), .B0(n1234), .C0(n1235), .Y(n2726)
         );
  OAI211XLTS U1070 ( .A0(n3760), .A1(n4027), .B0(n1232), .C0(n1233), .Y(n2727)
         );
  OAI211XLTS U1071 ( .A0(n3760), .A1(n4024), .B0(n1230), .C0(n1231), .Y(n2728)
         );
  OAI211XLTS U1072 ( .A0(n3761), .A1(n4021), .B0(n1228), .C0(n1229), .Y(n2729)
         );
  OAI211XLTS U1073 ( .A0(n3761), .A1(n4018), .B0(n1226), .C0(n1227), .Y(n2730)
         );
  OAI211XLTS U1074 ( .A0(n3761), .A1(n4012), .B0(n1222), .C0(n1223), .Y(n2732)
         );
  OAI211XLTS U1075 ( .A0(n3762), .A1(n4003), .B0(n1216), .C0(n1217), .Y(n2735)
         );
  OAI211XLTS U1076 ( .A0(n3766), .A1(n4069), .B0(n1260), .C0(n1261), .Y(n2713)
         );
  OAI211XLTS U1077 ( .A0(n3768), .A1(n4063), .B0(n1256), .C0(n1257), .Y(n2715)
         );
  OAI211XLTS U1078 ( .A0(n3758), .A1(n4054), .B0(n1250), .C0(n1251), .Y(n2718)
         );
  OAI211XLTS U1079 ( .A0(n3758), .A1(n4048), .B0(n1246), .C0(n1247), .Y(n2720)
         );
  OAI211XLTS U1080 ( .A0(n3759), .A1(n4039), .B0(n1240), .C0(n1241), .Y(n2723)
         );
  OAI211XLTS U1081 ( .A0(n3760), .A1(n4033), .B0(n1236), .C0(n1237), .Y(n2725)
         );
  OAI211XLTS U1082 ( .A0(n3762), .A1(n4009), .B0(n1220), .C0(n1221), .Y(n2733)
         );
  OAI211XLTS U1083 ( .A0(n3762), .A1(n4006), .B0(n1218), .C0(n1219), .Y(n2734)
         );
  OAI211XLTS U1084 ( .A0(n3762), .A1(n4000), .B0(n1214), .C0(n1215), .Y(n2736)
         );
  OAI211XLTS U1085 ( .A0(n3761), .A1(n4015), .B0(n1224), .C0(n1225), .Y(n2731)
         );
  OAI2BB1XLTS U1086 ( .A0N(n2278), .A1N(n2250), .B0(n2279), .Y(n2267) );
  AOI32XLTS U1087 ( .A0(n168), .A1(n825), .A2(n233), .B0(n169), .B1(n2280), 
        .Y(n2279) );
  XNOR2XLTS U1088 ( .A(n872), .B(n720), .Y(n2280) );
  AOI32XLTS U1089 ( .A0(n163), .A1(n1551), .A2(n1552), .B0(n591), .B1(n152), 
        .Y(n2570) );
  AOI22XLTS U1090 ( .A0(n3826), .A1(n1553), .B0(n3821), .B1(n1554), .Y(n1552)
         );
  AOI32XLTS U1091 ( .A0(n213), .A1(n1572), .A2(n1573), .B0(n3379), .B1(n151), 
        .Y(n2567) );
  AOI21XLTS U1092 ( .A0(n3833), .A1(n1574), .B0(n1575), .Y(n1573) );
  AOI32XLTS U1093 ( .A0(n212), .A1(n1558), .A2(n1559), .B0(n729), .B1(n28), 
        .Y(n2569) );
  NAND2XLTS U1094 ( .A(n3820), .B(n1563), .Y(n1558) );
  NAND2XLTS U1095 ( .A(n219), .B(selectBit_EAST), .Y(n1679) );
  AOI22XLTS U1096 ( .A0(n1599), .A1(n1600), .B0(n238), .B1(n583), .Y(n2563) );
  AOI31XLTS U1097 ( .A0(n1601), .A1(n215), .A2(readIn_SOUTH), .B0(n1603), .Y(
        n1600) );
  AOI21XLTS U1098 ( .A0(n3833), .A1(n1605), .B0(n498), .Y(n1599) );
  OAI32XLTS U1099 ( .A0(n3828), .A1(n518), .A2(n227), .B0(n1604), .B1(n3822), 
        .Y(n1603) );
  NAND3XLTS U1100 ( .A(n2251), .B(n718), .C(n170), .Y(n1813) );
  NAND3XLTS U1101 ( .A(n251), .B(n2250), .C(n254), .Y(n1812) );
  NAND4XLTS U1102 ( .A(n169), .B(n251), .C(n872), .D(n255), .Y(n1811) );
  NAND4XLTS U1103 ( .A(n168), .B(n251), .C(n255), .D(n825), .Y(n1815) );
  CLKBUFX2TS U1104 ( .A(n5323), .Y(n594) );
  CLKBUFX2TS U1105 ( .A(n5327), .Y(n595) );
  NOR3X1TS U1106 ( .A(n237), .B(n8), .C(n320), .Y(n1833) );
  OAI2BB2XLTS U1107 ( .B0(n620), .B1(n3610), .A0N(
        \requesterAddressbuffer[2][5] ), .A1N(n229), .Y(n1991) );
  OAI2BB2XLTS U1108 ( .B0(n619), .B1(n3610), .A0N(
        \requesterAddressbuffer[2][4] ), .A1N(n229), .Y(n1983) );
  OAI2BB2XLTS U1109 ( .B0(n617), .B1(n3609), .A0N(
        \requesterAddressbuffer[2][2] ), .A1N(n228), .Y(n1967) );
  OAI2BB2XLTS U1110 ( .B0(n616), .B1(n3609), .A0N(
        \requesterAddressbuffer[2][1] ), .A1N(n228), .Y(n1959) );
  OAI2BB2XLTS U1111 ( .B0(n618), .B1(n3609), .A0N(
        \requesterAddressbuffer[2][3] ), .A1N(n229), .Y(n1975) );
  OAI2BB2XLTS U1112 ( .B0(n615), .B1(n3609), .A0N(
        \requesterAddressbuffer[2][0] ), .A1N(n229), .Y(n1951) );
  NAND2X1TS U1113 ( .A(n10), .B(n319), .Y(n881) );
  CLKBUFX2TS U1114 ( .A(n3769), .Y(n3758) );
  CLKBUFX2TS U1115 ( .A(n3767), .Y(n3759) );
  CLKBUFX2TS U1116 ( .A(n3767), .Y(n3760) );
  CLKBUFX2TS U1117 ( .A(n3766), .Y(n3762) );
  CLKBUFX2TS U1118 ( .A(n3766), .Y(n3761) );
  CLKBUFX2TS U1119 ( .A(n3765), .Y(n3763) );
  CLKBUFX2TS U1120 ( .A(n3765), .Y(n3764) );
  CLKBUFX2TS U1121 ( .A(n3770), .Y(n3765) );
  CLKBUFX2TS U1122 ( .A(n3770), .Y(n3767) );
  CLKBUFX2TS U1123 ( .A(n3770), .Y(n3766) );
  CLKBUFX2TS U1124 ( .A(n3732), .Y(n3726) );
  CLKBUFX2TS U1125 ( .A(n3730), .Y(n3722) );
  CLKBUFX2TS U1126 ( .A(n3730), .Y(n3721) );
  CLKBUFX2TS U1127 ( .A(n3731), .Y(n3720) );
  CLKBUFX2TS U1128 ( .A(n3729), .Y(n3724) );
  CLKBUFX2TS U1129 ( .A(n3730), .Y(n3725) );
  CLKBUFX2TS U1130 ( .A(n3729), .Y(n3723) );
  CLKBUFX2TS U1131 ( .A(n3731), .Y(n3719) );
  CLKBUFX2TS U1132 ( .A(n3733), .Y(n3727) );
  CLKBUFX2TS U1133 ( .A(n3813), .Y(n3804) );
  CLKBUFX2TS U1134 ( .A(n3813), .Y(n3805) );
  CLKBUFX2TS U1135 ( .A(n3812), .Y(n3806) );
  CLKBUFX2TS U1136 ( .A(n3812), .Y(n3807) );
  CLKBUFX2TS U1137 ( .A(n3816), .Y(n3808) );
  CLKBUFX2TS U1138 ( .A(n3768), .Y(n3757) );
  CLKBUFX2TS U1139 ( .A(n3769), .Y(n3768) );
  CLKBUFX2TS U1140 ( .A(n3733), .Y(n3728) );
  CLKBUFX2TS U1141 ( .A(n3740), .Y(n3738) );
  CLKBUFX2TS U1142 ( .A(n3741), .Y(n3736) );
  CLKBUFX2TS U1143 ( .A(n3732), .Y(n3730) );
  CLKBUFX2TS U1144 ( .A(n3741), .Y(n3734) );
  CLKBUFX2TS U1145 ( .A(n4), .Y(n3718) );
  CLKBUFX2TS U1146 ( .A(n3732), .Y(n3729) );
  CLKBUFX2TS U1147 ( .A(n3740), .Y(n3737) );
  CLKBUFX2TS U1148 ( .A(n3732), .Y(n3731) );
  CLKBUFX2TS U1149 ( .A(n3741), .Y(n3735) );
  CLKBUFX2TS U1150 ( .A(n3815), .Y(n3813) );
  CLKBUFX2TS U1151 ( .A(n3815), .Y(n3812) );
  CLKBUFX2TS U1152 ( .A(n3816), .Y(n3811) );
  CLKBUFX2TS U1153 ( .A(n506), .Y(n3769) );
  CLKBUFX2TS U1154 ( .A(n506), .Y(n3770) );
  CLKBUFX2TS U1155 ( .A(n802), .Y(n788) );
  CLKBUFX2TS U1156 ( .A(n3397), .Y(n3383) );
  CLKBUFX2TS U1157 ( .A(n3397), .Y(n3384) );
  CLKBUFX2TS U1158 ( .A(n802), .Y(n789) );
  CLKBUFX2TS U1159 ( .A(n797), .Y(n795) );
  CLKBUFX2TS U1160 ( .A(n800), .Y(n793) );
  CLKBUFX2TS U1161 ( .A(n800), .Y(n792) );
  CLKBUFX2TS U1162 ( .A(n799), .Y(n794) );
  CLKBUFX2TS U1163 ( .A(n801), .Y(n791) );
  CLKBUFX2TS U1164 ( .A(n801), .Y(n790) );
  CLKBUFX2TS U1165 ( .A(n3394), .Y(n3390) );
  CLKBUFX2TS U1166 ( .A(n3395), .Y(n3388) );
  CLKBUFX2TS U1167 ( .A(n3395), .Y(n3387) );
  CLKBUFX2TS U1168 ( .A(n3394), .Y(n3389) );
  CLKBUFX2TS U1169 ( .A(n3396), .Y(n3386) );
  CLKBUFX2TS U1170 ( .A(n3396), .Y(n3385) );
  CLKBUFX2TS U1171 ( .A(n3508), .Y(n3505) );
  CLKBUFX2TS U1172 ( .A(n3509), .Y(n3504) );
  CLKBUFX2TS U1173 ( .A(n3510), .Y(n3502) );
  CLKBUFX2TS U1174 ( .A(n3510), .Y(n3501) );
  CLKBUFX2TS U1175 ( .A(n3511), .Y(n3500) );
  CLKBUFX2TS U1176 ( .A(n3511), .Y(n3499) );
  CLKBUFX2TS U1177 ( .A(n3512), .Y(n3498) );
  CLKBUFX2TS U1178 ( .A(n3512), .Y(n3497) );
  CLKBUFX2TS U1179 ( .A(n3509), .Y(n3503) );
  CLKBUFX2TS U1180 ( .A(n869), .Y(n855) );
  CLKBUFX2TS U1181 ( .A(n3752), .Y(n3743) );
  CLKBUFX2TS U1182 ( .A(n3798), .Y(n3790) );
  CLKBUFX2TS U1183 ( .A(n869), .Y(n856) );
  CLKBUFX2TS U1184 ( .A(n867), .Y(n859) );
  CLKBUFX2TS U1185 ( .A(n866), .Y(n861) );
  CLKBUFX2TS U1186 ( .A(n3796), .Y(n3795) );
  CLKBUFX2TS U1187 ( .A(n3796), .Y(n3794) );
  CLKBUFX2TS U1188 ( .A(n3797), .Y(n3793) );
  CLKBUFX2TS U1189 ( .A(n3797), .Y(n3792) );
  CLKBUFX2TS U1190 ( .A(n3798), .Y(n3791) );
  CLKBUFX2TS U1191 ( .A(n3748), .Y(n3747) );
  CLKBUFX2TS U1192 ( .A(n3751), .Y(n3746) );
  CLKBUFX2TS U1193 ( .A(n3751), .Y(n3745) );
  CLKBUFX2TS U1194 ( .A(n3752), .Y(n3744) );
  CLKBUFX2TS U1195 ( .A(n866), .Y(n862) );
  CLKBUFX2TS U1196 ( .A(n867), .Y(n860) );
  CLKBUFX2TS U1197 ( .A(n868), .Y(n858) );
  CLKBUFX2TS U1198 ( .A(n868), .Y(n857) );
  CLKBUFX2TS U1199 ( .A(n3740), .Y(n3739) );
  CLKBUFX2TS U1200 ( .A(n975), .Y(n863) );
  CLKBUFX2TS U1201 ( .A(n833), .Y(n819) );
  CLKBUFX2TS U1202 ( .A(n3428), .Y(n3414) );
  CLKBUFX2TS U1203 ( .A(n3362), .Y(n3349) );
  CLKBUFX2TS U1204 ( .A(n3428), .Y(n3415) );
  CLKBUFX2TS U1205 ( .A(n833), .Y(n820) );
  CLKBUFX2TS U1206 ( .A(n3283), .Y(n3269) );
  CLKBUFX2TS U1207 ( .A(n3283), .Y(n3270) );
  CLKBUFX2TS U1208 ( .A(n835), .Y(n827) );
  CLKBUFX2TS U1209 ( .A(n831), .Y(n824) );
  CLKBUFX2TS U1210 ( .A(n831), .Y(n823) );
  CLKBUFX2TS U1211 ( .A(n829), .Y(n826) );
  CLKBUFX2TS U1212 ( .A(n832), .Y(n822) );
  CLKBUFX2TS U1213 ( .A(n832), .Y(n821) );
  CLKBUFX2TS U1214 ( .A(n3359), .Y(n3354) );
  CLKBUFX2TS U1215 ( .A(n3361), .Y(n3351) );
  CLKBUFX2TS U1216 ( .A(n3423), .Y(n3420) );
  CLKBUFX2TS U1217 ( .A(n3426), .Y(n3419) );
  CLKBUFX2TS U1218 ( .A(n3426), .Y(n3418) );
  CLKBUFX2TS U1219 ( .A(n3427), .Y(n3417) );
  CLKBUFX2TS U1220 ( .A(n3427), .Y(n3416) );
  CLKBUFX2TS U1221 ( .A(n786), .Y(n770) );
  CLKBUFX2TS U1222 ( .A(n786), .Y(n771) );
  CLKBUFX2TS U1223 ( .A(n3202), .Y(n1669) );
  CLKBUFX2TS U1224 ( .A(n3202), .Y(n1728) );
  CLKBUFX2TS U1225 ( .A(n3360), .Y(n3353) );
  CLKBUFX2TS U1226 ( .A(n3360), .Y(n3352) );
  CLKBUFX2TS U1227 ( .A(n3361), .Y(n3350) );
  CLKBUFX2TS U1228 ( .A(n3508), .Y(n3506) );
  CLKBUFX2TS U1229 ( .A(n785), .Y(n772) );
  CLKBUFX2TS U1230 ( .A(n3282), .Y(n3271) );
  CLKBUFX2TS U1231 ( .A(n784), .Y(n775) );
  CLKBUFX2TS U1232 ( .A(n3200), .Y(n3192) );
  CLKBUFX2TS U1233 ( .A(n3279), .Y(n3278) );
  CLKBUFX2TS U1234 ( .A(n781), .Y(n779) );
  CLKBUFX2TS U1235 ( .A(n3198), .Y(n3196) );
  CLKBUFX2TS U1236 ( .A(n3200), .Y(n1894) );
  CLKBUFX2TS U1237 ( .A(n3279), .Y(n3277) );
  CLKBUFX2TS U1238 ( .A(n3280), .Y(n3276) );
  CLKBUFX2TS U1239 ( .A(n3280), .Y(n3275) );
  CLKBUFX2TS U1240 ( .A(n3281), .Y(n3274) );
  CLKBUFX2TS U1241 ( .A(n3282), .Y(n3272) );
  CLKBUFX2TS U1242 ( .A(n782), .Y(n777) );
  CLKBUFX2TS U1243 ( .A(n782), .Y(n776) );
  CLKBUFX2TS U1244 ( .A(n784), .Y(n774) );
  CLKBUFX2TS U1245 ( .A(n785), .Y(n773) );
  CLKBUFX2TS U1246 ( .A(n3198), .Y(n3195) );
  CLKBUFX2TS U1247 ( .A(n3199), .Y(n3193) );
  CLKBUFX2TS U1248 ( .A(n3199), .Y(n3194) );
  CLKBUFX2TS U1249 ( .A(n3201), .Y(n1822) );
  CLKBUFX2TS U1250 ( .A(n3281), .Y(n3273) );
  CLKBUFX2TS U1251 ( .A(n3331), .Y(n3317) );
  CLKBUFX2TS U1252 ( .A(n3331), .Y(n3318) );
  CLKBUFX2TS U1253 ( .A(n781), .Y(n780) );
  CLKBUFX2TS U1254 ( .A(n3198), .Y(n3197) );
  CLKBUFX2TS U1255 ( .A(n3785), .Y(n3775) );
  CLKBUFX2TS U1256 ( .A(n3782), .Y(n3781) );
  CLKBUFX2TS U1257 ( .A(n3784), .Y(n3778) );
  CLKBUFX2TS U1258 ( .A(n3328), .Y(n3323) );
  CLKBUFX2TS U1259 ( .A(n3329), .Y(n3322) );
  CLKBUFX2TS U1260 ( .A(n3782), .Y(n3780) );
  CLKBUFX2TS U1261 ( .A(n3788), .Y(n3779) );
  CLKBUFX2TS U1262 ( .A(n3784), .Y(n3777) );
  CLKBUFX2TS U1263 ( .A(n3785), .Y(n3776) );
  CLKBUFX2TS U1264 ( .A(n3328), .Y(n3324) );
  CLKBUFX2TS U1265 ( .A(n3329), .Y(n3321) );
  CLKBUFX2TS U1266 ( .A(n3814), .Y(n3803) );
  CLKBUFX2TS U1267 ( .A(n3815), .Y(n3814) );
  INVX2TS U1268 ( .A(n3264), .Y(n3261) );
  INVX2TS U1269 ( .A(n3265), .Y(n3260) );
  INVX2TS U1270 ( .A(n3263), .Y(n3262) );
  CLKBUFX2TS U1271 ( .A(n767), .Y(n756) );
  CLKBUFX2TS U1272 ( .A(n765), .Y(n758) );
  CLKBUFX2TS U1273 ( .A(n764), .Y(n759) );
  CLKBUFX2TS U1274 ( .A(n765), .Y(n757) );
  CLKBUFX2TS U1275 ( .A(n764), .Y(n760) );
  CLKBUFX2TS U1276 ( .A(n763), .Y(n761) );
  CLKBUFX2TS U1277 ( .A(n763), .Y(n762) );
  CLKBUFX2TS U1278 ( .A(n3268), .Y(n3263) );
  CLKBUFX2TS U1279 ( .A(n3268), .Y(n3264) );
  CLKBUFX2TS U1280 ( .A(n3268), .Y(n3265) );
  CLKBUFX2TS U1281 ( .A(n3220), .Y(n3215) );
  CLKBUFX2TS U1282 ( .A(n3220), .Y(n3217) );
  CLKBUFX2TS U1283 ( .A(n3220), .Y(n3216) );
  CLKBUFX2TS U1284 ( .A(n354), .Y(n3771) );
  CLKBUFX2TS U1285 ( .A(n1005), .Y(n781) );
  CLKBUFX2TS U1286 ( .A(n3203), .Y(n3200) );
  CLKBUFX2TS U1287 ( .A(n956), .Y(n3279) );
  CLKBUFX2TS U1288 ( .A(n3284), .Y(n3280) );
  CLKBUFX2TS U1289 ( .A(n3333), .Y(n3326) );
  CLKBUFX2TS U1290 ( .A(n3332), .Y(n3330) );
  CLKBUFX2TS U1291 ( .A(n1005), .Y(n782) );
  CLKBUFX2TS U1292 ( .A(n787), .Y(n783) );
  CLKBUFX2TS U1293 ( .A(n787), .Y(n784) );
  CLKBUFX2TS U1294 ( .A(n787), .Y(n785) );
  CLKBUFX2TS U1295 ( .A(n3788), .Y(n3782) );
  CLKBUFX2TS U1296 ( .A(n973), .Y(n3198) );
  CLKBUFX2TS U1297 ( .A(n3788), .Y(n3783) );
  CLKBUFX2TS U1298 ( .A(n973), .Y(n3199) );
  CLKBUFX2TS U1299 ( .A(n3787), .Y(n3784) );
  CLKBUFX2TS U1300 ( .A(n3203), .Y(n3201) );
  CLKBUFX2TS U1301 ( .A(n3787), .Y(n3785) );
  CLKBUFX2TS U1302 ( .A(n3284), .Y(n3283) );
  CLKBUFX2TS U1303 ( .A(n3284), .Y(n3282) );
  CLKBUFX2TS U1304 ( .A(n3284), .Y(n3281) );
  CLKBUFX2TS U1305 ( .A(n3332), .Y(n3331) );
  CLKBUFX2TS U1306 ( .A(n3333), .Y(n3327) );
  CLKBUFX2TS U1307 ( .A(n3333), .Y(n3328) );
  CLKBUFX2TS U1308 ( .A(n3332), .Y(n3329) );
  CLKBUFX2TS U1309 ( .A(n3430), .Y(n3423) );
  CLKBUFX2TS U1310 ( .A(n835), .Y(n830) );
  CLKBUFX2TS U1311 ( .A(n804), .Y(n797) );
  CLKBUFX2TS U1312 ( .A(n3801), .Y(n3796) );
  CLKBUFX2TS U1313 ( .A(n804), .Y(n798) );
  CLKBUFX2TS U1314 ( .A(n834), .Y(n831) );
  CLKBUFX2TS U1315 ( .A(n803), .Y(n800) );
  CLKBUFX2TS U1316 ( .A(n804), .Y(n799) );
  CLKBUFX2TS U1317 ( .A(n3800), .Y(n3797) );
  CLKBUFX2TS U1318 ( .A(n834), .Y(n832) );
  CLKBUFX2TS U1319 ( .A(n803), .Y(n801) );
  CLKBUFX2TS U1320 ( .A(n3364), .Y(n3358) );
  CLKBUFX2TS U1321 ( .A(n3364), .Y(n3359) );
  CLKBUFX2TS U1322 ( .A(n3363), .Y(n3362) );
  CLKBUFX2TS U1323 ( .A(n3399), .Y(n3392) );
  CLKBUFX2TS U1324 ( .A(n3755), .Y(n3748) );
  CLKBUFX2TS U1325 ( .A(n3430), .Y(n3424) );
  CLKBUFX2TS U1326 ( .A(n3399), .Y(n3393) );
  CLKBUFX2TS U1327 ( .A(n3755), .Y(n3749) );
  CLKBUFX2TS U1328 ( .A(n3755), .Y(n3750) );
  CLKBUFX2TS U1329 ( .A(n3429), .Y(n3426) );
  CLKBUFX2TS U1330 ( .A(n3398), .Y(n3395) );
  CLKBUFX2TS U1331 ( .A(n3430), .Y(n3425) );
  CLKBUFX2TS U1332 ( .A(n3399), .Y(n3394) );
  CLKBUFX2TS U1333 ( .A(n3754), .Y(n3751) );
  CLKBUFX2TS U1334 ( .A(n3429), .Y(n3427) );
  CLKBUFX2TS U1335 ( .A(n3398), .Y(n3396) );
  CLKBUFX2TS U1336 ( .A(n3754), .Y(n3752) );
  CLKBUFX2TS U1337 ( .A(n3429), .Y(n3428) );
  CLKBUFX2TS U1338 ( .A(n3398), .Y(n3397) );
  CLKBUFX2TS U1339 ( .A(n3508), .Y(n3510) );
  CLKBUFX2TS U1340 ( .A(n892), .Y(n3511) );
  CLKBUFX2TS U1341 ( .A(n3508), .Y(n3512) );
  CLKBUFX2TS U1342 ( .A(n892), .Y(n3509) );
  CLKBUFX2TS U1343 ( .A(n787), .Y(n786) );
  CLKBUFX2TS U1344 ( .A(n834), .Y(n833) );
  CLKBUFX2TS U1345 ( .A(n3800), .Y(n3798) );
  CLKBUFX2TS U1346 ( .A(n803), .Y(n802) );
  CLKBUFX2TS U1347 ( .A(n3203), .Y(n3202) );
  CLKBUFX2TS U1348 ( .A(n3363), .Y(n3360) );
  CLKBUFX2TS U1349 ( .A(n3363), .Y(n3361) );
  CLKBUFX2TS U1350 ( .A(n892), .Y(n3508) );
  CLKBUFX2TS U1351 ( .A(n868), .Y(n866) );
  CLKBUFX2TS U1352 ( .A(n870), .Y(n867) );
  CLKBUFX2TS U1353 ( .A(n870), .Y(n868) );
  CLKBUFX2TS U1354 ( .A(n870), .Y(n869) );
  CLKBUFX2TS U1355 ( .A(n497), .Y(n3815) );
  CLKBUFX2TS U1356 ( .A(n387), .Y(n3756) );
  CLKBUFX2TS U1357 ( .A(n175), .Y(n3740) );
  CLKBUFX2TS U1358 ( .A(n513), .Y(n3732) );
  CLKBUFX2TS U1359 ( .A(n3314), .Y(n3300) );
  CLKBUFX2TS U1360 ( .A(n3314), .Y(n3301) );
  CLKBUFX2TS U1361 ( .A(n3310), .Y(n3308) );
  CLKBUFX2TS U1362 ( .A(n3311), .Y(n3307) );
  CLKBUFX2TS U1363 ( .A(n3311), .Y(n3306) );
  CLKBUFX2TS U1364 ( .A(n3313), .Y(n3303) );
  CLKBUFX2TS U1365 ( .A(n3491), .Y(n3487) );
  CLKBUFX2TS U1366 ( .A(n3492), .Y(n3485) );
  CLKBUFX2TS U1367 ( .A(n3493), .Y(n3483) );
  CLKBUFX2TS U1368 ( .A(n3493), .Y(n3482) );
  CLKBUFX2TS U1369 ( .A(n3494), .Y(n3480) );
  CLKBUFX2TS U1370 ( .A(n3312), .Y(n3305) );
  CLKBUFX2TS U1371 ( .A(n3312), .Y(n3304) );
  CLKBUFX2TS U1372 ( .A(n3313), .Y(n3302) );
  CLKBUFX2TS U1373 ( .A(n3491), .Y(n3486) );
  CLKBUFX2TS U1374 ( .A(n3492), .Y(n3484) );
  CLKBUFX2TS U1375 ( .A(n3494), .Y(n3481) );
  CLKBUFX2TS U1376 ( .A(n3235), .Y(n3221) );
  CLKBUFX2TS U1377 ( .A(n3464), .Y(n3449) );
  CLKBUFX2TS U1378 ( .A(n3799), .Y(n3789) );
  CLKBUFX2TS U1379 ( .A(n3800), .Y(n3799) );
  CLKBUFX2TS U1380 ( .A(n3753), .Y(n3742) );
  CLKBUFX2TS U1381 ( .A(n3754), .Y(n3753) );
  CLKBUFX2TS U1382 ( .A(n3235), .Y(n3222) );
  CLKBUFX2TS U1383 ( .A(n751), .Y(n738) );
  CLKBUFX2TS U1384 ( .A(n751), .Y(n737) );
  CLKBUFX2TS U1385 ( .A(n752), .Y(n736) );
  CLKBUFX2TS U1386 ( .A(n748), .Y(n743) );
  CLKBUFX2TS U1387 ( .A(n749), .Y(n742) );
  CLKBUFX2TS U1388 ( .A(n3232), .Y(n3228) );
  CLKBUFX2TS U1389 ( .A(n3232), .Y(n3227) );
  CLKBUFX2TS U1390 ( .A(n3233), .Y(n3226) );
  CLKBUFX2TS U1391 ( .A(n3233), .Y(n3225) );
  CLKBUFX2TS U1392 ( .A(n3234), .Y(n3223) );
  CLKBUFX2TS U1393 ( .A(n749), .Y(n741) );
  CLKBUFX2TS U1394 ( .A(n750), .Y(n740) );
  CLKBUFX2TS U1395 ( .A(n750), .Y(n739) );
  CLKBUFX2TS U1396 ( .A(n752), .Y(n735) );
  CLKBUFX2TS U1397 ( .A(n3234), .Y(n3224) );
  CLKBUFX2TS U1398 ( .A(n3491), .Y(n3488) );
  CLKBUFX2TS U1399 ( .A(n803), .Y(n796) );
  CLKBUFX2TS U1400 ( .A(n3398), .Y(n3391) );
  CLKBUFX2TS U1401 ( .A(n3556), .Y(n3549) );
  CLKBUFX2TS U1402 ( .A(n3557), .Y(n3548) );
  CLKBUFX2TS U1403 ( .A(n3558), .Y(n3545) );
  CLKBUFX2TS U1404 ( .A(n3557), .Y(n3547) );
  CLKBUFX2TS U1405 ( .A(n3459), .Y(n3457) );
  CLKBUFX2TS U1406 ( .A(n3460), .Y(n3455) );
  CLKBUFX2TS U1407 ( .A(n3461), .Y(n3453) );
  CLKBUFX2TS U1408 ( .A(n3461), .Y(n3452) );
  CLKBUFX2TS U1409 ( .A(n3462), .Y(n3450) );
  CLKBUFX2TS U1410 ( .A(n3523), .Y(n3522) );
  CLKBUFX2TS U1411 ( .A(n3523), .Y(n3521) );
  CLKBUFX2TS U1412 ( .A(n3526), .Y(n3519) );
  CLKBUFX2TS U1413 ( .A(n3526), .Y(n3518) );
  CLKBUFX2TS U1414 ( .A(n3459), .Y(n3456) );
  CLKBUFX2TS U1415 ( .A(n3460), .Y(n3454) );
  CLKBUFX2TS U1416 ( .A(n3462), .Y(n3451) );
  CLKBUFX2TS U1417 ( .A(n3786), .Y(n3774) );
  CLKBUFX2TS U1418 ( .A(n3787), .Y(n3786) );
  INVX2TS U1419 ( .A(n3266), .Y(n3252) );
  INVX2TS U1420 ( .A(n3267), .Y(n3253) );
  INVX2TS U1421 ( .A(n3266), .Y(n3259) );
  CLKBUFX2TS U1422 ( .A(n3267), .Y(n3266) );
  INVX2TS U1423 ( .A(n3267), .Y(n3258) );
  INVX2TS U1424 ( .A(n3267), .Y(n3257) );
  INVX2TS U1425 ( .A(n3266), .Y(n3256) );
  INVX2TS U1426 ( .A(n3268), .Y(n3254) );
  INVX2TS U1427 ( .A(n3266), .Y(n3255) );
  INVX2TS U1428 ( .A(n3219), .Y(n3208) );
  INVX2TS U1429 ( .A(n3218), .Y(n3204) );
  INVX2TS U1430 ( .A(n3218), .Y(n3206) );
  INVX2TS U1431 ( .A(n3219), .Y(n3210) );
  INVX2TS U1432 ( .A(n3219), .Y(n3205) );
  INVX2TS U1433 ( .A(n3218), .Y(n3207) );
  INVX2TS U1434 ( .A(n3218), .Y(n3209) );
  INVX2TS U1435 ( .A(n3219), .Y(n3211) );
  INVX2TS U1436 ( .A(n3295), .Y(n3287) );
  INVX2TS U1437 ( .A(n3295), .Y(n3286) );
  INVX2TS U1438 ( .A(n3296), .Y(n3288) );
  INVX2TS U1439 ( .A(n3296), .Y(n3289) );
  INVX2TS U1440 ( .A(n3297), .Y(n3290) );
  INVX2TS U1441 ( .A(n3297), .Y(n3291) );
  INVX2TS U1442 ( .A(n3298), .Y(n3293) );
  INVX2TS U1443 ( .A(n3298), .Y(n3292) );
  INVX2TS U1444 ( .A(n3297), .Y(n3294) );
  INVX2TS U1445 ( .A(n732), .Y(n715) );
  INVX2TS U1446 ( .A(n732), .Y(n714) );
  INVX2TS U1447 ( .A(n717), .Y(n707) );
  INVX2TS U1448 ( .A(n717), .Y(n706) );
  INVX2TS U1449 ( .A(n727), .Y(n711) );
  INVX2TS U1450 ( .A(n733), .Y(n712) );
  INVX2TS U1451 ( .A(n727), .Y(n708) );
  INVX2TS U1452 ( .A(n717), .Y(n705) );
  INVX2TS U1453 ( .A(n3379), .Y(n3375) );
  INVX2TS U1454 ( .A(n851), .Y(n847) );
  INVX2TS U1455 ( .A(n851), .Y(n846) );
  INVX2TS U1456 ( .A(n851), .Y(n845) );
  INVX2TS U1457 ( .A(n3379), .Y(n3374) );
  INVX2TS U1458 ( .A(n3446), .Y(n3441) );
  INVX2TS U1459 ( .A(n3447), .Y(n3440) );
  INVX2TS U1460 ( .A(n3448), .Y(n3439) );
  INVX2TS U1461 ( .A(n3579), .Y(n3572) );
  INVX2TS U1462 ( .A(n3579), .Y(n3571) );
  INVX2TS U1463 ( .A(n3578), .Y(n3570) );
  INVX2TS U1464 ( .A(n3379), .Y(n3373) );
  INVX2TS U1465 ( .A(n590), .Y(n839) );
  INVX2TS U1466 ( .A(n3446), .Y(n3433) );
  INVX2TS U1467 ( .A(n3576), .Y(n3564) );
  INVX2TS U1468 ( .A(n3381), .Y(n3367) );
  INVX2TS U1469 ( .A(n854), .Y(n840) );
  INVX2TS U1470 ( .A(n3446), .Y(n3434) );
  INVX2TS U1471 ( .A(n3576), .Y(n3565) );
  INVX2TS U1472 ( .A(n3381), .Y(n3368) );
  INVX2TS U1473 ( .A(n852), .Y(n843) );
  INVX2TS U1474 ( .A(n852), .Y(n844) );
  INVX2TS U1475 ( .A(n852), .Y(n842) );
  INVX2TS U1476 ( .A(n3380), .Y(n3371) );
  INVX2TS U1477 ( .A(n3382), .Y(n3370) );
  INVX2TS U1478 ( .A(n3445), .Y(n3437) );
  INVX2TS U1479 ( .A(n3445), .Y(n3438) );
  INVX2TS U1480 ( .A(n3445), .Y(n3436) );
  INVX2TS U1481 ( .A(n3446), .Y(n3435) );
  INVX2TS U1482 ( .A(n3576), .Y(n3568) );
  INVX2TS U1483 ( .A(n3577), .Y(n3569) );
  INVX2TS U1484 ( .A(n3578), .Y(n3567) );
  INVX2TS U1485 ( .A(n3576), .Y(n3566) );
  INVX2TS U1486 ( .A(n590), .Y(n841) );
  INVX2TS U1487 ( .A(n3381), .Y(n3372) );
  INVX2TS U1488 ( .A(n584), .Y(n3369) );
  INVX2TS U1489 ( .A(n727), .Y(n716) );
  INVX2TS U1490 ( .A(n853), .Y(n837) );
  INVX2TS U1491 ( .A(n3447), .Y(n3431) );
  INVX2TS U1492 ( .A(n3380), .Y(n3365) );
  INVX2TS U1493 ( .A(n3577), .Y(n3562) );
  INVX2TS U1494 ( .A(n853), .Y(n838) );
  INVX2TS U1495 ( .A(n3380), .Y(n3366) );
  INVX2TS U1496 ( .A(n3447), .Y(n3432) );
  INVX2TS U1497 ( .A(n3577), .Y(n3563) );
  CLKBUFX2TS U1498 ( .A(n768), .Y(n767) );
  CLKBUFX2TS U1499 ( .A(n768), .Y(n766) );
  CLKBUFX2TS U1500 ( .A(n769), .Y(n765) );
  CLKBUFX2TS U1501 ( .A(n769), .Y(n764) );
  CLKBUFX2TS U1502 ( .A(n769), .Y(n763) );
  CLKBUFX2TS U1503 ( .A(n3249), .Y(n3238) );
  CLKBUFX2TS U1504 ( .A(n3248), .Y(n3240) );
  CLKBUFX2TS U1505 ( .A(n1585), .Y(n886) );
  CLKBUFX2TS U1506 ( .A(n3249), .Y(n3239) );
  CLKBUFX2TS U1507 ( .A(n1544), .Y(n919) );
  CLKBUFX2TS U1508 ( .A(n1531), .Y(n955) );
  CLKBUFX2TS U1509 ( .A(n1531), .Y(n957) );
  CLKBUFX2TS U1510 ( .A(n3251), .Y(n3244) );
  CLKBUFX2TS U1511 ( .A(n3247), .Y(n3243) );
  CLKBUFX2TS U1512 ( .A(n3248), .Y(n3241) );
  CLKBUFX2TS U1513 ( .A(n1544), .Y(n936) );
  CLKBUFX2TS U1514 ( .A(n1402), .Y(n970) );
  CLKBUFX2TS U1515 ( .A(n1402), .Y(n986) );
  CLKBUFX2TS U1516 ( .A(n3247), .Y(n3242) );
  CLKBUFX2TS U1517 ( .A(n3477), .Y(n3467) );
  CLKBUFX2TS U1518 ( .A(n816), .Y(n806) );
  CLKBUFX2TS U1519 ( .A(n815), .Y(n808) );
  CLKBUFX2TS U1520 ( .A(n816), .Y(n807) );
  CLKBUFX2TS U1521 ( .A(n815), .Y(n810) );
  CLKBUFX2TS U1522 ( .A(n3344), .Y(n3337) );
  CLKBUFX2TS U1523 ( .A(n3347), .Y(n3339) );
  CLKBUFX2TS U1524 ( .A(n3410), .Y(n3402) );
  CLKBUFX2TS U1525 ( .A(n3410), .Y(n3403) );
  CLKBUFX2TS U1526 ( .A(n3409), .Y(n3404) );
  CLKBUFX2TS U1527 ( .A(n3411), .Y(n3401) );
  CLKBUFX2TS U1528 ( .A(n3476), .Y(n3474) );
  CLKBUFX2TS U1529 ( .A(n3475), .Y(n3471) );
  CLKBUFX2TS U1530 ( .A(n3476), .Y(n3470) );
  CLKBUFX2TS U1531 ( .A(n3476), .Y(n3469) );
  CLKBUFX2TS U1532 ( .A(n3542), .Y(n3532) );
  CLKBUFX2TS U1533 ( .A(n3542), .Y(n3533) );
  CLKBUFX2TS U1534 ( .A(n3541), .Y(n3534) );
  CLKBUFX2TS U1535 ( .A(n3540), .Y(n3535) );
  CLKBUFX2TS U1536 ( .A(n3540), .Y(n3536) );
  CLKBUFX2TS U1537 ( .A(n3539), .Y(n3537) );
  CLKBUFX2TS U1538 ( .A(n3539), .Y(n3538) );
  CLKBUFX2TS U1539 ( .A(n815), .Y(n809) );
  CLKBUFX2TS U1540 ( .A(n3345), .Y(n3336) );
  CLKBUFX2TS U1541 ( .A(n3345), .Y(n3335) );
  CLKBUFX2TS U1542 ( .A(n3344), .Y(n3338) );
  CLKBUFX2TS U1543 ( .A(n3476), .Y(n3473) );
  CLKBUFX2TS U1544 ( .A(n3475), .Y(n3472) );
  CLKBUFX2TS U1545 ( .A(n3477), .Y(n3468) );
  CLKBUFX2TS U1546 ( .A(n3343), .Y(n3342) );
  CLKBUFX2TS U1547 ( .A(n3343), .Y(n3340) );
  CLKBUFX2TS U1548 ( .A(n814), .Y(n813) );
  CLKBUFX2TS U1549 ( .A(n990), .Y(n811) );
  CLKBUFX2TS U1550 ( .A(n814), .Y(n812) );
  CLKBUFX2TS U1551 ( .A(n3343), .Y(n3341) );
  CLKBUFX2TS U1552 ( .A(n3408), .Y(n3407) );
  CLKBUFX2TS U1553 ( .A(n3409), .Y(n3405) );
  CLKBUFX2TS U1554 ( .A(n3408), .Y(n3406) );
  CLKBUFX2TS U1555 ( .A(n3606), .Y(n3594) );
  CLKBUFX2TS U1556 ( .A(n3606), .Y(n3602) );
  CLKBUFX2TS U1557 ( .A(n3603), .Y(n3601) );
  CLKBUFX2TS U1558 ( .A(n3603), .Y(n3600) );
  CLKBUFX2TS U1559 ( .A(n3604), .Y(n3599) );
  CLKBUFX2TS U1560 ( .A(n3604), .Y(n3598) );
  CLKBUFX2TS U1561 ( .A(n3605), .Y(n3597) );
  CLKBUFX2TS U1562 ( .A(n3606), .Y(n3595) );
  CLKBUFX2TS U1563 ( .A(n3605), .Y(n3596) );
  CLKBUFX2TS U1564 ( .A(n3591), .Y(n3580) );
  CLKBUFX2TS U1565 ( .A(n3589), .Y(n3581) );
  CLKBUFX2TS U1566 ( .A(n3589), .Y(n3582) );
  CLKBUFX2TS U1567 ( .A(n3588), .Y(n3583) );
  CLKBUFX2TS U1568 ( .A(n3587), .Y(n3586) );
  CLKBUFX2TS U1569 ( .A(n3588), .Y(n3584) );
  CLKBUFX2TS U1570 ( .A(n3587), .Y(n3585) );
  CLKBUFX2TS U1571 ( .A(n3700), .Y(n3688) );
  CLKBUFX2TS U1572 ( .A(n3700), .Y(n3689) );
  CLKBUFX2TS U1573 ( .A(n3672), .Y(n3665) );
  CLKBUFX2TS U1574 ( .A(n3667), .Y(n3664) );
  CLKBUFX2TS U1575 ( .A(n3667), .Y(n3663) );
  CLKBUFX2TS U1576 ( .A(n3701), .Y(n3690) );
  CLKBUFX2TS U1577 ( .A(n3699), .Y(n3691) );
  CLKBUFX2TS U1578 ( .A(n3668), .Y(n3661) );
  CLKBUFX2TS U1579 ( .A(n3699), .Y(n3692) );
  CLKBUFX2TS U1580 ( .A(n3669), .Y(n3660) );
  CLKBUFX2TS U1581 ( .A(n3698), .Y(n3693) );
  CLKBUFX2TS U1582 ( .A(n3670), .Y(n3657) );
  CLKBUFX2TS U1583 ( .A(n3669), .Y(n3659) );
  CLKBUFX2TS U1584 ( .A(n3670), .Y(n3658) );
  CLKBUFX2TS U1585 ( .A(n3668), .Y(n3662) );
  CLKBUFX2TS U1586 ( .A(n3698), .Y(n3694) );
  CLKBUFX2TS U1587 ( .A(n3697), .Y(n3695) );
  CLKBUFX2TS U1588 ( .A(n3697), .Y(n3696) );
  CLKBUFX2TS U1589 ( .A(n504), .Y(n3773) );
  CLKBUFX2TS U1590 ( .A(n499), .Y(n3802) );
  CLKBUFX2TS U1591 ( .A(n3236), .Y(n3235) );
  CLKBUFX2TS U1592 ( .A(n3236), .Y(n3233) );
  CLKBUFX2TS U1593 ( .A(n3236), .Y(n3234) );
  CLKBUFX2TS U1594 ( .A(n3464), .Y(n3463) );
  CLKBUFX2TS U1595 ( .A(n3316), .Y(n3311) );
  CLKBUFX2TS U1596 ( .A(n3315), .Y(n3314) );
  CLKBUFX2TS U1597 ( .A(n3465), .Y(n3461) );
  CLKBUFX2TS U1598 ( .A(n3495), .Y(n3493) );
  CLKBUFX2TS U1599 ( .A(n3529), .Y(n3528) );
  CLKBUFX2TS U1600 ( .A(n3560), .Y(n3556) );
  CLKBUFX2TS U1601 ( .A(n3530), .Y(n3523) );
  CLKBUFX2TS U1602 ( .A(n3530), .Y(n3524) );
  CLKBUFX2TS U1603 ( .A(n3529), .Y(n3526) );
  CLKBUFX2TS U1604 ( .A(n3559), .Y(n3558) );
  CLKBUFX2TS U1605 ( .A(n3530), .Y(n3525) );
  CLKBUFX2TS U1606 ( .A(n3560), .Y(n3557) );
  CLKBUFX2TS U1607 ( .A(n3315), .Y(n3312) );
  CLKBUFX2TS U1608 ( .A(n3315), .Y(n3313) );
  CLKBUFX2TS U1609 ( .A(n3496), .Y(n3490) );
  CLKBUFX2TS U1610 ( .A(n3465), .Y(n3459) );
  CLKBUFX2TS U1611 ( .A(n3496), .Y(n3491) );
  CLKBUFX2TS U1612 ( .A(n3465), .Y(n3460) );
  CLKBUFX2TS U1613 ( .A(n3495), .Y(n3492) );
  CLKBUFX2TS U1614 ( .A(n3464), .Y(n3462) );
  CLKBUFX2TS U1615 ( .A(n3495), .Y(n3494) );
  CLKBUFX2TS U1616 ( .A(n3560), .Y(n3555) );
  CLKBUFX2TS U1617 ( .A(n3529), .Y(n3527) );
  CLKBUFX2TS U1618 ( .A(n754), .Y(n751) );
  CLKBUFX2TS U1619 ( .A(n3237), .Y(n3231) );
  CLKBUFX2TS U1620 ( .A(n956), .Y(n3285) );
  CLKBUFX2TS U1621 ( .A(n836), .Y(n829) );
  CLKBUFX2TS U1622 ( .A(n989), .Y(n836) );
  CLKBUFX2TS U1623 ( .A(n3237), .Y(n3232) );
  CLKBUFX2TS U1624 ( .A(n3513), .Y(n3507) );
  CLKBUFX2TS U1625 ( .A(n892), .Y(n3513) );
  CLKBUFX2TS U1626 ( .A(n754), .Y(n749) );
  CLKBUFX2TS U1627 ( .A(n753), .Y(n750) );
  CLKBUFX2TS U1628 ( .A(n754), .Y(n752) );
  CLKBUFX2TS U1629 ( .A(n754), .Y(n753) );
  CLKBUFX2TS U1630 ( .A(n975), .Y(n871) );
  CLKBUFX2TS U1631 ( .A(n975), .Y(n870) );
  CLKBUFX2TS U1632 ( .A(n956), .Y(n3284) );
  CLKBUFX2TS U1633 ( .A(n973), .Y(n3203) );
  CLKBUFX2TS U1634 ( .A(n941), .Y(n3333) );
  CLKBUFX2TS U1635 ( .A(n941), .Y(n3332) );
  CLKBUFX2TS U1636 ( .A(n939), .Y(n3364) );
  CLKBUFX2TS U1637 ( .A(n922), .Y(n3429) );
  CLKBUFX2TS U1638 ( .A(n925), .Y(n3398) );
  CLKBUFX2TS U1639 ( .A(n989), .Y(n834) );
  CLKBUFX2TS U1640 ( .A(n992), .Y(n803) );
  CLKBUFX2TS U1641 ( .A(n939), .Y(n3363) );
  CLKBUFX2TS U1642 ( .A(n1005), .Y(n787) );
  CLKBUFX2TS U1643 ( .A(n502), .Y(n3788) );
  CLKBUFX2TS U1644 ( .A(n502), .Y(n3787) );
  CLKBUFX2TS U1645 ( .A(n500), .Y(n3801) );
  CLKBUFX2TS U1646 ( .A(n510), .Y(n3755) );
  CLKBUFX2TS U1647 ( .A(n510), .Y(n3754) );
  CLKBUFX2TS U1648 ( .A(n500), .Y(n3800) );
  CLKBUFX2TS U1649 ( .A(n582), .Y(n3218) );
  CLKBUFX2TS U1650 ( .A(n582), .Y(n3219) );
  CLKBUFX2TS U1651 ( .A(n581), .Y(n3267) );
  CLKBUFX2TS U1652 ( .A(n581), .Y(n3268) );
  CLKBUFX2TS U1653 ( .A(n582), .Y(n3220) );
  CLKBUFX2TS U1654 ( .A(n732), .Y(n729) );
  CLKBUFX2TS U1655 ( .A(n3237), .Y(n3229) );
  CLKBUFX2TS U1656 ( .A(n3491), .Y(n3489) );
  CLKBUFX2TS U1657 ( .A(n908), .Y(n3458) );
  CLKBUFX2TS U1658 ( .A(n3299), .Y(n3295) );
  CLKBUFX2TS U1659 ( .A(n3299), .Y(n3296) );
  CLKBUFX2TS U1660 ( .A(n3299), .Y(n3297) );
  CLKBUFX2TS U1661 ( .A(n854), .Y(n853) );
  CLKBUFX2TS U1662 ( .A(n3448), .Y(n3447) );
  CLKBUFX2TS U1663 ( .A(n3381), .Y(n3380) );
  CLKBUFX2TS U1664 ( .A(n3578), .Y(n3577) );
  INVX2TS U1665 ( .A(n734), .Y(n702) );
  INVX2TS U1666 ( .A(n734), .Y(n703) );
  INVX2TS U1667 ( .A(n734), .Y(n704) );
  INVX2TS U1668 ( .A(n852), .Y(n849) );
  INVX2TS U1669 ( .A(n853), .Y(n848) );
  INVX2TS U1670 ( .A(n3447), .Y(n3443) );
  INVX2TS U1671 ( .A(n588), .Y(n3442) );
  INVX2TS U1672 ( .A(n3579), .Y(n3574) );
  INVX2TS U1673 ( .A(n3579), .Y(n3573) );
  CLKBUFX2TS U1674 ( .A(n1654), .Y(n1531) );
  CLKBUFX2TS U1675 ( .A(n818), .Y(n816) );
  CLKBUFX2TS U1676 ( .A(n990), .Y(n814) );
  CLKBUFX2TS U1677 ( .A(n1653), .Y(n1585) );
  CLKBUFX2TS U1678 ( .A(n3250), .Y(n3249) );
  CLKBUFX2TS U1679 ( .A(n3251), .Y(n3245) );
  CLKBUFX2TS U1680 ( .A(n3251), .Y(n3246) );
  CLKBUFX2TS U1681 ( .A(n3250), .Y(n3248) );
  CLKBUFX2TS U1682 ( .A(n3347), .Y(n3343) );
  CLKBUFX2TS U1683 ( .A(n3413), .Y(n3410) );
  CLKBUFX2TS U1684 ( .A(n3413), .Y(n3409) );
  CLKBUFX2TS U1685 ( .A(n3413), .Y(n3408) );
  CLKBUFX2TS U1686 ( .A(n3479), .Y(n3476) );
  CLKBUFX2TS U1687 ( .A(n3541), .Y(n3542) );
  CLKBUFX2TS U1688 ( .A(n3544), .Y(n3541) );
  CLKBUFX2TS U1689 ( .A(n3544), .Y(n3540) );
  CLKBUFX2TS U1690 ( .A(n3544), .Y(n3539) );
  CLKBUFX2TS U1691 ( .A(n818), .Y(n815) );
  CLKBUFX2TS U1692 ( .A(n1653), .Y(n1546) );
  CLKBUFX2TS U1693 ( .A(n1654), .Y(n1544) );
  CLKBUFX2TS U1694 ( .A(n1654), .Y(n1402) );
  CLKBUFX2TS U1695 ( .A(n3250), .Y(n3247) );
  CLKBUFX2TS U1696 ( .A(n940), .Y(n3345) );
  CLKBUFX2TS U1697 ( .A(n3347), .Y(n3344) );
  CLKBUFX2TS U1698 ( .A(n907), .Y(n3475) );
  CLKBUFX2TS U1699 ( .A(n3479), .Y(n3477) );
  CLKBUFX2TS U1700 ( .A(n1006), .Y(n768) );
  CLKBUFX2TS U1701 ( .A(n1006), .Y(n769) );
  INVX2TS U1702 ( .A(n700), .Y(n685) );
  INVX2TS U1703 ( .A(n701), .Y(n686) );
  INVX2TS U1704 ( .A(n699), .Y(n695) );
  INVX2TS U1705 ( .A(n699), .Y(n694) );
  INVX2TS U1706 ( .A(n696), .Y(n693) );
  INVX2TS U1707 ( .A(n696), .Y(n692) );
  INVX2TS U1708 ( .A(n696), .Y(n691) );
  INVX2TS U1709 ( .A(n700), .Y(n689) );
  INVX2TS U1710 ( .A(n700), .Y(n688) );
  INVX2TS U1711 ( .A(n700), .Y(n690) );
  INVX2TS U1712 ( .A(n696), .Y(n687) );
  CLKBUFX2TS U1713 ( .A(n3478), .Y(n3466) );
  CLKBUFX2TS U1714 ( .A(n3479), .Y(n3478) );
  CLKBUFX2TS U1715 ( .A(n817), .Y(n805) );
  CLKBUFX2TS U1716 ( .A(n818), .Y(n817) );
  CLKBUFX2TS U1717 ( .A(n3346), .Y(n3334) );
  CLKBUFX2TS U1718 ( .A(n940), .Y(n3346) );
  CLKBUFX2TS U1719 ( .A(n3411), .Y(n3400) );
  CLKBUFX2TS U1720 ( .A(n3412), .Y(n3411) );
  CLKBUFX2TS U1721 ( .A(n3543), .Y(n3531) );
  CLKBUFX2TS U1722 ( .A(n890), .Y(n3543) );
  CLKBUFX2TS U1723 ( .A(n664), .Y(n653) );
  CLKBUFX2TS U1724 ( .A(n660), .Y(n659) );
  CLKBUFX2TS U1725 ( .A(n660), .Y(n658) );
  CLKBUFX2TS U1726 ( .A(n661), .Y(n657) );
  CLKBUFX2TS U1727 ( .A(n664), .Y(n654) );
  CLKBUFX2TS U1728 ( .A(n663), .Y(n656) );
  CLKBUFX2TS U1729 ( .A(n663), .Y(n655) );
  INVX2TS U1730 ( .A(n631), .Y(n630) );
  INVX2TS U1731 ( .A(n632), .Y(n629) );
  INVX2TS U1732 ( .A(n633), .Y(n628) );
  CLKBUFX2TS U1733 ( .A(n3608), .Y(n3603) );
  CLKBUFX2TS U1734 ( .A(n3607), .Y(n3604) );
  CLKBUFX2TS U1735 ( .A(n3607), .Y(n3606) );
  CLKBUFX2TS U1736 ( .A(n3607), .Y(n3605) );
  CLKBUFX2TS U1737 ( .A(n3592), .Y(n3591) );
  CLKBUFX2TS U1738 ( .A(n3592), .Y(n3590) );
  CLKBUFX2TS U1739 ( .A(n3593), .Y(n3589) );
  CLKBUFX2TS U1740 ( .A(n3593), .Y(n3588) );
  CLKBUFX2TS U1741 ( .A(n3593), .Y(n3587) );
  CLKBUFX2TS U1742 ( .A(n607), .Y(n596) );
  CLKBUFX2TS U1743 ( .A(n605), .Y(n597) );
  CLKBUFX2TS U1744 ( .A(n605), .Y(n598) );
  CLKBUFX2TS U1745 ( .A(n604), .Y(n599) );
  CLKBUFX2TS U1746 ( .A(n603), .Y(n602) );
  CLKBUFX2TS U1747 ( .A(n604), .Y(n600) );
  CLKBUFX2TS U1748 ( .A(n603), .Y(n601) );
  CLKBUFX2TS U1749 ( .A(n648), .Y(n636) );
  CLKBUFX2TS U1750 ( .A(n648), .Y(n637) );
  CLKBUFX2TS U1751 ( .A(n646), .Y(n638) );
  CLKBUFX2TS U1752 ( .A(n646), .Y(n639) );
  CLKBUFX2TS U1753 ( .A(n645), .Y(n640) );
  CLKBUFX2TS U1754 ( .A(n644), .Y(n643) );
  CLKBUFX2TS U1755 ( .A(n645), .Y(n641) );
  CLKBUFX2TS U1756 ( .A(n644), .Y(n642) );
  INVX2TS U1757 ( .A(reset), .Y(n4392) );
  CLKBUFX2TS U1758 ( .A(n3638), .Y(n3626) );
  CLKBUFX2TS U1759 ( .A(n3682), .Y(n3679) );
  CLKBUFX2TS U1760 ( .A(n3638), .Y(n3627) );
  CLKBUFX2TS U1761 ( .A(n3716), .Y(n3703) );
  CLKBUFX2TS U1762 ( .A(n3683), .Y(n3678) );
  CLKBUFX2TS U1763 ( .A(n3683), .Y(n3677) );
  CLKBUFX2TS U1764 ( .A(n3712), .Y(n3704) );
  CLKBUFX2TS U1765 ( .A(n3639), .Y(n3628) );
  CLKBUFX2TS U1766 ( .A(n3684), .Y(n3676) );
  CLKBUFX2TS U1767 ( .A(n3713), .Y(n3705) );
  CLKBUFX2TS U1768 ( .A(n3637), .Y(n3629) );
  CLKBUFX2TS U1769 ( .A(n3684), .Y(n3675) );
  CLKBUFX2TS U1770 ( .A(n3713), .Y(n3706) );
  CLKBUFX2TS U1771 ( .A(n3637), .Y(n3630) );
  CLKBUFX2TS U1772 ( .A(n3685), .Y(n3674) );
  CLKBUFX2TS U1773 ( .A(n3712), .Y(n3707) );
  CLKBUFX2TS U1774 ( .A(n3636), .Y(n3631) );
  CLKBUFX2TS U1775 ( .A(n3685), .Y(n3673) );
  CLKBUFX2TS U1776 ( .A(n3623), .Y(n3609) );
  CLKBUFX2TS U1777 ( .A(n3623), .Y(n3610) );
  CLKBUFX2TS U1778 ( .A(n3652), .Y(n3642) );
  CLKBUFX2TS U1779 ( .A(n3625), .Y(n3617) );
  CLKBUFX2TS U1780 ( .A(n3620), .Y(n3616) );
  CLKBUFX2TS U1781 ( .A(n3620), .Y(n3615) );
  CLKBUFX2TS U1782 ( .A(n3650), .Y(n3646) );
  CLKBUFX2TS U1783 ( .A(n3621), .Y(n3614) );
  CLKBUFX2TS U1784 ( .A(n3650), .Y(n3645) );
  CLKBUFX2TS U1785 ( .A(n3621), .Y(n3613) );
  CLKBUFX2TS U1786 ( .A(n3651), .Y(n3644) );
  CLKBUFX2TS U1787 ( .A(n3622), .Y(n3612) );
  CLKBUFX2TS U1788 ( .A(n3651), .Y(n3643) );
  CLKBUFX2TS U1789 ( .A(n3622), .Y(n3611) );
  CLKBUFX2TS U1790 ( .A(n3636), .Y(n3632) );
  CLKBUFX2TS U1791 ( .A(n3712), .Y(n3708) );
  CLKBUFX2TS U1792 ( .A(n3635), .Y(n3634) );
  CLKBUFX2TS U1793 ( .A(n3701), .Y(n3700) );
  CLKBUFX2TS U1794 ( .A(n3672), .Y(n3667) );
  CLKBUFX2TS U1795 ( .A(n3702), .Y(n3699) );
  CLKBUFX2TS U1796 ( .A(n3702), .Y(n3698) );
  CLKBUFX2TS U1797 ( .A(n3671), .Y(n3669) );
  CLKBUFX2TS U1798 ( .A(n3671), .Y(n3670) );
  CLKBUFX2TS U1799 ( .A(n3671), .Y(n3668) );
  CLKBUFX2TS U1800 ( .A(n3702), .Y(n3697) );
  CLKBUFX2TS U1801 ( .A(n549), .Y(n3666) );
  CLKBUFX2TS U1802 ( .A(n3635), .Y(n3633) );
  CLKBUFX2TS U1803 ( .A(n3682), .Y(n3680) );
  CLKBUFX2TS U1804 ( .A(n3711), .Y(n3709) );
  CLKBUFX2TS U1805 ( .A(n3684), .Y(n3681) );
  CLKBUFX2TS U1806 ( .A(n3711), .Y(n3710) );
  NOR2X1TS U1807 ( .A(n1581), .B(n216), .Y(n956) );
  NOR2X1TS U1808 ( .A(n1604), .B(n498), .Y(n1005) );
  AND2X2TS U1809 ( .A(n1554), .B(n163), .Y(n892) );
  AND2X2TS U1810 ( .A(n1564), .B(n523), .Y(n925) );
  AND2X2TS U1811 ( .A(n1593), .B(n520), .Y(n989) );
  INVX2TS U1812 ( .A(n1547), .Y(n499) );
  CLKBUFX2TS U1813 ( .A(n959), .Y(n3236) );
  CLKBUFX2TS U1814 ( .A(n589), .Y(n732) );
  CLKBUFX2TS U1815 ( .A(n589), .Y(n733) );
  CLKBUFX2TS U1816 ( .A(n1007), .Y(n755) );
  INVX2TS U1817 ( .A(n1577), .Y(n526) );
  CLKBUFX2TS U1818 ( .A(n942), .Y(n3316) );
  CLKBUFX2TS U1819 ( .A(n942), .Y(n3315) );
  CLKBUFX2TS U1820 ( .A(n908), .Y(n3464) );
  CLKBUFX2TS U1821 ( .A(n889), .Y(n3559) );
  CLKBUFX2TS U1822 ( .A(n891), .Y(n3530) );
  CLKBUFX2TS U1823 ( .A(n906), .Y(n3496) );
  CLKBUFX2TS U1824 ( .A(n908), .Y(n3465) );
  CLKBUFX2TS U1825 ( .A(n906), .Y(n3495) );
  CLKBUFX2TS U1826 ( .A(n889), .Y(n3560) );
  CLKBUFX2TS U1827 ( .A(n891), .Y(n3529) );
  CLKBUFX2TS U1828 ( .A(n958), .Y(n3251) );
  INVX2TS U1829 ( .A(n1604), .Y(n518) );
  CLKBUFX2TS U1830 ( .A(n435), .Y(n3298) );
  CLKBUFX2TS U1831 ( .A(n1007), .Y(n754) );
  INVX2TS U1832 ( .A(n2), .Y(n510) );
  INVX2TS U1833 ( .A(n444), .Y(n500) );
  INVX2TS U1834 ( .A(n1582), .Y(n521) );
  CLKBUFX2TS U1835 ( .A(n3561), .Y(n3554) );
  CLKBUFX2TS U1836 ( .A(n889), .Y(n3561) );
  INVX2TS U1837 ( .A(n1581), .Y(n522) );
  CLKBUFX2TS U1838 ( .A(n588), .Y(n3448) );
  CLKBUFX2TS U1839 ( .A(n591), .Y(n3579) );
  CLKBUFX2TS U1840 ( .A(n590), .Y(n854) );
  CLKBUFX2TS U1841 ( .A(n584), .Y(n3382) );
  CLKBUFX2TS U1842 ( .A(n584), .Y(n3381) );
  CLKBUFX2TS U1843 ( .A(n591), .Y(n3578) );
  CLKBUFX2TS U1844 ( .A(n435), .Y(n3299) );
  CLKBUFX2TS U1845 ( .A(n635), .Y(n631) );
  CLKBUFX2TS U1846 ( .A(n635), .Y(n632) );
  CLKBUFX2TS U1847 ( .A(n635), .Y(n633) );
  AND2X2TS U1848 ( .A(n1644), .B(n1763), .Y(n1006) );
  CLKBUFX2TS U1849 ( .A(n667), .Y(n660) );
  CLKBUFX2TS U1850 ( .A(n667), .Y(n661) );
  CLKBUFX2TS U1851 ( .A(n667), .Y(n662) );
  CLKBUFX2TS U1852 ( .A(n666), .Y(n664) );
  CLKBUFX2TS U1853 ( .A(n666), .Y(n663) );
  CLKBUFX2TS U1854 ( .A(n923), .Y(n3412) );
  CLKBUFX2TS U1855 ( .A(n923), .Y(n3413) );
  CLKBUFX2TS U1856 ( .A(n890), .Y(n3544) );
  CLKBUFX2TS U1857 ( .A(n990), .Y(n818) );
  CLKBUFX2TS U1858 ( .A(n974), .Y(n1653) );
  CLKBUFX2TS U1859 ( .A(n974), .Y(n1654) );
  CLKBUFX2TS U1860 ( .A(n958), .Y(n3250) );
  CLKBUFX2TS U1861 ( .A(n940), .Y(n3347) );
  CLKBUFX2TS U1862 ( .A(n907), .Y(n3479) );
  CLKBUFX2TS U1863 ( .A(n699), .Y(n697) );
  CLKBUFX2TS U1864 ( .A(n699), .Y(n698) );
  CLKBUFX2TS U1865 ( .A(n665), .Y(n652) );
  CLKBUFX2TS U1866 ( .A(n666), .Y(n665) );
  INVX2TS U1867 ( .A(n633), .Y(n610) );
  INVX2TS U1868 ( .A(n634), .Y(n611) );
  CLKBUFX2TS U1869 ( .A(n592), .Y(n634) );
  INVX2TS U1870 ( .A(n634), .Y(n612) );
  INVX2TS U1871 ( .A(n634), .Y(n613) );
  INVX2TS U1872 ( .A(n635), .Y(n614) );
  INVX2TS U1873 ( .A(n592), .Y(n622) );
  INVX2TS U1874 ( .A(n634), .Y(n623) );
  INVX2TS U1875 ( .A(n592), .Y(n624) );
  CLKBUFX2TS U1876 ( .A(n650), .Y(n648) );
  CLKBUFX2TS U1877 ( .A(n608), .Y(n607) );
  CLKBUFX2TS U1878 ( .A(n650), .Y(n647) );
  CLKBUFX2TS U1879 ( .A(n608), .Y(n606) );
  CLKBUFX2TS U1880 ( .A(n651), .Y(n646) );
  CLKBUFX2TS U1881 ( .A(n609), .Y(n605) );
  CLKBUFX2TS U1882 ( .A(n651), .Y(n645) );
  CLKBUFX2TS U1883 ( .A(n609), .Y(n604) );
  CLKBUFX2TS U1884 ( .A(n651), .Y(n644) );
  CLKBUFX2TS U1885 ( .A(n609), .Y(n603) );
  CLKBUFX2TS U1886 ( .A(n709), .Y(n3608) );
  CLKBUFX2TS U1887 ( .A(n709), .Y(n3607) );
  CLKBUFX2TS U1888 ( .A(n1837), .Y(n3592) );
  CLKBUFX2TS U1889 ( .A(n1837), .Y(n3593) );
  CLKBUFX2TS U1890 ( .A(n650), .Y(n649) );
  CLKBUFX2TS U1891 ( .A(n4280), .Y(n4281) );
  CLKBUFX2TS U1892 ( .A(n4283), .Y(n4284) );
  CLKBUFX2TS U1893 ( .A(n4280), .Y(n4282) );
  CLKBUFX2TS U1894 ( .A(n4283), .Y(n4285) );
  INVX2TS U1895 ( .A(n3828), .Y(n3826) );
  CLKBUFX2TS U1896 ( .A(n3716), .Y(n3715) );
  CLKBUFX2TS U1897 ( .A(n3687), .Y(n3682) );
  CLKBUFX2TS U1898 ( .A(n3639), .Y(n3638) );
  CLKBUFX2TS U1899 ( .A(n3716), .Y(n3714) );
  CLKBUFX2TS U1900 ( .A(n552), .Y(n3620) );
  CLKBUFX2TS U1901 ( .A(n3686), .Y(n3683) );
  CLKBUFX2TS U1902 ( .A(n3655), .Y(n3650) );
  CLKBUFX2TS U1903 ( .A(n3624), .Y(n3621) );
  CLKBUFX2TS U1904 ( .A(n3686), .Y(n3684) );
  CLKBUFX2TS U1905 ( .A(n3717), .Y(n3713) );
  CLKBUFX2TS U1906 ( .A(n3640), .Y(n3637) );
  CLKBUFX2TS U1907 ( .A(n3654), .Y(n3651) );
  CLKBUFX2TS U1908 ( .A(n3717), .Y(n3712) );
  CLKBUFX2TS U1909 ( .A(n3640), .Y(n3636) );
  CLKBUFX2TS U1910 ( .A(n3624), .Y(n3622) );
  CLKBUFX2TS U1911 ( .A(n3686), .Y(n3685) );
  CLKBUFX2TS U1912 ( .A(n3654), .Y(n3652) );
  CLKBUFX2TS U1913 ( .A(n3624), .Y(n3623) );
  CLKBUFX2TS U1914 ( .A(n3640), .Y(n3635) );
  CLKBUFX2TS U1915 ( .A(n684), .Y(n676) );
  CLKBUFX2TS U1916 ( .A(n680), .Y(n675) );
  CLKBUFX2TS U1917 ( .A(n680), .Y(n674) );
  CLKBUFX2TS U1918 ( .A(n680), .Y(n673) );
  CLKBUFX2TS U1919 ( .A(n683), .Y(n672) );
  CLKBUFX2TS U1920 ( .A(n681), .Y(n671) );
  CLKBUFX2TS U1921 ( .A(n681), .Y(n670) );
  CLKBUFX2TS U1922 ( .A(n682), .Y(n669) );
  CLKBUFX2TS U1923 ( .A(n682), .Y(n668) );
  CLKBUFX2TS U1924 ( .A(n3653), .Y(n3641) );
  CLKBUFX2TS U1925 ( .A(n3654), .Y(n3653) );
  INVX2TS U1926 ( .A(n1763), .Y(n542) );
  CLKBUFX2TS U1927 ( .A(n3717), .Y(n3711) );
  CLKBUFX2TS U1928 ( .A(n547), .Y(n3701) );
  CLKBUFX2TS U1929 ( .A(n547), .Y(n3702) );
  CLKBUFX2TS U1930 ( .A(n549), .Y(n3672) );
  CLKBUFX2TS U1931 ( .A(n549), .Y(n3671) );
  CLKBUFX2TS U1932 ( .A(n3649), .Y(n3647) );
  CLKBUFX2TS U1933 ( .A(n3649), .Y(n3648) );
  CLKBUFX2TS U1934 ( .A(n3619), .Y(n3618) );
  OAI21X1TS U1935 ( .A0(n531), .A1(n226), .B0(n257), .Y(n1750) );
  NOR2X1TS U1936 ( .A(n226), .B(n1729), .Y(n1580) );
  NOR2X1TS U1937 ( .A(n2264), .B(n538), .Y(n2259) );
  OAI2BB1X1TS U1938 ( .A0N(n1797), .A1N(n1798), .B0(n1799), .Y(n1796) );
  OAI21X1TS U1939 ( .A0(n1798), .A1(n1797), .B0(n316), .Y(n1799) );
  NOR2X1TS U1940 ( .A(n1723), .B(n576), .Y(n958) );
  INVX2TS U1941 ( .A(n2265), .Y(n538) );
  INVX2TS U1942 ( .A(n1678), .Y(n532) );
  OR2X2TS U1943 ( .A(n2259), .B(n2260), .Y(n2258) );
  INVX2TS U1944 ( .A(n1555), .Y(n533) );
  AOI21X1TS U1945 ( .A0(n223), .A1(n532), .B0(n521), .Y(n1724) );
  XNOR2X1TS U1946 ( .A(n553), .B(n873), .Y(n2261) );
  NAND2X1TS U1947 ( .A(n223), .B(n1628), .Y(n1723) );
  NOR2BX1TS U1948 ( .AN(n220), .B(n253), .Y(n1644) );
  AND2X2TS U1949 ( .A(n1644), .B(n223), .Y(n974) );
  AND2X2TS U1950 ( .A(n1618), .B(n241), .Y(n890) );
  AND2X2TS U1951 ( .A(n1618), .B(n239), .Y(n990) );
  AND2X2TS U1952 ( .A(n1644), .B(n1619), .Y(n907) );
  AND2X2TS U1953 ( .A(n1618), .B(n224), .Y(n923) );
  AND2X2TS U1954 ( .A(n1644), .B(n224), .Y(n940) );
  CLKBUFX2TS U1955 ( .A(n701), .Y(n700) );
  CLKBUFX2TS U1956 ( .A(n701), .Y(n699) );
  CLKBUFX2TS U1957 ( .A(n1838), .Y(n667) );
  CLKBUFX2TS U1958 ( .A(n1838), .Y(n666) );
  CLKBUFX2TS U1959 ( .A(n592), .Y(n635) );
  NAND2X1TS U1960 ( .A(n578), .B(n4392), .Y(n875) );
  CLKBUFX2TS U1961 ( .A(n3829), .Y(n3828) );
  CLKBUFX2TS U1962 ( .A(destinationAddressIn_SOUTH[6]), .Y(n4280) );
  CLKBUFX2TS U1963 ( .A(destinationAddressIn_SOUTH[7]), .Y(n4283) );
  CLKBUFX2TS U1964 ( .A(n1839), .Y(n650) );
  CLKBUFX2TS U1965 ( .A(n1839), .Y(n651) );
  CLKBUFX2TS U1966 ( .A(n1903), .Y(n608) );
  CLKBUFX2TS U1967 ( .A(n1903), .Y(n609) );
  CLKBUFX2TS U1968 ( .A(n4306), .Y(n4307) );
  CLKBUFX2TS U1969 ( .A(n4380), .Y(n4381) );
  CLKBUFX2TS U1970 ( .A(dataIn_NORTH[29]), .Y(n4362) );
  CLKBUFX2TS U1971 ( .A(n4350), .Y(n4351) );
  CLKBUFX2TS U1972 ( .A(n4346), .Y(n4347) );
  CLKBUFX2TS U1973 ( .A(dataIn_NORTH[20]), .Y(n4344) );
  CLKBUFX2TS U1974 ( .A(n4330), .Y(n4331) );
  CLKBUFX2TS U1975 ( .A(n4328), .Y(n4329) );
  CLKBUFX2TS U1976 ( .A(n4324), .Y(n4325) );
  CLKBUFX2TS U1977 ( .A(n4316), .Y(n4317) );
  CLKBUFX2TS U1978 ( .A(n4366), .Y(n4367) );
  CLKBUFX2TS U1979 ( .A(n4364), .Y(n4365) );
  CLKBUFX2TS U1980 ( .A(n4360), .Y(n4361) );
  CLKBUFX2TS U1981 ( .A(n4358), .Y(n4359) );
  CLKBUFX2TS U1982 ( .A(dataIn_NORTH[26]), .Y(n4356) );
  CLKBUFX2TS U1983 ( .A(n4352), .Y(n4353) );
  CLKBUFX2TS U1984 ( .A(n4348), .Y(n4349) );
  CLKBUFX2TS U1985 ( .A(n4342), .Y(n4343) );
  CLKBUFX2TS U1986 ( .A(n4336), .Y(n4337) );
  CLKBUFX2TS U1987 ( .A(n4326), .Y(n4327) );
  CLKBUFX2TS U1988 ( .A(n4322), .Y(n4323) );
  CLKBUFX2TS U1989 ( .A(n4320), .Y(n4321) );
  CLKBUFX2TS U1990 ( .A(n4318), .Y(n4319) );
  CLKBUFX2TS U1991 ( .A(dataIn_NORTH[5]), .Y(n4314) );
  CLKBUFX2TS U1992 ( .A(n4308), .Y(n4309) );
  CLKBUFX2TS U1993 ( .A(destinationAddressIn_NORTH[5]), .Y(n4390) );
  CLKBUFX2TS U1994 ( .A(destinationAddressIn_NORTH[3]), .Y(n4386) );
  CLKBUFX2TS U1995 ( .A(n4384), .Y(n4385) );
  CLKBUFX2TS U1996 ( .A(n4382), .Y(n4383) );
  CLKBUFX2TS U1997 ( .A(dataIn_NORTH[0]), .Y(n4304) );
  CLKBUFX2TS U1998 ( .A(n4338), .Y(n4339) );
  CLKBUFX2TS U1999 ( .A(n4334), .Y(n4335) );
  CLKBUFX2TS U2000 ( .A(dataIn_NORTH[14]), .Y(n4332) );
  CLKBUFX2TS U2001 ( .A(dataIn_NORTH[3]), .Y(n4310) );
  CLKBUFX2TS U2002 ( .A(n4388), .Y(n4389) );
  CLKBUFX2TS U2003 ( .A(n4354), .Y(n4355) );
  CLKBUFX2TS U2004 ( .A(n4340), .Y(n4341) );
  CLKBUFX2TS U2005 ( .A(n4312), .Y(n4313) );
  CLKBUFX2TS U2006 ( .A(requesterAddressIn_NORTH[5]), .Y(n4378) );
  CLKBUFX2TS U2007 ( .A(n4376), .Y(n4377) );
  CLKBUFX2TS U2008 ( .A(requesterAddressIn_NORTH[2]), .Y(n4372) );
  CLKBUFX2TS U2009 ( .A(n4374), .Y(n4375) );
  CLKBUFX2TS U2010 ( .A(n4370), .Y(n4371) );
  CLKBUFX2TS U2011 ( .A(n4368), .Y(n4369) );
  INVX2TS U2012 ( .A(n3931), .Y(n3929) );
  INVX2TS U2013 ( .A(n3928), .Y(n3926) );
  INVX2TS U2014 ( .A(n3925), .Y(n3923) );
  INVX2TS U2015 ( .A(n3922), .Y(n3920) );
  INVX2TS U2016 ( .A(n3919), .Y(n3917) );
  INVX2TS U2017 ( .A(n3916), .Y(n3914) );
  INVX2TS U2018 ( .A(n3913), .Y(n3911) );
  INVX2TS U2019 ( .A(n3910), .Y(n3908) );
  INVX2TS U2020 ( .A(n3907), .Y(n3905) );
  INVX2TS U2021 ( .A(n3904), .Y(n3902) );
  INVX2TS U2022 ( .A(n3901), .Y(n3899) );
  INVX2TS U2023 ( .A(n3898), .Y(n3896) );
  INVX2TS U2024 ( .A(n3895), .Y(n3893) );
  INVX2TS U2025 ( .A(n3892), .Y(n3890) );
  INVX2TS U2026 ( .A(n3889), .Y(n3887) );
  INVX2TS U2027 ( .A(n3886), .Y(n3884) );
  INVX2TS U2028 ( .A(n3883), .Y(n3881) );
  INVX2TS U2029 ( .A(n3880), .Y(n3878) );
  INVX2TS U2030 ( .A(n3877), .Y(n3875) );
  INVX2TS U2031 ( .A(n3874), .Y(n3872) );
  INVX2TS U2032 ( .A(n3871), .Y(n3869) );
  INVX2TS U2033 ( .A(n3868), .Y(n3866) );
  INVX2TS U2034 ( .A(n3865), .Y(n3863) );
  INVX2TS U2035 ( .A(n3862), .Y(n3860) );
  INVX2TS U2036 ( .A(n3859), .Y(n3857) );
  INVX2TS U2037 ( .A(n3856), .Y(n3854) );
  INVX2TS U2038 ( .A(n3853), .Y(n3851) );
  INVX2TS U2039 ( .A(n3850), .Y(n3848) );
  INVX2TS U2040 ( .A(n3847), .Y(n3845) );
  INVX2TS U2041 ( .A(n3844), .Y(n3842) );
  INVX2TS U2042 ( .A(n3841), .Y(n3839) );
  INVX2TS U2043 ( .A(n3838), .Y(n3836) );
  INVX2TS U2044 ( .A(n3952), .Y(n3950) );
  INVX2TS U2045 ( .A(n3967), .Y(n3965) );
  INVX2TS U2046 ( .A(n3961), .Y(n3959) );
  INVX2TS U2047 ( .A(n3958), .Y(n3956) );
  INVX2TS U2048 ( .A(n3955), .Y(n3953) );
  INVX2TS U2049 ( .A(n3964), .Y(n3962) );
  INVX2TS U2050 ( .A(n3949), .Y(n3947) );
  INVX2TS U2051 ( .A(n3946), .Y(n3944) );
  INVX2TS U2052 ( .A(n3940), .Y(n3938) );
  INVX2TS U2053 ( .A(n3943), .Y(n3941) );
  INVX2TS U2054 ( .A(n3937), .Y(n3935) );
  INVX2TS U2055 ( .A(n3934), .Y(n3932) );
  INVX2TS U2056 ( .A(n885), .Y(n709) );
  INVX2TS U2057 ( .A(n4102), .Y(n4100) );
  INVX2TS U2058 ( .A(n4105), .Y(n4103) );
  INVX2TS U2059 ( .A(n4096), .Y(n4094) );
  INVX2TS U2060 ( .A(n4099), .Y(n4097) );
  INVX2TS U2061 ( .A(n4093), .Y(n4091) );
  INVX2TS U2062 ( .A(n4090), .Y(n4088) );
  INVX2TS U2063 ( .A(n4255), .Y(n4253) );
  INVX2TS U2064 ( .A(n4252), .Y(n4250) );
  INVX2TS U2065 ( .A(n4249), .Y(n4247) );
  INVX2TS U2066 ( .A(n4246), .Y(n4244) );
  INVX2TS U2067 ( .A(n4261), .Y(n4259) );
  INVX2TS U2068 ( .A(n4258), .Y(n4256) );
  INVX2TS U2069 ( .A(n3822), .Y(n3821) );
  CLKBUFX2TS U2070 ( .A(destinationAddressIn_NORTH[5]), .Y(n4391) );
  CLKBUFX2TS U2071 ( .A(destinationAddressIn_NORTH[3]), .Y(n4387) );
  CLKBUFX2TS U2072 ( .A(dataIn_NORTH[29]), .Y(n4363) );
  CLKBUFX2TS U2073 ( .A(dataIn_NORTH[26]), .Y(n4357) );
  CLKBUFX2TS U2074 ( .A(dataIn_NORTH[14]), .Y(n4333) );
  CLKBUFX2TS U2075 ( .A(dataIn_NORTH[3]), .Y(n4311) );
  CLKBUFX2TS U2076 ( .A(dataIn_NORTH[20]), .Y(n4345) );
  CLKBUFX2TS U2077 ( .A(dataIn_NORTH[5]), .Y(n4315) );
  CLKBUFX2TS U2078 ( .A(dataIn_NORTH[0]), .Y(n4305) );
  INVX2TS U2079 ( .A(n4027), .Y(n4025) );
  INVX2TS U2080 ( .A(n3997), .Y(n3995) );
  INVX2TS U2081 ( .A(n4084), .Y(n4082) );
  INVX2TS U2082 ( .A(n4081), .Y(n4079) );
  INVX2TS U2083 ( .A(n4078), .Y(n4076) );
  INVX2TS U2084 ( .A(n4075), .Y(n4073) );
  INVX2TS U2085 ( .A(n4072), .Y(n4070) );
  INVX2TS U2086 ( .A(n4069), .Y(n4067) );
  INVX2TS U2087 ( .A(n4063), .Y(n4061) );
  INVX2TS U2088 ( .A(n4057), .Y(n4055) );
  INVX2TS U2089 ( .A(n4054), .Y(n4052) );
  INVX2TS U2090 ( .A(n4051), .Y(n4049) );
  INVX2TS U2091 ( .A(n4048), .Y(n4046) );
  INVX2TS U2092 ( .A(n4033), .Y(n4031) );
  INVX2TS U2093 ( .A(n4030), .Y(n4028) );
  INVX2TS U2094 ( .A(n4024), .Y(n4022) );
  INVX2TS U2095 ( .A(n4021), .Y(n4019) );
  INVX2TS U2096 ( .A(n4018), .Y(n4016) );
  INVX2TS U2097 ( .A(n4015), .Y(n4013) );
  INVX2TS U2098 ( .A(n4009), .Y(n4007) );
  INVX2TS U2099 ( .A(n4006), .Y(n4004) );
  INVX2TS U2100 ( .A(n4087), .Y(n4085) );
  INVX2TS U2101 ( .A(n4066), .Y(n4064) );
  INVX2TS U2102 ( .A(n4060), .Y(n4058) );
  INVX2TS U2103 ( .A(n4042), .Y(n4040) );
  INVX2TS U2104 ( .A(n4012), .Y(n4010) );
  INVX2TS U2105 ( .A(n4000), .Y(n3998) );
  INVX2TS U2106 ( .A(n3994), .Y(n3992) );
  INVX2TS U2107 ( .A(n4045), .Y(n4043) );
  INVX2TS U2108 ( .A(n4039), .Y(n4037) );
  INVX2TS U2109 ( .A(n4036), .Y(n4034) );
  INVX2TS U2110 ( .A(n4003), .Y(n4001) );
  INVX2TS U2111 ( .A(n4123), .Y(n4121) );
  INVX2TS U2112 ( .A(n4120), .Y(n4118) );
  INVX2TS U2113 ( .A(n4117), .Y(n4115) );
  INVX2TS U2114 ( .A(n4114), .Y(n4112) );
  INVX2TS U2115 ( .A(n4111), .Y(n4109) );
  INVX2TS U2116 ( .A(n4108), .Y(n4106) );
  INVX2TS U2117 ( .A(n3835), .Y(n3833) );
  CLKBUFX2TS U2118 ( .A(n3986), .Y(n3987) );
  CLKBUFX2TS U2119 ( .A(n3974), .Y(n3975) );
  CLKBUFX2TS U2120 ( .A(n3968), .Y(n3969) );
  CLKBUFX2TS U2121 ( .A(n3983), .Y(n3984) );
  CLKBUFX2TS U2122 ( .A(n3977), .Y(n3978) );
  CLKBUFX2TS U2123 ( .A(n3989), .Y(n3990) );
  CLKBUFX2TS U2124 ( .A(n3980), .Y(n3981) );
  CLKBUFX2TS U2125 ( .A(n3971), .Y(n3972) );
  CLKBUFX2TS U2126 ( .A(n4298), .Y(n4299) );
  CLKBUFX2TS U2127 ( .A(n4292), .Y(n4293) );
  CLKBUFX2TS U2128 ( .A(n4289), .Y(n4290) );
  CLKBUFX2TS U2129 ( .A(n4301), .Y(n4302) );
  CLKBUFX2TS U2130 ( .A(n4295), .Y(n4296) );
  CLKBUFX2TS U2131 ( .A(n4286), .Y(n4287) );
  CLKBUFX2TS U2132 ( .A(n4145), .Y(n4146) );
  CLKBUFX2TS U2133 ( .A(n4142), .Y(n4143) );
  CLKBUFX2TS U2134 ( .A(n4136), .Y(n4137) );
  CLKBUFX2TS U2135 ( .A(n4130), .Y(n4131) );
  CLKBUFX2TS U2136 ( .A(n4124), .Y(n4125) );
  CLKBUFX2TS U2137 ( .A(n4139), .Y(n4140) );
  CLKBUFX2TS U2138 ( .A(n4133), .Y(n4134) );
  CLKBUFX2TS U2139 ( .A(n4127), .Y(n4128) );
  CLKBUFX2TS U2140 ( .A(n4142), .Y(n4144) );
  CLKBUFX2TS U2141 ( .A(n4124), .Y(n4126) );
  CLKBUFX2TS U2142 ( .A(n3986), .Y(n3988) );
  CLKBUFX2TS U2143 ( .A(n3980), .Y(n3982) );
  CLKBUFX2TS U2144 ( .A(n3968), .Y(n3970) );
  CLKBUFX2TS U2145 ( .A(n4136), .Y(n4138) );
  CLKBUFX2TS U2146 ( .A(n4133), .Y(n4135) );
  CLKBUFX2TS U2147 ( .A(n3977), .Y(n3979) );
  CLKBUFX2TS U2148 ( .A(n3989), .Y(n3991) );
  CLKBUFX2TS U2149 ( .A(n4145), .Y(n4147) );
  CLKBUFX2TS U2150 ( .A(n3983), .Y(n3985) );
  CLKBUFX2TS U2151 ( .A(n4139), .Y(n4141) );
  CLKBUFX2TS U2152 ( .A(n3974), .Y(n3976) );
  CLKBUFX2TS U2153 ( .A(n4130), .Y(n4132) );
  CLKBUFX2TS U2154 ( .A(n3971), .Y(n3973) );
  CLKBUFX2TS U2155 ( .A(n4127), .Y(n4129) );
  CLKBUFX2TS U2156 ( .A(n4298), .Y(n4300) );
  CLKBUFX2TS U2157 ( .A(n4286), .Y(n4288) );
  CLKBUFX2TS U2158 ( .A(n4295), .Y(n4297) );
  CLKBUFX2TS U2159 ( .A(n4289), .Y(n4291) );
  CLKBUFX2TS U2160 ( .A(n4301), .Y(n4303) );
  CLKBUFX2TS U2161 ( .A(n4292), .Y(n4294) );
  CLKBUFX2TS U2162 ( .A(requesterAddressIn_NORTH[5]), .Y(n4379) );
  CLKBUFX2TS U2163 ( .A(requesterAddressIn_NORTH[2]), .Y(n4373) );
  INVX2TS U2164 ( .A(n3819), .Y(n3817) );
  INVX2TS U2165 ( .A(n3832), .Y(n3830) );
  INVX2TS U2166 ( .A(n3825), .Y(n3823) );
  INVX2TS U2167 ( .A(n3877), .Y(n3876) );
  INVX2TS U2168 ( .A(n3925), .Y(n3924) );
  INVX2TS U2169 ( .A(n3901), .Y(n3900) );
  INVX2TS U2170 ( .A(n3874), .Y(n3873) );
  INVX2TS U2171 ( .A(n3868), .Y(n3867) );
  INVX2TS U2172 ( .A(n3856), .Y(n3855) );
  INVX2TS U2173 ( .A(n3931), .Y(n3930) );
  INVX2TS U2174 ( .A(n3928), .Y(n3927) );
  INVX2TS U2175 ( .A(n3916), .Y(n3915) );
  INVX2TS U2176 ( .A(n3910), .Y(n3909) );
  INVX2TS U2177 ( .A(n3904), .Y(n3903) );
  INVX2TS U2178 ( .A(n3895), .Y(n3894) );
  INVX2TS U2179 ( .A(n3886), .Y(n3885) );
  INVX2TS U2180 ( .A(n3871), .Y(n3870) );
  INVX2TS U2181 ( .A(n3862), .Y(n3861) );
  INVX2TS U2182 ( .A(n3922), .Y(n3921) );
  INVX2TS U2183 ( .A(n3919), .Y(n3918) );
  INVX2TS U2184 ( .A(n3907), .Y(n3906) );
  INVX2TS U2185 ( .A(n3898), .Y(n3897) );
  INVX2TS U2186 ( .A(n3865), .Y(n3864) );
  INVX2TS U2187 ( .A(n3853), .Y(n3852) );
  INVX2TS U2188 ( .A(n3844), .Y(n3843) );
  INVX2TS U2189 ( .A(n3841), .Y(n3840) );
  INVX2TS U2190 ( .A(n3838), .Y(n3837) );
  INVX2TS U2191 ( .A(n3859), .Y(n3858) );
  INVX2TS U2192 ( .A(n3889), .Y(n3888) );
  INVX2TS U2193 ( .A(n3883), .Y(n3882) );
  INVX2TS U2194 ( .A(n3880), .Y(n3879) );
  INVX2TS U2195 ( .A(n3847), .Y(n3846) );
  INVX2TS U2196 ( .A(n3913), .Y(n3912) );
  INVX2TS U2197 ( .A(n3892), .Y(n3891) );
  INVX2TS U2198 ( .A(n3850), .Y(n3849) );
  INVX2TS U2199 ( .A(n3967), .Y(n3966) );
  INVX2TS U2200 ( .A(n3964), .Y(n3963) );
  INVX2TS U2201 ( .A(n3961), .Y(n3960) );
  INVX2TS U2202 ( .A(n3955), .Y(n3954) );
  INVX2TS U2203 ( .A(n3952), .Y(n3951) );
  INVX2TS U2204 ( .A(n3958), .Y(n3957) );
  INVX2TS U2205 ( .A(n3819), .Y(n3818) );
  INVX2TS U2206 ( .A(n4276), .Y(n4275) );
  INVX2TS U2207 ( .A(n4264), .Y(n4263) );
  INVX2TS U2208 ( .A(n4279), .Y(n4278) );
  INVX2TS U2209 ( .A(n4273), .Y(n4272) );
  INVX2TS U2210 ( .A(n4270), .Y(n4269) );
  INVX2TS U2211 ( .A(n4267), .Y(n4266) );
  INVX2TS U2212 ( .A(n4240), .Y(n4239) );
  INVX2TS U2213 ( .A(n4237), .Y(n4236) );
  INVX2TS U2214 ( .A(n4234), .Y(n4233) );
  INVX2TS U2215 ( .A(n4231), .Y(n4230) );
  INVX2TS U2216 ( .A(n4228), .Y(n4227) );
  INVX2TS U2217 ( .A(n4225), .Y(n4224) );
  INVX2TS U2218 ( .A(n4219), .Y(n4218) );
  INVX2TS U2219 ( .A(n4213), .Y(n4212) );
  INVX2TS U2220 ( .A(n4210), .Y(n4209) );
  INVX2TS U2221 ( .A(n4207), .Y(n4206) );
  INVX2TS U2222 ( .A(n4204), .Y(n4203) );
  INVX2TS U2223 ( .A(n4201), .Y(n4200) );
  INVX2TS U2224 ( .A(n4195), .Y(n4194) );
  INVX2TS U2225 ( .A(n4192), .Y(n4191) );
  INVX2TS U2226 ( .A(n4189), .Y(n4188) );
  INVX2TS U2227 ( .A(n4186), .Y(n4185) );
  INVX2TS U2228 ( .A(n4183), .Y(n4182) );
  INVX2TS U2229 ( .A(n4180), .Y(n4179) );
  INVX2TS U2230 ( .A(n4177), .Y(n4176) );
  INVX2TS U2231 ( .A(n4174), .Y(n4173) );
  INVX2TS U2232 ( .A(n4171), .Y(n4170) );
  INVX2TS U2233 ( .A(n4165), .Y(n4164) );
  INVX2TS U2234 ( .A(n4162), .Y(n4161) );
  INVX2TS U2235 ( .A(n4159), .Y(n4158) );
  INVX2TS U2236 ( .A(n4153), .Y(n4152) );
  INVX2TS U2237 ( .A(n4243), .Y(n4242) );
  INVX2TS U2238 ( .A(n4222), .Y(n4221) );
  INVX2TS U2239 ( .A(n4216), .Y(n4215) );
  INVX2TS U2240 ( .A(n4198), .Y(n4197) );
  INVX2TS U2241 ( .A(n4168), .Y(n4167) );
  INVX2TS U2242 ( .A(n4156), .Y(n4155) );
  INVX2TS U2243 ( .A(n4150), .Y(n4149) );
  INVX2TS U2244 ( .A(n3832), .Y(n3831) );
  INVX2TS U2245 ( .A(n4261), .Y(n4260) );
  INVX2TS U2246 ( .A(n4258), .Y(n4257) );
  INVX2TS U2247 ( .A(n4252), .Y(n4251) );
  INVX2TS U2248 ( .A(n4255), .Y(n4254) );
  INVX2TS U2249 ( .A(n4249), .Y(n4248) );
  INVX2TS U2250 ( .A(n4246), .Y(n4245) );
  INVX2TS U2251 ( .A(n3825), .Y(n3824) );
  INVX2TS U2252 ( .A(n4087), .Y(n4086) );
  INVX2TS U2253 ( .A(n4084), .Y(n4083) );
  INVX2TS U2254 ( .A(n4081), .Y(n4080) );
  INVX2TS U2255 ( .A(n4078), .Y(n4077) );
  INVX2TS U2256 ( .A(n4075), .Y(n4074) );
  INVX2TS U2257 ( .A(n4072), .Y(n4071) );
  INVX2TS U2258 ( .A(n4066), .Y(n4065) );
  INVX2TS U2259 ( .A(n4063), .Y(n4062) );
  INVX2TS U2260 ( .A(n4060), .Y(n4059) );
  INVX2TS U2261 ( .A(n4057), .Y(n4056) );
  INVX2TS U2262 ( .A(n4054), .Y(n4053) );
  INVX2TS U2263 ( .A(n4051), .Y(n4050) );
  INVX2TS U2264 ( .A(n4045), .Y(n4044) );
  INVX2TS U2265 ( .A(n4042), .Y(n4041) );
  INVX2TS U2266 ( .A(n4039), .Y(n4038) );
  INVX2TS U2267 ( .A(n4036), .Y(n4035) );
  INVX2TS U2268 ( .A(n4033), .Y(n4032) );
  INVX2TS U2269 ( .A(n4030), .Y(n4029) );
  INVX2TS U2270 ( .A(n4027), .Y(n4026) );
  INVX2TS U2271 ( .A(n4024), .Y(n4023) );
  INVX2TS U2272 ( .A(n4021), .Y(n4020) );
  INVX2TS U2273 ( .A(n4018), .Y(n4017) );
  INVX2TS U2274 ( .A(n4015), .Y(n4014) );
  INVX2TS U2275 ( .A(n4012), .Y(n4011) );
  INVX2TS U2276 ( .A(n4009), .Y(n4008) );
  INVX2TS U2277 ( .A(n4003), .Y(n4002) );
  INVX2TS U2278 ( .A(n4000), .Y(n3999) );
  INVX2TS U2279 ( .A(n3997), .Y(n3996) );
  INVX2TS U2280 ( .A(n3994), .Y(n3993) );
  INVX2TS U2281 ( .A(n4069), .Y(n4068) );
  INVX2TS U2282 ( .A(n4048), .Y(n4047) );
  INVX2TS U2283 ( .A(n4006), .Y(n4005) );
  INVX2TS U2284 ( .A(n4108), .Y(n4107) );
  INVX2TS U2285 ( .A(n4123), .Y(n4122) );
  INVX2TS U2286 ( .A(n4117), .Y(n4116) );
  INVX2TS U2287 ( .A(n4114), .Y(n4113) );
  INVX2TS U2288 ( .A(n4111), .Y(n4110) );
  INVX2TS U2289 ( .A(n4120), .Y(n4119) );
  INVX2TS U2290 ( .A(n4105), .Y(n4104) );
  INVX2TS U2291 ( .A(n4102), .Y(n4101) );
  INVX2TS U2292 ( .A(n4099), .Y(n4098) );
  INVX2TS U2293 ( .A(n4096), .Y(n4095) );
  INVX2TS U2294 ( .A(n4093), .Y(n4092) );
  INVX2TS U2295 ( .A(n4090), .Y(n4089) );
  INVX2TS U2296 ( .A(n3943), .Y(n3942) );
  INVX2TS U2297 ( .A(n3940), .Y(n3939) );
  INVX2TS U2298 ( .A(n3937), .Y(n3936) );
  INVX2TS U2299 ( .A(n3934), .Y(n3933) );
  INVX2TS U2300 ( .A(n3949), .Y(n3948) );
  INVX2TS U2301 ( .A(n3946), .Y(n3945) );
  INVX2TS U2302 ( .A(n3835), .Y(n3834) );
  INVX2TS U2303 ( .A(n3822), .Y(n3820) );
  INVX2TS U2304 ( .A(n4279), .Y(n4277) );
  INVX2TS U2305 ( .A(n4273), .Y(n4271) );
  INVX2TS U2306 ( .A(n4267), .Y(n4265) );
  INVX2TS U2307 ( .A(n4264), .Y(n4262) );
  INVX2TS U2308 ( .A(n4270), .Y(n4268) );
  INVX2TS U2309 ( .A(n4189), .Y(n4187) );
  INVX2TS U2310 ( .A(n4237), .Y(n4235) );
  INVX2TS U2311 ( .A(n4213), .Y(n4211) );
  INVX2TS U2312 ( .A(n4186), .Y(n4184) );
  INVX2TS U2313 ( .A(n4180), .Y(n4178) );
  INVX2TS U2314 ( .A(n4168), .Y(n4166) );
  INVX2TS U2315 ( .A(n4243), .Y(n4241) );
  INVX2TS U2316 ( .A(n4240), .Y(n4238) );
  INVX2TS U2317 ( .A(n4228), .Y(n4226) );
  INVX2TS U2318 ( .A(n4222), .Y(n4220) );
  INVX2TS U2319 ( .A(n4216), .Y(n4214) );
  INVX2TS U2320 ( .A(n4207), .Y(n4205) );
  INVX2TS U2321 ( .A(n4198), .Y(n4196) );
  INVX2TS U2322 ( .A(n4183), .Y(n4181) );
  INVX2TS U2323 ( .A(n4174), .Y(n4172) );
  INVX2TS U2324 ( .A(n4234), .Y(n4232) );
  INVX2TS U2325 ( .A(n4231), .Y(n4229) );
  INVX2TS U2326 ( .A(n4219), .Y(n4217) );
  INVX2TS U2327 ( .A(n4210), .Y(n4208) );
  INVX2TS U2328 ( .A(n4177), .Y(n4175) );
  INVX2TS U2329 ( .A(n4165), .Y(n4163) );
  INVX2TS U2330 ( .A(n4156), .Y(n4154) );
  INVX2TS U2331 ( .A(n4153), .Y(n4151) );
  INVX2TS U2332 ( .A(n4150), .Y(n4148) );
  INVX2TS U2333 ( .A(n4171), .Y(n4169) );
  INVX2TS U2334 ( .A(n4201), .Y(n4199) );
  INVX2TS U2335 ( .A(n4195), .Y(n4193) );
  INVX2TS U2336 ( .A(n4192), .Y(n4190) );
  INVX2TS U2337 ( .A(n4159), .Y(n4157) );
  INVX2TS U2338 ( .A(n4276), .Y(n4274) );
  INVX2TS U2339 ( .A(n4225), .Y(n4223) );
  INVX2TS U2340 ( .A(n4204), .Y(n4202) );
  INVX2TS U2341 ( .A(n4162), .Y(n4160) );
  INVX2TS U2342 ( .A(n2273), .Y(n539) );
  INVX2TS U2343 ( .A(n2276), .Y(n540) );
  CLKBUFX2TS U2344 ( .A(n683), .Y(n680) );
  CLKBUFX2TS U2345 ( .A(n683), .Y(n681) );
  CLKBUFX2TS U2346 ( .A(n683), .Y(n682) );
  CLKBUFX2TS U2347 ( .A(n15), .Y(n3716) );
  CLKBUFX2TS U2348 ( .A(n275), .Y(n3639) );
  CLKBUFX2TS U2349 ( .A(n275), .Y(n3640) );
  CLKBUFX2TS U2350 ( .A(n550), .Y(n3655) );
  CLKBUFX2TS U2351 ( .A(n15), .Y(n3717) );
  CLKBUFX2TS U2352 ( .A(n3), .Y(n3687) );
  CLKBUFX2TS U2353 ( .A(n3), .Y(n3686) );
  CLKBUFX2TS U2354 ( .A(n550), .Y(n3654) );
  CLKBUFX2TS U2355 ( .A(n552), .Y(n3624) );
  INVX2TS U2356 ( .A(n1834), .Y(n547) );
  CLKBUFX2TS U2357 ( .A(n3656), .Y(n3649) );
  CLKBUFX2TS U2358 ( .A(n550), .Y(n3656) );
  CLKBUFX2TS U2359 ( .A(n3625), .Y(n3619) );
  CLKBUFX2TS U2360 ( .A(n552), .Y(n3625) );
  INVX2TS U2361 ( .A(n1821), .Y(n549) );
  CLKBUFX2TS U2362 ( .A(n679), .Y(n677) );
  CLKBUFX2TS U2363 ( .A(n679), .Y(n678) );
  XNOR2X1TS U2364 ( .A(n2263), .B(n2259), .Y(n876) );
  XNOR2X1TS U2365 ( .A(n2260), .B(n5323), .Y(n2263) );
  XNOR2X1TS U2366 ( .A(n206), .B(n876), .Y(n2262) );
  NOR2X1TS U2367 ( .A(n594), .B(n1802), .Y(n1801) );
  NOR3X1TS U2368 ( .A(n538), .B(n318), .C(n719), .Y(n2260) );
  OAI211X1TS U2369 ( .A0(n2268), .A1(n2269), .B0(n2270), .C0(n2271), .Y(n2265)
         );
  NAND3BX1TS U2370 ( .AN(n880), .B(n882), .C(n2273), .Y(n2270) );
  OAI21X1TS U2371 ( .A0(n207), .A1(n2256), .B0(n2272), .Y(n2271) );
  OAI32X1TS U2372 ( .A0(n2272), .A1(n207), .A2(n2256), .B0(n880), .B1(n2264), 
        .Y(n2269) );
  XOR2X1TS U2373 ( .A(n2256), .B(n208), .Y(n2264) );
  XOR2X1TS U2374 ( .A(n2254), .B(n2255), .Y(n877) );
  NOR3X1TS U2375 ( .A(n2256), .B(n538), .C(n207), .Y(n2255) );
  XNOR2X1TS U2376 ( .A(n5326), .B(n2257), .Y(n2254) );
  AOI22X1TS U2377 ( .A0(n2258), .A1(n6), .B0(n2259), .B1(n2260), .Y(n2257) );
  INVX2TS U2378 ( .A(n2278), .Y(n720) );
  INVX2TS U2379 ( .A(n1802), .Y(n531) );
  INVX2TS U2380 ( .A(n2267), .Y(n719) );
  OAI221XLTS U2381 ( .A0(n2), .A1(n291), .B0(n3431), .B1(n21), .C0(n1536), .Y(
        n2576) );
  AOI222XLTS U2382 ( .A0(n3817), .A1(n3399), .B0(n3831), .B1(n359), .C0(n3823), 
        .C1(n3421), .Y(n1536) );
  OAI221XLTS U2383 ( .A0(n449), .A1(n291), .B0(n3562), .B1(n558), .C0(n1532), 
        .Y(n2578) );
  AOI222XLTS U2384 ( .A0(n3817), .A1(n3506), .B0(n3831), .B1(n3516), .C0(n3824), .C1(n3552), .Y(n1532) );
  AOI211X1TS U2385 ( .A0(n880), .A1(n2264), .B0(n539), .C0(n719), .Y(n2268) );
  NOR2X1TS U2386 ( .A(n529), .B(n5326), .Y(n1561) );
  XOR2X1TS U2387 ( .A(n2266), .B(n13), .Y(n873) );
  NAND2X1TS U2388 ( .A(n2267), .B(n2265), .Y(n2266) );
  OAI33XLTS U2389 ( .A0(n744), .A1(n530), .A2(n1576), .B0(n3829), .B1(n519), 
        .B2(n1577), .Y(n1575) );
  NAND2X1TS U2390 ( .A(n3820), .B(n520), .Y(n1594) );
  INVX2TS U2391 ( .A(n3828), .Y(n3827) );
  NAND2X1TS U2392 ( .A(n3820), .B(n523), .Y(n1565) );
  NOR2X1TS U2393 ( .A(n1811), .B(n713), .Y(n1839) );
  NOR2X1TS U2394 ( .A(n1812), .B(n713), .Y(n1838) );
  OAI2BB2XLTS U2395 ( .B0(n1598), .B1(n744), .A0N(n1598), .A1N(n3833), .Y(
        n1570) );
  INVX2TS U2396 ( .A(n1805), .Y(n701) );
  NAND4X1TS U2397 ( .A(n1811), .B(n1813), .C(n1815), .D(n2248), .Y(n1805) );
  AND3X2TS U2398 ( .A(n1825), .B(n1812), .C(n1814), .Y(n2248) );
  OAI222X1TS U2399 ( .A0(n3822), .A1(n1811), .B0(n3828), .B1(n1812), .C0(n235), 
        .C1(n1813), .Y(n1810) );
  OR2X2TS U2400 ( .A(n1814), .B(n713), .Y(n592) );
  OAI211X1TS U2401 ( .A0(n3835), .A1(n1814), .B0(n1815), .C0(n710), .Y(n1809)
         );
  INVX2TS U2402 ( .A(n1825), .Y(n713) );
  NOR2X1TS U2403 ( .A(n710), .B(reset), .Y(n885) );
  NOR2X1TS U2404 ( .A(n1815), .B(n465), .Y(n1903) );
  INVX2TS U2405 ( .A(readIn_NORTH), .Y(n3835) );
  INVX2TS U2406 ( .A(writeIn_SOUTH), .Y(n3832) );
  INVX2TS U2407 ( .A(writeIn_WEST), .Y(n3819) );
  OAI221XLTS U2408 ( .A0(n290), .A1(n1814), .B0(n3825), .B1(n1812), .C0(n710), 
        .Y(n1826) );
  INVX2TS U2409 ( .A(readIn_WEST), .Y(n3822) );
  INVX2TS U2410 ( .A(requesterAddressIn_EAST[5]), .Y(n4105) );
  INVX2TS U2411 ( .A(requesterAddressIn_EAST[3]), .Y(n4099) );
  INVX2TS U2412 ( .A(requesterAddressIn_EAST[4]), .Y(n4102) );
  INVX2TS U2413 ( .A(requesterAddressIn_EAST[2]), .Y(n4096) );
  INVX2TS U2414 ( .A(requesterAddressIn_EAST[1]), .Y(n4093) );
  INVX2TS U2415 ( .A(requesterAddressIn_EAST[0]), .Y(n4090) );
  INVX2TS U2416 ( .A(dataIn_EAST[31]), .Y(n4087) );
  INVX2TS U2417 ( .A(dataIn_EAST[30]), .Y(n4084) );
  INVX2TS U2418 ( .A(dataIn_EAST[29]), .Y(n4081) );
  INVX2TS U2419 ( .A(dataIn_EAST[26]), .Y(n4072) );
  INVX2TS U2420 ( .A(dataIn_EAST[24]), .Y(n4066) );
  INVX2TS U2421 ( .A(dataIn_EAST[22]), .Y(n4060) );
  INVX2TS U2422 ( .A(dataIn_EAST[21]), .Y(n4057) );
  INVX2TS U2423 ( .A(dataIn_EAST[19]), .Y(n4051) );
  INVX2TS U2424 ( .A(dataIn_EAST[17]), .Y(n4045) );
  INVX2TS U2425 ( .A(dataIn_EAST[16]), .Y(n4042) );
  INVX2TS U2426 ( .A(dataIn_EAST[14]), .Y(n4036) );
  INVX2TS U2427 ( .A(dataIn_EAST[12]), .Y(n4030) );
  INVX2TS U2428 ( .A(dataIn_EAST[11]), .Y(n4027) );
  INVX2TS U2429 ( .A(dataIn_EAST[10]), .Y(n4024) );
  INVX2TS U2430 ( .A(dataIn_EAST[8]), .Y(n4018) );
  INVX2TS U2431 ( .A(dataIn_EAST[6]), .Y(n4012) );
  INVX2TS U2432 ( .A(dataIn_EAST[3]), .Y(n4003) );
  INVX2TS U2433 ( .A(dataIn_EAST[25]), .Y(n4069) );
  INVX2TS U2434 ( .A(dataIn_EAST[18]), .Y(n4048) );
  INVX2TS U2435 ( .A(dataIn_EAST[15]), .Y(n4039) );
  INVX2TS U2436 ( .A(dataIn_EAST[13]), .Y(n4033) );
  INVX2TS U2437 ( .A(dataIn_EAST[4]), .Y(n4006) );
  INVX2TS U2438 ( .A(dataIn_EAST[28]), .Y(n4078) );
  INVX2TS U2439 ( .A(dataIn_EAST[27]), .Y(n4075) );
  INVX2TS U2440 ( .A(dataIn_EAST[23]), .Y(n4063) );
  INVX2TS U2441 ( .A(dataIn_EAST[20]), .Y(n4054) );
  INVX2TS U2442 ( .A(dataIn_EAST[9]), .Y(n4021) );
  INVX2TS U2443 ( .A(dataIn_EAST[5]), .Y(n4009) );
  INVX2TS U2444 ( .A(dataIn_EAST[2]), .Y(n4000) );
  INVX2TS U2445 ( .A(dataIn_EAST[1]), .Y(n3997) );
  INVX2TS U2446 ( .A(dataIn_EAST[0]), .Y(n3994) );
  INVX2TS U2447 ( .A(dataIn_EAST[7]), .Y(n4015) );
  INVX2TS U2448 ( .A(requesterAddressIn_WEST[4]), .Y(n3946) );
  INVX2TS U2449 ( .A(requesterAddressIn_WEST[1]), .Y(n3937) );
  INVX2TS U2450 ( .A(requesterAddressIn_WEST[0]), .Y(n3934) );
  INVX2TS U2451 ( .A(requesterAddressIn_WEST[5]), .Y(n3949) );
  INVX2TS U2452 ( .A(requesterAddressIn_WEST[3]), .Y(n3943) );
  INVX2TS U2453 ( .A(requesterAddressIn_WEST[2]), .Y(n3940) );
  INVX2TS U2454 ( .A(destinationAddressIn_EAST[5]), .Y(n4123) );
  INVX2TS U2455 ( .A(destinationAddressIn_EAST[3]), .Y(n4117) );
  INVX2TS U2456 ( .A(destinationAddressIn_EAST[1]), .Y(n4111) );
  INVX2TS U2457 ( .A(destinationAddressIn_EAST[4]), .Y(n4120) );
  INVX2TS U2458 ( .A(destinationAddressIn_EAST[0]), .Y(n4108) );
  INVX2TS U2459 ( .A(destinationAddressIn_EAST[2]), .Y(n4114) );
  INVX2TS U2460 ( .A(writeIn_EAST), .Y(n3825) );
  INVX2TS U2461 ( .A(destinationAddressIn_SOUTH[0]), .Y(n4264) );
  INVX2TS U2462 ( .A(requesterAddressIn_SOUTH[5]), .Y(n4261) );
  INVX2TS U2463 ( .A(requesterAddressIn_SOUTH[4]), .Y(n4258) );
  INVX2TS U2464 ( .A(requesterAddressIn_SOUTH[2]), .Y(n4252) );
  INVX2TS U2465 ( .A(destinationAddressIn_SOUTH[5]), .Y(n4279) );
  INVX2TS U2466 ( .A(destinationAddressIn_SOUTH[3]), .Y(n4273) );
  INVX2TS U2467 ( .A(destinationAddressIn_SOUTH[2]), .Y(n4270) );
  INVX2TS U2468 ( .A(destinationAddressIn_SOUTH[1]), .Y(n4267) );
  INVX2TS U2469 ( .A(dataIn_SOUTH[30]), .Y(n4240) );
  INVX2TS U2470 ( .A(dataIn_SOUTH[29]), .Y(n4237) );
  INVX2TS U2471 ( .A(dataIn_SOUTH[26]), .Y(n4228) );
  INVX2TS U2472 ( .A(dataIn_SOUTH[21]), .Y(n4213) );
  INVX2TS U2473 ( .A(dataIn_SOUTH[19]), .Y(n4207) );
  INVX2TS U2474 ( .A(dataIn_SOUTH[13]), .Y(n4189) );
  INVX2TS U2475 ( .A(dataIn_SOUTH[12]), .Y(n4186) );
  INVX2TS U2476 ( .A(dataIn_SOUTH[11]), .Y(n4183) );
  INVX2TS U2477 ( .A(dataIn_SOUTH[10]), .Y(n4180) );
  INVX2TS U2478 ( .A(dataIn_SOUTH[8]), .Y(n4174) );
  INVX2TS U2479 ( .A(requesterAddressIn_SOUTH[3]), .Y(n4255) );
  INVX2TS U2480 ( .A(requesterAddressIn_SOUTH[1]), .Y(n4249) );
  INVX2TS U2481 ( .A(requesterAddressIn_SOUTH[0]), .Y(n4246) );
  INVX2TS U2482 ( .A(dataIn_SOUTH[28]), .Y(n4234) );
  INVX2TS U2483 ( .A(dataIn_SOUTH[27]), .Y(n4231) );
  INVX2TS U2484 ( .A(dataIn_SOUTH[23]), .Y(n4219) );
  INVX2TS U2485 ( .A(dataIn_SOUTH[20]), .Y(n4210) );
  INVX2TS U2486 ( .A(dataIn_SOUTH[9]), .Y(n4177) );
  INVX2TS U2487 ( .A(dataIn_SOUTH[5]), .Y(n4165) );
  INVX2TS U2488 ( .A(dataIn_SOUTH[1]), .Y(n4153) );
  INVX2TS U2489 ( .A(dataIn_SOUTH[31]), .Y(n4243) );
  INVX2TS U2490 ( .A(dataIn_SOUTH[24]), .Y(n4222) );
  INVX2TS U2491 ( .A(dataIn_SOUTH[22]), .Y(n4216) );
  INVX2TS U2492 ( .A(dataIn_SOUTH[16]), .Y(n4198) );
  INVX2TS U2493 ( .A(dataIn_SOUTH[6]), .Y(n4168) );
  INVX2TS U2494 ( .A(dataIn_SOUTH[2]), .Y(n4156) );
  INVX2TS U2495 ( .A(dataIn_SOUTH[0]), .Y(n4150) );
  INVX2TS U2496 ( .A(dataIn_SOUTH[7]), .Y(n4171) );
  INVX2TS U2497 ( .A(dataIn_SOUTH[17]), .Y(n4201) );
  INVX2TS U2498 ( .A(dataIn_SOUTH[15]), .Y(n4195) );
  INVX2TS U2499 ( .A(dataIn_SOUTH[14]), .Y(n4192) );
  INVX2TS U2500 ( .A(dataIn_SOUTH[3]), .Y(n4159) );
  INVX2TS U2501 ( .A(destinationAddressIn_SOUTH[4]), .Y(n4276) );
  INVX2TS U2502 ( .A(dataIn_SOUTH[25]), .Y(n4225) );
  INVX2TS U2503 ( .A(dataIn_SOUTH[18]), .Y(n4204) );
  INVX2TS U2504 ( .A(dataIn_SOUTH[4]), .Y(n4162) );
  INVX2TS U2505 ( .A(dataIn_WEST[31]), .Y(n3931) );
  INVX2TS U2506 ( .A(dataIn_WEST[30]), .Y(n3928) );
  INVX2TS U2507 ( .A(dataIn_WEST[29]), .Y(n3925) );
  INVX2TS U2508 ( .A(dataIn_WEST[26]), .Y(n3916) );
  INVX2TS U2509 ( .A(dataIn_WEST[24]), .Y(n3910) );
  INVX2TS U2510 ( .A(dataIn_WEST[22]), .Y(n3904) );
  INVX2TS U2511 ( .A(dataIn_WEST[21]), .Y(n3901) );
  INVX2TS U2512 ( .A(dataIn_WEST[19]), .Y(n3895) );
  INVX2TS U2513 ( .A(dataIn_WEST[16]), .Y(n3886) );
  INVX2TS U2514 ( .A(dataIn_WEST[13]), .Y(n3877) );
  INVX2TS U2515 ( .A(dataIn_WEST[12]), .Y(n3874) );
  INVX2TS U2516 ( .A(dataIn_WEST[11]), .Y(n3871) );
  INVX2TS U2517 ( .A(dataIn_WEST[10]), .Y(n3868) );
  INVX2TS U2518 ( .A(dataIn_WEST[8]), .Y(n3862) );
  INVX2TS U2519 ( .A(dataIn_WEST[6]), .Y(n3856) );
  INVX2TS U2520 ( .A(dataIn_WEST[28]), .Y(n3922) );
  INVX2TS U2521 ( .A(dataIn_WEST[27]), .Y(n3919) );
  INVX2TS U2522 ( .A(dataIn_WEST[23]), .Y(n3907) );
  INVX2TS U2523 ( .A(dataIn_WEST[20]), .Y(n3898) );
  INVX2TS U2524 ( .A(dataIn_WEST[9]), .Y(n3865) );
  INVX2TS U2525 ( .A(dataIn_WEST[5]), .Y(n3853) );
  INVX2TS U2526 ( .A(dataIn_WEST[2]), .Y(n3844) );
  INVX2TS U2527 ( .A(dataIn_WEST[1]), .Y(n3841) );
  INVX2TS U2528 ( .A(dataIn_WEST[0]), .Y(n3838) );
  INVX2TS U2529 ( .A(dataIn_WEST[7]), .Y(n3859) );
  INVX2TS U2530 ( .A(dataIn_WEST[17]), .Y(n3889) );
  INVX2TS U2531 ( .A(dataIn_WEST[15]), .Y(n3883) );
  INVX2TS U2532 ( .A(dataIn_WEST[14]), .Y(n3880) );
  INVX2TS U2533 ( .A(dataIn_WEST[3]), .Y(n3847) );
  INVX2TS U2534 ( .A(dataIn_WEST[25]), .Y(n3913) );
  INVX2TS U2535 ( .A(dataIn_WEST[18]), .Y(n3892) );
  INVX2TS U2536 ( .A(dataIn_WEST[4]), .Y(n3850) );
  INVX2TS U2537 ( .A(destinationAddressIn_WEST[0]), .Y(n3952) );
  INVX2TS U2538 ( .A(destinationAddressIn_WEST[5]), .Y(n3967) );
  INVX2TS U2539 ( .A(destinationAddressIn_WEST[3]), .Y(n3961) );
  INVX2TS U2540 ( .A(destinationAddressIn_WEST[2]), .Y(n3958) );
  INVX2TS U2541 ( .A(destinationAddressIn_WEST[1]), .Y(n3955) );
  INVX2TS U2542 ( .A(destinationAddressIn_WEST[4]), .Y(n3964) );
  NOR2BX1TS U2543 ( .AN(n457), .B(n878), .Y(n2885) );
  AOI31X1TS U2544 ( .A0(n879), .A1(n539), .A2(n880), .B0(n3607), .Y(n878) );
  XNOR2X1TS U2545 ( .A(n881), .B(n882), .Y(n879) );
  CLKBUFX2TS U2546 ( .A(destinationAddressIn_EAST[6]), .Y(n4124) );
  CLKBUFX2TS U2547 ( .A(destinationAddressIn_WEST[6]), .Y(n3968) );
  CLKBUFX2TS U2548 ( .A(destinationAddressIn_EAST[10]), .Y(n4136) );
  CLKBUFX2TS U2549 ( .A(destinationAddressIn_SOUTH[10]), .Y(n4292) );
  CLKBUFX2TS U2550 ( .A(destinationAddressIn_WEST[10]), .Y(n3980) );
  CLKBUFX2TS U2551 ( .A(destinationAddressIn_NORTH[0]), .Y(n4380) );
  CLKBUFX2TS U2552 ( .A(requesterAddressIn_NORTH[4]), .Y(n4376) );
  CLKBUFX2TS U2553 ( .A(destinationAddressIn_EAST[12]), .Y(n4142) );
  CLKBUFX2TS U2554 ( .A(destinationAddressIn_NORTH[2]), .Y(n4384) );
  CLKBUFX2TS U2555 ( .A(destinationAddressIn_NORTH[1]), .Y(n4382) );
  CLKBUFX2TS U2556 ( .A(dataIn_NORTH[30]), .Y(n4364) );
  CLKBUFX2TS U2557 ( .A(dataIn_NORTH[21]), .Y(n4346) );
  CLKBUFX2TS U2558 ( .A(dataIn_NORTH[19]), .Y(n4342) );
  CLKBUFX2TS U2559 ( .A(dataIn_NORTH[13]), .Y(n4330) );
  CLKBUFX2TS U2560 ( .A(dataIn_NORTH[12]), .Y(n4328) );
  CLKBUFX2TS U2561 ( .A(dataIn_NORTH[11]), .Y(n4326) );
  CLKBUFX2TS U2562 ( .A(dataIn_NORTH[10]), .Y(n4324) );
  CLKBUFX2TS U2563 ( .A(dataIn_NORTH[8]), .Y(n4320) );
  CLKBUFX2TS U2564 ( .A(requesterAddressIn_NORTH[3]), .Y(n4374) );
  CLKBUFX2TS U2565 ( .A(requesterAddressIn_NORTH[1]), .Y(n4370) );
  CLKBUFX2TS U2566 ( .A(requesterAddressIn_NORTH[0]), .Y(n4368) );
  CLKBUFX2TS U2567 ( .A(dataIn_NORTH[28]), .Y(n4360) );
  CLKBUFX2TS U2568 ( .A(dataIn_NORTH[27]), .Y(n4358) );
  CLKBUFX2TS U2569 ( .A(dataIn_NORTH[23]), .Y(n4350) );
  CLKBUFX2TS U2570 ( .A(dataIn_NORTH[9]), .Y(n4322) );
  CLKBUFX2TS U2571 ( .A(dataIn_NORTH[1]), .Y(n4306) );
  CLKBUFX2TS U2572 ( .A(destinationAddressIn_WEST[12]), .Y(n3986) );
  CLKBUFX2TS U2573 ( .A(destinationAddressIn_SOUTH[12]), .Y(n4298) );
  CLKBUFX2TS U2574 ( .A(dataIn_NORTH[31]), .Y(n4366) );
  CLKBUFX2TS U2575 ( .A(dataIn_NORTH[24]), .Y(n4352) );
  CLKBUFX2TS U2576 ( .A(dataIn_NORTH[22]), .Y(n4348) );
  CLKBUFX2TS U2577 ( .A(dataIn_NORTH[16]), .Y(n4336) );
  CLKBUFX2TS U2578 ( .A(dataIn_NORTH[6]), .Y(n4316) );
  CLKBUFX2TS U2579 ( .A(dataIn_NORTH[2]), .Y(n4308) );
  CLKBUFX2TS U2580 ( .A(dataIn_NORTH[7]), .Y(n4318) );
  CLKBUFX2TS U2581 ( .A(destinationAddressIn_EAST[9]), .Y(n4133) );
  CLKBUFX2TS U2582 ( .A(destinationAddressIn_WEST[9]), .Y(n3977) );
  CLKBUFX2TS U2583 ( .A(destinationAddressIn_SOUTH[9]), .Y(n4289) );
  CLKBUFX2TS U2584 ( .A(dataIn_NORTH[17]), .Y(n4338) );
  CLKBUFX2TS U2585 ( .A(dataIn_NORTH[15]), .Y(n4334) );
  CLKBUFX2TS U2586 ( .A(destinationAddressIn_WEST[13]), .Y(n3989) );
  CLKBUFX2TS U2587 ( .A(destinationAddressIn_EAST[13]), .Y(n4145) );
  CLKBUFX2TS U2588 ( .A(destinationAddressIn_SOUTH[13]), .Y(n4301) );
  CLKBUFX2TS U2589 ( .A(destinationAddressIn_WEST[11]), .Y(n3983) );
  CLKBUFX2TS U2590 ( .A(destinationAddressIn_EAST[11]), .Y(n4139) );
  CLKBUFX2TS U2591 ( .A(destinationAddressIn_SOUTH[11]), .Y(n4295) );
  CLKBUFX2TS U2592 ( .A(destinationAddressIn_WEST[8]), .Y(n3974) );
  CLKBUFX2TS U2593 ( .A(destinationAddressIn_EAST[8]), .Y(n4130) );
  CLKBUFX2TS U2594 ( .A(destinationAddressIn_SOUTH[8]), .Y(n4286) );
  CLKBUFX2TS U2595 ( .A(destinationAddressIn_WEST[7]), .Y(n3971) );
  CLKBUFX2TS U2596 ( .A(destinationAddressIn_EAST[7]), .Y(n4127) );
  CLKBUFX2TS U2597 ( .A(destinationAddressIn_NORTH[4]), .Y(n4388) );
  CLKBUFX2TS U2598 ( .A(dataIn_NORTH[25]), .Y(n4354) );
  CLKBUFX2TS U2599 ( .A(dataIn_NORTH[18]), .Y(n4340) );
  CLKBUFX2TS U2600 ( .A(dataIn_NORTH[4]), .Y(n4312) );
  INVX2TS U2601 ( .A(readIn_EAST), .Y(n3829) );
  OAI21X1TS U2602 ( .A0(n710), .A1(n881), .B0(n4392), .Y(n883) );
  OAI22X1TS U2603 ( .A0(n3594), .A1(n3677), .B0(n205), .B1(n883), .Y(n2884) );
  XNOR2X1TS U2604 ( .A(n279), .B(n205), .Y(n882) );
  AOI21X1TS U2605 ( .A0(n9), .A1(n5327), .B0(n2276), .Y(n2273) );
  XNOR2X1TS U2606 ( .A(n882), .B(n2274), .Y(n2272) );
  AOI21X1TS U2607 ( .A0(n594), .A1(n540), .B0(n2275), .Y(n2274) );
  AOI21X1TS U2608 ( .A0(n2276), .A1(n6), .B0(n206), .Y(n2275) );
  OAI22X1TS U2609 ( .A0(n22), .A1(n671), .B0(n627), .B1(n3660), .Y(n1990) );
  OAI22X1TS U2610 ( .A0(n23), .A1(n670), .B0(n626), .B1(n3659), .Y(n1982) );
  OAI22X1TS U2611 ( .A0(n24), .A1(n670), .B0(n625), .B1(n3659), .Y(n1966) );
  OAI22X1TS U2612 ( .A0(n25), .A1(n670), .B0(n586), .B1(n3659), .Y(n1958) );
  OAI22X1TS U2613 ( .A0(n26), .A1(n670), .B0(n587), .B1(n3659), .Y(n1974) );
  OAI22X1TS U2614 ( .A0(n27), .A1(n669), .B0(n585), .B1(n3658), .Y(n1950) );
  CLKBUFX2TS U2615 ( .A(n1818), .Y(n683) );
  INVX2TS U2616 ( .A(n1820), .Y(n550) );
  INVX2TS U2617 ( .A(n1831), .Y(n552) );
  NOR2X1TS U2618 ( .A(n881), .B(n205), .Y(n1821) );
  INVX2TS U2619 ( .A(n319), .Y(n553) );
  CLKBUFX2TS U2620 ( .A(n684), .Y(n679) );
  CLKBUFX2TS U2621 ( .A(n1818), .Y(n684) );
  NOR2X1TS U2622 ( .A(selectBit_SOUTH), .B(selectBit_NORTH), .Y(n2249) );
  AOI222XLTS U2623 ( .A0(n3987), .A1(n770), .B0(n4300), .B1(n746), .C0(n4143), 
        .C1(n1549), .Y(n1793) );
  AOI222XLTS U2624 ( .A0(n3975), .A1(n771), .B0(n4288), .B1(n745), .C0(n4131), 
        .C1(n575), .Y(n1789) );
  AOI222XLTS U2625 ( .A0(n4302), .A1(n1669), .B0(destinationAddressIn_EAST[13]), .B1(n870), .C0(n3991), .C1(n3215), .Y(n1749) );
  AOI222XLTS U2626 ( .A0(n3981), .A1(n770), .B0(n4294), .B1(n746), .C0(n4137), 
        .C1(n574), .Y(n1791) );
  AOI222XLTS U2627 ( .A0(n3969), .A1(n771), .B0(n4282), .B1(n745), .C0(n4125), 
        .C1(n575), .Y(n1787) );
  AOI222XLTS U2628 ( .A0(n3817), .A1(n772), .B0(n3830), .B1(n745), .C0(n3823), 
        .C1(n574), .Y(n1548) );
  AOI222XLTS U2629 ( .A0(n4290), .A1(n1728), .B0(destinationAddressIn_EAST[9]), 
        .B1(n864), .C0(n3979), .C1(n3216), .Y(n1745) );
  AOI222XLTS U2630 ( .A0(n4284), .A1(n1728), .B0(destinationAddressIn_EAST[7]), 
        .B1(n863), .C0(n3973), .C1(n3217), .Y(n1743) );
  AOI222XLTS U2631 ( .A0(n3830), .A1(n1817), .B0(n3824), .B1(n863), .C0(n3818), 
        .C1(n3217), .Y(n1543) );
  AOI222XLTS U2632 ( .A0(n3984), .A1(n770), .B0(n4297), .B1(n746), .C0(n4140), 
        .C1(n575), .Y(n1792) );
  AOI222XLTS U2633 ( .A0(n3978), .A1(n771), .B0(n4291), .B1(n746), .C0(n4134), 
        .C1(n574), .Y(n1790) );
  AOI222XLTS U2634 ( .A0(n3972), .A1(n771), .B0(n4285), .B1(n745), .C0(n4128), 
        .C1(n575), .Y(n1788) );
  AOI222XLTS U2635 ( .A0(n4299), .A1(n1669), .B0(destinationAddressIn_EAST[12]), .B1(n864), .C0(n3988), .C1(n3215), .Y(n1748) );
  AOI222XLTS U2636 ( .A0(n4293), .A1(n1669), .B0(destinationAddressIn_EAST[10]), .B1(n864), .C0(n3982), .C1(n3216), .Y(n1746) );
  AOI222XLTS U2637 ( .A0(n4287), .A1(n1728), .B0(destinationAddressIn_EAST[8]), 
        .B1(n863), .C0(n3976), .C1(n3216), .Y(n1744) );
  AOI222XLTS U2638 ( .A0(n4281), .A1(n1728), .B0(destinationAddressIn_EAST[6]), 
        .B1(n863), .C0(n3970), .C1(n3217), .Y(n1742) );
  NOR2X1TS U2639 ( .A(selectBit_WEST), .B(readReady), .Y(n2250) );
  INVX2TS U2640 ( .A(selectBit_EAST), .Y(n778) );
  OAI22X1TS U2641 ( .A0(n877), .A1(n458), .B0(n5326), .B1(n875), .Y(n2886) );
  INVX2TS U2642 ( .A(readReady), .Y(n872) );
  OAI32X1TS U2643 ( .A0(n2252), .A1(n458), .A2(n2253), .B0(n465), .B1(n150), 
        .Y(N4718) );
  NAND2X1TS U2644 ( .A(n2261), .B(n2262), .Y(n2252) );
  XNOR2X1TS U2645 ( .A(n236), .B(n877), .Y(n2253) );
  OAI221XLTS U2646 ( .A0(n204), .A1(n299), .B0(n2340), .B1(n702), .C0(n1651), 
        .Y(n2536) );
  AOI222XLTS U2647 ( .A0(n4299), .A1(n3490), .B0(n4144), .B1(n908), .C0(n3988), 
        .C1(n3728), .Y(n1651) );
  OAI221XLTS U2648 ( .A0(n1533), .A1(n302), .B0(n2328), .B1(n703), .C0(n1649), 
        .Y(n2538) );
  AOI222XLTS U2649 ( .A0(n4293), .A1(n3490), .B0(n4138), .B1(n3462), .C0(n3982), .C1(n3727), .Y(n1649) );
  OAI221XLTS U2650 ( .A0(n1533), .A1(n305), .B0(n2320), .B1(n703), .C0(n1648), 
        .Y(n2539) );
  AOI222XLTS U2651 ( .A0(n4290), .A1(n3494), .B0(n4135), .B1(n3463), .C0(n3979), .C1(n3727), .Y(n1648) );
  OAI221XLTS U2652 ( .A0(n453), .A1(n293), .B0(n2296), .B1(n704), .C0(n1645), 
        .Y(n2542) );
  AOI222XLTS U2653 ( .A0(n4281), .A1(n3496), .B0(n4126), .B1(n3463), .C0(n3970), .C1(n3728), .Y(n1645) );
  OAI221XLTS U2654 ( .A0(n453), .A1(n311), .B0(n2330), .B1(n702), .C0(n1650), 
        .Y(n2537) );
  AOI222XLTS U2655 ( .A0(n4296), .A1(n906), .B0(n4141), .B1(n3459), .C0(n3985), 
        .C1(n3728), .Y(n1650) );
  OAI221XLTS U2656 ( .A0(n453), .A1(n314), .B0(n2306), .B1(n703), .C0(n1647), 
        .Y(n2540) );
  AOI222XLTS U2657 ( .A0(n4287), .A1(n3490), .B0(n4132), .B1(n3463), .C0(n3976), .C1(n3727), .Y(n1647) );
  OAI221XLTS U2658 ( .A0(n1533), .A1(n295), .B0(n2300), .B1(n703), .C0(n1646), 
        .Y(n2541) );
  AOI222XLTS U2659 ( .A0(n4284), .A1(n3494), .B0(n4129), .B1(n3460), .C0(n3973), .C1(n3727), .Y(n1646) );
  OAI221XLTS U2660 ( .A0(n446), .A1(n309), .B0(n2351), .B1(n839), .C0(n1772), 
        .Y(n2465) );
  OAI221XLTS U2661 ( .A0(n445), .A1(n299), .B0(n2343), .B1(n838), .C0(n1771), 
        .Y(n2466) );
  AOI222XLTS U2662 ( .A0(n4143), .A1(n796), .B0(destinationAddressIn_SOUTH[12]), .B1(n266), .C0(n3988), .C1(n828), .Y(n1771) );
  OAI221XLTS U2663 ( .A0(n446), .A1(n311), .B0(n2333), .B1(n839), .C0(n1770), 
        .Y(n2467) );
  AOI222XLTS U2664 ( .A0(n4140), .A1(n796), .B0(destinationAddressIn_SOUTH[11]), .B1(n269), .C0(n3985), .C1(n828), .Y(n1770) );
  OAI221XLTS U2665 ( .A0(n445), .A1(n302), .B0(n2327), .B1(n839), .C0(n1769), 
        .Y(n2468) );
  AOI222XLTS U2666 ( .A0(n4137), .A1(n796), .B0(destinationAddressIn_SOUTH[10]), .B1(n378), .C0(n3982), .C1(n828), .Y(n1769) );
  OAI221XLTS U2667 ( .A0(n446), .A1(n305), .B0(n2315), .B1(n840), .C0(n1768), 
        .Y(n2469) );
  AOI222XLTS U2668 ( .A0(n4134), .A1(n796), .B0(destinationAddressIn_SOUTH[9]), 
        .B1(n378), .C0(n3979), .C1(n828), .Y(n1768) );
  OAI221XLTS U2669 ( .A0(n445), .A1(n314), .B0(n2311), .B1(n840), .C0(n1767), 
        .Y(n2470) );
  AOI222XLTS U2670 ( .A0(n4131), .A1(n797), .B0(destinationAddressIn_SOUTH[8]), 
        .B1(n269), .C0(n3976), .C1(n830), .Y(n1767) );
  OAI221XLTS U2671 ( .A0(n446), .A1(n295), .B0(n2303), .B1(n840), .C0(n1766), 
        .Y(n2471) );
  AOI222XLTS U2672 ( .A0(n4128), .A1(n992), .B0(n4283), .B1(n382), .C0(n3973), 
        .C1(n832), .Y(n1766) );
  OAI221XLTS U2673 ( .A0(n445), .A1(n293), .B0(n2291), .B1(n839), .C0(n1765), 
        .Y(n2472) );
  AOI222XLTS U2674 ( .A0(n4125), .A1(n797), .B0(n4280), .B1(n266), .C0(n3970), 
        .C1(n830), .Y(n1765) );
  OAI221XLTS U2675 ( .A0(n444), .A1(n730), .B0(n837), .B1(n621), .C0(n1545), 
        .Y(n2572) );
  AOI222XLTS U2676 ( .A0(n3823), .A1(n797), .B0(n3831), .B1(n378), .C0(n3818), 
        .C1(n830), .Y(n1545) );
  OAI221XLTS U2677 ( .A0(n453), .A1(n308), .B0(n2350), .B1(n702), .C0(n1652), 
        .Y(n2535) );
  AOI222XLTS U2678 ( .A0(n4302), .A1(n3488), .B0(n4147), .B1(n3460), .C0(n3991), .C1(n3728), .Y(n1652) );
  OAI221XLTS U2679 ( .A0(n203), .A1(n291), .B0(n702), .B1(n154), .C0(n1534), 
        .Y(n2577) );
  AOI222XLTS U2680 ( .A0(n3830), .A1(n3488), .B0(n3824), .B1(n3459), .C0(n3818), .C1(n3733), .Y(n1534) );
  OAI221XLTS U2681 ( .A0(n3265), .A1(n291), .B0(n3295), .B1(n157), .C0(n1539), 
        .Y(n2574) );
  AOI222XLTS U2682 ( .A0(n3817), .A1(n3271), .B0(n3831), .B1(n3230), .C0(n3824), .C1(n572), .Y(n1539) );
  OAI221XLTS U2683 ( .A0(n1537), .A1(n730), .B0(n3365), .B1(n155), .C0(n1538), 
        .Y(n2575) );
  AOI222XLTS U2684 ( .A0(n3830), .A1(n3309), .B0(n3818), .B1(n3319), .C0(n3823), .C1(n3357), .Y(n1538) );
  OAI221XLTS U2685 ( .A0(n3263), .A1(n311), .B0(n2334), .B1(n3295), .C0(n1720), 
        .Y(n2495) );
  AOI222XLTS U2686 ( .A0(n3984), .A1(n3269), .B0(n4297), .B1(n3229), .C0(n4141), .C1(n572), .Y(n1720) );
  OAI221XLTS U2687 ( .A0(n3265), .A1(n293), .B0(n2294), .B1(n3297), .C0(n1715), 
        .Y(n2500) );
  AOI222XLTS U2688 ( .A0(n3969), .A1(n3270), .B0(n4282), .B1(n3230), .C0(n4126), .C1(n572), .Y(n1715) );
  OAI221XLTS U2689 ( .A0(n451), .A1(n299), .B0(n2342), .B1(n3366), .C0(n1699), 
        .Y(n2508) );
  AOI222XLTS U2690 ( .A0(n4299), .A1(n3310), .B0(n3988), .B1(n3317), .C0(n4144), .C1(n3356), .Y(n1699) );
  OAI221XLTS U2691 ( .A0(n451), .A1(n312), .B0(n2336), .B1(n3367), .C0(n1698), 
        .Y(n2509) );
  AOI222XLTS U2692 ( .A0(n4296), .A1(n3311), .B0(n3985), .B1(n3317), .C0(n4141), .C1(n3356), .Y(n1698) );
  OAI221XLTS U2693 ( .A0(n329), .A1(n302), .B0(n2326), .B1(n3367), .C0(n1697), 
        .Y(n2510) );
  AOI222XLTS U2694 ( .A0(n4293), .A1(n3314), .B0(n3982), .B1(n3317), .C0(n4138), .C1(n3356), .Y(n1697) );
  OAI221XLTS U2695 ( .A0(n333), .A1(n314), .B0(n2308), .B1(n3368), .C0(n1695), 
        .Y(n2512) );
  AOI222XLTS U2696 ( .A0(n4287), .A1(n3309), .B0(n3976), .B1(n3318), .C0(n4132), .C1(n3364), .Y(n1695) );
  OAI221XLTS U2697 ( .A0(n451), .A1(n296), .B0(n2304), .B1(n3368), .C0(n1694), 
        .Y(n2513) );
  AOI222XLTS U2698 ( .A0(n4284), .A1(n3309), .B0(n3973), .B1(n3318), .C0(n4129), .C1(n3357), .Y(n1694) );
  OAI221XLTS U2699 ( .A0(n451), .A1(n294), .B0(n2292), .B1(n3367), .C0(n1693), 
        .Y(n2514) );
  AOI222XLTS U2700 ( .A0(n4281), .A1(n3309), .B0(n3970), .B1(n3318), .C0(n4126), .C1(n3357), .Y(n1693) );
  OAI221XLTS U2701 ( .A0(n3263), .A1(n300), .B0(n2341), .B1(n436), .C0(n1721), 
        .Y(n2494) );
  AOI222XLTS U2702 ( .A0(n3987), .A1(n3269), .B0(n4300), .B1(n3229), .C0(n4144), .C1(n572), .Y(n1721) );
  OAI221XLTS U2703 ( .A0(n3264), .A1(n305), .B0(n2319), .B1(n3296), .C0(n1718), 
        .Y(n2497) );
  AOI222XLTS U2704 ( .A0(n3978), .A1(n3270), .B0(n4291), .B1(n3229), .C0(n4135), .C1(n1540), .Y(n1718) );
  OAI221XLTS U2705 ( .A0(n3264), .A1(n315), .B0(n2305), .B1(n436), .C0(n1717), 
        .Y(n2498) );
  AOI222XLTS U2706 ( .A0(n3975), .A1(n3270), .B0(n4288), .B1(n3230), .C0(n4132), .C1(n573), .Y(n1717) );
  OAI221XLTS U2707 ( .A0(n440), .A1(n721), .B0(n2347), .B1(n3433), .C0(n1677), 
        .Y(n2521) );
  OAI221XLTS U2708 ( .A0(n439), .A1(n299), .B0(n2337), .B1(n3432), .C0(n1676), 
        .Y(n2522) );
  AOI222XLTS U2709 ( .A0(n3987), .A1(n3391), .B0(n4300), .B1(n359), .C0(n4143), 
        .C1(n3422), .Y(n1676) );
  OAI221XLTS U2710 ( .A0(n440), .A1(n311), .B0(n2331), .B1(n3433), .C0(n1675), 
        .Y(n2523) );
  AOI222XLTS U2711 ( .A0(n3984), .A1(n3391), .B0(n4297), .B1(n360), .C0(n4140), 
        .C1(n3422), .Y(n1675) );
  OAI221XLTS U2712 ( .A0(n439), .A1(n303), .B0(n2321), .B1(n3433), .C0(n1674), 
        .Y(n2524) );
  AOI222XLTS U2713 ( .A0(n3981), .A1(n3391), .B0(n4294), .B1(n284), .C0(n4137), 
        .C1(n3422), .Y(n1674) );
  OAI221XLTS U2714 ( .A0(n440), .A1(n306), .B0(n2317), .B1(n3434), .C0(n1673), 
        .Y(n2525) );
  AOI222XLTS U2715 ( .A0(n3978), .A1(n3391), .B0(n4291), .B1(n284), .C0(n4134), 
        .C1(n3422), .Y(n1673) );
  OAI221XLTS U2716 ( .A0(n439), .A1(n314), .B0(n2307), .B1(n3434), .C0(n1672), 
        .Y(n2526) );
  AOI222XLTS U2717 ( .A0(n3975), .A1(n3392), .B0(n4288), .B1(n360), .C0(n4131), 
        .C1(n3421), .Y(n1672) );
  OAI221XLTS U2718 ( .A0(n440), .A1(n297), .B0(n2301), .B1(n3434), .C0(n1671), 
        .Y(n2527) );
  AOI222XLTS U2719 ( .A0(n3972), .A1(n3392), .B0(n4285), .B1(n358), .C0(n4128), 
        .C1(n3421), .Y(n1671) );
  OAI221XLTS U2720 ( .A0(n439), .A1(n293), .B0(n2295), .B1(n3433), .C0(n1670), 
        .Y(n2528) );
  AOI222XLTS U2721 ( .A0(n3969), .A1(n3394), .B0(n4282), .B1(n283), .C0(n4125), 
        .C1(n3421), .Y(n1670) );
  OAI221XLTS U2722 ( .A0(n3263), .A1(n309), .B0(n2348), .B1(n436), .C0(n1722), 
        .Y(n2493) );
  AOI222XLTS U2723 ( .A0(n3990), .A1(n3269), .B0(n4303), .B1(n3236), .C0(n4147), .C1(n573), .Y(n1722) );
  OAI221XLTS U2724 ( .A0(n3264), .A1(n302), .B0(n2322), .B1(n435), .C0(n1719), 
        .Y(n2496) );
  AOI222XLTS U2725 ( .A0(n3981), .A1(n3269), .B0(n4294), .B1(n3229), .C0(n4138), .C1(n573), .Y(n1719) );
  OAI221XLTS U2726 ( .A0(n3265), .A1(n295), .B0(n2298), .B1(n436), .C0(n1716), 
        .Y(n2499) );
  AOI222XLTS U2727 ( .A0(n3972), .A1(n3270), .B0(n4285), .B1(n3232), .C0(n4129), .C1(n573), .Y(n1716) );
  OAI221XLTS U2728 ( .A0(n1537), .A1(n308), .B0(n2346), .B1(n3367), .C0(n1700), 
        .Y(n2507) );
  AOI222XLTS U2729 ( .A0(n4302), .A1(n3315), .B0(n3991), .B1(n3317), .C0(n4147), .C1(n3360), .Y(n1700) );
  OAI221XLTS U2730 ( .A0(n337), .A1(n305), .B0(n2314), .B1(n3368), .C0(n1696), 
        .Y(n2511) );
  AOI222XLTS U2731 ( .A0(n4290), .A1(n3312), .B0(n3979), .B1(n3318), .C0(n4135), .C1(n3356), .Y(n1696) );
  OAI221XLTS U2732 ( .A0(n450), .A1(n725), .B0(n2316), .B1(n3565), .C0(n1623), 
        .Y(n2553) );
  AOI222XLTS U2733 ( .A0(n3978), .A1(n3513), .B0(n4291), .B1(n3515), .C0(n4135), .C1(n3553), .Y(n1623) );
  OAI221XLTS U2734 ( .A0(n450), .A1(n308), .B0(n2349), .B1(n3564), .C0(n1627), 
        .Y(n2549) );
  AOI222XLTS U2735 ( .A0(n3990), .A1(n3510), .B0(n4303), .B1(n3514), .C0(n4147), .C1(n3554), .Y(n1627) );
  OAI221XLTS U2736 ( .A0(n448), .A1(n722), .B0(n2339), .B1(n3563), .C0(n1626), 
        .Y(n2550) );
  OAI221XLTS U2737 ( .A0(n450), .A1(n723), .B0(n2335), .B1(n3564), .C0(n1625), 
        .Y(n2551) );
  AOI222XLTS U2738 ( .A0(n3984), .A1(n3513), .B0(n4297), .B1(n3514), .C0(n4141), .C1(n3553), .Y(n1625) );
  OAI221XLTS U2739 ( .A0(n448), .A1(n724), .B0(n2325), .B1(n3564), .C0(n1624), 
        .Y(n2552) );
  OAI221XLTS U2740 ( .A0(n450), .A1(n726), .B0(n2309), .B1(n3565), .C0(n1622), 
        .Y(n2554) );
  AOI222XLTS U2741 ( .A0(n3975), .A1(n3506), .B0(n4288), .B1(n3515), .C0(n4132), .C1(n3552), .Y(n1622) );
  OAI221XLTS U2742 ( .A0(n448), .A1(n296), .B0(n2299), .B1(n3565), .C0(n1621), 
        .Y(n2555) );
  AOI222XLTS U2743 ( .A0(n3972), .A1(n3506), .B0(n4285), .B1(n3515), .C0(n4129), .C1(n3552), .Y(n1621) );
  OAI221XLTS U2744 ( .A0(n448), .A1(n728), .B0(n2293), .B1(n3564), .C0(n1620), 
        .Y(n2556) );
  AOI222XLTS U2745 ( .A0(n3969), .A1(n3506), .B0(n4282), .B1(n3515), .C0(n4126), .C1(n3552), .Y(n1620) );
  AOI22X1TS U2746 ( .A0(n3300), .A1(n4253), .B0(n335), .B1(n4375), .Y(n947) );
  AOI222XLTS U2747 ( .A0(n3348), .A1(n4098), .B0(n3340), .B1(n192), .C0(n3319), 
        .C1(n3942), .Y(n948) );
  AOI22X1TS U2748 ( .A0(n3300), .A1(n4250), .B0(n339), .B1(n4372), .Y(n945) );
  AOI222XLTS U2749 ( .A0(n3348), .A1(n4095), .B0(n3340), .B1(n188), .C0(n3319), 
        .C1(n3939), .Y(n946) );
  AOI22X1TS U2750 ( .A0(n3300), .A1(n4247), .B0(n331), .B1(n4371), .Y(n943) );
  AOI222XLTS U2751 ( .A0(n3348), .A1(n4092), .B0(n3340), .B1(n184), .C0(n3319), 
        .C1(n3936), .Y(n944) );
  AOI22X1TS U2752 ( .A0(n3301), .A1(n4244), .B0(n334), .B1(n4369), .Y(n937) );
  AOI222XLTS U2753 ( .A0(n3349), .A1(n4089), .B0(n3341), .B1(n179), .C0(n3320), 
        .C1(n3933), .Y(n938) );
  AOI22X1TS U2754 ( .A0(n3301), .A1(n4259), .B0(n338), .B1(n4378), .Y(n951) );
  AOI222XLTS U2755 ( .A0(n3349), .A1(n4104), .B0(n3341), .B1(n200), .C0(n3320), 
        .C1(n3948), .Y(n952) );
  AOI22X1TS U2756 ( .A0(n3300), .A1(n4256), .B0(n330), .B1(n4377), .Y(n949) );
  AOI22X1TS U2757 ( .A0(n3384), .A1(n3947), .B0(n3743), .B1(n4378), .Y(n934)
         );
  AOI222XLTS U2758 ( .A0(n3415), .A1(n4104), .B0(n3406), .B1(n201), .C0(n284), 
        .C1(n4260), .Y(n935) );
  AOI22X1TS U2759 ( .A0(n3383), .A1(n3944), .B0(n3743), .B1(n4377), .Y(n932)
         );
  AOI222XLTS U2760 ( .A0(n3414), .A1(n4101), .B0(n3406), .B1(n195), .C0(n283), 
        .C1(n4257), .Y(n933) );
  AOI22X1TS U2761 ( .A0(n3383), .A1(n3941), .B0(n3742), .B1(n4375), .Y(n930)
         );
  AOI222XLTS U2762 ( .A0(n3414), .A1(n4098), .B0(n3405), .B1(n191), .C0(n283), 
        .C1(n4254), .Y(n931) );
  AOI22X1TS U2763 ( .A0(n3383), .A1(n3938), .B0(n3742), .B1(n4372), .Y(n928)
         );
  AOI222XLTS U2764 ( .A0(n3414), .A1(n4095), .B0(n3405), .B1(n187), .C0(n358), 
        .C1(n4251), .Y(n929) );
  AOI22X1TS U2765 ( .A0(n3383), .A1(n3935), .B0(n3742), .B1(n4371), .Y(n926)
         );
  AOI222XLTS U2766 ( .A0(n3414), .A1(n4092), .B0(n3405), .B1(n183), .C0(n359), 
        .C1(n4248), .Y(n927) );
  AOI22X1TS U2767 ( .A0(n3384), .A1(n3932), .B0(n3742), .B1(n4369), .Y(n920)
         );
  AOI222XLTS U2768 ( .A0(n3415), .A1(n4089), .B0(n3406), .B1(n180), .C0(n358), 
        .C1(n4245), .Y(n921) );
  AOI22X1TS U2769 ( .A0(n3240), .A1(n199), .B0(n3222), .B1(n4259), .Y(n968) );
  AOI222XLTS U2770 ( .A0(\requesterAddressbuffer[3][5] ), .A1(n3294), .B0(
        n3283), .B1(n3948), .C0(n3253), .C1(n4379), .Y(n969) );
  AOI22X1TS U2771 ( .A0(n3240), .A1(n195), .B0(n3221), .B1(n4256), .Y(n966) );
  AOI222XLTS U2772 ( .A0(\requesterAddressbuffer[3][4] ), .A1(n3287), .B0(
        n3285), .B1(n3945), .C0(n3253), .C1(n4376), .Y(n967) );
  AOI22X1TS U2773 ( .A0(n3240), .A1(n191), .B0(n3221), .B1(n4253), .Y(n964) );
  AOI222XLTS U2774 ( .A0(\requesterAddressbuffer[3][3] ), .A1(n3286), .B0(
        n3285), .B1(n3942), .C0(n3252), .C1(n4374), .Y(n965) );
  AOI22X1TS U2775 ( .A0(n3239), .A1(n187), .B0(n3221), .B1(n4250), .Y(n962) );
  AOI222XLTS U2776 ( .A0(\requesterAddressbuffer[3][2] ), .A1(n3288), .B0(
        n3279), .B1(n3939), .C0(n3252), .C1(n4373), .Y(n963) );
  AOI22X1TS U2777 ( .A0(n3238), .A1(n183), .B0(n3221), .B1(n4247), .Y(n960) );
  AOI222XLTS U2778 ( .A0(\requesterAddressbuffer[3][1] ), .A1(n3289), .B0(
        n3279), .B1(n3936), .C0(n3252), .C1(n4370), .Y(n961) );
  AOI22X1TS U2779 ( .A0(n3240), .A1(n178), .B0(n3222), .B1(n4244), .Y(n953) );
  AOI222XLTS U2780 ( .A0(\requesterAddressbuffer[3][0] ), .A1(n3290), .B0(
        n3280), .B1(n3933), .C0(n3252), .C1(n4368), .Y(n954) );
  AOI22X1TS U2781 ( .A0(n789), .A1(n4103), .B0(n3790), .B1(n4378), .Y(n1001)
         );
  AOI222XLTS U2782 ( .A0(n820), .A1(n3947), .B0(n812), .B1(n199), .C0(n379), 
        .C1(n4260), .Y(n1002) );
  AOI22X1TS U2783 ( .A0(n788), .A1(n4100), .B0(n3790), .B1(n4377), .Y(n999) );
  AOI222XLTS U2784 ( .A0(n819), .A1(n3944), .B0(n812), .B1(n167), .C0(n266), 
        .C1(n4257), .Y(n1000) );
  AOI22X1TS U2785 ( .A0(n788), .A1(n4097), .B0(n3789), .B1(n4375), .Y(n997) );
  AOI222XLTS U2786 ( .A0(n819), .A1(n3941), .B0(n811), .B1(n190), .C0(n266), 
        .C1(n4254), .Y(n998) );
  AOI22X1TS U2787 ( .A0(n788), .A1(n4094), .B0(n3789), .B1(n4372), .Y(n995) );
  AOI222XLTS U2788 ( .A0(n819), .A1(n3938), .B0(n811), .B1(n186), .C0(n260), 
        .C1(n4251), .Y(n996) );
  AOI22X1TS U2789 ( .A0(n788), .A1(n4091), .B0(n3789), .B1(n4371), .Y(n993) );
  AOI222XLTS U2790 ( .A0(n819), .A1(n3935), .B0(n811), .B1(n182), .C0(n259), 
        .C1(n4248), .Y(n994) );
  AOI22X1TS U2791 ( .A0(n789), .A1(n4088), .B0(n3789), .B1(n4369), .Y(n987) );
  AOI222XLTS U2792 ( .A0(n820), .A1(n3932), .B0(n812), .B1(n179), .C0(n269), 
        .C1(n4245), .Y(n988) );
  AOI222XLTS U2793 ( .A0(\requesterAddressbuffer[6][5] ), .A1(n727), .B0(n3490), .B1(n4259), .C0(n172), .C1(n4379), .Y(n918) );
  AOI22X1TS U2794 ( .A0(n3467), .A1(n194), .B0(n3449), .B1(n4100), .Y(n915) );
  AOI222XLTS U2795 ( .A0(\requesterAddressbuffer[6][4] ), .A1(n717), .B0(n3489), .B1(n4256), .C0(n172), .C1(n4376), .Y(n916) );
  AOI22X1TS U2796 ( .A0(n3466), .A1(n186), .B0(n3449), .B1(n4094), .Y(n911) );
  AOI222XLTS U2797 ( .A0(\requesterAddressbuffer[6][2] ), .A1(n732), .B0(n3489), .B1(n4250), .C0(n202), .C1(n4373), .Y(n912) );
  AOI22X1TS U2798 ( .A0(n4277), .A1(n3308), .B0(n4391), .B1(n387), .Y(n1691)
         );
  AOI22X1TS U2799 ( .A0(n4274), .A1(n3308), .B0(n4388), .B1(n340), .Y(n1689)
         );
  AOI222XLTS U2800 ( .A0(n4118), .A1(n3355), .B0(n3342), .B1(n194), .C0(n3963), 
        .C1(n3333), .Y(n1690) );
  AOI22X1TS U2801 ( .A0(n4271), .A1(n3308), .B0(n4387), .B1(n336), .Y(n1687)
         );
  AOI222XLTS U2802 ( .A0(n4115), .A1(n3355), .B0(n3342), .B1(n190), .C0(n3960), 
        .C1(n3325), .Y(n1688) );
  AOI22X1TS U2803 ( .A0(n4268), .A1(n3308), .B0(n4384), .B1(n388), .Y(n1685)
         );
  AOI222XLTS U2804 ( .A0(n4112), .A1(n3355), .B0(n3342), .B1(n186), .C0(n3957), 
        .C1(n3325), .Y(n1686) );
  AOI22X1TS U2805 ( .A0(n4265), .A1(n3314), .B0(n4382), .B1(n332), .Y(n1683)
         );
  AOI222XLTS U2806 ( .A0(n4109), .A1(n3358), .B0(n3342), .B1(n182), .C0(n3954), 
        .C1(n3325), .Y(n1684) );
  AOI22X1TS U2807 ( .A0(n4262), .A1(n3310), .B0(n4380), .B1(n388), .Y(n1681)
         );
  AOI222XLTS U2808 ( .A0(n4106), .A1(n3360), .B0(n3341), .B1(n177), .C0(n3951), 
        .C1(n3325), .Y(n1682) );
  AOI22X1TS U2809 ( .A0(n4238), .A1(n3312), .B0(n4365), .B1(n388), .Y(n1334)
         );
  AOI22X1TS U2810 ( .A0(n4232), .A1(n3313), .B0(n4361), .B1(n387), .Y(n1330)
         );
  AOI22X1TS U2811 ( .A0(n4229), .A1(n3311), .B0(n4359), .B1(n330), .Y(n1328)
         );
  AOI22X1TS U2812 ( .A0(n4226), .A1(n942), .B0(n4356), .B1(n388), .Y(n1326) );
  AOI22X1TS U2813 ( .A0(n4223), .A1(n3307), .B0(n4355), .B1(n339), .Y(n1324)
         );
  AOI22X1TS U2814 ( .A0(n4220), .A1(n3307), .B0(n4353), .B1(n331), .Y(n1322)
         );
  AOI22X1TS U2815 ( .A0(n4217), .A1(n3307), .B0(n4351), .B1(n334), .Y(n1320)
         );
  AOI22X1TS U2816 ( .A0(n4202), .A1(n3305), .B0(n4341), .B1(n336), .Y(n1310)
         );
  AOI22X1TS U2817 ( .A0(n4187), .A1(n3304), .B0(n4331), .B1(n340), .Y(n1300)
         );
  AOI22X1TS U2818 ( .A0(n4175), .A1(n3306), .B0(n4323), .B1(n334), .Y(n1292)
         );
  AOI22X1TS U2819 ( .A0(n4169), .A1(n3303), .B0(n4319), .B1(n338), .Y(n1288)
         );
  AOI22X1TS U2820 ( .A0(n4163), .A1(n3302), .B0(n4314), .B1(n332), .Y(n1284)
         );
  AOI22X1TS U2821 ( .A0(n4160), .A1(n3302), .B0(n4313), .B1(n335), .Y(n1282)
         );
  AOI22X1TS U2822 ( .A0(n4154), .A1(n3302), .B0(n4309), .B1(n339), .Y(n1278)
         );
  AOI22X1TS U2823 ( .A0(n3929), .A1(n3397), .B0(n4367), .B1(n3748), .Y(n1400)
         );
  AOI22X1TS U2824 ( .A0(n3884), .A1(n3388), .B0(n4337), .B1(n3753), .Y(n1370)
         );
  AOI22X1TS U2825 ( .A0(n3881), .A1(n3388), .B0(n4335), .B1(n3753), .Y(n1368)
         );
  AOI22X1TS U2826 ( .A0(n3869), .A1(n3387), .B0(n4327), .B1(n3746), .Y(n1360)
         );
  AOI22X1TS U2827 ( .A0(n3839), .A1(n3384), .B0(n4307), .B1(n3743), .Y(n1340)
         );
  AOI22X1TS U2828 ( .A0(n4241), .A1(n3316), .B0(n4367), .B1(n387), .Y(n1336)
         );
  AOI22X1TS U2829 ( .A0(n4235), .A1(n3313), .B0(n4362), .B1(n3756), .Y(n1332)
         );
  AOI22X1TS U2830 ( .A0(n4214), .A1(n3307), .B0(n4349), .B1(n338), .Y(n1318)
         );
  AOI22X1TS U2831 ( .A0(n4211), .A1(n3306), .B0(n4347), .B1(n340), .Y(n1316)
         );
  AOI22X1TS U2832 ( .A0(n4208), .A1(n3306), .B0(n4344), .B1(n332), .Y(n1314)
         );
  AOI22X1TS U2833 ( .A0(n4205), .A1(n3306), .B0(n4343), .B1(n335), .Y(n1312)
         );
  AOI22X1TS U2834 ( .A0(n4196), .A1(n3305), .B0(n4337), .B1(n331), .Y(n1306)
         );
  AOI22X1TS U2835 ( .A0(n4184), .A1(n3304), .B0(n4329), .B1(n332), .Y(n1298)
         );
  AOI22X1TS U2836 ( .A0(n4181), .A1(n3304), .B0(n4327), .B1(n335), .Y(n1296)
         );
  AOI22X1TS U2837 ( .A0(n4178), .A1(n3303), .B0(n4325), .B1(n339), .Y(n1294)
         );
  AOI22X1TS U2838 ( .A0(n4172), .A1(n3303), .B0(n4321), .B1(n330), .Y(n1290)
         );
  AOI22X1TS U2839 ( .A0(n4166), .A1(n3303), .B0(n4317), .B1(n336), .Y(n1286)
         );
  AOI22X1TS U2840 ( .A0(n4151), .A1(n3301), .B0(n4307), .B1(n336), .Y(n1276)
         );
  AOI22X1TS U2841 ( .A0(n4148), .A1(n3301), .B0(n4304), .B1(n340), .Y(n1274)
         );
  AOI22X1TS U2842 ( .A0(n3965), .A1(n3395), .B0(n4390), .B1(n3747), .Y(n1667)
         );
  AOI222XLTS U2843 ( .A0(n4121), .A1(n3420), .B0(n3405), .B1(
        readRequesterAddress[5]), .C0(n4278), .C1(n375), .Y(n1668) );
  AOI22X1TS U2844 ( .A0(n3962), .A1(n3396), .B0(n4389), .B1(n3747), .Y(n1665)
         );
  AOI222XLTS U2845 ( .A0(n4118), .A1(n3420), .B0(n3407), .B1(n196), .C0(n4275), 
        .C1(n357), .Y(n1666) );
  AOI22X1TS U2846 ( .A0(n3959), .A1(n3392), .B0(n4386), .B1(n3747), .Y(n1663)
         );
  AOI222XLTS U2847 ( .A0(n4115), .A1(n3420), .B0(n3407), .B1(n192), .C0(n4272), 
        .C1(n360), .Y(n1664) );
  AOI22X1TS U2848 ( .A0(n3956), .A1(n3392), .B0(n4385), .B1(n3747), .Y(n1661)
         );
  AOI222XLTS U2849 ( .A0(n4112), .A1(n3420), .B0(n3407), .B1(n188), .C0(n4269), 
        .C1(n357), .Y(n1662) );
  AOI22X1TS U2850 ( .A0(n3953), .A1(n3393), .B0(n4383), .B1(n3753), .Y(n1659)
         );
  AOI222XLTS U2851 ( .A0(n4109), .A1(n3424), .B0(n3407), .B1(n184), .C0(n4266), 
        .C1(n357), .Y(n1660) );
  AOI22X1TS U2852 ( .A0(n3950), .A1(n3393), .B0(n4381), .B1(n3748), .Y(n1657)
         );
  AOI222XLTS U2853 ( .A0(n4106), .A1(n3424), .B0(n3406), .B1(
        readRequesterAddress[0]), .C0(n4263), .C1(n357), .Y(n1658) );
  AOI22X1TS U2854 ( .A0(n3926), .A1(n3397), .B0(n4365), .B1(n510), .Y(n1398)
         );
  AOI22X1TS U2855 ( .A0(n3923), .A1(n3395), .B0(n4362), .B1(n3751), .Y(n1396)
         );
  AOI22X1TS U2856 ( .A0(n3920), .A1(n3393), .B0(n4361), .B1(n3749), .Y(n1394)
         );
  AOI22X1TS U2857 ( .A0(n3917), .A1(n3396), .B0(n4359), .B1(n3748), .Y(n1392)
         );
  AOI22X1TS U2858 ( .A0(n3914), .A1(n3393), .B0(n4356), .B1(n3749), .Y(n1390)
         );
  AOI22X1TS U2859 ( .A0(n3911), .A1(n3390), .B0(n4355), .B1(n3752), .Y(n1388)
         );
  AOI22X1TS U2860 ( .A0(n3908), .A1(n3390), .B0(n4353), .B1(n3749), .Y(n1386)
         );
  AOI22X1TS U2861 ( .A0(n3905), .A1(n3390), .B0(n4351), .B1(n3752), .Y(n1384)
         );
  AOI22X1TS U2862 ( .A0(n3902), .A1(n3390), .B0(n4349), .B1(n3749), .Y(n1382)
         );
  AOI22X1TS U2863 ( .A0(n3899), .A1(n3389), .B0(n4347), .B1(n3750), .Y(n1380)
         );
  AOI22X1TS U2864 ( .A0(n3896), .A1(n3389), .B0(n4344), .B1(n3755), .Y(n1378)
         );
  AOI22X1TS U2865 ( .A0(n3893), .A1(n3389), .B0(n4343), .B1(n3750), .Y(n1376)
         );
  AOI22X1TS U2866 ( .A0(n3890), .A1(n3388), .B0(n4341), .B1(n3751), .Y(n1374)
         );
  AOI22X1TS U2867 ( .A0(n3887), .A1(n3388), .B0(n4339), .B1(n3750), .Y(n1372)
         );
  AOI22X1TS U2868 ( .A0(n3878), .A1(n3387), .B0(n4332), .B1(n3750), .Y(n1366)
         );
  AOI22X1TS U2869 ( .A0(n3875), .A1(n3387), .B0(n4331), .B1(n3746), .Y(n1364)
         );
  AOI22X1TS U2870 ( .A0(n3872), .A1(n3387), .B0(n4329), .B1(n3746), .Y(n1362)
         );
  AOI22X1TS U2871 ( .A0(n3866), .A1(n3386), .B0(n4325), .B1(n3746), .Y(n1358)
         );
  AOI22X1TS U2872 ( .A0(n3863), .A1(n3389), .B0(n4323), .B1(n3745), .Y(n1356)
         );
  AOI22X1TS U2873 ( .A0(n3860), .A1(n3386), .B0(n4321), .B1(n3745), .Y(n1354)
         );
  AOI22X1TS U2874 ( .A0(n3857), .A1(n3386), .B0(n4319), .B1(n3745), .Y(n1352)
         );
  AOI22X1TS U2875 ( .A0(n3854), .A1(n3386), .B0(n4317), .B1(n3745), .Y(n1350)
         );
  AOI22X1TS U2876 ( .A0(n3851), .A1(n3385), .B0(n4314), .B1(n3744), .Y(n1348)
         );
  AOI22X1TS U2877 ( .A0(n3848), .A1(n3385), .B0(n4313), .B1(n3744), .Y(n1346)
         );
  AOI22X1TS U2878 ( .A0(n3845), .A1(n3385), .B0(n4310), .B1(n3744), .Y(n1344)
         );
  AOI22X1TS U2879 ( .A0(n3842), .A1(n3385), .B0(n4309), .B1(n3744), .Y(n1342)
         );
  AOI22X1TS U2880 ( .A0(n3836), .A1(n3384), .B0(n4304), .B1(n3743), .Y(n1338)
         );
  AOI22X1TS U2881 ( .A0(n4199), .A1(n3305), .B0(n4339), .B1(n334), .Y(n1308)
         );
  AOI22X1TS U2882 ( .A0(n4193), .A1(n3305), .B0(n4335), .B1(n338), .Y(n1304)
         );
  AOI22X1TS U2883 ( .A0(n4190), .A1(n3304), .B0(n4332), .B1(n330), .Y(n1302)
         );
  AOI22X1TS U2884 ( .A0(n4157), .A1(n3302), .B0(n4310), .B1(n331), .Y(n1280)
         );
  AOI22X1TS U2885 ( .A0(n4073), .A1(n802), .B0(n4359), .B1(n3801), .Y(n1136)
         );
  AOI222XLTS U2886 ( .A0(n3917), .A1(n829), .B0(cacheDataOut[27]), .B1(n805), 
        .C0(n4230), .C1(n258), .Y(n1137) );
  AOI22X1TS U2887 ( .A0(n4058), .A1(n799), .B0(n4349), .B1(n3797), .Y(n1126)
         );
  AOI222XLTS U2888 ( .A0(n3902), .A1(n827), .B0(cacheDataOut[22]), .B1(n808), 
        .C0(n4215), .C1(n258), .Y(n1127) );
  AOI22X1TS U2889 ( .A0(n4052), .A1(n794), .B0(n4344), .B1(n3799), .Y(n1122)
         );
  AOI222XLTS U2890 ( .A0(n3896), .A1(n826), .B0(cacheDataOut[20]), .B1(n808), 
        .C0(n4209), .C1(n258), .Y(n1123) );
  AOI22X1TS U2891 ( .A0(n4049), .A1(n794), .B0(n4343), .B1(n500), .Y(n1120) );
  AOI222XLTS U2892 ( .A0(n3893), .A1(n826), .B0(cacheDataOut[19]), .B1(n809), 
        .C0(n4206), .C1(n262), .Y(n1121) );
  AOI22X1TS U2893 ( .A0(n4022), .A1(n791), .B0(n4325), .B1(n3793), .Y(n1102)
         );
  AOI222XLTS U2894 ( .A0(n3866), .A1(n822), .B0(cacheDataOut[10]), .B1(n814), 
        .C0(n4179), .C1(n380), .Y(n1103) );
  AOI22X1TS U2895 ( .A0(n4016), .A1(n791), .B0(n4321), .B1(n3792), .Y(n1098)
         );
  AOI222XLTS U2896 ( .A0(n3860), .A1(n822), .B0(cacheDataOut[8]), .B1(n817), 
        .C0(n4173), .C1(n262), .Y(n1099) );
  AOI22X1TS U2897 ( .A0(n4007), .A1(n790), .B0(n4314), .B1(n3791), .Y(n1092)
         );
  AOI222XLTS U2898 ( .A0(n3851), .A1(n821), .B0(cacheDataOut[5]), .B1(n810), 
        .C0(n4164), .C1(n379), .Y(n1093) );
  AOI22X1TS U2899 ( .A0(n3998), .A1(n790), .B0(n4309), .B1(n3791), .Y(n1086)
         );
  AOI222XLTS U2900 ( .A0(n3842), .A1(n821), .B0(cacheDataOut[2]), .B1(n810), 
        .C0(n4155), .C1(n262), .Y(n1087) );
  AOI22X1TS U2901 ( .A0(n4277), .A1(n3486), .B0(n4390), .B1(n174), .Y(n1642)
         );
  AOI222XLTS U2902 ( .A0(n3965), .A1(n513), .B0(n3478), .B1(n200), .C0(n4122), 
        .C1(n3463), .Y(n1643) );
  AOI22X1TS U2903 ( .A0(n4271), .A1(n3488), .B0(n4386), .B1(n3737), .Y(n1638)
         );
  AOI222XLTS U2904 ( .A0(n3959), .A1(n3730), .B0(n3478), .B1(n166), .C0(n4116), 
        .C1(n3458), .Y(n1639) );
  AOI22X1TS U2905 ( .A0(n4268), .A1(n3493), .B0(n4385), .B1(n172), .Y(n1636)
         );
  AOI222XLTS U2906 ( .A0(n3956), .A1(n3729), .B0(n3478), .B1(n165), .C0(n4113), 
        .C1(n3458), .Y(n1637) );
  AOI22X1TS U2907 ( .A0(n4265), .A1(n3492), .B0(n4383), .B1(n173), .Y(n1634)
         );
  AOI222XLTS U2908 ( .A0(n3953), .A1(n3731), .B0(n907), .B1(n164), .C0(n4110), 
        .C1(n3458), .Y(n1635) );
  AOI22X1TS U2909 ( .A0(n4262), .A1(n3493), .B0(n4381), .B1(n3736), .Y(n1632)
         );
  AOI222XLTS U2910 ( .A0(n3950), .A1(n3731), .B0(n3479), .B1(n177), .C0(n4107), 
        .C1(n3458), .Y(n1633) );
  AOI22X1TS U2911 ( .A0(n4235), .A1(n3487), .B0(n4362), .B1(n3739), .Y(n1461)
         );
  AOI22X1TS U2912 ( .A0(n4217), .A1(n3485), .B0(n4351), .B1(n175), .Y(n1449)
         );
  AOI22X1TS U2913 ( .A0(n4211), .A1(n3485), .B0(n4347), .B1(n3738), .Y(n1445)
         );
  AOI22X1TS U2914 ( .A0(n4208), .A1(n3485), .B0(n4344), .B1(n3737), .Y(n1443)
         );
  AOI22X1TS U2915 ( .A0(n4187), .A1(n3483), .B0(n4331), .B1(n175), .Y(n1429)
         );
  AOI22X1TS U2916 ( .A0(n4184), .A1(n3483), .B0(n4329), .B1(n3739), .Y(n1427)
         );
  AOI22X1TS U2917 ( .A0(n4178), .A1(n3482), .B0(n4325), .B1(n3736), .Y(n1423)
         );
  AOI22X1TS U2918 ( .A0(n4166), .A1(n3481), .B0(n4317), .B1(n175), .Y(n1415)
         );
  AOI22X1TS U2919 ( .A0(n3962), .A1(n3505), .B0(n4389), .B1(n367), .Y(n1614)
         );
  AOI222XLTS U2920 ( .A0(n4119), .A1(n3551), .B0(n195), .B1(n3531), .C0(n4275), 
        .C1(n3523), .Y(n1615) );
  AOI22X1TS U2921 ( .A0(n3950), .A1(n3512), .B0(n4381), .B1(n367), .Y(n1606)
         );
  AOI222XLTS U2922 ( .A0(n4107), .A1(n3550), .B0(n180), .B1(n890), .C0(n4263), 
        .C1(n3524), .Y(n1607) );
  AOI22X1TS U2923 ( .A0(n4121), .A1(n795), .B0(n4390), .B1(n3795), .Y(n1761)
         );
  OAI211X1TS U2924 ( .A0(n2395), .A1(n850), .B0(n1759), .C0(n1760), .Y(n2474)
         );
  INVX2TS U2925 ( .A(n853), .Y(n850) );
  AOI22X1TS U2926 ( .A0(n4118), .A1(n795), .B0(n4389), .B1(n3795), .Y(n1759)
         );
  AOI222XLTS U2927 ( .A0(n3963), .A1(n833), .B0(n813), .B1(n167), .C0(n4275), 
        .C1(n269), .Y(n1760) );
  AOI22X1TS U2928 ( .A0(n4115), .A1(n795), .B0(n4386), .B1(n3795), .Y(n1757)
         );
  AOI222XLTS U2929 ( .A0(n3960), .A1(n830), .B0(n813), .B1(n166), .C0(n4272), 
        .C1(n380), .Y(n1758) );
  AOI22X1TS U2930 ( .A0(n4112), .A1(n795), .B0(n4385), .B1(n3795), .Y(n1755)
         );
  AOI222XLTS U2931 ( .A0(n3957), .A1(n831), .B0(n813), .B1(n165), .C0(n4269), 
        .C1(n379), .Y(n1756) );
  AOI22X1TS U2932 ( .A0(n4109), .A1(n798), .B0(n4383), .B1(n11), .Y(n1753) );
  AOI222XLTS U2933 ( .A0(n3954), .A1(n832), .B0(n813), .B1(n164), .C0(n4266), 
        .C1(n382), .Y(n1754) );
  AOI22X1TS U2934 ( .A0(n4106), .A1(n798), .B0(n4381), .B1(n3796), .Y(n1751)
         );
  AOI222XLTS U2935 ( .A0(n3951), .A1(n834), .B0(n812), .B1(n178), .C0(n4263), 
        .C1(n268), .Y(n1752) );
  AOI22X1TS U2936 ( .A0(n4085), .A1(n801), .B0(n4367), .B1(n3800), .Y(n1144)
         );
  AOI222XLTS U2937 ( .A0(n3929), .A1(n989), .B0(cacheDataOut[31]), .B1(n806), 
        .C0(n4242), .C1(n259), .Y(n1145) );
  AOI22X1TS U2938 ( .A0(n4082), .A1(n798), .B0(n4365), .B1(n500), .Y(n1142) );
  AOI222XLTS U2939 ( .A0(n3926), .A1(n831), .B0(cacheDataOut[30]), .B1(n805), 
        .C0(n4239), .C1(n260), .Y(n1143) );
  AOI22X1TS U2940 ( .A0(n4079), .A1(n799), .B0(n4362), .B1(n3801), .Y(n1140)
         );
  AOI222XLTS U2941 ( .A0(n3923), .A1(n833), .B0(cacheDataOut[29]), .B1(n806), 
        .C0(n4236), .C1(n383), .Y(n1141) );
  AOI22X1TS U2942 ( .A0(n4076), .A1(n800), .B0(n4361), .B1(n3799), .Y(n1138)
         );
  AOI222XLTS U2943 ( .A0(n3920), .A1(n836), .B0(cacheDataOut[28]), .B1(n805), 
        .C0(n4233), .C1(n381), .Y(n1139) );
  AOI22X1TS U2944 ( .A0(n4070), .A1(n802), .B0(n4356), .B1(n3796), .Y(n1134)
         );
  AOI222XLTS U2945 ( .A0(n3914), .A1(n836), .B0(cacheDataOut[26]), .B1(n807), 
        .C0(n4227), .C1(n260), .Y(n1135) );
  AOI22X1TS U2946 ( .A0(n4067), .A1(n799), .B0(n4355), .B1(n3798), .Y(n1132)
         );
  AOI222XLTS U2947 ( .A0(n3911), .A1(n827), .B0(cacheDataOut[25]), .B1(n807), 
        .C0(n4224), .C1(n383), .Y(n1133) );
  AOI22X1TS U2948 ( .A0(n4064), .A1(n800), .B0(n4353), .B1(n3797), .Y(n1130)
         );
  AOI222XLTS U2949 ( .A0(n3908), .A1(n827), .B0(cacheDataOut[24]), .B1(n806), 
        .C0(n4221), .C1(n381), .Y(n1131) );
  AOI22X1TS U2950 ( .A0(n4061), .A1(n801), .B0(n4351), .B1(n3798), .Y(n1128)
         );
  AOI222XLTS U2951 ( .A0(n3905), .A1(n827), .B0(cacheDataOut[23]), .B1(n808), 
        .C0(n4218), .C1(n383), .Y(n1129) );
  AOI22X1TS U2952 ( .A0(n4055), .A1(n794), .B0(n4347), .B1(n3799), .Y(n1124)
         );
  AOI222XLTS U2953 ( .A0(n3899), .A1(n826), .B0(cacheDataOut[21]), .B1(n806), 
        .C0(n4212), .C1(n381), .Y(n1125) );
  AOI22X1TS U2954 ( .A0(n4046), .A1(n793), .B0(n4341), .B1(n3801), .Y(n1118)
         );
  AOI222XLTS U2955 ( .A0(n3890), .A1(n824), .B0(cacheDataOut[18]), .B1(n807), 
        .C0(n4203), .C1(n259), .Y(n1119) );
  AOI22X1TS U2956 ( .A0(n4043), .A1(n793), .B0(n4339), .B1(n3794), .Y(n1116)
         );
  AOI222XLTS U2957 ( .A0(n3887), .A1(n824), .B0(cacheDataOut[17]), .B1(n809), 
        .C0(n4200), .C1(n265), .Y(n1117) );
  AOI22X1TS U2958 ( .A0(n4040), .A1(n793), .B0(n4337), .B1(n3794), .Y(n1114)
         );
  AOI222XLTS U2959 ( .A0(n3884), .A1(n824), .B0(cacheDataOut[16]), .B1(n805), 
        .C0(n4197), .C1(n268), .Y(n1115) );
  AOI22X1TS U2960 ( .A0(n4037), .A1(n793), .B0(n4335), .B1(n3794), .Y(n1112)
         );
  AOI222XLTS U2961 ( .A0(n3881), .A1(n824), .B0(cacheDataOut[15]), .B1(n808), 
        .C0(n4194), .C1(n378), .Y(n1113) );
  AOI22X1TS U2962 ( .A0(n4034), .A1(n792), .B0(n4332), .B1(n3794), .Y(n1110)
         );
  AOI222XLTS U2963 ( .A0(n3878), .A1(n823), .B0(cacheDataOut[14]), .B1(n807), 
        .C0(n4191), .C1(n262), .Y(n1111) );
  AOI22X1TS U2964 ( .A0(n4031), .A1(n792), .B0(n4331), .B1(n3793), .Y(n1108)
         );
  AOI222XLTS U2965 ( .A0(n3875), .A1(n823), .B0(cacheDataOut[13]), .B1(n990), 
        .C0(n4188), .C1(n382), .Y(n1109) );
  AOI22X1TS U2966 ( .A0(n4028), .A1(n792), .B0(n4329), .B1(n3793), .Y(n1106)
         );
  AOI222XLTS U2967 ( .A0(n3872), .A1(n823), .B0(cacheDataOut[12]), .B1(n809), 
        .C0(n4185), .C1(n379), .Y(n1107) );
  AOI22X1TS U2968 ( .A0(n4025), .A1(n792), .B0(n4327), .B1(n3793), .Y(n1104)
         );
  AOI222XLTS U2969 ( .A0(n3869), .A1(n823), .B0(cacheDataOut[11]), .B1(n814), 
        .C0(n4182), .C1(n268), .Y(n1105) );
  AOI22X1TS U2970 ( .A0(n4019), .A1(n794), .B0(n4323), .B1(n3792), .Y(n1100)
         );
  AOI222XLTS U2971 ( .A0(n3863), .A1(n826), .B0(cacheDataOut[9]), .B1(n817), 
        .C0(n4176), .C1(n383), .Y(n1101) );
  AOI22X1TS U2972 ( .A0(n4013), .A1(n791), .B0(n4319), .B1(n3792), .Y(n1096)
         );
  AOI222XLTS U2973 ( .A0(n3857), .A1(n822), .B0(cacheDataOut[7]), .B1(n815), 
        .C0(n4170), .C1(n265), .Y(n1097) );
  AOI22X1TS U2974 ( .A0(n4010), .A1(n791), .B0(n4317), .B1(n3792), .Y(n1094)
         );
  AOI222XLTS U2975 ( .A0(n3854), .A1(n822), .B0(cacheDataOut[6]), .B1(n818), 
        .C0(n4167), .C1(n265), .Y(n1095) );
  AOI22X1TS U2976 ( .A0(n4004), .A1(n790), .B0(n4313), .B1(n3791), .Y(n1090)
         );
  AOI222XLTS U2977 ( .A0(n3848), .A1(n821), .B0(cacheDataOut[4]), .B1(n810), 
        .C0(n4161), .C1(n268), .Y(n1091) );
  AOI22X1TS U2978 ( .A0(n4001), .A1(n790), .B0(n4310), .B1(n3791), .Y(n1088)
         );
  AOI222XLTS U2979 ( .A0(n3845), .A1(n821), .B0(cacheDataOut[3]), .B1(n817), 
        .C0(n4158), .C1(n380), .Y(n1089) );
  AOI22X1TS U2980 ( .A0(n3995), .A1(n789), .B0(n4307), .B1(n3790), .Y(n1084)
         );
  AOI222XLTS U2981 ( .A0(n3839), .A1(n820), .B0(cacheDataOut[1]), .B1(n810), 
        .C0(n4152), .C1(n265), .Y(n1085) );
  AOI22X1TS U2982 ( .A0(n4241), .A1(n3492), .B0(n4367), .B1(n3735), .Y(n1465)
         );
  AOI22X1TS U2983 ( .A0(n4238), .A1(n3487), .B0(n4365), .B1(n3741), .Y(n1463)
         );
  AOI22X1TS U2984 ( .A0(n4232), .A1(n3487), .B0(n4361), .B1(n3738), .Y(n1459)
         );
  AOI22X1TS U2985 ( .A0(n4229), .A1(n3487), .B0(n4359), .B1(n173), .Y(n1457)
         );
  AOI22X1TS U2986 ( .A0(n4226), .A1(n3486), .B0(n4356), .B1(n174), .Y(n1455)
         );
  AOI22X1TS U2987 ( .A0(n4220), .A1(n3486), .B0(n4353), .B1(n3734), .Y(n1451)
         );
  AOI22X1TS U2988 ( .A0(n4214), .A1(n3485), .B0(n4349), .B1(n3735), .Y(n1447)
         );
  AOI22X1TS U2989 ( .A0(n4205), .A1(n3484), .B0(n4343), .B1(n3738), .Y(n1441)
         );
  AOI22X1TS U2990 ( .A0(n4199), .A1(n3484), .B0(n4339), .B1(n3737), .Y(n1437)
         );
  AOI22X1TS U2991 ( .A0(n4196), .A1(n3484), .B0(n4337), .B1(n3735), .Y(n1435)
         );
  AOI22X1TS U2992 ( .A0(n4193), .A1(n3483), .B0(n4335), .B1(n3734), .Y(n1433)
         );
  AOI22X1TS U2993 ( .A0(n4190), .A1(n3483), .B0(n4332), .B1(n173), .Y(n1431)
         );
  AOI22X1TS U2994 ( .A0(n4181), .A1(n3482), .B0(n4327), .B1(n3735), .Y(n1425)
         );
  AOI22X1TS U2995 ( .A0(n4175), .A1(n3482), .B0(n4323), .B1(n3739), .Y(n1421)
         );
  AOI22X1TS U2996 ( .A0(n4172), .A1(n3482), .B0(n4321), .B1(n3738), .Y(n1419)
         );
  AOI22X1TS U2997 ( .A0(n4169), .A1(n3481), .B0(n4319), .B1(n173), .Y(n1417)
         );
  AOI22X1TS U2998 ( .A0(n4163), .A1(n3481), .B0(n4314), .B1(n3734), .Y(n1413)
         );
  AOI22X1TS U2999 ( .A0(n4157), .A1(n3480), .B0(n4310), .B1(n174), .Y(n1409)
         );
  AOI22X1TS U3000 ( .A0(n4154), .A1(n3480), .B0(n4309), .B1(n3737), .Y(n1407)
         );
  AOI22X1TS U3001 ( .A0(n3965), .A1(n3505), .B0(n4390), .B1(n366), .Y(n1616)
         );
  AOI22X1TS U3002 ( .A0(n3959), .A1(n3505), .B0(n4386), .B1(n3718), .Y(n1612)
         );
  AOI222XLTS U3003 ( .A0(n4116), .A1(n3551), .B0(n191), .B1(n3531), .C0(n4272), 
        .C1(n3528), .Y(n1613) );
  AOI22X1TS U3004 ( .A0(n3956), .A1(n3505), .B0(n4385), .B1(n368), .Y(n1610)
         );
  AOI222XLTS U3005 ( .A0(n4113), .A1(n3551), .B0(n187), .B1(n3531), .C0(n4269), 
        .C1(n891), .Y(n1611) );
  AOI22X1TS U3006 ( .A0(n3953), .A1(n3512), .B0(n4383), .B1(n366), .Y(n1608)
         );
  AOI222XLTS U3007 ( .A0(n4110), .A1(n3550), .B0(n184), .B1(n890), .C0(n4266), 
        .C1(n3524), .Y(n1609) );
  AOI22X1TS U3008 ( .A0(n3929), .A1(n3510), .B0(n4366), .B1(n366), .Y(n1529)
         );
  AOI22X1TS U3009 ( .A0(n3926), .A1(n3511), .B0(n4364), .B1(n365), .Y(n1527)
         );
  AOI22X1TS U3010 ( .A0(n3923), .A1(n3513), .B0(n4363), .B1(n362), .Y(n1525)
         );
  AOI22X1TS U3011 ( .A0(n3920), .A1(n3509), .B0(n4360), .B1(n371), .Y(n1523)
         );
  AOI22X1TS U3012 ( .A0(n3917), .A1(n3511), .B0(n4358), .B1(n368), .Y(n1521)
         );
  AOI22X1TS U3013 ( .A0(n3914), .A1(n3509), .B0(n4357), .B1(n367), .Y(n1519)
         );
  AOI22X1TS U3014 ( .A0(n3911), .A1(n3504), .B0(n4354), .B1(n364), .Y(n1517)
         );
  AOI22X1TS U3015 ( .A0(n3908), .A1(n3504), .B0(n4352), .B1(n373), .Y(n1515)
         );
  AOI22X1TS U3016 ( .A0(n3905), .A1(n3504), .B0(n4350), .B1(n363), .Y(n1513)
         );
  AOI22X1TS U3017 ( .A0(n3902), .A1(n3504), .B0(n4348), .B1(n372), .Y(n1511)
         );
  AOI22X1TS U3018 ( .A0(n3899), .A1(n3503), .B0(n4346), .B1(n362), .Y(n1509)
         );
  AOI22X1TS U3019 ( .A0(n3896), .A1(n3503), .B0(n4345), .B1(n371), .Y(n1507)
         );
  AOI22X1TS U3020 ( .A0(n3893), .A1(n3503), .B0(n4342), .B1(n365), .Y(n1505)
         );
  AOI22X1TS U3021 ( .A0(n3890), .A1(n3502), .B0(n4340), .B1(n370), .Y(n1503)
         );
  AOI22X1TS U3022 ( .A0(n3887), .A1(n3502), .B0(n4338), .B1(n364), .Y(n1501)
         );
  AOI22X1TS U3023 ( .A0(n3884), .A1(n3502), .B0(n4336), .B1(n373), .Y(n1499)
         );
  AOI22X1TS U3024 ( .A0(n3881), .A1(n3502), .B0(n4334), .B1(n363), .Y(n1497)
         );
  AOI22X1TS U3025 ( .A0(n3878), .A1(n3501), .B0(n4333), .B1(n372), .Y(n1495)
         );
  AOI22X1TS U3026 ( .A0(n3875), .A1(n3501), .B0(n4330), .B1(n362), .Y(n1493)
         );
  AOI22X1TS U3027 ( .A0(n3872), .A1(n3501), .B0(n4328), .B1(n371), .Y(n1491)
         );
  AOI22X1TS U3028 ( .A0(n3869), .A1(n3501), .B0(n4326), .B1(n365), .Y(n1489)
         );
  AOI22X1TS U3029 ( .A0(n3866), .A1(n3500), .B0(n4324), .B1(n370), .Y(n1487)
         );
  AOI22X1TS U3030 ( .A0(n3863), .A1(n3500), .B0(n4322), .B1(n364), .Y(n1485)
         );
  AOI22X1TS U3031 ( .A0(n3860), .A1(n3500), .B0(n4320), .B1(n373), .Y(n1483)
         );
  AOI22X1TS U3032 ( .A0(n3857), .A1(n3500), .B0(n4318), .B1(n363), .Y(n1481)
         );
  AOI22X1TS U3033 ( .A0(n3854), .A1(n3499), .B0(n4316), .B1(n372), .Y(n1479)
         );
  AOI22X1TS U3034 ( .A0(n3851), .A1(n3499), .B0(n4315), .B1(n362), .Y(n1477)
         );
  AOI22X1TS U3035 ( .A0(n3848), .A1(n3499), .B0(n4312), .B1(n371), .Y(n1475)
         );
  AOI22X1TS U3036 ( .A0(n3845), .A1(n3499), .B0(n4311), .B1(n365), .Y(n1473)
         );
  AOI22X1TS U3037 ( .A0(n3842), .A1(n3498), .B0(n4308), .B1(n370), .Y(n1471)
         );
  AOI22X1TS U3038 ( .A0(n3839), .A1(n3498), .B0(n4306), .B1(n363), .Y(n1469)
         );
  AOI22X1TS U3039 ( .A0(n3836), .A1(n3498), .B0(n4305), .B1(n372), .Y(n1467)
         );
  AOI22X1TS U3040 ( .A0(n3992), .A1(n789), .B0(n4304), .B1(n3790), .Y(n1082)
         );
  AOI222XLTS U3041 ( .A0(n3836), .A1(n820), .B0(cacheDataOut[0]), .B1(n809), 
        .C0(n4149), .C1(n382), .Y(n1083) );
  AOI22X1TS U3042 ( .A0(n4274), .A1(n3488), .B0(n4389), .B1(n3734), .Y(n1640)
         );
  AOI222XLTS U3043 ( .A0(n3962), .A1(n513), .B0(n907), .B1(n194), .C0(n4119), 
        .C1(n3465), .Y(n1641) );
  AOI22X1TS U3044 ( .A0(n4223), .A1(n3486), .B0(n4355), .B1(n3740), .Y(n1453)
         );
  AOI22X1TS U3045 ( .A0(n4202), .A1(n3484), .B0(n4341), .B1(n3736), .Y(n1439)
         );
  AOI22X1TS U3046 ( .A0(n4160), .A1(n3481), .B0(n4313), .B1(n3736), .Y(n1411)
         );
  AOI22X1TS U3047 ( .A0(n974), .A1(n164), .B0(n855), .B1(n4091), .Y(n976) );
  AOI222XLTS U3048 ( .A0(\requesterAddressbuffer[2][1] ), .A1(n432), .B0(n3198), .B1(n4248), .C0(n3774), .C1(n4370), .Y(n977) );
  AOI22X1TS U3049 ( .A0(n1653), .A1(readRequesterAddress[0]), .B0(n856), .B1(
        n4088), .Y(n971) );
  AOI222XLTS U3050 ( .A0(\requesterAddressbuffer[2][0] ), .A1(n433), .B0(n3200), .B1(n4245), .C0(n3774), .C1(requesterAddressIn_NORTH[0]), .Y(n972) );
  AOI22X1TS U3051 ( .A0(n1546), .A1(n166), .B0(n855), .B1(n4097), .Y(n980) );
  AOI222XLTS U3052 ( .A0(\requesterAddressbuffer[2][3] ), .A1(n273), .B0(n3203), .B1(n4254), .C0(n3774), .C1(n4374), .Y(n981) );
  AOI22X1TS U3053 ( .A0(n1653), .A1(n165), .B0(n855), .B1(n4094), .Y(n978) );
  AOI222XLTS U3054 ( .A0(\requesterAddressbuffer[2][2] ), .A1(n355), .B0(n3201), .B1(n4251), .C0(n3774), .C1(n4373), .Y(n979) );
  AOI22X1TS U3055 ( .A0(n1585), .A1(n167), .B0(n855), .B1(n4100), .Y(n982) );
  AOI222XLTS U3056 ( .A0(\requesterAddressbuffer[2][4] ), .A1(n350), .B0(n3199), .B1(n4257), .C0(n3775), .C1(n4376), .Y(n983) );
  AOI22X1TS U3057 ( .A0(n1544), .A1(readRequesterAddress[5]), .B0(n856), .B1(
        n4103), .Y(n984) );
  AOI222XLTS U3058 ( .A0(\requesterAddressbuffer[2][5] ), .A1(n352), .B0(n3197), .B1(n4260), .C0(n3775), .C1(n4379), .Y(n985) );
  AOI22X1TS U3059 ( .A0(n767), .A1(n200), .B0(n752), .B1(n4259), .Y(n1016) );
  AOI22X1TS U3060 ( .A0(n766), .A1(n166), .B0(n748), .B1(n4253), .Y(n1012) );
  AOI222XLTS U3061 ( .A0(\requesterAddressbuffer[0][3] ), .A1(n385), .B0(n781), 
        .B1(n3942), .C0(n245), .C1(requesterAddressIn_NORTH[3]), .Y(n1013) );
  AOI22X1TS U3062 ( .A0(n768), .A1(n167), .B0(n748), .B1(n4256), .Y(n1014) );
  AOI222XLTS U3063 ( .A0(\requesterAddressbuffer[0][4] ), .A1(n3802), .B0(n781), .B1(n3945), .C0(n246), .C1(requesterAddressIn_NORTH[4]), .Y(n1015) );
  AOI22X1TS U3064 ( .A0(n768), .A1(readRequesterAddress[2]), .B0(n749), .B1(
        n4250), .Y(n1010) );
  AOI222XLTS U3065 ( .A0(\requesterAddressbuffer[0][2] ), .A1(n326), .B0(n782), 
        .B1(n3939), .C0(n246), .C1(n4373), .Y(n1011) );
  AOI22X1TS U3066 ( .A0(n1006), .A1(readRequesterAddress[1]), .B0(n750), .B1(
        n4247), .Y(n1008) );
  AOI222XLTS U3067 ( .A0(\requesterAddressbuffer[0][1] ), .A1(n286), .B0(n782), 
        .B1(n3936), .C0(n245), .C1(requesterAddressIn_NORTH[1]), .Y(n1009) );
  AOI22X1TS U3068 ( .A0(n765), .A1(n180), .B0(n752), .B1(n4244), .Y(n1003) );
  AOI222XLTS U3069 ( .A0(\requesterAddressbuffer[0][0] ), .A1(n238), .B0(n786), 
        .B1(n3933), .C0(n343), .C1(n4368), .Y(n1004) );
  AOI22X1TS U3070 ( .A0(n3466), .A1(n190), .B0(n3449), .B1(n4097), .Y(n913) );
  AOI222XLTS U3071 ( .A0(\requesterAddressbuffer[6][3] ), .A1(n729), .B0(n3489), .B1(n4253), .C0(n202), .C1(n4374), .Y(n914) );
  AOI22X1TS U3072 ( .A0(n3466), .A1(n182), .B0(n3449), .B1(n4091), .Y(n909) );
  AOI222XLTS U3073 ( .A0(\requesterAddressbuffer[6][1] ), .A1(n729), .B0(n3489), .B1(n4247), .C0(n202), .C1(n4370), .Y(n910) );
  AOI222XLTS U3074 ( .A0(\requesterAddressbuffer[6][0] ), .A1(n729), .B0(n3495), .B1(n4244), .C0(n202), .C1(n4368), .Y(n905) );
  AOI22X1TS U3075 ( .A0(n767), .A1(n199), .B0(n4277), .B1(n743), .Y(n1785) );
  AOI222XLTS U3076 ( .A0(n323), .A1(n36), .B0(n3966), .B1(n772), .C0(n4391), 
        .C1(n391), .Y(n1786) );
  AOI22X1TS U3077 ( .A0(n756), .A1(n190), .B0(n4271), .B1(n743), .Y(n1781) );
  AOI222XLTS U3078 ( .A0(n328), .A1(n37), .B0(n3960), .B1(n780), .C0(n4387), 
        .C1(n246), .Y(n1782) );
  AOI22X1TS U3079 ( .A0(n756), .A1(n188), .B0(n4268), .B1(n743), .Y(n1779) );
  AOI222XLTS U3080 ( .A0(n322), .A1(n38), .B0(n3957), .B1(n780), .C0(
        destinationAddressIn_NORTH[2]), .C1(n271), .Y(n1780) );
  AOI22X1TS U3081 ( .A0(n1006), .A1(n184), .B0(n4265), .B1(n742), .Y(n1777) );
  AOI222XLTS U3082 ( .A0(n385), .A1(n39), .B0(n3954), .B1(n779), .C0(
        destinationAddressIn_NORTH[1]), .C1(n346), .Y(n1778) );
  AOI22X1TS U3083 ( .A0(n467), .A1(n762), .B0(n4241), .B1(n742), .Y(n1080) );
  AOI222XLTS U3084 ( .A0(n323), .A1(n40), .B0(n3930), .B1(n779), .C0(
        dataIn_NORTH[31]), .C1(n391), .Y(n1081) );
  AOI22X1TS U3085 ( .A0(n469), .A1(n766), .B0(n4238), .B1(n742), .Y(n1078) );
  AOI222XLTS U3086 ( .A0(n288), .A1(n41), .B0(n3927), .B1(n779), .C0(
        dataIn_NORTH[30]), .C1(n342), .Y(n1079) );
  AOI22X1TS U3087 ( .A0(n471), .A1(n766), .B0(n4235), .B1(n741), .Y(n1076) );
  AOI222XLTS U3088 ( .A0(n323), .A1(n42), .B0(n3924), .B1(n777), .C0(n4363), 
        .C1(n344), .Y(n1077) );
  AOI22X1TS U3089 ( .A0(n477), .A1(n759), .B0(n4226), .B1(n741), .Y(n1070) );
  AOI222XLTS U3090 ( .A0(n326), .A1(n43), .B0(n3915), .B1(n777), .C0(n4357), 
        .C1(n343), .Y(n1071) );
  AOI22X1TS U3091 ( .A0(n479), .A1(n763), .B0(n4223), .B1(n740), .Y(n1068) );
  AOI222XLTS U3092 ( .A0(n327), .A1(n44), .B0(n3912), .B1(n776), .C0(
        dataIn_NORTH[25]), .C1(n344), .Y(n1069) );
  AOI22X1TS U3093 ( .A0(n481), .A1(n769), .B0(n4220), .B1(n740), .Y(n1066) );
  AOI222XLTS U3094 ( .A0(n287), .A1(n45), .B0(n3909), .B1(n776), .C0(
        dataIn_NORTH[24]), .C1(n346), .Y(n1067) );
  AOI22X1TS U3095 ( .A0(n485), .A1(n766), .B0(n4214), .B1(n740), .Y(n1062) );
  AOI222XLTS U3096 ( .A0(n327), .A1(n46), .B0(n3903), .B1(n776), .C0(
        dataIn_NORTH[22]), .C1(n246), .Y(n1063) );
  AOI22X1TS U3097 ( .A0(n487), .A1(n757), .B0(n4211), .B1(n739), .Y(n1060) );
  AOI222XLTS U3098 ( .A0(n286), .A1(n47), .B0(n3900), .B1(n786), .C0(
        dataIn_NORTH[21]), .C1(n391), .Y(n1061) );
  AOI22X1TS U3099 ( .A0(n491), .A1(n757), .B0(n4205), .B1(n739), .Y(n1056) );
  AOI222XLTS U3100 ( .A0(n288), .A1(n48), .B0(n3894), .B1(n783), .C0(
        dataIn_NORTH[19]), .C1(n344), .Y(n1057) );
  AOI22X1TS U3101 ( .A0(n493), .A1(n758), .B0(n4202), .B1(n738), .Y(n1054) );
  AOI222XLTS U3102 ( .A0(n287), .A1(n49), .B0(n3891), .B1(n783), .C0(
        dataIn_NORTH[18]), .C1(n346), .Y(n1055) );
  AOI22X1TS U3103 ( .A0(n495), .A1(n757), .B0(n4199), .B1(n738), .Y(n1052) );
  AOI222XLTS U3104 ( .A0(n324), .A1(n50), .B0(n3888), .B1(n783), .C0(
        dataIn_NORTH[17]), .C1(n347), .Y(n1053) );
  AOI22X1TS U3105 ( .A0(n503), .A1(n758), .B0(n4196), .B1(n738), .Y(n1050) );
  AOI222XLTS U3106 ( .A0(n326), .A1(n51), .B0(n3885), .B1(n785), .C0(
        dataIn_NORTH[16]), .C1(n271), .Y(n1051) );
  AOI22X1TS U3107 ( .A0(n507), .A1(n759), .B0(n4193), .B1(n738), .Y(n1048) );
  AOI222XLTS U3108 ( .A0(n499), .A1(n52), .B0(n3882), .B1(n785), .C0(
        dataIn_NORTH[15]), .C1(n343), .Y(n1049) );
  AOI22X1TS U3109 ( .A0(n509), .A1(n758), .B0(n4190), .B1(n737), .Y(n1046) );
  AOI222XLTS U3110 ( .A0(n324), .A1(n53), .B0(n3879), .B1(n775), .C0(n4333), 
        .C1(n348), .Y(n1047) );
  AOI22X1TS U3111 ( .A0(n512), .A1(n758), .B0(n4187), .B1(n737), .Y(n1044) );
  AOI222XLTS U3112 ( .A0(n288), .A1(n54), .B0(n3876), .B1(n775), .C0(
        dataIn_NORTH[13]), .C1(n391), .Y(n1045) );
  AOI22X1TS U3113 ( .A0(n515), .A1(n759), .B0(n4184), .B1(n737), .Y(n1042) );
  AOI222XLTS U3114 ( .A0(n326), .A1(n55), .B0(n3873), .B1(n775), .C0(
        dataIn_NORTH[12]), .C1(n245), .Y(n1043) );
  AOI22X1TS U3115 ( .A0(n536), .A1(n759), .B0(n4181), .B1(n737), .Y(n1040) );
  AOI222XLTS U3116 ( .A0(n385), .A1(n56), .B0(n3870), .B1(n775), .C0(
        dataIn_NORTH[11]), .C1(n271), .Y(n1041) );
  AOI22X1TS U3117 ( .A0(n541), .A1(n762), .B0(n4178), .B1(n736), .Y(n1038) );
  AOI222XLTS U3118 ( .A0(n287), .A1(n57), .B0(n3867), .B1(n774), .C0(
        dataIn_NORTH[10]), .C1(n346), .Y(n1039) );
  AOI22X1TS U3119 ( .A0(n546), .A1(n760), .B0(n4172), .B1(n736), .Y(n1034) );
  AOI222XLTS U3120 ( .A0(n327), .A1(n58), .B0(n3861), .B1(n774), .C0(
        dataIn_NORTH[8]), .C1(n392), .Y(n1035) );
  AOI22X1TS U3121 ( .A0(n551), .A1(n760), .B0(n4169), .B1(n736), .Y(n1032) );
  AOI222XLTS U3122 ( .A0(n287), .A1(n59), .B0(n3858), .B1(n774), .C0(
        dataIn_NORTH[7]), .C1(n342), .Y(n1033) );
  AOI22X1TS U3123 ( .A0(n555), .A1(n761), .B0(n4166), .B1(n736), .Y(n1030) );
  AOI222XLTS U3124 ( .A0(n324), .A1(n60), .B0(n3855), .B1(n783), .C0(
        dataIn_NORTH[6]), .C1(n347), .Y(n1031) );
  AOI22X1TS U3125 ( .A0(n560), .A1(n761), .B0(n4160), .B1(n735), .Y(n1026) );
  AOI222XLTS U3126 ( .A0(n286), .A1(n61), .B0(n3849), .B1(n773), .C0(
        dataIn_NORTH[4]), .C1(n343), .Y(n1027) );
  AOI22X1TS U3127 ( .A0(n562), .A1(n762), .B0(n4157), .B1(n735), .Y(n1024) );
  AOI222XLTS U3128 ( .A0(n288), .A1(n62), .B0(n3846), .B1(n773), .C0(n4311), 
        .C1(n348), .Y(n1025) );
  AOI22X1TS U3129 ( .A0(n3238), .A1(n200), .B0(n4277), .B1(n3233), .Y(n1713)
         );
  AOI222XLTS U3130 ( .A0(n3287), .A1(n63), .B0(n3966), .B1(n3271), .C0(n4391), 
        .C1(n3262), .Y(n1714) );
  AOI22X1TS U3131 ( .A0(n3238), .A1(n194), .B0(n4274), .B1(n3234), .Y(n1711)
         );
  AOI222XLTS U3132 ( .A0(n3286), .A1(n64), .B0(n3963), .B1(n3285), .C0(n4388), 
        .C1(n3262), .Y(n1712) );
  AOI22X1TS U3133 ( .A0(n3238), .A1(readRequesterAddress[3]), .B0(n4271), .B1(
        n3235), .Y(n1709) );
  AOI222XLTS U3134 ( .A0(n3288), .A1(n65), .B0(n3960), .B1(n3285), .C0(n4387), 
        .C1(n3262), .Y(n1710) );
  AOI22X1TS U3135 ( .A0(n3239), .A1(n182), .B0(n4265), .B1(n3231), .Y(n1705)
         );
  AOI222XLTS U3136 ( .A0(n3290), .A1(n66), .B0(n3954), .B1(n3282), .C0(n4382), 
        .C1(n3261), .Y(n1706) );
  AOI22X1TS U3137 ( .A0(n3239), .A1(n177), .B0(n4262), .B1(n3231), .Y(n1703)
         );
  AOI222XLTS U3138 ( .A0(n3293), .A1(n67), .B0(n3951), .B1(n3282), .C0(
        destinationAddressIn_NORTH[0]), .C1(n3261), .Y(n1704) );
  AOI22X1TS U3139 ( .A0(n468), .A1(n3244), .B0(n4241), .B1(n3234), .Y(n1272)
         );
  AOI222XLTS U3140 ( .A0(n3292), .A1(n68), .B0(n3930), .B1(n956), .C0(n4366), 
        .C1(n3261), .Y(n1273) );
  AOI22X1TS U3141 ( .A0(n470), .A1(n3244), .B0(n4238), .B1(n3235), .Y(n1270)
         );
  AOI222XLTS U3142 ( .A0(n3291), .A1(n69), .B0(n3927), .B1(n3281), .C0(n4364), 
        .C1(n3261), .Y(n1271) );
  AOI22X1TS U3143 ( .A0(n472), .A1(n3244), .B0(n4235), .B1(n3231), .Y(n1268)
         );
  AOI222XLTS U3144 ( .A0(n3293), .A1(n70), .B0(n3924), .B1(n3278), .C0(n4363), 
        .C1(n3260), .Y(n1269) );
  AOI22X1TS U3145 ( .A0(n473), .A1(n3246), .B0(n4232), .B1(n3231), .Y(n1266)
         );
  AOI222XLTS U3146 ( .A0(n280), .A1(n71), .B0(n3921), .B1(n3278), .C0(
        dataIn_NORTH[28]), .C1(n3260), .Y(n1267) );
  AOI22X1TS U3147 ( .A0(n475), .A1(n3244), .B0(n4229), .B1(n3232), .Y(n1264)
         );
  AOI222XLTS U3148 ( .A0(n281), .A1(n72), .B0(n3918), .B1(n3278), .C0(
        dataIn_NORTH[27]), .C1(n3260), .Y(n1265) );
  AOI22X1TS U3149 ( .A0(n478), .A1(n3245), .B0(n4226), .B1(n3233), .Y(n1262)
         );
  AOI222XLTS U3150 ( .A0(n3294), .A1(n73), .B0(n3915), .B1(n3278), .C0(n4357), 
        .C1(n3260), .Y(n1263) );
  AOI22X1TS U3151 ( .A0(n482), .A1(n3248), .B0(n4220), .B1(n3228), .Y(n1258)
         );
  AOI222XLTS U3152 ( .A0(n3290), .A1(n74), .B0(n3909), .B1(n3277), .C0(n4352), 
        .C1(n3259), .Y(n1259) );
  AOI22X1TS U3153 ( .A0(n486), .A1(n3248), .B0(n4214), .B1(n3228), .Y(n1254)
         );
  AOI222XLTS U3154 ( .A0(n3293), .A1(n75), .B0(n3903), .B1(n3277), .C0(n4348), 
        .C1(n3259), .Y(n1255) );
  AOI22X1TS U3155 ( .A0(n488), .A1(n3247), .B0(n4211), .B1(n3227), .Y(n1252)
         );
  AOI222XLTS U3156 ( .A0(n3287), .A1(n76), .B0(n3900), .B1(n3276), .C0(n4346), 
        .C1(n3258), .Y(n1253) );
  AOI22X1TS U3157 ( .A0(n492), .A1(n3245), .B0(n4205), .B1(n3227), .Y(n1248)
         );
  AOI222XLTS U3158 ( .A0(n3286), .A1(n77), .B0(n3894), .B1(n3276), .C0(n4342), 
        .C1(n3258), .Y(n1249) );
  AOI22X1TS U3159 ( .A0(n501), .A1(n3246), .B0(n4199), .B1(n3226), .Y(n1244)
         );
  AOI222XLTS U3160 ( .A0(n3294), .A1(n78), .B0(n3888), .B1(n3275), .C0(n4338), 
        .C1(n3257), .Y(n1245) );
  AOI22X1TS U3161 ( .A0(n505), .A1(n3246), .B0(n4196), .B1(n3226), .Y(n1242)
         );
  AOI222XLTS U3162 ( .A0(n3287), .A1(n79), .B0(n3885), .B1(n3275), .C0(n4336), 
        .C1(n3257), .Y(n1243) );
  AOI22X1TS U3163 ( .A0(n511), .A1(n3249), .B0(n4190), .B1(n3225), .Y(n1238)
         );
  AOI222XLTS U3164 ( .A0(n3286), .A1(n80), .B0(n3879), .B1(n3274), .C0(n4333), 
        .C1(n3257), .Y(n1239) );
  AOI22X1TS U3165 ( .A0(n516), .A1(n3250), .B0(n4184), .B1(n3225), .Y(n1234)
         );
  AOI222XLTS U3166 ( .A0(n281), .A1(n81), .B0(n3873), .B1(n3274), .C0(n4328), 
        .C1(n3256), .Y(n1235) );
  AOI22X1TS U3167 ( .A0(n537), .A1(n3243), .B0(n4181), .B1(n3225), .Y(n1232)
         );
  AOI222XLTS U3168 ( .A0(n280), .A1(n82), .B0(n3870), .B1(n3274), .C0(n4326), 
        .C1(n3256), .Y(n1233) );
  AOI22X1TS U3169 ( .A0(n543), .A1(n3243), .B0(n4178), .B1(n3224), .Y(n1230)
         );
  AOI222XLTS U3170 ( .A0(n281), .A1(n83), .B0(n3867), .B1(n3273), .C0(n4324), 
        .C1(n3256), .Y(n1231) );
  AOI22X1TS U3171 ( .A0(n544), .A1(n3243), .B0(n4175), .B1(n3227), .Y(n1228)
         );
  AOI222XLTS U3172 ( .A0(n3289), .A1(n84), .B0(n3864), .B1(n3273), .C0(
        dataIn_NORTH[9]), .C1(n3255), .Y(n1229) );
  AOI22X1TS U3173 ( .A0(n548), .A1(n3243), .B0(n4172), .B1(n3224), .Y(n1226)
         );
  AOI222XLTS U3174 ( .A0(n3290), .A1(n85), .B0(n3861), .B1(n3273), .C0(n4320), 
        .C1(n3255), .Y(n1227) );
  AOI22X1TS U3175 ( .A0(n556), .A1(n3242), .B0(n4166), .B1(n3224), .Y(n1222)
         );
  AOI222XLTS U3176 ( .A0(n3293), .A1(n86), .B0(n3855), .B1(n3276), .C0(n4316), 
        .C1(n3255), .Y(n1223) );
  AOI22X1TS U3177 ( .A0(n563), .A1(n3241), .B0(n4157), .B1(n3223), .Y(n1216)
         );
  AOI222XLTS U3178 ( .A0(n3291), .A1(n87), .B0(n3846), .B1(n3272), .C0(n4311), 
        .C1(n3254), .Y(n1217) );
  AOI22X1TS U3179 ( .A0(n566), .A1(n3241), .B0(n4151), .B1(n3222), .Y(n1212)
         );
  AOI222XLTS U3180 ( .A0(n3291), .A1(n88), .B0(n3840), .B1(n3271), .C0(
        dataIn_NORTH[1]), .C1(n3253), .Y(n1213) );
  AOI22X1TS U3181 ( .A0(n568), .A1(n3241), .B0(n4148), .B1(n3222), .Y(n1210)
         );
  AOI222XLTS U3182 ( .A0(n280), .A1(n89), .B0(n3837), .B1(n3271), .C0(n4305), 
        .C1(n3253), .Y(n1211) );
  AOI22X1TS U3183 ( .A0(n756), .A1(readRequesterAddress[4]), .B0(n4274), .B1(
        n743), .Y(n1783) );
  AOI222XLTS U3184 ( .A0(n327), .A1(n90), .B0(n3963), .B1(n780), .C0(
        destinationAddressIn_NORTH[4]), .C1(n392), .Y(n1784) );
  AOI22X1TS U3185 ( .A0(n756), .A1(n178), .B0(n4262), .B1(n742), .Y(n1775) );
  AOI222XLTS U3186 ( .A0(n323), .A1(n91), .B0(n3951), .B1(n779), .C0(n4380), 
        .C1(n347), .Y(n1776) );
  AOI22X1TS U3187 ( .A0(n3239), .A1(n186), .B0(n4268), .B1(n3230), .Y(n1707)
         );
  AOI222XLTS U3188 ( .A0(n3289), .A1(n92), .B0(n3957), .B1(n3283), .C0(n4384), 
        .C1(n3262), .Y(n1708) );
  AOI22X1TS U3189 ( .A0(n480), .A1(n3247), .B0(n4223), .B1(n3228), .Y(n1260)
         );
  AOI222XLTS U3190 ( .A0(n3292), .A1(n93), .B0(n3912), .B1(n3277), .C0(n4354), 
        .C1(n3259), .Y(n1261) );
  AOI22X1TS U3191 ( .A0(n483), .A1(n958), .B0(n4217), .B1(n3228), .Y(n1256) );
  AOI222XLTS U3192 ( .A0(n3291), .A1(n94), .B0(n3906), .B1(n3277), .C0(
        dataIn_NORTH[23]), .C1(n3259), .Y(n1257) );
  AOI22X1TS U3193 ( .A0(n489), .A1(n3249), .B0(n4208), .B1(n3227), .Y(n1250)
         );
  AOI222XLTS U3194 ( .A0(n3288), .A1(n95), .B0(n3897), .B1(n3276), .C0(n4345), 
        .C1(n3258), .Y(n1251) );
  AOI22X1TS U3195 ( .A0(n494), .A1(n3246), .B0(n4202), .B1(n3226), .Y(n1246)
         );
  AOI222XLTS U3196 ( .A0(n3289), .A1(n96), .B0(n3891), .B1(n3275), .C0(n4340), 
        .C1(n3258), .Y(n1247) );
  AOI22X1TS U3197 ( .A0(n508), .A1(n3245), .B0(n4193), .B1(n3226), .Y(n1240)
         );
  AOI222XLTS U3198 ( .A0(n3288), .A1(n97), .B0(n3882), .B1(n3275), .C0(n4334), 
        .C1(n3257), .Y(n1241) );
  AOI22X1TS U3199 ( .A0(n514), .A1(n3245), .B0(n4187), .B1(n3225), .Y(n1236)
         );
  AOI222XLTS U3200 ( .A0(n280), .A1(n98), .B0(n3876), .B1(n3274), .C0(n4330), 
        .C1(n3256), .Y(n1237) );
  AOI22X1TS U3201 ( .A0(n557), .A1(n3242), .B0(n4163), .B1(n3223), .Y(n1220)
         );
  AOI222XLTS U3202 ( .A0(n3292), .A1(n99), .B0(n3852), .B1(n3272), .C0(n4315), 
        .C1(n3254), .Y(n1221) );
  AOI22X1TS U3203 ( .A0(n561), .A1(n3242), .B0(n4160), .B1(n3223), .Y(n1218)
         );
  AOI222XLTS U3204 ( .A0(n281), .A1(n100), .B0(n3849), .B1(n3272), .C0(n4312), 
        .C1(n3254), .Y(n1219) );
  AOI22X1TS U3205 ( .A0(n564), .A1(n3241), .B0(n4154), .B1(n3223), .Y(n1214)
         );
  AOI222XLTS U3206 ( .A0(n3294), .A1(n101), .B0(n3843), .B1(n3272), .C0(
        dataIn_NORTH[2]), .C1(n3254), .Y(n1215) );
  AOI22X1TS U3207 ( .A0(n474), .A1(n767), .B0(n4232), .B1(n741), .Y(n1074) );
  AOI222XLTS U3208 ( .A0(n286), .A1(n102), .B0(n3921), .B1(n777), .C0(n4360), 
        .C1(n348), .Y(n1075) );
  AOI22X1TS U3209 ( .A0(n476), .A1(n765), .B0(n4229), .B1(n741), .Y(n1072) );
  AOI222XLTS U3210 ( .A0(n328), .A1(n103), .B0(n3918), .B1(n777), .C0(n4358), 
        .C1(n392), .Y(n1073) );
  AOI22X1TS U3211 ( .A0(n484), .A1(n764), .B0(n4217), .B1(n740), .Y(n1064) );
  AOI222XLTS U3212 ( .A0(n328), .A1(n104), .B0(n3906), .B1(n776), .C0(n4350), 
        .C1(n342), .Y(n1065) );
  AOI22X1TS U3213 ( .A0(n490), .A1(n757), .B0(n4208), .B1(n739), .Y(n1058) );
  AOI222XLTS U3214 ( .A0(n322), .A1(n105), .B0(n3897), .B1(n784), .C0(n4345), 
        .C1(n342), .Y(n1059) );
  AOI22X1TS U3215 ( .A0(n545), .A1(n760), .B0(n4175), .B1(n739), .Y(n1036) );
  AOI222XLTS U3216 ( .A0(n322), .A1(n106), .B0(n3864), .B1(n774), .C0(n4322), 
        .C1(n271), .Y(n1037) );
  AOI22X1TS U3217 ( .A0(n559), .A1(n760), .B0(n4163), .B1(n735), .Y(n1028) );
  AOI222XLTS U3218 ( .A0(n322), .A1(n107), .B0(n3852), .B1(n773), .C0(n4315), 
        .C1(n392), .Y(n1029) );
  AOI22X1TS U3219 ( .A0(n565), .A1(n761), .B0(n4154), .B1(n735), .Y(n1022) );
  AOI222XLTS U3220 ( .A0(n324), .A1(n108), .B0(n3843), .B1(n773), .C0(n4308), 
        .C1(n344), .Y(n1023) );
  AOI22X1TS U3221 ( .A0(n567), .A1(n761), .B0(n4151), .B1(n751), .Y(n1020) );
  AOI222XLTS U3222 ( .A0(n385), .A1(n109), .B0(n3840), .B1(n772), .C0(n4306), 
        .C1(n245), .Y(n1021) );
  AOI22X1TS U3223 ( .A0(n569), .A1(n762), .B0(n4148), .B1(n751), .Y(n1018) );
  AOI222XLTS U3224 ( .A0(n328), .A1(n110), .B0(n3837), .B1(n772), .C0(n4305), 
        .C1(n348), .Y(n1019) );
  AOI22X1TS U3225 ( .A0(n554), .A1(n3242), .B0(n4169), .B1(n3224), .Y(n1224)
         );
  AOI222XLTS U3226 ( .A0(n3292), .A1(n111), .B0(n3858), .B1(n3273), .C0(n4318), 
        .C1(n3255), .Y(n1225) );
  AOI22X1TS U3227 ( .A0(n886), .A1(readRequesterAddress[2]), .B0(n4112), .B1(
        n869), .Y(n1734) );
  AOI222XLTS U3228 ( .A0(n3773), .A1(n112), .B0(n4269), .B1(n3197), .C0(n4384), 
        .C1(n3781), .Y(n1735) );
  AOI22X1TS U3229 ( .A0(n469), .A1(n1546), .B0(n4082), .B1(n867), .Y(n1206) );
  AOI222XLTS U3230 ( .A0(n350), .A1(n113), .B0(n4239), .B1(n973), .C0(n4364), 
        .C1(n3780), .Y(n1207) );
  AOI22X1TS U3231 ( .A0(n471), .A1(n1546), .B0(n4079), .B1(n871), .Y(n1204) );
  AOI222XLTS U3232 ( .A0(n3772), .A1(n114), .B0(n4236), .B1(n3196), .C0(n4363), 
        .C1(n3783), .Y(n1205) );
  AOI22X1TS U3233 ( .A0(n473), .A1(n1531), .B0(n4076), .B1(n865), .Y(n1202) );
  AOI222XLTS U3234 ( .A0(n274), .A1(n115), .B0(n4233), .B1(n3196), .C0(n4360), 
        .C1(n3783), .Y(n1203) );
  AOI22X1TS U3235 ( .A0(n477), .A1(n955), .B0(n4070), .B1(n975), .Y(n1198) );
  AOI222XLTS U3236 ( .A0(n351), .A1(n116), .B0(n4227), .B1(n3196), .C0(n4357), 
        .C1(n3783), .Y(n1199) );
  AOI22X1TS U3237 ( .A0(n479), .A1(n1402), .B0(n4067), .B1(n862), .Y(n1196) );
  AOI222XLTS U3238 ( .A0(n354), .A1(n117), .B0(n4224), .B1(n3195), .C0(n4354), 
        .C1(n3784), .Y(n1197) );
  AOI22X1TS U3239 ( .A0(n483), .A1(n1654), .B0(n4061), .B1(n862), .Y(n1192) );
  AOI222XLTS U3240 ( .A0(n351), .A1(n118), .B0(n4218), .B1(n3195), .C0(n4350), 
        .C1(n3783), .Y(n1193) );
  AOI22X1TS U3241 ( .A0(n487), .A1(n919), .B0(n4055), .B1(n861), .Y(n1188) );
  AOI222XLTS U3242 ( .A0(n3772), .A1(n119), .B0(n4212), .B1(n3194), .C0(n4346), 
        .C1(n3788), .Y(n1189) );
  AOI22X1TS U3243 ( .A0(n489), .A1(n919), .B0(n4052), .B1(n861), .Y(n1186) );
  AOI222XLTS U3244 ( .A0(n432), .A1(n120), .B0(n4209), .B1(n3194), .C0(n4345), 
        .C1(n3786), .Y(n1187) );
  AOI22X1TS U3245 ( .A0(n491), .A1(n919), .B0(n4049), .B1(n861), .Y(n1184) );
  AOI222XLTS U3246 ( .A0(n3771), .A1(n121), .B0(n4206), .B1(n3194), .C0(n4342), 
        .C1(n502), .Y(n1185) );
  AOI22X1TS U3247 ( .A0(n493), .A1(n936), .B0(n4046), .B1(n860), .Y(n1182) );
  AOI222XLTS U3248 ( .A0(n354), .A1(n122), .B0(n4203), .B1(n3193), .C0(n4340), 
        .C1(n502), .Y(n1183) );
  AOI22X1TS U3249 ( .A0(n495), .A1(n919), .B0(n4043), .B1(n860), .Y(n1180) );
  AOI222XLTS U3250 ( .A0(n433), .A1(n123), .B0(n4200), .B1(n3193), .C0(n4338), 
        .C1(n3779), .Y(n1181) );
  AOI22X1TS U3251 ( .A0(n507), .A1(n955), .B0(n4037), .B1(n860), .Y(n1176) );
  AOI222XLTS U3252 ( .A0(n273), .A1(n124), .B0(n4194), .B1(n3193), .C0(n4334), 
        .C1(n3779), .Y(n1177) );
  AOI22X1TS U3253 ( .A0(n509), .A1(n936), .B0(n4034), .B1(n859), .Y(n1174) );
  AOI222XLTS U3254 ( .A0(n356), .A1(n125), .B0(n4191), .B1(n3192), .C0(n4333), 
        .C1(n3779), .Y(n1175) );
  AOI22X1TS U3255 ( .A0(n512), .A1(n936), .B0(n4031), .B1(n859), .Y(n1172) );
  AOI222XLTS U3256 ( .A0(n3772), .A1(n126), .B0(n4188), .B1(n3192), .C0(n4330), 
        .C1(n3778), .Y(n1173) );
  AOI22X1TS U3257 ( .A0(n515), .A1(n955), .B0(n4028), .B1(n859), .Y(n1170) );
  AOI222XLTS U3258 ( .A0(n273), .A1(n127), .B0(n4185), .B1(n3192), .C0(n4328), 
        .C1(n3778), .Y(n1171) );
  AOI22X1TS U3259 ( .A0(n536), .A1(n955), .B0(n4025), .B1(n859), .Y(n1168) );
  AOI222XLTS U3260 ( .A0(n356), .A1(n128), .B0(n4182), .B1(n3192), .C0(n4326), 
        .C1(n3778), .Y(n1169) );
  AOI22X1TS U3261 ( .A0(n544), .A1(n957), .B0(n4019), .B1(n861), .Y(n1164) );
  AOI222XLTS U3262 ( .A0(n351), .A1(n129), .B0(n4176), .B1(n1894), .C0(n4322), 
        .C1(n3777), .Y(n1165) );
  AOI22X1TS U3263 ( .A0(n546), .A1(n957), .B0(n4016), .B1(n858), .Y(n1162) );
  AOI222XLTS U3264 ( .A0(n273), .A1(n130), .B0(n4173), .B1(n1894), .C0(n4320), 
        .C1(n3777), .Y(n1163) );
  AOI22X1TS U3265 ( .A0(n551), .A1(n957), .B0(n4013), .B1(n858), .Y(n1160) );
  AOI222XLTS U3266 ( .A0(n3772), .A1(n131), .B0(n4170), .B1(n1894), .C0(n4318), 
        .C1(n3777), .Y(n1161) );
  AOI22X1TS U3267 ( .A0(n557), .A1(n957), .B0(n4007), .B1(n857), .Y(n1156) );
  AOI222XLTS U3268 ( .A0(n352), .A1(n132), .B0(n4164), .B1(n1822), .C0(n4315), 
        .C1(n3776), .Y(n1157) );
  AOI22X1TS U3269 ( .A0(n560), .A1(n970), .B0(n4004), .B1(n857), .Y(n1154) );
  AOI222XLTS U3270 ( .A0(n274), .A1(n133), .B0(n4161), .B1(n1822), .C0(n4312), 
        .C1(n3776), .Y(n1155) );
  AOI22X1TS U3271 ( .A0(n562), .A1(n986), .B0(n4001), .B1(n857), .Y(n1152) );
  AOI222XLTS U3272 ( .A0(n355), .A1(n134), .B0(n4158), .B1(n1822), .C0(n4311), 
        .C1(n3776), .Y(n1153) );
  AOI22X1TS U3273 ( .A0(n1585), .A1(n201), .B0(n4121), .B1(n866), .Y(n1740) );
  AOI222XLTS U3274 ( .A0(n350), .A1(n135), .B0(n4278), .B1(n1817), .C0(n4391), 
        .C1(n3781), .Y(n1741) );
  AOI22X1TS U3275 ( .A0(n886), .A1(readRequesterAddress[4]), .B0(n4118), .B1(
        n871), .Y(n1738) );
  AOI222XLTS U3276 ( .A0(n274), .A1(n136), .B0(n4275), .B1(n3197), .C0(n4388), 
        .C1(n3781), .Y(n1739) );
  AOI22X1TS U3277 ( .A0(n886), .A1(readRequesterAddress[3]), .B0(n4115), .B1(
        n866), .Y(n1736) );
  AOI222XLTS U3278 ( .A0(n3773), .A1(n137), .B0(n4272), .B1(n3197), .C0(n4387), 
        .C1(n3781), .Y(n1737) );
  AOI22X1TS U3279 ( .A0(n1544), .A1(readRequesterAddress[1]), .B0(n4109), .B1(
        n867), .Y(n1732) );
  AOI222XLTS U3280 ( .A0(n355), .A1(n138), .B0(n4266), .B1(n3199), .C0(n4382), 
        .C1(n3780), .Y(n1733) );
  AOI22X1TS U3281 ( .A0(n886), .A1(n179), .B0(n4106), .B1(n869), .Y(n1730) );
  AOI222XLTS U3282 ( .A0(n355), .A1(n139), .B0(n4263), .B1(n3202), .C0(n4380), 
        .C1(n3780), .Y(n1731) );
  AOI22X1TS U3283 ( .A0(n475), .A1(n974), .B0(n4073), .B1(n871), .Y(n1200) );
  AOI222XLTS U3284 ( .A0(n354), .A1(n140), .B0(n4230), .B1(n3196), .C0(n4358), 
        .C1(n3782), .Y(n1201) );
  AOI22X1TS U3285 ( .A0(n541), .A1(n986), .B0(n4022), .B1(n858), .Y(n1166) );
  AOI222XLTS U3286 ( .A0(n352), .A1(n141), .B0(n4179), .B1(n1894), .C0(n4324), 
        .C1(n3778), .Y(n1167) );
  AOI22X1TS U3287 ( .A0(n566), .A1(n970), .B0(n3995), .B1(n856), .Y(n1148) );
  AOI222XLTS U3288 ( .A0(n432), .A1(n142), .B0(n4152), .B1(n1817), .C0(n4306), 
        .C1(n3775), .Y(n1149) );
  AOI22X1TS U3289 ( .A0(n467), .A1(n986), .B0(n4085), .B1(n868), .Y(n1208) );
  AOI222XLTS U3290 ( .A0(n356), .A1(n143), .B0(n4242), .B1(n3202), .C0(n4366), 
        .C1(n3780), .Y(n1209) );
  AOI22X1TS U3291 ( .A0(n481), .A1(n1546), .B0(n4064), .B1(n862), .Y(n1194) );
  AOI222XLTS U3292 ( .A0(n274), .A1(n144), .B0(n4221), .B1(n3195), .C0(n4352), 
        .C1(n3785), .Y(n1195) );
  AOI22X1TS U3293 ( .A0(n485), .A1(n1585), .B0(n4058), .B1(n862), .Y(n1190) );
  AOI222XLTS U3294 ( .A0(n352), .A1(n145), .B0(n4215), .B1(n3195), .C0(n4348), 
        .C1(n3787), .Y(n1191) );
  AOI22X1TS U3295 ( .A0(n503), .A1(n936), .B0(n4040), .B1(n860), .Y(n1178) );
  AOI222XLTS U3296 ( .A0(n350), .A1(n146), .B0(n4197), .B1(n3193), .C0(n4336), 
        .C1(n3779), .Y(n1179) );
  AOI22X1TS U3297 ( .A0(n555), .A1(n970), .B0(n4010), .B1(n858), .Y(n1158) );
  AOI222XLTS U3298 ( .A0(n433), .A1(n147), .B0(n4167), .B1(n3194), .C0(n4316), 
        .C1(n3777), .Y(n1159) );
  AOI22X1TS U3299 ( .A0(n564), .A1(n970), .B0(n3998), .B1(n857), .Y(n1150) );
  AOI222XLTS U3300 ( .A0(n356), .A1(n148), .B0(n4155), .B1(n1822), .C0(n4308), 
        .C1(n3776), .Y(n1151) );
  AOI22X1TS U3301 ( .A0(n568), .A1(n986), .B0(n3992), .B1(n856), .Y(n1146) );
  AOI222XLTS U3302 ( .A0(n3771), .A1(n149), .B0(n4149), .B1(n1817), .C0(n4305), 
        .C1(n3775), .Y(n1147) );
  AOI22X1TS U3303 ( .A0(n3947), .A1(n3498), .B0(n4378), .B1(n367), .Y(n901) );
  AOI22X1TS U3304 ( .A0(n3944), .A1(n3497), .B0(n4377), .B1(n366), .Y(n899) );
  AOI22X1TS U3305 ( .A0(n3938), .A1(n3497), .B0(n4372), .B1(n3718), .Y(n895)
         );
  AOI22X1TS U3306 ( .A0(n3941), .A1(n3497), .B0(n4375), .B1(n368), .Y(n897) );
  AOI22X1TS U3307 ( .A0(n3935), .A1(n3497), .B0(n4371), .B1(n368), .Y(n893) );
  AOI222XLTS U3308 ( .A0(n4091), .A1(n3545), .B0(n183), .B1(n3538), .C0(n4248), 
        .C1(n3516), .Y(n894) );
  AOI22X1TS U3309 ( .A0(n3932), .A1(n3503), .B0(n4369), .B1(n370), .Y(n887) );
  AOI222XLTS U3310 ( .A0(n3826), .A1(n1560), .B0(readIn_SOUTH), .B1(n1561), 
        .C0(n3834), .C1(n1562), .Y(n1559) );
  AOI2BB2X1TS U3311 ( .B0(n1578), .B1(n1579), .A0N(n3296), .A1N(
        readOutbuffer[3]), .Y(n2566) );
  OAI22X1TS U3312 ( .A0(n458), .A1(n876), .B0(n594), .B1(n875), .Y(n2887) );
  OAI22X1TS U3313 ( .A0(n873), .A1(n458), .B0(n595), .B1(n875), .Y(n2888) );
  NAND2X1TS U3314 ( .A(n3820), .B(n519), .Y(n1572) );
  OAI22X1TS U3315 ( .A0(n686), .A1(n2903), .B0(n1987), .B1(n3597), .Y(n1986)
         );
  NOR4XLTS U3316 ( .A(n1988), .B(n1989), .C(n1990), .D(n1991), .Y(n1987) );
  AO22X1TS U3317 ( .A0(n230), .A1(\requesterAddressbuffer[3][5] ), .B0(
        \requesterAddressbuffer[6][5] ), .B1(n1834), .Y(n1989) );
  OAI2BB2XLTS U3318 ( .B0(n30), .B1(n3642), .A0N(
        \requesterAddressbuffer[0][5] ), .A1N(n276), .Y(n1988) );
  OAI22X1TS U3319 ( .A0(n686), .A1(n2902), .B0(n1979), .B1(n3597), .Y(n1978)
         );
  NOR4XLTS U3320 ( .A(n1980), .B(n1981), .C(n1982), .D(n1983), .Y(n1979) );
  AO22X1TS U3321 ( .A0(n282), .A1(\requesterAddressbuffer[3][4] ), .B0(
        \requesterAddressbuffer[6][4] ), .B1(n1834), .Y(n1981) );
  OAI2BB2XLTS U3322 ( .B0(n31), .B1(n3642), .A0N(
        \requesterAddressbuffer[0][4] ), .A1N(n1833), .Y(n1980) );
  OAI22X1TS U3323 ( .A0(n685), .A1(n2901), .B0(n1963), .B1(n3596), .Y(n1962)
         );
  NOR4XLTS U3324 ( .A(n1964), .B(n1965), .C(n1966), .D(n1967), .Y(n1963) );
  AO22X1TS U3325 ( .A0(n230), .A1(\requesterAddressbuffer[3][2] ), .B0(
        \requesterAddressbuffer[6][2] ), .B1(n1834), .Y(n1965) );
  OAI2BB2XLTS U3326 ( .B0(n32), .B1(n3641), .A0N(
        \requesterAddressbuffer[0][2] ), .A1N(n276), .Y(n1964) );
  OAI22X1TS U3327 ( .A0(n685), .A1(n2900), .B0(n1955), .B1(n3596), .Y(n1954)
         );
  NOR4XLTS U3328 ( .A(n1956), .B(n1957), .C(n1958), .D(n1959), .Y(n1955) );
  AO22X1TS U3329 ( .A0(n282), .A1(\requesterAddressbuffer[3][1] ), .B0(
        \requesterAddressbuffer[6][1] ), .B1(n466), .Y(n1957) );
  OAI2BB2XLTS U3330 ( .B0(n33), .B1(n3641), .A0N(
        \requesterAddressbuffer[0][1] ), .A1N(n1833), .Y(n1956) );
  OAI22X1TS U3331 ( .A0(n685), .A1(n2283), .B0(n1971), .B1(n3596), .Y(n1970)
         );
  NOR4XLTS U3332 ( .A(n1972), .B(n1973), .C(n1974), .D(n1975), .Y(n1971) );
  AO22X1TS U3333 ( .A0(n230), .A1(\requesterAddressbuffer[3][3] ), .B0(
        \requesterAddressbuffer[6][3] ), .B1(n466), .Y(n1973) );
  OAI2BB2XLTS U3334 ( .B0(n34), .B1(n3641), .A0N(
        \requesterAddressbuffer[0][3] ), .A1N(n276), .Y(n1972) );
  OAI22X1TS U3335 ( .A0(n685), .A1(n2284), .B0(n1947), .B1(n3596), .Y(n1946)
         );
  NOR4XLTS U3336 ( .A(n1948), .B(n1949), .C(n1950), .D(n1951), .Y(n1947) );
  AO22X1TS U3337 ( .A0(n282), .A1(\requesterAddressbuffer[3][0] ), .B0(
        \requesterAddressbuffer[6][0] ), .B1(n466), .Y(n1949) );
  OAI2BB2XLTS U3338 ( .B0(n35), .B1(n3641), .A0N(
        \requesterAddressbuffer[0][0] ), .A1N(n1833), .Y(n1948) );
  OAI22X1TS U3339 ( .A0(n3191), .A1(n686), .B0(n2243), .B1(n3594), .Y(n2242)
         );
  NOR4XLTS U3340 ( .A(n2244), .B(n2245), .C(n2246), .D(n2247), .Y(n2243) );
  OAI22X1TS U3341 ( .A0(n3190), .A1(n3626), .B0(n3189), .B1(n3645), .Y(n2244)
         );
  OAI22X1TS U3342 ( .A0(n3188), .A1(n3673), .B0(n3187), .B1(n3688), .Y(n2245)
         );
  OAI22X1TS U3343 ( .A0(n3182), .A1(n695), .B0(n2235), .B1(n3608), .Y(n2234)
         );
  NOR4XLTS U3344 ( .A(n2236), .B(n2237), .C(n2238), .D(n2239), .Y(n2235) );
  OAI22X1TS U3345 ( .A0(n3177), .A1(n3626), .B0(n3181), .B1(n3655), .Y(n2236)
         );
  OAI22X1TS U3346 ( .A0(n3175), .A1(n3682), .B0(n3176), .B1(n3688), .Y(n2237)
         );
  OAI22X1TS U3347 ( .A0(n3173), .A1(n695), .B0(n2227), .B1(n3606), .Y(n2226)
         );
  NOR4XLTS U3348 ( .A(n2228), .B(n2229), .C(n2230), .D(n2231), .Y(n2227) );
  OAI22X1TS U3349 ( .A0(n3166), .A1(n3626), .B0(n3165), .B1(n550), .Y(n2228)
         );
  OAI22X1TS U3350 ( .A0(n3170), .A1(n3687), .B0(n3168), .B1(n3688), .Y(n2229)
         );
  OAI22X1TS U3351 ( .A0(n3164), .A1(n695), .B0(n2219), .B1(n3603), .Y(n2218)
         );
  NOR4XLTS U3352 ( .A(n2220), .B(n2221), .C(n2222), .D(n2223), .Y(n2219) );
  OAI22X1TS U3353 ( .A0(n3157), .A1(n3626), .B0(n3163), .B1(n3652), .Y(n2220)
         );
  OAI22X1TS U3354 ( .A0(n3159), .A1(n3687), .B0(n3160), .B1(n3688), .Y(n2221)
         );
  OAI22X1TS U3355 ( .A0(n3155), .A1(n695), .B0(n2211), .B1(n3603), .Y(n2210)
         );
  NOR4XLTS U3356 ( .A(n2212), .B(n2213), .C(n2214), .D(n2215), .Y(n2211) );
  OAI22X1TS U3357 ( .A0(n3148), .A1(n3627), .B0(n3152), .B1(n3651), .Y(n2212)
         );
  OAI22X1TS U3358 ( .A0(n3150), .A1(n3679), .B0(n3151), .B1(n3689), .Y(n2213)
         );
  OAI22X1TS U3359 ( .A0(n3146), .A1(n694), .B0(n2203), .B1(n3608), .Y(n2202)
         );
  NOR4XLTS U3360 ( .A(n2204), .B(n2205), .C(n2206), .D(n2207), .Y(n2203) );
  OAI22X1TS U3361 ( .A0(n3141), .A1(n3627), .B0(n3145), .B1(n3654), .Y(n2204)
         );
  OAI22X1TS U3362 ( .A0(n3139), .A1(n3679), .B0(n3140), .B1(n3689), .Y(n2205)
         );
  OAI22X1TS U3363 ( .A0(n3137), .A1(n694), .B0(n2195), .B1(n3604), .Y(n2194)
         );
  NOR4XLTS U3364 ( .A(n2196), .B(n2197), .C(n2198), .D(n2199), .Y(n2195) );
  OAI22X1TS U3365 ( .A0(n3134), .A1(n3627), .B0(n3132), .B1(n3650), .Y(n2196)
         );
  OAI22X1TS U3366 ( .A0(n3135), .A1(n3679), .B0(n3130), .B1(n3689), .Y(n2197)
         );
  OAI22X1TS U3367 ( .A0(n3128), .A1(n694), .B0(n2187), .B1(n3605), .Y(n2186)
         );
  NOR4XLTS U3368 ( .A(n2188), .B(n2189), .C(n2190), .D(n2191), .Y(n2187) );
  OAI22X1TS U3369 ( .A0(n3125), .A1(n3627), .B0(n3127), .B1(n3655), .Y(n2188)
         );
  OAI22X1TS U3370 ( .A0(n3123), .A1(n3679), .B0(n3120), .B1(n3689), .Y(n2189)
         );
  OAI22X1TS U3371 ( .A0(n3119), .A1(n694), .B0(n2179), .B1(n3605), .Y(n2178)
         );
  NOR4XLTS U3372 ( .A(n2180), .B(n2181), .C(n2182), .D(n2183), .Y(n2179) );
  OAI22X1TS U3373 ( .A0(n3112), .A1(n3639), .B0(n3116), .B1(n3655), .Y(n2180)
         );
  OAI22X1TS U3374 ( .A0(n3111), .A1(n3684), .B0(n3118), .B1(n3701), .Y(n2181)
         );
  OAI22X1TS U3375 ( .A0(n3110), .A1(n693), .B0(n2171), .B1(n3608), .Y(n2170)
         );
  NOR4XLTS U3376 ( .A(n2172), .B(n2173), .C(n2174), .D(n2175), .Y(n2171) );
  OAI22X1TS U3377 ( .A0(n3109), .A1(n3636), .B0(n3106), .B1(n3649), .Y(n2172)
         );
  OAI22X1TS U3378 ( .A0(n3107), .A1(n3685), .B0(n3102), .B1(n3698), .Y(n2173)
         );
  OAI22X1TS U3379 ( .A0(n3101), .A1(n693), .B0(n2163), .B1(n3604), .Y(n2162)
         );
  NOR4XLTS U3380 ( .A(n2164), .B(n2165), .C(n2166), .D(n2167), .Y(n2163) );
  OAI22X1TS U3381 ( .A0(n3094), .A1(n3637), .B0(n3095), .B1(n3653), .Y(n2164)
         );
  OAI22X1TS U3382 ( .A0(n3096), .A1(n3685), .B0(n3098), .B1(n3700), .Y(n2165)
         );
  OAI22X1TS U3383 ( .A0(n3092), .A1(n693), .B0(n2155), .B1(n3602), .Y(n2154)
         );
  NOR4XLTS U3384 ( .A(n2156), .B(n2157), .C(n2158), .D(n2159), .Y(n2155) );
  OAI22X1TS U3385 ( .A0(n3085), .A1(n3634), .B0(n3086), .B1(n3653), .Y(n2156)
         );
  OAI22X1TS U3386 ( .A0(n3084), .A1(n3683), .B0(n3091), .B1(n3696), .Y(n2157)
         );
  OAI22X1TS U3387 ( .A0(n3083), .A1(n693), .B0(n2147), .B1(n3602), .Y(n2146)
         );
  NOR4XLTS U3388 ( .A(n2148), .B(n2149), .C(n2150), .D(n2151), .Y(n2147) );
  OAI22X1TS U3389 ( .A0(n3080), .A1(n3638), .B0(n3081), .B1(n3653), .Y(n2148)
         );
  OAI22X1TS U3390 ( .A0(n3076), .A1(n3681), .B0(n3079), .B1(n3699), .Y(n2149)
         );
  OAI22X1TS U3391 ( .A0(n3074), .A1(n692), .B0(n2139), .B1(n3602), .Y(n2138)
         );
  NOR4XLTS U3392 ( .A(n2140), .B(n2141), .C(n2142), .D(n2143), .Y(n2139) );
  OAI22X1TS U3393 ( .A0(n3071), .A1(n3636), .B0(n3073), .B1(n3656), .Y(n2140)
         );
  OAI22X1TS U3394 ( .A0(n3068), .A1(n3683), .B0(n3067), .B1(n547), .Y(n2141)
         );
  OAI22X1TS U3395 ( .A0(n3065), .A1(n692), .B0(n2131), .B1(n3602), .Y(n2130)
         );
  NOR4XLTS U3396 ( .A(n2132), .B(n2133), .C(n2134), .D(n2135), .Y(n2131) );
  OAI22X1TS U3397 ( .A0(n3062), .A1(n3638), .B0(n3058), .B1(n3656), .Y(n2132)
         );
  OAI22X1TS U3398 ( .A0(n3064), .A1(n3686), .B0(n3057), .B1(n3698), .Y(n2133)
         );
  OAI22X1TS U3399 ( .A0(n3056), .A1(n692), .B0(n2123), .B1(n3601), .Y(n2122)
         );
  NOR4XLTS U3400 ( .A(n2124), .B(n2125), .C(n2126), .D(n2127), .Y(n2123) );
  OAI22X1TS U3401 ( .A0(n3053), .A1(n3637), .B0(n3054), .B1(n3656), .Y(n2124)
         );
  OAI22X1TS U3402 ( .A0(n3055), .A1(n3682), .B0(n3052), .B1(n3699), .Y(n2125)
         );
  OAI22X1TS U3403 ( .A0(n3047), .A1(n692), .B0(n2115), .B1(n3601), .Y(n2114)
         );
  NOR4XLTS U3404 ( .A(n2116), .B(n2117), .C(n2118), .D(n2119), .Y(n2115) );
  OAI22X1TS U3405 ( .A0(n3042), .A1(n3635), .B0(n3040), .B1(n3649), .Y(n2116)
         );
  OAI22X1TS U3406 ( .A0(n3043), .A1(n3678), .B0(n3039), .B1(n3697), .Y(n2117)
         );
  OAI22X1TS U3407 ( .A0(n3038), .A1(n691), .B0(n2107), .B1(n3601), .Y(n2106)
         );
  NOR4XLTS U3408 ( .A(n2108), .B(n2109), .C(n2110), .D(n2111), .Y(n2107) );
  OAI22X1TS U3409 ( .A0(n3035), .A1(n3635), .B0(n3031), .B1(n3646), .Y(n2108)
         );
  OAI22X1TS U3410 ( .A0(n3033), .A1(n3678), .B0(n3032), .B1(n3697), .Y(n2109)
         );
  OAI22X1TS U3411 ( .A0(n3029), .A1(n691), .B0(n2099), .B1(n3601), .Y(n2098)
         );
  NOR4XLTS U3412 ( .A(n2100), .B(n2101), .C(n2102), .D(n2103), .Y(n2099) );
  OAI22X1TS U3413 ( .A0(n3022), .A1(n3639), .B0(n3028), .B1(n3646), .Y(n2100)
         );
  OAI22X1TS U3414 ( .A0(n3025), .A1(n3678), .B0(n3024), .B1(n3700), .Y(n2101)
         );
  OAI22X1TS U3415 ( .A0(n3020), .A1(n691), .B0(n2091), .B1(n3600), .Y(n2090)
         );
  NOR4XLTS U3416 ( .A(n2092), .B(n2093), .C(n2094), .D(n2095), .Y(n2091) );
  OAI22X1TS U3417 ( .A0(n3015), .A1(n3640), .B0(n3016), .B1(n3646), .Y(n2092)
         );
  OAI22X1TS U3418 ( .A0(n3017), .A1(n3678), .B0(n3013), .B1(n3701), .Y(n2093)
         );
  OAI22X1TS U3419 ( .A0(n3011), .A1(n691), .B0(n2083), .B1(n3600), .Y(n2082)
         );
  NOR4XLTS U3420 ( .A(n2084), .B(n2085), .C(n2086), .D(n2087), .Y(n2083) );
  OAI22X1TS U3421 ( .A0(n3010), .A1(n3628), .B0(n3005), .B1(n3646), .Y(n2084)
         );
  OAI22X1TS U3422 ( .A0(n3006), .A1(n3677), .B0(n3003), .B1(n3690), .Y(n2085)
         );
  OAI22X1TS U3423 ( .A0(n3002), .A1(n690), .B0(n2075), .B1(n3600), .Y(n2074)
         );
  NOR4XLTS U3424 ( .A(n2076), .B(n2077), .C(n2078), .D(n2079), .Y(n2075) );
  OAI22X1TS U3425 ( .A0(n2997), .A1(n3628), .B0(n2998), .B1(n3645), .Y(n2076)
         );
  OAI22X1TS U3426 ( .A0(n2999), .A1(n3677), .B0(n3001), .B1(n3690), .Y(n2077)
         );
  OAI22X1TS U3427 ( .A0(n2993), .A1(n690), .B0(n2067), .B1(n3600), .Y(n2066)
         );
  NOR4XLTS U3428 ( .A(n2068), .B(n2069), .C(n2070), .D(n2071), .Y(n2067) );
  OAI22X1TS U3429 ( .A0(n2986), .A1(n3628), .B0(n2988), .B1(n3645), .Y(n2068)
         );
  OAI22X1TS U3430 ( .A0(n2990), .A1(n3677), .B0(n2987), .B1(n3690), .Y(n2069)
         );
  OAI22X1TS U3431 ( .A0(n2984), .A1(n690), .B0(n2059), .B1(n3599), .Y(n2058)
         );
  NOR4XLTS U3432 ( .A(n2060), .B(n2061), .C(n2062), .D(n2063), .Y(n2059) );
  OAI22X1TS U3433 ( .A0(n2977), .A1(n3628), .B0(n2982), .B1(n3645), .Y(n2060)
         );
  OAI22X1TS U3434 ( .A0(n2983), .A1(n3676), .B0(n2976), .B1(n3690), .Y(n2061)
         );
  OAI22X1TS U3435 ( .A0(n2975), .A1(n689), .B0(n2051), .B1(n3599), .Y(n2050)
         );
  NOR4XLTS U3436 ( .A(n2052), .B(n2053), .C(n2054), .D(n2055), .Y(n2051) );
  OAI22X1TS U3437 ( .A0(n2972), .A1(n3629), .B0(n2970), .B1(n3644), .Y(n2052)
         );
  OAI22X1TS U3438 ( .A0(n2968), .A1(n3676), .B0(n2971), .B1(n3691), .Y(n2053)
         );
  OAI22X1TS U3439 ( .A0(n2966), .A1(n689), .B0(n2043), .B1(n3599), .Y(n2042)
         );
  NOR4XLTS U3440 ( .A(n2044), .B(n2045), .C(n2046), .D(n2047), .Y(n2043) );
  OAI22X1TS U3441 ( .A0(n2963), .A1(n3629), .B0(n2960), .B1(n3644), .Y(n2044)
         );
  OAI22X1TS U3442 ( .A0(n2961), .A1(n3676), .B0(n2965), .B1(n3691), .Y(n2045)
         );
  OAI22X1TS U3443 ( .A0(n2957), .A1(n689), .B0(n2035), .B1(n3598), .Y(n2034)
         );
  NOR4XLTS U3444 ( .A(n2036), .B(n2037), .C(n2038), .D(n2039), .Y(n2035) );
  OAI22X1TS U3445 ( .A0(n2950), .A1(n3629), .B0(n2954), .B1(n3644), .Y(n2036)
         );
  OAI22X1TS U3446 ( .A0(n2951), .A1(n3676), .B0(n2953), .B1(n3691), .Y(n2037)
         );
  OAI22X1TS U3447 ( .A0(n2948), .A1(n689), .B0(n2027), .B1(n3598), .Y(n2026)
         );
  NOR4XLTS U3448 ( .A(n2028), .B(n2029), .C(n2030), .D(n2031), .Y(n2027) );
  OAI22X1TS U3449 ( .A0(n2947), .A1(n3629), .B0(n2943), .B1(n3644), .Y(n2028)
         );
  OAI22X1TS U3450 ( .A0(n2944), .A1(n3675), .B0(n2941), .B1(n3691), .Y(n2029)
         );
  OAI22X1TS U3451 ( .A0(n2939), .A1(n688), .B0(n2019), .B1(n3598), .Y(n2018)
         );
  NOR4XLTS U3452 ( .A(n2020), .B(n2021), .C(n2022), .D(n2023), .Y(n2019) );
  OAI22X1TS U3453 ( .A0(n2936), .A1(n3630), .B0(n2932), .B1(n3643), .Y(n2020)
         );
  OAI22X1TS U3454 ( .A0(n2934), .A1(n3675), .B0(n2937), .B1(n3692), .Y(n2021)
         );
  OAI22X1TS U3455 ( .A0(n2930), .A1(n688), .B0(n2011), .B1(n3598), .Y(n2010)
         );
  NOR4XLTS U3456 ( .A(n2012), .B(n2013), .C(n2014), .D(n2015), .Y(n2011) );
  OAI22X1TS U3457 ( .A0(n2923), .A1(n3630), .B0(n2927), .B1(n3643), .Y(n2012)
         );
  OAI22X1TS U3458 ( .A0(n2924), .A1(n3675), .B0(n2922), .B1(n3692), .Y(n2013)
         );
  OAI22X1TS U3459 ( .A0(n2921), .A1(n688), .B0(n2003), .B1(n3597), .Y(n2002)
         );
  NOR4XLTS U3460 ( .A(n2004), .B(n2005), .C(n2006), .D(n2007), .Y(n2003) );
  OAI22X1TS U3461 ( .A0(n2914), .A1(n3630), .B0(n2919), .B1(n3643), .Y(n2004)
         );
  OAI22X1TS U3462 ( .A0(n2920), .A1(n3675), .B0(n2918), .B1(n3692), .Y(n2005)
         );
  OAI22X1TS U3463 ( .A0(n2912), .A1(n688), .B0(n1995), .B1(n3597), .Y(n1994)
         );
  NOR4XLTS U3464 ( .A(n1996), .B(n1997), .C(n1998), .D(n1999), .Y(n1995) );
  OAI22X1TS U3465 ( .A0(n2907), .A1(n3630), .B0(n2908), .B1(n3643), .Y(n1996)
         );
  OAI22X1TS U3466 ( .A0(n2911), .A1(n3674), .B0(n2906), .B1(n3692), .Y(n1997)
         );
  OAI22X1TS U3467 ( .A0(n2899), .A1(n687), .B0(n1939), .B1(n3595), .Y(n1938)
         );
  NOR4XLTS U3468 ( .A(n1940), .B(n1941), .C(n1942), .D(n1943), .Y(n1939) );
  OAI22X1TS U3469 ( .A0(n2898), .A1(n3631), .B0(n2896), .B1(n3652), .Y(n1940)
         );
  OAI22X1TS U3470 ( .A0(n2892), .A1(n3674), .B0(n2894), .B1(n3693), .Y(n1941)
         );
  OAI22X1TS U3471 ( .A0(n2890), .A1(n687), .B0(n1931), .B1(n3595), .Y(n1930)
         );
  NOR4XLTS U3472 ( .A(n1932), .B(n1933), .C(n1934), .D(n1935), .Y(n1931) );
  OAI22X1TS U3473 ( .A0(n2393), .A1(n3631), .B0(n2392), .B1(n3652), .Y(n1932)
         );
  OAI22X1TS U3474 ( .A0(n2394), .A1(n3674), .B0(n2390), .B1(n3693), .Y(n1933)
         );
  OAI22X1TS U3475 ( .A0(n2388), .A1(n690), .B0(n1923), .B1(n3595), .Y(n1922)
         );
  NOR4XLTS U3476 ( .A(n1924), .B(n1925), .C(n1926), .D(n1927), .Y(n1923) );
  OAI22X1TS U3477 ( .A0(n2385), .A1(n3631), .B0(n2383), .B1(n3651), .Y(n1924)
         );
  OAI22X1TS U3478 ( .A0(n2381), .A1(n3674), .B0(n2387), .B1(n3693), .Y(n1925)
         );
  OAI22X1TS U3479 ( .A0(n2379), .A1(n687), .B0(n1915), .B1(n3595), .Y(n1914)
         );
  NOR4XLTS U3480 ( .A(n1916), .B(n1917), .C(n1918), .D(n1919), .Y(n1915) );
  OAI22X1TS U3481 ( .A0(n2374), .A1(n3631), .B0(n2378), .B1(n3642), .Y(n1916)
         );
  OAI22X1TS U3482 ( .A0(n2377), .A1(n3673), .B0(n2376), .B1(n3693), .Y(n1917)
         );
  OAI22X1TS U3483 ( .A0(n2370), .A1(n686), .B0(n1907), .B1(n3594), .Y(n1906)
         );
  NOR4XLTS U3484 ( .A(n1908), .B(n1909), .C(n1910), .D(n1911), .Y(n1907) );
  OAI22X1TS U3485 ( .A0(n2369), .A1(n3632), .B0(n2365), .B1(n3650), .Y(n1908)
         );
  OAI22X1TS U3486 ( .A0(n2363), .A1(n3673), .B0(n2367), .B1(n3694), .Y(n1909)
         );
  OAI22X1TS U3487 ( .A0(n2361), .A1(n687), .B0(n1898), .B1(n3594), .Y(n1897)
         );
  NOR4XLTS U3488 ( .A(n1899), .B(n1900), .C(n1901), .D(n1902), .Y(n1898) );
  OAI22X1TS U3489 ( .A0(n2355), .A1(n3632), .B0(n2360), .B1(n3642), .Y(n1899)
         );
  OAI22X1TS U3490 ( .A0(n2356), .A1(n3673), .B0(n2358), .B1(n3694), .Y(n1900)
         );
  OAI221XLTS U3491 ( .A0(n1807), .A1(n1808), .B0(n1809), .B1(n1810), .C0(n4392), .Y(n1806) );
  OAI211X1TS U3492 ( .A0(n3625), .A1(n20), .B0(n2287), .C0(n1816), .Y(n1808)
         );
  OAI221XLTS U3493 ( .A0(n3634), .A1(n583), .B0(n3696), .B1(n28), .C0(n1819), 
        .Y(n1807) );
  OAI211X1TS U3494 ( .A0(n309), .A1(n631), .B0(n1887), .C0(n1888), .Y(n2441)
         );
  AOI22X1TS U3495 ( .A0(n570), .A1(n1889), .B0(n697), .B1(
        destinationAddressOut[13]), .Y(n1887) );
  AOI222XLTS U3496 ( .A0(n462), .A1(n4302), .B0(n653), .B1(n4146), .C0(n644), 
        .C1(destinationAddressIn_WEST[13]), .Y(n1888) );
  NAND4X1TS U3497 ( .A(n1890), .B(n1891), .C(n1892), .D(n1893), .Y(n1889) );
  OAI211X1TS U3498 ( .A0(n300), .A1(n631), .B0(n1880), .C0(n1881), .Y(n2442)
         );
  AOI22X1TS U3499 ( .A0(n571), .A1(n1882), .B0(n697), .B1(
        destinationAddressOut[12]), .Y(n1880) );
  AOI222XLTS U3500 ( .A0(n461), .A1(n4299), .B0(n653), .B1(n4143), .C0(n648), 
        .C1(destinationAddressIn_WEST[12]), .Y(n1881) );
  NAND4X1TS U3501 ( .A(n1883), .B(n1884), .C(n1885), .D(n1886), .Y(n1882) );
  OAI211X1TS U3502 ( .A0(n312), .A1(n631), .B0(n1873), .C0(n1874), .Y(n2443)
         );
  AOI22X1TS U3503 ( .A0(n571), .A1(n1875), .B0(n697), .B1(
        destinationAddressOut[11]), .Y(n1873) );
  AOI222XLTS U3504 ( .A0(n462), .A1(n4296), .B0(n653), .B1(n4140), .C0(n647), 
        .C1(destinationAddressIn_WEST[11]), .Y(n1874) );
  NAND4X1TS U3505 ( .A(n1876), .B(n1877), .C(n1878), .D(n1879), .Y(n1875) );
  OAI211X1TS U3506 ( .A0(n303), .A1(n632), .B0(n1866), .C0(n1867), .Y(n2444)
         );
  AOI22X1TS U3507 ( .A0(n570), .A1(n1868), .B0(n697), .B1(
        destinationAddressOut[10]), .Y(n1866) );
  AOI222XLTS U3508 ( .A0(n461), .A1(n4293), .B0(n653), .B1(n4137), .C0(n646), 
        .C1(destinationAddressIn_WEST[10]), .Y(n1867) );
  NAND4X1TS U3509 ( .A(n1869), .B(n1870), .C(n1871), .D(n1872), .Y(n1868) );
  OAI211X1TS U3510 ( .A0(n306), .A1(n632), .B0(n1859), .C0(n1860), .Y(n2445)
         );
  AOI22X1TS U3511 ( .A0(n571), .A1(n1861), .B0(n698), .B1(
        destinationAddressOut[9]), .Y(n1859) );
  AOI222XLTS U3512 ( .A0(n462), .A1(n4290), .B0(n652), .B1(n4134), .C0(n651), 
        .C1(destinationAddressIn_WEST[9]), .Y(n1860) );
  NAND4X1TS U3513 ( .A(n1862), .B(n1863), .C(n1864), .D(n1865), .Y(n1861) );
  OAI211X1TS U3514 ( .A0(n315), .A1(n632), .B0(n1852), .C0(n1853), .Y(n2446)
         );
  AOI22X1TS U3515 ( .A0(n570), .A1(n1854), .B0(n698), .B1(
        destinationAddressOut[8]), .Y(n1852) );
  AOI222XLTS U3516 ( .A0(n461), .A1(n4287), .B0(n652), .B1(n4131), .C0(n650), 
        .C1(destinationAddressIn_WEST[8]), .Y(n1853) );
  NAND4X1TS U3517 ( .A(n1855), .B(n1856), .C(n1857), .D(n1858), .Y(n1854) );
  OAI211X1TS U3518 ( .A0(n297), .A1(n633), .B0(n1845), .C0(n1846), .Y(n2447)
         );
  AOI22X1TS U3519 ( .A0(n570), .A1(n1847), .B0(n698), .B1(
        destinationAddressOut[7]), .Y(n1845) );
  AOI222XLTS U3520 ( .A0(n462), .A1(n4284), .B0(n652), .B1(n4128), .C0(n649), 
        .C1(destinationAddressIn_WEST[7]), .Y(n1846) );
  NAND4X1TS U3521 ( .A(n1848), .B(n1849), .C(n1850), .D(n1851), .Y(n1847) );
  OAI211X1TS U3522 ( .A0(n294), .A1(n633), .B0(n1835), .C0(n1836), .Y(n2448)
         );
  AOI22X1TS U3523 ( .A0(n571), .A1(n1840), .B0(n698), .B1(
        destinationAddressOut[6]), .Y(n1835) );
  AOI222XLTS U3524 ( .A0(n461), .A1(n4281), .B0(n652), .B1(n4125), .C0(n645), 
        .C1(destinationAddressIn_WEST[6]), .Y(n1836) );
  NAND4X1TS U3525 ( .A(n1841), .B(n1842), .C(n1843), .D(n1844), .Y(n1840) );
  OAI211X1TS U3526 ( .A0(n4243), .A1(n3592), .B0(n2240), .C0(n2241), .Y(n2397)
         );
  AOI22X1TS U3527 ( .A0(n606), .A1(n468), .B0(n649), .B1(n3929), .Y(n2240) );
  AOI221X1TS U3528 ( .A0(n610), .A1(dataIn_NORTH[31]), .B0(n661), .B1(n4086), 
        .C0(n2242), .Y(n2241) );
  OAI211X1TS U3529 ( .A0(n4240), .A1(n3592), .B0(n2232), .C0(n2233), .Y(n2398)
         );
  AOI22X1TS U3530 ( .A0(n607), .A1(n470), .B0(n649), .B1(n3926), .Y(n2232) );
  AOI221X1TS U3531 ( .A0(n610), .A1(dataIn_NORTH[30]), .B0(n663), .B1(n4083), 
        .C0(n2234), .Y(n2233) );
  OAI211X1TS U3532 ( .A0(n4237), .A1(n3593), .B0(n2224), .C0(n2225), .Y(n2399)
         );
  AOI22X1TS U3533 ( .A0(n608), .A1(n472), .B0(n649), .B1(n3923), .Y(n2224) );
  AOI221X1TS U3534 ( .A0(n610), .A1(dataIn_NORTH[29]), .B0(n663), .B1(n4080), 
        .C0(n2226), .Y(n2225) );
  OAI211X1TS U3535 ( .A0(n4234), .A1(n3589), .B0(n2216), .C0(n2217), .Y(n2400)
         );
  AOI22X1TS U3536 ( .A0(n609), .A1(n474), .B0(n645), .B1(n3920), .Y(n2216) );
  AOI221X1TS U3537 ( .A0(n610), .A1(dataIn_NORTH[28]), .B0(n660), .B1(n4077), 
        .C0(n2218), .Y(n2217) );
  OAI211X1TS U3538 ( .A0(n4231), .A1(n3580), .B0(n2208), .C0(n2209), .Y(n2401)
         );
  AOI22X1TS U3539 ( .A0(n596), .A1(n476), .B0(n636), .B1(n3917), .Y(n2208) );
  AOI221X1TS U3540 ( .A0(n611), .A1(dataIn_NORTH[27]), .B0(n662), .B1(n4074), 
        .C0(n2210), .Y(n2209) );
  OAI211X1TS U3541 ( .A0(n4228), .A1(n3580), .B0(n2200), .C0(n2201), .Y(n2402)
         );
  AOI22X1TS U3542 ( .A0(n596), .A1(n478), .B0(n636), .B1(n3914), .Y(n2200) );
  AOI221X1TS U3543 ( .A0(n611), .A1(dataIn_NORTH[26]), .B0(n661), .B1(n4071), 
        .C0(n2202), .Y(n2201) );
  OAI211X1TS U3544 ( .A0(n4225), .A1(n3580), .B0(n2192), .C0(n2193), .Y(n2403)
         );
  AOI22X1TS U3545 ( .A0(n596), .A1(n480), .B0(n636), .B1(n3911), .Y(n2192) );
  AOI221X1TS U3546 ( .A0(n611), .A1(dataIn_NORTH[25]), .B0(n662), .B1(n4068), 
        .C0(n2194), .Y(n2193) );
  OAI211X1TS U3547 ( .A0(n4222), .A1(n3580), .B0(n2184), .C0(n2185), .Y(n2404)
         );
  AOI22X1TS U3548 ( .A0(n596), .A1(n482), .B0(n636), .B1(n3908), .Y(n2184) );
  AOI221X1TS U3549 ( .A0(n611), .A1(dataIn_NORTH[24]), .B0(n667), .B1(n4065), 
        .C0(n2186), .Y(n2185) );
  OAI211X1TS U3550 ( .A0(n4219), .A1(n3589), .B0(n2176), .C0(n2177), .Y(n2405)
         );
  AOI22X1TS U3551 ( .A0(n607), .A1(n484), .B0(n637), .B1(n3905), .Y(n2176) );
  AOI221X1TS U3552 ( .A0(n612), .A1(dataIn_NORTH[23]), .B0(n659), .B1(n4062), 
        .C0(n2178), .Y(n2177) );
  OAI211X1TS U3553 ( .A0(n4216), .A1(n3588), .B0(n2168), .C0(n2169), .Y(n2406)
         );
  AOI22X1TS U3554 ( .A0(n603), .A1(n486), .B0(n637), .B1(n3902), .Y(n2168) );
  AOI221X1TS U3555 ( .A0(n612), .A1(dataIn_NORTH[22]), .B0(n659), .B1(n4059), 
        .C0(n2170), .Y(n2169) );
  OAI211X1TS U3556 ( .A0(n4213), .A1(n3587), .B0(n2160), .C0(n2161), .Y(n2407)
         );
  AOI22X1TS U3557 ( .A0(n605), .A1(n488), .B0(n637), .B1(n3899), .Y(n2160) );
  AOI221X1TS U3558 ( .A0(n612), .A1(dataIn_NORTH[21]), .B0(n659), .B1(n4056), 
        .C0(n2162), .Y(n2161) );
  OAI211X1TS U3559 ( .A0(n4210), .A1(n3591), .B0(n2152), .C0(n2153), .Y(n2408)
         );
  AOI22X1TS U3560 ( .A0(n607), .A1(n490), .B0(n637), .B1(n3896), .Y(n2152) );
  AOI221X1TS U3561 ( .A0(n612), .A1(dataIn_NORTH[20]), .B0(n659), .B1(n4053), 
        .C0(n2154), .Y(n2153) );
  OAI211X1TS U3562 ( .A0(n4207), .A1(n3590), .B0(n2144), .C0(n2145), .Y(n2409)
         );
  AOI22X1TS U3563 ( .A0(n606), .A1(n492), .B0(n646), .B1(n3893), .Y(n2144) );
  AOI221X1TS U3564 ( .A0(n613), .A1(dataIn_NORTH[19]), .B0(n658), .B1(n4050), 
        .C0(n2146), .Y(n2145) );
  OAI211X1TS U3565 ( .A0(n4204), .A1(n3590), .B0(n2136), .C0(n2137), .Y(n2410)
         );
  AOI22X1TS U3566 ( .A0(n606), .A1(n494), .B0(n647), .B1(n3890), .Y(n2136) );
  AOI221X1TS U3567 ( .A0(n613), .A1(dataIn_NORTH[18]), .B0(n658), .B1(n4047), 
        .C0(n2138), .Y(n2137) );
  OAI211X1TS U3568 ( .A0(n4201), .A1(n3591), .B0(n2128), .C0(n2129), .Y(n2411)
         );
  AOI22X1TS U3569 ( .A0(n608), .A1(n501), .B0(n1839), .B1(n3887), .Y(n2128) );
  AOI221X1TS U3570 ( .A0(n613), .A1(dataIn_NORTH[17]), .B0(n658), .B1(n4044), 
        .C0(n2130), .Y(n2129) );
  OAI211X1TS U3571 ( .A0(n4198), .A1(n3591), .B0(n2120), .C0(n2121), .Y(n2412)
         );
  AOI22X1TS U3572 ( .A0(n604), .A1(n505), .B0(n1839), .B1(n3884), .Y(n2120) );
  AOI221X1TS U3573 ( .A0(n613), .A1(dataIn_NORTH[16]), .B0(n658), .B1(n4041), 
        .C0(n2122), .Y(n2121) );
  OAI211X1TS U3574 ( .A0(n4195), .A1(n3590), .B0(n2112), .C0(n2113), .Y(n2413)
         );
  AOI22X1TS U3575 ( .A0(n606), .A1(n508), .B0(n647), .B1(n3881), .Y(n2112) );
  AOI221X1TS U3576 ( .A0(n614), .A1(dataIn_NORTH[15]), .B0(n657), .B1(n4038), 
        .C0(n2114), .Y(n2113) );
  OAI211X1TS U3577 ( .A0(n4192), .A1(n3588), .B0(n2104), .C0(n2105), .Y(n2414)
         );
  AOI22X1TS U3578 ( .A0(n604), .A1(n511), .B0(n647), .B1(n3878), .Y(n2104) );
  AOI221X1TS U3579 ( .A0(n614), .A1(dataIn_NORTH[14]), .B0(n657), .B1(n4035), 
        .C0(n2106), .Y(n2105) );
  OAI211X1TS U3580 ( .A0(n4189), .A1(n3587), .B0(n2096), .C0(n2097), .Y(n2415)
         );
  AOI22X1TS U3581 ( .A0(n603), .A1(n514), .B0(n644), .B1(n3875), .Y(n2096) );
  AOI221X1TS U3582 ( .A0(n614), .A1(dataIn_NORTH[13]), .B0(n657), .B1(n4032), 
        .C0(n2098), .Y(n2097) );
  OAI211X1TS U3583 ( .A0(n4186), .A1(n3590), .B0(n2088), .C0(n2089), .Y(n2416)
         );
  AOI22X1TS U3584 ( .A0(n605), .A1(n516), .B0(n648), .B1(n3872), .Y(n2088) );
  AOI221X1TS U3585 ( .A0(n614), .A1(dataIn_NORTH[12]), .B0(n657), .B1(n4029), 
        .C0(n2090), .Y(n2089) );
  OAI211X1TS U3586 ( .A0(n4183), .A1(n3581), .B0(n2080), .C0(n2081), .Y(n2417)
         );
  AOI22X1TS U3587 ( .A0(n597), .A1(n537), .B0(n638), .B1(n3869), .Y(n2080) );
  AOI221X1TS U3588 ( .A0(n622), .A1(dataIn_NORTH[11]), .B0(n661), .B1(n4026), 
        .C0(n2082), .Y(n2081) );
  OAI211X1TS U3589 ( .A0(n4180), .A1(n3581), .B0(n2072), .C0(n2073), .Y(n2418)
         );
  AOI22X1TS U3590 ( .A0(n597), .A1(n543), .B0(n638), .B1(n3866), .Y(n2072) );
  AOI221X1TS U3591 ( .A0(n622), .A1(dataIn_NORTH[10]), .B0(n664), .B1(n4023), 
        .C0(n2074), .Y(n2073) );
  OAI211X1TS U3592 ( .A0(n4177), .A1(n3581), .B0(n2064), .C0(n2065), .Y(n2419)
         );
  AOI22X1TS U3593 ( .A0(n597), .A1(n545), .B0(n638), .B1(n3863), .Y(n2064) );
  AOI221X1TS U3594 ( .A0(n622), .A1(dataIn_NORTH[9]), .B0(n665), .B1(n4020), 
        .C0(n2066), .Y(n2065) );
  OAI211X1TS U3595 ( .A0(n4174), .A1(n3581), .B0(n2056), .C0(n2057), .Y(n2420)
         );
  AOI22X1TS U3596 ( .A0(n597), .A1(n548), .B0(n638), .B1(n3860), .Y(n2056) );
  AOI221X1TS U3597 ( .A0(n622), .A1(dataIn_NORTH[8]), .B0(n1838), .B1(n4017), 
        .C0(n2058), .Y(n2057) );
  OAI211X1TS U3598 ( .A0(n4171), .A1(n3582), .B0(n2048), .C0(n2049), .Y(n2421)
         );
  AOI22X1TS U3599 ( .A0(n598), .A1(n554), .B0(n639), .B1(n3857), .Y(n2048) );
  AOI221X1TS U3600 ( .A0(n623), .A1(dataIn_NORTH[7]), .B0(n662), .B1(n4014), 
        .C0(n2050), .Y(n2049) );
  OAI211X1TS U3601 ( .A0(n4168), .A1(n3582), .B0(n2040), .C0(n2041), .Y(n2422)
         );
  AOI22X1TS U3602 ( .A0(n598), .A1(n556), .B0(n639), .B1(n3854), .Y(n2040) );
  AOI221X1TS U3603 ( .A0(n623), .A1(dataIn_NORTH[6]), .B0(n664), .B1(n4011), 
        .C0(n2042), .Y(n2041) );
  OAI211X1TS U3604 ( .A0(n4165), .A1(n3582), .B0(n2032), .C0(n2033), .Y(n2423)
         );
  AOI22X1TS U3605 ( .A0(n598), .A1(n559), .B0(n639), .B1(n3851), .Y(n2032) );
  AOI221X1TS U3606 ( .A0(n623), .A1(dataIn_NORTH[5]), .B0(n665), .B1(n4008), 
        .C0(n2034), .Y(n2033) );
  OAI211X1TS U3607 ( .A0(n4162), .A1(n3582), .B0(n2024), .C0(n2025), .Y(n2424)
         );
  AOI22X1TS U3608 ( .A0(n598), .A1(n561), .B0(n639), .B1(n3848), .Y(n2024) );
  AOI221X1TS U3609 ( .A0(n623), .A1(dataIn_NORTH[4]), .B0(n1838), .B1(n4005), 
        .C0(n2026), .Y(n2025) );
  OAI211X1TS U3610 ( .A0(n4159), .A1(n3583), .B0(n2016), .C0(n2017), .Y(n2425)
         );
  AOI22X1TS U3611 ( .A0(n599), .A1(n563), .B0(n640), .B1(n3845), .Y(n2016) );
  AOI221X1TS U3612 ( .A0(n624), .A1(dataIn_NORTH[3]), .B0(n660), .B1(n4002), 
        .C0(n2018), .Y(n2017) );
  OAI211X1TS U3613 ( .A0(n4156), .A1(n3583), .B0(n2008), .C0(n2009), .Y(n2426)
         );
  AOI22X1TS U3614 ( .A0(n599), .A1(n565), .B0(n640), .B1(n3842), .Y(n2008) );
  AOI221X1TS U3615 ( .A0(n624), .A1(dataIn_NORTH[2]), .B0(n662), .B1(n3999), 
        .C0(n2010), .Y(n2009) );
  OAI211X1TS U3616 ( .A0(n4153), .A1(n3583), .B0(n2000), .C0(n2001), .Y(n2427)
         );
  AOI22X1TS U3617 ( .A0(n599), .A1(n567), .B0(n640), .B1(n3839), .Y(n2000) );
  AOI221X1TS U3618 ( .A0(n624), .A1(dataIn_NORTH[1]), .B0(n665), .B1(n3996), 
        .C0(n2002), .Y(n2001) );
  OAI211X1TS U3619 ( .A0(n4150), .A1(n3583), .B0(n1992), .C0(n1993), .Y(n2428)
         );
  AOI22X1TS U3620 ( .A0(n599), .A1(n569), .B0(n640), .B1(n3836), .Y(n1992) );
  AOI221X1TS U3621 ( .A0(n624), .A1(dataIn_NORTH[0]), .B0(n666), .B1(n3993), 
        .C0(n1994), .Y(n1993) );
  OAI211X1TS U3622 ( .A0(n4261), .A1(n3584), .B0(n1984), .C0(n1985), .Y(n2429)
         );
  AOI22X1TS U3623 ( .A0(n600), .A1(n201), .B0(n641), .B1(n3947), .Y(n1984) );
  AOI221X1TS U3624 ( .A0(n628), .A1(requesterAddressIn_NORTH[5]), .B0(n656), 
        .B1(n4104), .C0(n1986), .Y(n1985) );
  OAI211X1TS U3625 ( .A0(n4258), .A1(n3584), .B0(n1976), .C0(n1977), .Y(n2430)
         );
  AOI22X1TS U3626 ( .A0(n600), .A1(n196), .B0(n641), .B1(n3944), .Y(n1976) );
  AOI221X1TS U3627 ( .A0(n628), .A1(requesterAddressIn_NORTH[4]), .B0(n656), 
        .B1(n4101), .C0(n1978), .Y(n1977) );
  OAI211X1TS U3628 ( .A0(n4252), .A1(n3584), .B0(n1960), .C0(n1961), .Y(n2432)
         );
  AOI22X1TS U3629 ( .A0(n600), .A1(n165), .B0(n641), .B1(n3938), .Y(n1960) );
  AOI221X1TS U3630 ( .A0(n628), .A1(requesterAddressIn_NORTH[2]), .B0(n656), 
        .B1(n4095), .C0(n1962), .Y(n1961) );
  OAI211X1TS U3631 ( .A0(n4249), .A1(n3585), .B0(n1952), .C0(n1953), .Y(n2433)
         );
  AOI22X1TS U3632 ( .A0(n601), .A1(n164), .B0(n642), .B1(n3935), .Y(n1952) );
  AOI221X1TS U3633 ( .A0(n629), .A1(requesterAddressIn_NORTH[1]), .B0(n655), 
        .B1(n4092), .C0(n1954), .Y(n1953) );
  OAI211X1TS U3634 ( .A0(n4279), .A1(n3585), .B0(n1936), .C0(n1937), .Y(n2435)
         );
  AOI22X1TS U3635 ( .A0(n601), .A1(n198), .B0(n642), .B1(n3965), .Y(n1936) );
  AOI221X1TS U3636 ( .A0(n629), .A1(destinationAddressIn_NORTH[5]), .B0(n655), 
        .B1(n4122), .C0(n1938), .Y(n1937) );
  OAI211X1TS U3637 ( .A0(n4276), .A1(n3585), .B0(n1928), .C0(n1929), .Y(n2436)
         );
  AOI22X1TS U3638 ( .A0(n601), .A1(n195), .B0(n642), .B1(n3962), .Y(n1928) );
  AOI221X1TS U3639 ( .A0(n629), .A1(destinationAddressIn_NORTH[4]), .B0(n655), 
        .B1(n4119), .C0(n1930), .Y(n1929) );
  OAI211X1TS U3640 ( .A0(n4273), .A1(n3586), .B0(n1920), .C0(n1921), .Y(n2437)
         );
  AOI22X1TS U3641 ( .A0(n602), .A1(n192), .B0(n643), .B1(n3959), .Y(n1920) );
  AOI221X1TS U3642 ( .A0(n630), .A1(destinationAddressIn_NORTH[3]), .B0(n654), 
        .B1(n4116), .C0(n1922), .Y(n1921) );
  OAI211X1TS U3643 ( .A0(n4270), .A1(n3586), .B0(n1912), .C0(n1913), .Y(n2438)
         );
  AOI22X1TS U3644 ( .A0(n602), .A1(n187), .B0(n643), .B1(n3956), .Y(n1912) );
  AOI221X1TS U3645 ( .A0(n630), .A1(destinationAddressIn_NORTH[2]), .B0(n654), 
        .B1(n4113), .C0(n1914), .Y(n1913) );
  OAI211X1TS U3646 ( .A0(n4267), .A1(n3586), .B0(n1904), .C0(n1905), .Y(n2439)
         );
  AOI22X1TS U3647 ( .A0(n602), .A1(n183), .B0(n643), .B1(n3953), .Y(n1904) );
  AOI221X1TS U3648 ( .A0(n630), .A1(destinationAddressIn_NORTH[1]), .B0(n654), 
        .B1(n4110), .C0(n1906), .Y(n1905) );
  OAI211X1TS U3649 ( .A0(n4264), .A1(n3586), .B0(n1895), .C0(n1896), .Y(n2440)
         );
  AOI22X1TS U3650 ( .A0(n602), .A1(n179), .B0(n643), .B1(n3950), .Y(n1895) );
  AOI221X1TS U3651 ( .A0(n630), .A1(destinationAddressIn_NORTH[0]), .B0(n654), 
        .B1(n4107), .C0(n1897), .Y(n1896) );
  OAI211X1TS U3652 ( .A0(n4255), .A1(n3584), .B0(n1968), .C0(n1969), .Y(n2431)
         );
  AOI22X1TS U3653 ( .A0(n600), .A1(n191), .B0(n641), .B1(n3941), .Y(n1968) );
  AOI221X1TS U3654 ( .A0(n628), .A1(requesterAddressIn_NORTH[3]), .B0(n656), 
        .B1(n4098), .C0(n1970), .Y(n1969) );
  OAI211X1TS U3655 ( .A0(n4246), .A1(n3585), .B0(n1944), .C0(n1945), .Y(n2434)
         );
  AOI22X1TS U3656 ( .A0(n601), .A1(n180), .B0(n642), .B1(n3932), .Y(n1944) );
  AOI221X1TS U3657 ( .A0(n629), .A1(requesterAddressIn_NORTH[0]), .B0(n655), 
        .B1(n4089), .C0(n1946), .Y(n1945) );
  NOR2X1TS U3658 ( .A(reset), .B(n2287), .Y(n1825) );
  INVX2TS U3659 ( .A(readIn_SOUTH), .Y(n744) );
  INVX2TS U3660 ( .A(writeIn_NORTH), .Y(n730) );
  OAI22X1TS U3661 ( .A0(n1824), .A1(n1825), .B0(n1826), .B1(n1827), .Y(n1823)
         );
  AOI31X1TS U3662 ( .A0(n1828), .A1(n1829), .A2(n1830), .B0(reset), .Y(n1824)
         );
  OAI22X1TS U3663 ( .A0(n3832), .A1(n1813), .B0(n3819), .B1(n1811), .Y(n1827)
         );
  OAI22X1TS U3664 ( .A0(n465), .A1(n553), .B0(n9), .B1(n3599), .Y(n2889) );
  INVX2TS U3665 ( .A(destinationAddressIn_NORTH[6]), .Y(n728) );
  INVX2TS U3666 ( .A(destinationAddressIn_NORTH[12]), .Y(n722) );
  INVX2TS U3667 ( .A(destinationAddressIn_NORTH[10]), .Y(n724) );
  INVX2TS U3668 ( .A(destinationAddressIn_NORTH[9]), .Y(n725) );
  INVX2TS U3669 ( .A(destinationAddressIn_NORTH[13]), .Y(n721) );
  INVX2TS U3670 ( .A(destinationAddressIn_NORTH[11]), .Y(n723) );
  INVX2TS U3671 ( .A(destinationAddressIn_NORTH[8]), .Y(n726) );
  NOR2X1TS U3672 ( .A(n884), .B(n883), .Y(n2883) );
  AOI21X1TS U3673 ( .A0(n319), .A1(n885), .B0(n10), .Y(n884) );
  XNOR2X1TS U3674 ( .A(n2277), .B(n540), .Y(n880) );
  XNOR2X1TS U3675 ( .A(n237), .B(n317), .Y(n2277) );
  OAI22X1TS U3676 ( .A0(n3184), .A1(n3715), .B0(n3183), .B1(n3614), .Y(n2247)
         );
  OAI22X1TS U3677 ( .A0(n3179), .A1(n3715), .B0(n3174), .B1(n3623), .Y(n2239)
         );
  OAI22X1TS U3678 ( .A0(n3172), .A1(n3715), .B0(n3169), .B1(n3621), .Y(n2231)
         );
  OAI22X1TS U3679 ( .A0(n3161), .A1(n3710), .B0(n3162), .B1(n552), .Y(n2223)
         );
  OAI22X1TS U3680 ( .A0(n3147), .A1(n3715), .B0(n3154), .B1(n3622), .Y(n2215)
         );
  OAI22X1TS U3681 ( .A0(n3143), .A1(n3712), .B0(n3138), .B1(n3617), .Y(n2207)
         );
  OAI22X1TS U3682 ( .A0(n3136), .A1(n3710), .B0(n3131), .B1(n3617), .Y(n2199)
         );
  OAI22X1TS U3683 ( .A0(n3121), .A1(n3713), .B0(n3126), .B1(n3617), .Y(n2191)
         );
  OAI22X1TS U3684 ( .A0(n3114), .A1(n3714), .B0(n3117), .B1(n3617), .Y(n2183)
         );
  OAI22X1TS U3685 ( .A0(n3103), .A1(n3714), .B0(n3105), .B1(n3620), .Y(n2175)
         );
  OAI22X1TS U3686 ( .A0(n3100), .A1(n3714), .B0(n3099), .B1(n3620), .Y(n2167)
         );
  OAI22X1TS U3687 ( .A0(n3087), .A1(n3716), .B0(n3089), .B1(n3625), .Y(n2159)
         );
  OAI22X1TS U3688 ( .A0(n3082), .A1(n3711), .B0(n3078), .B1(n3623), .Y(n2151)
         );
  OAI22X1TS U3689 ( .A0(n3069), .A1(n3711), .B0(n3066), .B1(n3616), .Y(n2143)
         );
  OAI22X1TS U3690 ( .A0(n3060), .A1(n3714), .B0(n3063), .B1(n3616), .Y(n2135)
         );
  OAI22X1TS U3691 ( .A0(n3049), .A1(n3717), .B0(n3048), .B1(n3616), .Y(n2127)
         );
  OAI22X1TS U3692 ( .A0(n3044), .A1(n3703), .B0(n3041), .B1(n3616), .Y(n2119)
         );
  OAI22X1TS U3693 ( .A0(n3037), .A1(n3703), .B0(n3034), .B1(n3615), .Y(n2111)
         );
  OAI22X1TS U3694 ( .A0(n3026), .A1(n3703), .B0(n3021), .B1(n3615), .Y(n2103)
         );
  OAI22X1TS U3695 ( .A0(n3019), .A1(n3703), .B0(n3012), .B1(n3615), .Y(n2095)
         );
  OAI22X1TS U3696 ( .A0(n3004), .A1(n3704), .B0(n3009), .B1(n3615), .Y(n2087)
         );
  OAI22X1TS U3697 ( .A0(n2996), .A1(n3704), .B0(n2995), .B1(n3614), .Y(n2079)
         );
  OAI22X1TS U3698 ( .A0(n2992), .A1(n3704), .B0(n2991), .B1(n3614), .Y(n2071)
         );
  OAI22X1TS U3699 ( .A0(n2979), .A1(n3704), .B0(n2981), .B1(n3614), .Y(n2063)
         );
  OAI22X1TS U3700 ( .A0(n2974), .A1(n3705), .B0(n2967), .B1(n3613), .Y(n2055)
         );
  OAI22X1TS U3701 ( .A0(n2959), .A1(n3705), .B0(n2964), .B1(n3613), .Y(n2047)
         );
  OAI22X1TS U3702 ( .A0(n2952), .A1(n3705), .B0(n2956), .B1(n3613), .Y(n2039)
         );
  OAI22X1TS U3703 ( .A0(n2945), .A1(n3705), .B0(n2940), .B1(n3613), .Y(n2031)
         );
  OAI22X1TS U3704 ( .A0(n2938), .A1(n3706), .B0(n2935), .B1(n3612), .Y(n2023)
         );
  OAI22X1TS U3705 ( .A0(n2925), .A1(n3706), .B0(n2929), .B1(n3612), .Y(n2015)
         );
  OAI22X1TS U3706 ( .A0(n2913), .A1(n3706), .B0(n2917), .B1(n3612), .Y(n2007)
         );
  OAI22X1TS U3707 ( .A0(n2909), .A1(n3706), .B0(n2905), .B1(n3612), .Y(n1999)
         );
  OAI22X1TS U3708 ( .A0(n2895), .A1(n3707), .B0(n2897), .B1(n3611), .Y(n1943)
         );
  OAI22X1TS U3709 ( .A0(n2389), .A1(n3707), .B0(n2395), .B1(n3611), .Y(n1935)
         );
  OAI22X1TS U3710 ( .A0(n2380), .A1(n3707), .B0(n2384), .B1(n3611), .Y(n1927)
         );
  OAI22X1TS U3711 ( .A0(n2372), .A1(n3707), .B0(n2371), .B1(n3610), .Y(n1919)
         );
  OAI22X1TS U3712 ( .A0(n2366), .A1(n3708), .B0(n2362), .B1(n3611), .Y(n1911)
         );
  OAI22X1TS U3713 ( .A0(n2359), .A1(n3708), .B0(n2353), .B1(n3610), .Y(n1902)
         );
  OAI22X1TS U3714 ( .A0(n3186), .A1(n673), .B0(n3185), .B1(n3657), .Y(n2246)
         );
  OAI22X1TS U3715 ( .A0(n3178), .A1(n679), .B0(n3180), .B1(n3669), .Y(n2238)
         );
  OAI22X1TS U3716 ( .A0(n3167), .A1(n676), .B0(n3171), .B1(n3672), .Y(n2230)
         );
  OAI22X1TS U3717 ( .A0(n3156), .A1(n676), .B0(n3158), .B1(n3668), .Y(n2222)
         );
  OAI22X1TS U3718 ( .A0(n3153), .A1(n676), .B0(n3149), .B1(n3670), .Y(n2214)
         );
  OAI22X1TS U3719 ( .A0(n3144), .A1(n676), .B0(n3142), .B1(n3667), .Y(n2206)
         );
  OAI22X1TS U3720 ( .A0(n3129), .A1(n684), .B0(n3133), .B1(n3668), .Y(n2198)
         );
  OAI22X1TS U3721 ( .A0(n3122), .A1(n681), .B0(n3124), .B1(n549), .Y(n2190) );
  OAI22X1TS U3722 ( .A0(n3115), .A1(n681), .B0(n3113), .B1(n3671), .Y(n2182)
         );
  OAI22X1TS U3723 ( .A0(n3104), .A1(n1818), .B0(n3108), .B1(n3672), .Y(n2174)
         );
  OAI22X1TS U3724 ( .A0(n3097), .A1(n684), .B0(n3093), .B1(n3665), .Y(n2166)
         );
  OAI22X1TS U3725 ( .A0(n3090), .A1(n682), .B0(n3088), .B1(n3665), .Y(n2158)
         );
  OAI22X1TS U3726 ( .A0(n3077), .A1(n682), .B0(n3075), .B1(n3665), .Y(n2150)
         );
  OAI22X1TS U3727 ( .A0(n3070), .A1(n680), .B0(n3072), .B1(n3665), .Y(n2142)
         );
  OAI22X1TS U3728 ( .A0(n3059), .A1(n675), .B0(n3061), .B1(n3664), .Y(n2134)
         );
  OAI22X1TS U3729 ( .A0(n3051), .A1(n675), .B0(n3050), .B1(n3664), .Y(n2126)
         );
  OAI22X1TS U3730 ( .A0(n3046), .A1(n675), .B0(n3045), .B1(n3664), .Y(n2118)
         );
  OAI22X1TS U3731 ( .A0(n3036), .A1(n675), .B0(n3030), .B1(n3664), .Y(n2110)
         );
  OAI22X1TS U3732 ( .A0(n3023), .A1(n674), .B0(n3027), .B1(n3663), .Y(n2102)
         );
  OAI22X1TS U3733 ( .A0(n3014), .A1(n674), .B0(n3018), .B1(n3663), .Y(n2094)
         );
  OAI22X1TS U3734 ( .A0(n3008), .A1(n674), .B0(n3007), .B1(n3663), .Y(n2086)
         );
  OAI22X1TS U3735 ( .A0(n3000), .A1(n674), .B0(n2994), .B1(n3663), .Y(n2078)
         );
  OAI22X1TS U3736 ( .A0(n2989), .A1(n673), .B0(n2985), .B1(n3662), .Y(n2070)
         );
  OAI22X1TS U3737 ( .A0(n2978), .A1(n673), .B0(n2980), .B1(n3662), .Y(n2062)
         );
  OAI22X1TS U3738 ( .A0(n2969), .A1(n673), .B0(n2973), .B1(n3662), .Y(n2054)
         );
  OAI22X1TS U3739 ( .A0(n2962), .A1(n672), .B0(n2958), .B1(n3661), .Y(n2046)
         );
  OAI22X1TS U3740 ( .A0(n2949), .A1(n672), .B0(n2955), .B1(n3661), .Y(n2038)
         );
  OAI22X1TS U3741 ( .A0(n2942), .A1(n672), .B0(n2946), .B1(n3661), .Y(n2030)
         );
  OAI22X1TS U3742 ( .A0(n2931), .A1(n672), .B0(n2933), .B1(n3661), .Y(n2022)
         );
  OAI22X1TS U3743 ( .A0(n2926), .A1(n671), .B0(n2928), .B1(n3660), .Y(n2014)
         );
  OAI22X1TS U3744 ( .A0(n2916), .A1(n671), .B0(n2915), .B1(n3660), .Y(n2006)
         );
  OAI22X1TS U3745 ( .A0(n2904), .A1(n671), .B0(n2910), .B1(n3660), .Y(n1998)
         );
  OAI22X1TS U3746 ( .A0(n2893), .A1(n669), .B0(n2891), .B1(n3658), .Y(n1942)
         );
  OAI22X1TS U3747 ( .A0(n2391), .A1(n669), .B0(n2396), .B1(n3658), .Y(n1934)
         );
  OAI22X1TS U3748 ( .A0(n2382), .A1(n669), .B0(n2386), .B1(n3658), .Y(n1926)
         );
  OAI22X1TS U3749 ( .A0(n2373), .A1(n668), .B0(n2375), .B1(n3657), .Y(n1918)
         );
  OAI22X1TS U3750 ( .A0(n2364), .A1(n668), .B0(n2368), .B1(n3657), .Y(n1910)
         );
  OAI22X1TS U3751 ( .A0(n2357), .A1(n668), .B0(n2354), .B1(n3657), .Y(n1901)
         );
  NOR3X1TS U3752 ( .A(n9), .B(n237), .C(n205), .Y(n1820) );
  NOR3X1TS U3753 ( .A(n10), .B(n236), .C(n553), .Y(n1831) );
  NAND3X1TS U3754 ( .A(n320), .B(n459), .C(n8), .Y(n1818) );
  AOI2BB2X1TS U3755 ( .B0(readOutbuffer[3]), .B1(n282), .A0N(n29), .A1N(n678), 
        .Y(n1816) );
  AOI222XLTS U3756 ( .A0(readOutbuffer[4]), .A1(n1820), .B0(readOutbuffer[7]), 
        .B1(n1821), .C0(readOutbuffer[2]), .C1(n228), .Y(n1819) );
  AOI221X1TS U3757 ( .A0(n1831), .A1(writeOutbuffer[1]), .B0(n228), .B1(
        writeOutbuffer[2]), .C0(n1832), .Y(n1830) );
  OAI22X1TS U3758 ( .A0(n21), .A1(n668), .B0(n558), .B1(n3662), .Y(n1832) );
  OA22X1TS U3759 ( .A0(n3619), .A1(n2351), .B0(n3708), .B1(n2352), .Y(n1890)
         );
  OA22X1TS U3760 ( .A0(n3619), .A1(n2343), .B0(n3708), .B1(n2338), .Y(n1883)
         );
  OA22X1TS U3761 ( .A0(n3619), .A1(n2333), .B0(n3709), .B1(n2329), .Y(n1876)
         );
  OA22X1TS U3762 ( .A0(n3624), .A1(n2327), .B0(n3709), .B1(n2324), .Y(n1869)
         );
  OA22X1TS U3763 ( .A0(n3618), .A1(n2315), .B0(n3709), .B1(n2313), .Y(n1862)
         );
  OA22X1TS U3764 ( .A0(n3618), .A1(n2311), .B0(n3709), .B1(n2310), .Y(n1855)
         );
  OA22X1TS U3765 ( .A0(n3618), .A1(n2303), .B0(n3710), .B1(n2297), .Y(n1848)
         );
  OA22X1TS U3766 ( .A0(n3618), .A1(n2291), .B0(n3710), .B1(n2290), .Y(n1841)
         );
  OA22X1TS U3767 ( .A0(n3647), .A1(n2346), .B0(n3632), .B1(n2345), .Y(n1893)
         );
  OA22X1TS U3768 ( .A0(n3647), .A1(n2342), .B0(n3632), .B1(n2344), .Y(n1886)
         );
  OA22X1TS U3769 ( .A0(n3647), .A1(n2336), .B0(n3633), .B1(n2332), .Y(n1879)
         );
  OA22X1TS U3770 ( .A0(n3647), .A1(n2326), .B0(n3633), .B1(n2323), .Y(n1872)
         );
  OA22X1TS U3771 ( .A0(n3648), .A1(n2314), .B0(n3633), .B1(n2318), .Y(n1865)
         );
  OA22X1TS U3772 ( .A0(n3648), .A1(n2308), .B0(n3633), .B1(n2312), .Y(n1858)
         );
  OA22X1TS U3773 ( .A0(n3648), .A1(n2304), .B0(n3634), .B1(n2302), .Y(n1851)
         );
  OA22X1TS U3774 ( .A0(n3648), .A1(n2292), .B0(n3634), .B1(n2289), .Y(n1844)
         );
  OA22X1TS U3775 ( .A0(n3670), .A1(n2349), .B0(n678), .B1(n2347), .Y(n1891) );
  OA22X1TS U3776 ( .A0(n3667), .A1(n2339), .B0(n677), .B1(n2337), .Y(n1884) );
  OA22X1TS U3777 ( .A0(n3669), .A1(n2335), .B0(n679), .B1(n2331), .Y(n1877) );
  AOI2BB2X1TS U3778 ( .B0(n1821), .B1(n593), .A0N(n678), .A1N(n2321), .Y(n1870) );
  OA22X1TS U3779 ( .A0(n3666), .A1(n2316), .B0(n677), .B1(n2317), .Y(n1863) );
  OA22X1TS U3780 ( .A0(n3666), .A1(n2309), .B0(n677), .B1(n2307), .Y(n1856) );
  OA22X1TS U3781 ( .A0(n3666), .A1(n2299), .B0(n677), .B1(n2301), .Y(n1849) );
  OA22X1TS U3782 ( .A0(n3666), .A1(n2293), .B0(n678), .B1(n2295), .Y(n1842) );
  OA22X1TS U3783 ( .A0(n3694), .A1(n2350), .B0(n3), .B1(n2348), .Y(n1892) );
  OA22X1TS U3784 ( .A0(n3694), .A1(n2340), .B0(n3680), .B1(n2341), .Y(n1885)
         );
  OA22X1TS U3785 ( .A0(n3695), .A1(n2330), .B0(n3680), .B1(n2334), .Y(n1878)
         );
  OA22X1TS U3786 ( .A0(n3695), .A1(n2328), .B0(n3681), .B1(n2322), .Y(n1871)
         );
  OA22X1TS U3787 ( .A0(n3695), .A1(n2320), .B0(n3680), .B1(n2319), .Y(n1864)
         );
  OA22X1TS U3788 ( .A0(n3695), .A1(n2306), .B0(n3680), .B1(n2305), .Y(n1857)
         );
  OA22X1TS U3789 ( .A0(n3696), .A1(n2300), .B0(n3681), .B1(n2298), .Y(n1850)
         );
  OA22X1TS U3790 ( .A0(n3696), .A1(n2296), .B0(n3681), .B1(n2294), .Y(n1843)
         );
  AOI22X1TS U3791 ( .A0(n466), .A1(writeOutbuffer[6]), .B0(writeOutbuffer[3]), 
        .B1(n230), .Y(n1828) );
  AOI22X1TS U3792 ( .A0(n1820), .A1(writeOutbuffer[4]), .B0(n276), .B1(
        writeOutbuffer[0]), .Y(n1829) );
  AOI32XLTS U3793 ( .A0(n210), .A1(n1587), .A2(n1588), .B0(n351), .B1(n153), 
        .Y(n2565) );
  AOI21XLTS U3794 ( .A0(n3833), .A1(n1589), .B0(n1590), .Y(n1588) );
  AOI21XLTS U3795 ( .A0(n3821), .A1(n522), .B0(n217), .Y(n1578) );
  OAI221XLTS U3796 ( .A0(n5), .A1(n290), .B0(n321), .B1(n158), .C0(n1548), .Y(
        n2571) );
  OAI221XLTS U3797 ( .A0(n389), .A1(n728), .B0(n2289), .B1(n434), .C0(n1787), 
        .Y(n2458) );
  OAI221XLTS U3798 ( .A0(n270), .A1(n296), .B0(n2302), .B1(n1547), .C0(n1788), 
        .Y(n2457) );
  OAI221XLTS U3799 ( .A0(n270), .A1(n726), .B0(n2312), .B1(n325), .C0(n1789), 
        .Y(n2456) );
  OAI221XLTS U3800 ( .A0(n244), .A1(n725), .B0(n2318), .B1(n1547), .C0(n1790), 
        .Y(n2455) );
  OAI221XLTS U3801 ( .A0(n5), .A1(n724), .B0(n2323), .B1(n434), .C0(n1791), 
        .Y(n2454) );
  OAI221XLTS U3802 ( .A0(n244), .A1(n723), .B0(n2332), .B1(n285), .C0(n1792), 
        .Y(n2453) );
  OAI221XLTS U3803 ( .A0(n341), .A1(n722), .B0(n2344), .B1(n434), .C0(n1793), 
        .Y(n2452) );
  OAI221XLTS U3804 ( .A0(n5), .A1(n721), .B0(n2345), .B1(n1547), .C0(n1794), 
        .Y(n2451) );
  OAI221XLTS U3805 ( .A0(n232), .A1(n290), .B0(n1542), .B1(n156), .C0(n1543), 
        .Y(n2573) );
  OAI221XLTS U3806 ( .A0(n1541), .A1(n294), .B0(n2290), .B1(n438), .C0(n1742), 
        .Y(n2486) );
  OAI221XLTS U3807 ( .A0(n1541), .A1(n297), .B0(n2297), .B1(n1542), .C0(n1743), 
        .Y(n2485) );
  OAI221XLTS U3808 ( .A0(n1541), .A1(n315), .B0(n2310), .B1(n438), .C0(n1744), 
        .Y(n2484) );
  OAI221XLTS U3809 ( .A0(n232), .A1(n306), .B0(n2313), .B1(n272), .C0(n1745), 
        .Y(n2483) );
  OAI221XLTS U3810 ( .A0(n231), .A1(n303), .B0(n2324), .B1(n272), .C0(n1746), 
        .Y(n2482) );
  OAI221XLTS U3811 ( .A0(n231), .A1(n312), .B0(n2329), .B1(n438), .C0(n1747), 
        .Y(n2481) );
  OAI221XLTS U3812 ( .A0(n232), .A1(n300), .B0(n2338), .B1(n438), .C0(n1748), 
        .Y(n2480) );
  OAI221XLTS U3813 ( .A0(n231), .A1(n308), .B0(n2352), .B1(n1542), .C0(n1749), 
        .Y(n2479) );
endmodule


module incomingPortHandler_1 ( clk, reset, localRouterAddress, 
        destinationAddressIn, requesterAddressIn, readIn, writeIn, 
        outputPortSelect, memRead, memWrite );
  input [5:0] localRouterAddress;
  input [13:0] destinationAddressIn;
  input [5:0] requesterAddressIn;
  output [3:0] outputPortSelect;
  input clk, reset, readIn, writeIn;
  output memRead, memWrite;
  wire   n70, n45, n44, n43, n42, n3, n34, n35, n36, n37, n38, n39, n40, n41,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69;

  DFFQX1TS memRead_reg ( .D(n68), .CK(clk), .Q(memRead) );
  DFFQX1TS memWrite_reg ( .D(n69), .CK(clk), .Q(n70) );
  DFFQX1TS \outputPortSelect_reg[1]  ( .D(n43), .CK(clk), .Q(
        outputPortSelect[1]) );
  DFFQX1TS \outputPortSelect_reg[3]  ( .D(n45), .CK(clk), .Q(
        outputPortSelect[3]) );
  DFFQX1TS \outputPortSelect_reg[2]  ( .D(n44), .CK(clk), .Q(
        outputPortSelect[2]) );
  DFFQX1TS \outputPortSelect_reg[0]  ( .D(n42), .CK(clk), .Q(
        outputPortSelect[0]) );
  OAI211X1TS U1 ( .A0(localRouterAddress[4]), .A1(n62), .B0(n61), .C0(
        localRouterAddress[3]), .Y(n39) );
  INVXLTS U2 ( .A(n70), .Y(n3) );
  INVXLTS U3 ( .A(n3), .Y(memWrite) );
  NAND2XLTS U4 ( .A(localRouterAddress[5]), .B(n63), .Y(n46) );
  INVXLTS U5 ( .A(destinationAddressIn[13]), .Y(n63) );
  NOR3BXLTS U6 ( .AN(n34), .B(writeIn), .C(readIn), .Y(n57) );
  NAND2XLTS U7 ( .A(localRouterAddress[2]), .B(n60), .Y(n52) );
  AOI2BB2XLTS U8 ( .B0(n59), .B1(localRouterAddress[1]), .A0N(
        destinationAddressIn[8]), .A1N(n64), .Y(n54) );
  INVX2TS U9 ( .A(reset), .Y(n34) );
  NOR2BX1TS U10 ( .AN(n56), .B(n55), .Y(n45) );
  NOR2X1TS U11 ( .A(n55), .B(n56), .Y(n44) );
  INVX2TS U12 ( .A(n49), .Y(n67) );
  OAI21X1TS U13 ( .A0(n54), .A1(n53), .B0(n52), .Y(n56) );
  NAND3BX1TS U14 ( .AN(n51), .B(n50), .C(n49), .Y(n55) );
  OAI22XLTS U15 ( .A0(localRouterAddress[1]), .A1(n59), .B0(
        localRouterAddress[2]), .B1(n60), .Y(n53) );
  AOI2BB1XLTS U16 ( .A0N(localRouterAddress[4]), .A1N(n62), .B0(n38), .Y(n48)
         );
  OAI21XLTS U17 ( .A0(readIn), .A1(writeIn), .B0(n34), .Y(n51) );
  NAND3X1TS U18 ( .A(n54), .B(n50), .C(n36), .Y(n49) );
  AOI211XLTS U19 ( .A0(destinationAddressIn[8]), .A1(n64), .B0(n53), .C0(n65), 
        .Y(n36) );
  INVX2TS U20 ( .A(n52), .Y(n65) );
  AND4X1TS U21 ( .A(n35), .B(n48), .C(n41), .D(n46), .Y(n50) );
  XNOR2XLTS U22 ( .A(destinationAddressIn[11]), .B(localRouterAddress[3]), .Y(
        n35) );
  INVXLTS U23 ( .A(destinationAddressIn[10]), .Y(n60) );
  AOI211X1TS U24 ( .A0(n40), .A1(n39), .B0(n51), .C0(n38), .Y(n42) );
  AND2X2TS U25 ( .A(n41), .B(n46), .Y(n40) );
  INVXLTS U26 ( .A(destinationAddressIn[11]), .Y(n61) );
  AOI211X1TS U27 ( .A0(n48), .A1(n47), .B0(n51), .C0(n66), .Y(n43) );
  INVX2TS U28 ( .A(n46), .Y(n66) );
  NAND3BXLTS U29 ( .AN(localRouterAddress[3]), .B(n41), .C(
        destinationAddressIn[11]), .Y(n47) );
  INVXLTS U30 ( .A(destinationAddressIn[12]), .Y(n62) );
  INVX2TS U31 ( .A(n58), .Y(n68) );
  AOI32XLTS U32 ( .A0(n67), .A1(n34), .A2(readIn), .B0(memRead), .B1(n57), .Y(
        n58) );
  INVX2TS U33 ( .A(n37), .Y(n69) );
  AOI32XLTS U34 ( .A0(n67), .A1(n34), .A2(writeIn), .B0(n70), .B1(n57), .Y(n37) );
  NAND2XLTS U35 ( .A(localRouterAddress[4]), .B(n62), .Y(n41) );
  NOR2XLTS U36 ( .A(n63), .B(localRouterAddress[5]), .Y(n38) );
  INVXLTS U37 ( .A(destinationAddressIn[9]), .Y(n59) );
  INVXLTS U38 ( .A(localRouterAddress[0]), .Y(n64) );
endmodule


module incomingPortHandler_2 ( clk, reset, localRouterAddress, 
        destinationAddressIn, requesterAddressIn, readIn, writeIn, 
        outputPortSelect, memRead, memWrite );
  input [5:0] localRouterAddress;
  input [13:0] destinationAddressIn;
  input [5:0] requesterAddressIn;
  output [3:0] outputPortSelect;
  input clk, reset, readIn, writeIn;
  output memRead, memWrite;
  wire   n69, n45, n44, n43, n42, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68;

  DFFQX1TS memRead_reg ( .D(n67), .CK(clk), .Q(memRead) );
  DFFQX1TS \outputPortSelect_reg[0]  ( .D(n42), .CK(clk), .Q(
        outputPortSelect[0]) );
  DFFQX1TS \outputPortSelect_reg[1]  ( .D(n43), .CK(clk), .Q(
        outputPortSelect[1]) );
  DFFQX4TS \outputPortSelect_reg[2]  ( .D(n44), .CK(clk), .Q(
        outputPortSelect[2]) );
  DFFQX4TS \outputPortSelect_reg[3]  ( .D(n45), .CK(clk), .Q(
        outputPortSelect[3]) );
  DFFQX1TS memWrite_reg ( .D(n68), .CK(clk), .Q(n69) );
  OAI211X1TS U1 ( .A0(localRouterAddress[4]), .A1(n61), .B0(n60), .C0(
        localRouterAddress[3]), .Y(n38) );
  CLKBUFX2TS U2 ( .A(n69), .Y(memWrite) );
  NAND2XLTS U3 ( .A(localRouterAddress[5]), .B(n62), .Y(n41) );
  INVXLTS U4 ( .A(destinationAddressIn[13]), .Y(n62) );
  NOR3BXLTS U5 ( .AN(n33), .B(writeIn), .C(readIn), .Y(n56) );
  NAND2XLTS U6 ( .A(localRouterAddress[2]), .B(n59), .Y(n51) );
  AOI2BB2XLTS U7 ( .B0(n58), .B1(localRouterAddress[1]), .A0N(
        destinationAddressIn[8]), .A1N(n63), .Y(n53) );
  INVX2TS U8 ( .A(reset), .Y(n33) );
  NOR2BX1TS U9 ( .AN(n55), .B(n54), .Y(n45) );
  NOR2X1TS U10 ( .A(n54), .B(n55), .Y(n44) );
  INVX2TS U11 ( .A(n48), .Y(n66) );
  OAI21X1TS U12 ( .A0(n53), .A1(n52), .B0(n51), .Y(n55) );
  NAND3BX1TS U13 ( .AN(n50), .B(n49), .C(n48), .Y(n54) );
  OAI22XLTS U14 ( .A0(localRouterAddress[1]), .A1(n58), .B0(
        localRouterAddress[2]), .B1(n59), .Y(n52) );
  AOI2BB1XLTS U15 ( .A0N(localRouterAddress[4]), .A1N(n61), .B0(n37), .Y(n47)
         );
  OAI21XLTS U16 ( .A0(readIn), .A1(writeIn), .B0(n33), .Y(n50) );
  NAND3X1TS U17 ( .A(n53), .B(n49), .C(n35), .Y(n48) );
  AOI211XLTS U18 ( .A0(destinationAddressIn[8]), .A1(n63), .B0(n52), .C0(n64), 
        .Y(n35) );
  INVX2TS U19 ( .A(n51), .Y(n64) );
  AND4X1TS U20 ( .A(n34), .B(n47), .C(n40), .D(n41), .Y(n49) );
  XNOR2XLTS U21 ( .A(destinationAddressIn[11]), .B(localRouterAddress[3]), .Y(
        n34) );
  INVXLTS U22 ( .A(destinationAddressIn[10]), .Y(n59) );
  AOI211X1TS U23 ( .A0(n39), .A1(n38), .B0(n50), .C0(n37), .Y(n42) );
  AND2X2TS U24 ( .A(n40), .B(n41), .Y(n39) );
  INVXLTS U25 ( .A(destinationAddressIn[11]), .Y(n60) );
  AOI211X1TS U26 ( .A0(n47), .A1(n46), .B0(n50), .C0(n65), .Y(n43) );
  INVX2TS U27 ( .A(n41), .Y(n65) );
  NAND3BXLTS U28 ( .AN(localRouterAddress[3]), .B(n40), .C(
        destinationAddressIn[11]), .Y(n46) );
  INVXLTS U29 ( .A(destinationAddressIn[12]), .Y(n61) );
  INVX2TS U30 ( .A(n57), .Y(n67) );
  AOI32XLTS U31 ( .A0(n66), .A1(n33), .A2(readIn), .B0(memRead), .B1(n56), .Y(
        n57) );
  INVX2TS U32 ( .A(n36), .Y(n68) );
  AOI32XLTS U33 ( .A0(n66), .A1(n33), .A2(writeIn), .B0(n69), .B1(n56), .Y(n36) );
  NAND2XLTS U34 ( .A(localRouterAddress[4]), .B(n61), .Y(n40) );
  NOR2XLTS U35 ( .A(n62), .B(localRouterAddress[5]), .Y(n37) );
  INVXLTS U36 ( .A(destinationAddressIn[9]), .Y(n58) );
  INVXLTS U37 ( .A(localRouterAddress[0]), .Y(n63) );
endmodule


module incomingPortHandler_3 ( clk, reset, localRouterAddress, 
        destinationAddressIn, requesterAddressIn, readIn, writeIn, 
        outputPortSelect, memRead, memWrite );
  input [5:0] localRouterAddress;
  input [13:0] destinationAddressIn;
  input [5:0] requesterAddressIn;
  output [3:0] outputPortSelect;
  input clk, reset, readIn, writeIn;
  output memRead, memWrite;
  wire   n45, n44, n43, n42, n3, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67;

  DFFQX1TS memWrite_reg ( .D(n67), .CK(clk), .Q(memWrite) );
  DFFQX1TS memRead_reg ( .D(n66), .CK(clk), .Q(memRead) );
  DFFQX1TS \outputPortSelect_reg[2]  ( .D(n44), .CK(clk), .Q(
        outputPortSelect[2]) );
  DFFHQX1TS \outputPortSelect_reg[0]  ( .D(n42), .CK(clk), .Q(
        outputPortSelect[0]) );
  DFFQX4TS \outputPortSelect_reg[1]  ( .D(n43), .CK(clk), .Q(
        outputPortSelect[1]) );
  DFFHQX1TS \outputPortSelect_reg[3]  ( .D(n45), .CK(clk), .Q(
        outputPortSelect[3]) );
  OAI211X1TS U1 ( .A0(localRouterAddress[4]), .A1(n60), .B0(n59), .C0(
        localRouterAddress[3]), .Y(n37) );
  NAND2XLTS U2 ( .A(localRouterAddress[5]), .B(n61), .Y(n40) );
  INVXLTS U3 ( .A(destinationAddressIn[13]), .Y(n61) );
  NOR3BXLTS U4 ( .AN(n3), .B(writeIn), .C(readIn), .Y(n55) );
  NAND2XLTS U5 ( .A(localRouterAddress[2]), .B(n58), .Y(n50) );
  AOI2BB2XLTS U6 ( .B0(n57), .B1(localRouterAddress[1]), .A0N(
        destinationAddressIn[8]), .A1N(n62), .Y(n52) );
  INVX2TS U7 ( .A(reset), .Y(n3) );
  NOR2BX1TS U8 ( .AN(n54), .B(n53), .Y(n45) );
  NOR2X1TS U9 ( .A(n53), .B(n54), .Y(n44) );
  INVX2TS U10 ( .A(n47), .Y(n65) );
  OAI21X1TS U11 ( .A0(n52), .A1(n51), .B0(n50), .Y(n54) );
  NAND3BX1TS U12 ( .AN(n49), .B(n48), .C(n47), .Y(n53) );
  OAI22XLTS U13 ( .A0(localRouterAddress[1]), .A1(n57), .B0(
        localRouterAddress[2]), .B1(n58), .Y(n51) );
  AOI2BB1XLTS U14 ( .A0N(localRouterAddress[4]), .A1N(n60), .B0(n36), .Y(n46)
         );
  OAI21XLTS U15 ( .A0(readIn), .A1(writeIn), .B0(n3), .Y(n49) );
  NAND3X1TS U16 ( .A(n52), .B(n48), .C(n34), .Y(n47) );
  AOI211XLTS U17 ( .A0(destinationAddressIn[8]), .A1(n62), .B0(n51), .C0(n63), 
        .Y(n34) );
  INVX2TS U18 ( .A(n50), .Y(n63) );
  AND4X1TS U19 ( .A(n33), .B(n46), .C(n39), .D(n40), .Y(n48) );
  XNOR2XLTS U20 ( .A(destinationAddressIn[11]), .B(localRouterAddress[3]), .Y(
        n33) );
  INVXLTS U21 ( .A(destinationAddressIn[10]), .Y(n58) );
  AOI211X1TS U22 ( .A0(n38), .A1(n37), .B0(n49), .C0(n36), .Y(n42) );
  AND2X2TS U23 ( .A(n39), .B(n40), .Y(n38) );
  INVXLTS U24 ( .A(destinationAddressIn[11]), .Y(n59) );
  AOI211X1TS U25 ( .A0(n46), .A1(n41), .B0(n49), .C0(n64), .Y(n43) );
  INVX2TS U26 ( .A(n40), .Y(n64) );
  NAND3BXLTS U27 ( .AN(localRouterAddress[3]), .B(n39), .C(
        destinationAddressIn[11]), .Y(n41) );
  INVXLTS U28 ( .A(destinationAddressIn[12]), .Y(n60) );
  INVX2TS U29 ( .A(n56), .Y(n66) );
  AOI32XLTS U30 ( .A0(n65), .A1(n3), .A2(readIn), .B0(memRead), .B1(n55), .Y(
        n56) );
  INVX2TS U31 ( .A(n35), .Y(n67) );
  AOI32XLTS U32 ( .A0(n65), .A1(n3), .A2(writeIn), .B0(memWrite), .B1(n55), 
        .Y(n35) );
  NAND2XLTS U33 ( .A(localRouterAddress[4]), .B(n60), .Y(n39) );
  NOR2XLTS U34 ( .A(n61), .B(localRouterAddress[5]), .Y(n36) );
  INVXLTS U35 ( .A(destinationAddressIn[9]), .Y(n57) );
  INVXLTS U36 ( .A(localRouterAddress[0]), .Y(n62) );
endmodule


module outputPortArbiter_1 ( clk, reset, selectBit_NORTH, 
        destinationAddressIn_NORTH, requesterAddressIn_NORTH, readIn_NORTH, 
        writeIn_NORTH, dataIn_NORTH, selectBit_SOUTH, 
        destinationAddressIn_SOUTH, requesterAddressIn_SOUTH, readIn_SOUTH, 
        writeIn_SOUTH, dataIn_SOUTH, selectBit_EAST, destinationAddressIn_EAST, 
        requesterAddressIn_EAST, readIn_EAST, writeIn_EAST, dataIn_EAST, 
        selectBit_WEST, destinationAddressIn_WEST, requesterAddressIn_WEST, 
        readIn_WEST, writeIn_WEST, dataIn_WEST, readReady, 
        readRequesterAddress, cacheDataOut, destinationAddressOut, 
        requesterAddressOut, readOut, writeOut, dataOut );
  input [13:0] destinationAddressIn_NORTH;
  input [5:0] requesterAddressIn_NORTH;
  input [31:0] dataIn_NORTH;
  input [13:0] destinationAddressIn_SOUTH;
  input [5:0] requesterAddressIn_SOUTH;
  input [31:0] dataIn_SOUTH;
  input [13:0] destinationAddressIn_EAST;
  input [5:0] requesterAddressIn_EAST;
  input [31:0] dataIn_EAST;
  input [13:0] destinationAddressIn_WEST;
  input [5:0] requesterAddressIn_WEST;
  input [31:0] dataIn_WEST;
  input [5:0] readRequesterAddress;
  input [31:0] cacheDataOut;
  output [13:0] destinationAddressOut;
  output [5:0] requesterAddressOut;
  output [31:0] dataOut;
  input clk, reset, selectBit_NORTH, readIn_NORTH, writeIn_NORTH,
         selectBit_SOUTH, readIn_SOUTH, writeIn_SOUTH, selectBit_EAST,
         readIn_EAST, writeIn_EAST, selectBit_WEST, readIn_WEST, writeIn_WEST,
         readReady;
  output readOut, writeOut;
  wire   N4718, n2888, n5327, n2886, n5326, n2889, n2883, n2887, n5323, n2569,
         n2567, n2566, n2578, n2638, n2624, n2617, n2577, n2544, n2541, n2540,
         n2537, n2535, n2703, n2692, n2691, n2689, n2511, n2507, n2731, n2574,
         n2499, n2496, n2493, n2770, n2768, n2764, n2754, n2748, n2746, n2739,
         n2486, n2484, n2482, n2480, n2802, n2834, n2833, n2832, n2829, n2825,
         n2814, n2811, n2807, n2806, n2457, n2455, n2453, n2570, n2565, n2573,
         n2568, n2564, n2563, n2575, n2882, n2881, n2879, n2610, n2609, n2608,
         n2607, n2606, n2605, n2604, n2603, n2602, n2601, n2600, n2599, n2598,
         n2597, n2596, n2595, n2594, n2593, n2592, n2591, n2590, n2589, n2588,
         n2587, n2586, n2585, n2584, n2583, n2582, n2581, n2580, n2579, n2561,
         n2560, n2559, n2557, n2556, n2555, n2554, n2552, n2551, n2550, n2549,
         n2642, n2640, n2639, n2637, n2635, n2634, n2633, n2631, n2628, n2627,
         n2626, n2625, n2623, n2620, n2618, n2616, n2615, n2614, n2612, n2611,
         n2870, n2869, n2868, n2867, n2866, n2865, n2674, n2672, n2671, n2670,
         n2669, n2668, n2667, n2666, n2665, n2664, n2662, n2661, n2660, n2657,
         n2656, n2655, n2654, n2653, n2652, n2651, n2650, n2649, n2648, n2647,
         n2646, n2645, n2644, n2576, n2534, n2533, n2532, n2531, n2530, n2529,
         n2528, n2527, n2526, n2525, n2524, n2523, n2522, n2521, n2860, n2859,
         n2706, n2705, n2700, n2698, n2696, n2695, n2694, n2690, n2687, n2686,
         n2685, n2684, n2677, n2675, n2736, n2734, n2733, n2725, n2723, n2720,
         n2718, n2715, n2713, n2504, n2498, n2497, n2494, n2850,
         \requesterAddressbuffer[2][2] , n2849, \requesterAddressbuffer[2][3] ,
         n2847, \requesterAddressbuffer[2][5] , n2769, n2760, n2743, n2492,
         n2491, n2489, n2488, n2487, n2485, n2483, n2481, n2846, n2845, n2844,
         n2843, n2842, n2841, n2801, n2799, n2798, n2796, n2795, n2793, n2791,
         n2790, n2789, n2788, n2787, n2786, n2785, n2784, n2781, n2779, n2778,
         n2777, n2776, n2774, n2773, n2772, n2771, n2572, n2478, n2477, n2476,
         n2475, n2474, n2473, n2472, n2471, n2470, n2469, n2468, n2467, n2466,
         n2465, n2840, \requesterAddressbuffer[0][0] , n2839,
         \requesterAddressbuffer[0][1] , n2838, \requesterAddressbuffer[0][2] ,
         n2836, \requesterAddressbuffer[0][4] , n2571, n2464, n2460, n2458,
         n2454, n2451, n2880, n2878, n2877, n2562, n2558, n2553, n2876,
         \requesterAddressbuffer[6][0] , n2875, \requesterAddressbuffer[6][1] ,
         n2874, \requesterAddressbuffer[6][2] , n2873,
         \requesterAddressbuffer[6][3] , n2872, \requesterAddressbuffer[6][4] ,
         n2871, \requesterAddressbuffer[6][5] , n2641, n2636, n2632, n2630,
         n2629, n2622, n2621, n2619, n2613, n2548, n2547, n2546, n2545, n2543,
         n2542, n2539, n2538, n2536, n2673, n2663, n2659, n2658, n2643, n2864,
         n2863, n2862, n2861, n2704, n2702, n2701, n2699, n2697, n2693, n2688,
         n2683, n2682, n2681, n2680, n2679, n2678, n2676, n2520, n2519, n2518,
         n2517, n2516, n2515, n2514, n2513, n2512, n2510, n2509, n2508, n2858,
         \requesterAddressbuffer[3][0] , n2857, \requesterAddressbuffer[3][1] ,
         n2856, \requesterAddressbuffer[3][2] , n2855,
         \requesterAddressbuffer[3][3] , n2854, \requesterAddressbuffer[3][4] ,
         n2853, \requesterAddressbuffer[3][5] , n2738, n2737, n2735, n2732,
         n2730, n2729, n2728, n2727, n2726, n2724, n2722, n2721, n2719, n2717,
         n2716, n2714, n2712, n2711, n2710, n2709, n2708, n2707, n2506, n2505,
         n2503, n2502, n2501, n2500, n2495, n2852,
         \requesterAddressbuffer[2][0] , n2851, \requesterAddressbuffer[2][1] ,
         n2848, \requesterAddressbuffer[2][4] , n2767, n2766, n2765, n2763,
         n2762, n2761, n2759, n2758, n2757, n2756, n2755, n2753, n2752, n2751,
         n2750, n2749, n2747, n2745, n2744, n2742, n2741, n2740, n2490, n2479,
         n2800, n2797, n2794, n2792, n2783, n2782, n2780, n2775, n2837,
         \requesterAddressbuffer[0][3] , n2835, \requesterAddressbuffer[0][5] ,
         n2831, n2830, n2828, n2827, n2826, n2824, n2823, n2822, n2821, n2820,
         n2819, n2818, n2817, n2816, n2815, n2813, n2812, n2810, n2809, n2808,
         n2805, n2804, n2803, n2463, n2462, n2461, n2459, n2456, n2452, n2885,
         n2449, n2434, n2431, n2450, n2448, n2447, n2446, n2445, n2444, n2443,
         n2442, n2441, n2440, n2439, n2438, n2437, n2436, n2435, n2433, n2432,
         n2430, n2429, n2428, n2427, n2426, n2425, n2424, n2423, n2422, n2421,
         n2420, n2419, n2418, n2417, n2416, n2415, n2414, n2413, n2412, n2411,
         n2410, n2409, n2408, n2407, n2406, n2405, n2404, n2403, n2402, n2401,
         n2400, n2399, n2398, n2397, n2884, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n501, n503, n505, n507, n508, n509, n510, n511, n512, n514,
         n515, n516, n526, n531, n536, n537, n541, n543, n544, n545, n546,
         n548, n551, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n621,
         n622, n623, n624, n625, n626, n627, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n711, n712, n714, n715, n716,
         n728, n729, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n886, n919, n936, n955,
         n957, n959, n970, n986, n1402, n1533, n1535, n1571, n1598, n1602,
         n1653, n1654, n1728, n1797, n1817, n1822, n1894, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5324, n5325,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311;
  wire   [0:7] readOutbuffer;
  wire   [0:7] writeOutbuffer;

  DFFNSRX2TS \destinationAddressbuffer_reg[2][6]  ( .D(n2486), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4839) );
  DFFNSRX2TS \destinationAddressbuffer_reg[2][8]  ( .D(n2484), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4819) );
  DFFNSRX2TS \destinationAddressbuffer_reg[2][10]  ( .D(n2482), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4805) );
  DFFNSRX2TS \destinationAddressbuffer_reg[2][12]  ( .D(n2480), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4791) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][7]  ( .D(n2457), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4827) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][9]  ( .D(n2455), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4811) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][11]  ( .D(n2453), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4797) );
  DFFNSRX2TS \destinationAddressbuffer_reg[2][7]  ( .D(n2485), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4832) );
  DFFNSRX2TS \destinationAddressbuffer_reg[2][9]  ( .D(n2483), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4816) );
  DFFNSRX2TS \destinationAddressbuffer_reg[2][11]  ( .D(n2481), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4800) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][6]  ( .D(n2458), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4840) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][10]  ( .D(n2454), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4806) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][13]  ( .D(n2451), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4784) );
  DFFNSRX2TS \destinationAddressbuffer_reg[2][13]  ( .D(n2479), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4777) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][8]  ( .D(n2456), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4817) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][12]  ( .D(n2452), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4785) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][7]  ( .D(n2499), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4831) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][10]  ( .D(n2496), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4807) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][13]  ( .D(n2493), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4781) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][8]  ( .D(n2498), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4824) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][9]  ( .D(n2497), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4810) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][12]  ( .D(n2494), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4788) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][6]  ( .D(n2500), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4835) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][11]  ( .D(n2495), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4795) );
  DFFNSRX2TS \destinationAddressbuffer_reg[6][7]  ( .D(n2541), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4829) );
  DFFNSRX2TS \destinationAddressbuffer_reg[6][8]  ( .D(n2540), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4823) );
  DFFNSRX2TS \destinationAddressbuffer_reg[6][11]  ( .D(n2537), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4799) );
  DFFNSRX2TS \destinationAddressbuffer_reg[6][13]  ( .D(n2535), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4779) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][9]  ( .D(n2511), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4815) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][13]  ( .D(n2507), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4783) );
  DFFNSRX2TS \destinationAddressbuffer_reg[7][6]  ( .D(n2556), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4836) );
  DFFNSRX2TS \destinationAddressbuffer_reg[7][7]  ( .D(n2555), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4830) );
  DFFNSRX2TS \destinationAddressbuffer_reg[7][8]  ( .D(n2554), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4820) );
  DFFNSRX2TS \destinationAddressbuffer_reg[7][10]  ( .D(n2552), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n567), .QN(n4804) );
  DFFNSRX2TS \destinationAddressbuffer_reg[7][11]  ( .D(n2551), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4794) );
  DFFNSRX2TS \destinationAddressbuffer_reg[7][12]  ( .D(n2550), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4790) );
  DFFNSRX2TS \destinationAddressbuffer_reg[7][13]  ( .D(n2549), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4780) );
  DFFNSRX2TS \destinationAddressbuffer_reg[1][6]  ( .D(n2472), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4838) );
  DFFNSRX2TS \destinationAddressbuffer_reg[1][7]  ( .D(n2471), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4826) );
  DFFNSRX2TS \destinationAddressbuffer_reg[1][8]  ( .D(n2470), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4818) );
  DFFNSRX2TS \destinationAddressbuffer_reg[1][9]  ( .D(n2469), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4814) );
  DFFNSRX2TS \destinationAddressbuffer_reg[1][10]  ( .D(n2468), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4802) );
  DFFNSRX2TS \destinationAddressbuffer_reg[1][11]  ( .D(n2467), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4796) );
  DFFNSRX2TS \destinationAddressbuffer_reg[1][12]  ( .D(n2466), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4786) );
  DFFNSRX2TS \destinationAddressbuffer_reg[1][13]  ( .D(n2465), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4778) );
  DFFNSRX2TS \destinationAddressbuffer_reg[7][9]  ( .D(n2553), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4813) );
  DFFNSRX2TS \destinationAddressbuffer_reg[6][6]  ( .D(n2542), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4833) );
  DFFNSRX2TS \destinationAddressbuffer_reg[6][9]  ( .D(n2539), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4809) );
  DFFNSRX2TS \destinationAddressbuffer_reg[6][10]  ( .D(n2538), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4801) );
  DFFNSRX2TS \destinationAddressbuffer_reg[6][12]  ( .D(n2536), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4789) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][10]  ( .D(n2510), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4803) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][11]  ( .D(n2509), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4793) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][12]  ( .D(n2508), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4787) );
  DFFNSRX2TS \dataoutbuffer_reg[6][4]  ( .D(n2638), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4681) );
  DFFNSRX2TS \dataoutbuffer_reg[6][18]  ( .D(n2624), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4555) );
  DFFNSRX2TS \dataoutbuffer_reg[6][25]  ( .D(n2617), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4492) );
  DFFNSRX2TS \dataoutbuffer_reg[7][0]  ( .D(n2610), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4712) );
  DFFNSRX2TS \dataoutbuffer_reg[7][1]  ( .D(n2609), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4707) );
  DFFNSRX2TS \dataoutbuffer_reg[7][2]  ( .D(n2608), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4694) );
  DFFNSRX2TS \dataoutbuffer_reg[7][3]  ( .D(n2607), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4689) );
  DFFNSRX2TS \dataoutbuffer_reg[7][4]  ( .D(n2606), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4676) );
  DFFNSRX2TS \dataoutbuffer_reg[7][5]  ( .D(n2605), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4667) );
  DFFNSRX2TS \dataoutbuffer_reg[7][6]  ( .D(n2604), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4664) );
  DFFNSRX2TS \dataoutbuffer_reg[7][7]  ( .D(n2603), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4649) );
  DFFNSRX2TS \dataoutbuffer_reg[7][8]  ( .D(n2602), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4642) );
  DFFNSRX2TS \dataoutbuffer_reg[7][9]  ( .D(n2601), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4637) );
  DFFNSRX2TS \dataoutbuffer_reg[7][10]  ( .D(n2600), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4628) );
  DFFNSRX2TS \dataoutbuffer_reg[7][11]  ( .D(n2599), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4615) );
  DFFNSRX2TS \dataoutbuffer_reg[7][12]  ( .D(n2598), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4604) );
  DFFNSRX2TS \dataoutbuffer_reg[7][13]  ( .D(n2597), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4595) );
  DFFNSRX2TS \dataoutbuffer_reg[7][14]  ( .D(n2596), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4592) );
  DFFNSRX2TS \dataoutbuffer_reg[7][15]  ( .D(n2595), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4577) );
  DFFNSRX2TS \dataoutbuffer_reg[7][16]  ( .D(n2594), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4572) );
  DFFNSRX2TS \dataoutbuffer_reg[7][17]  ( .D(n2593), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4561) );
  DFFNSRX2TS \dataoutbuffer_reg[7][18]  ( .D(n2592), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4550) );
  DFFNSRX2TS \dataoutbuffer_reg[7][19]  ( .D(n2591), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4547) );
  DFFNSRX2TS \dataoutbuffer_reg[7][20]  ( .D(n2590), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4534) );
  DFFNSRX2TS \dataoutbuffer_reg[7][21]  ( .D(n2589), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4529) );
  DFFNSRX2TS \dataoutbuffer_reg[7][22]  ( .D(n2588), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4514) );
  DFFNSRX2TS \dataoutbuffer_reg[7][23]  ( .D(n2587), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4509) );
  DFFNSRX2TS \dataoutbuffer_reg[7][24]  ( .D(n2586), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4498) );
  DFFNSRX2TS \dataoutbuffer_reg[7][25]  ( .D(n2585), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4489) );
  DFFNSRX2TS \dataoutbuffer_reg[7][26]  ( .D(n2584), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4480) );
  DFFNSRX2TS \dataoutbuffer_reg[7][27]  ( .D(n2583), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4473) );
  DFFNSRX2TS \dataoutbuffer_reg[7][28]  ( .D(n2582), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4464) );
  DFFNSRX2TS \dataoutbuffer_reg[7][29]  ( .D(n2581), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4451) );
  DFFNSRX2TS \dataoutbuffer_reg[7][30]  ( .D(n2580), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4442) );
  DFFNSRX2TS \dataoutbuffer_reg[7][31]  ( .D(n2579), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4437) );
  DFFNSRX2TS \destinationAddressbuffer_reg[7][1]  ( .D(n2561), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4761) );
  DFFNSRX2TS \destinationAddressbuffer_reg[7][2]  ( .D(n2560), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4754) );
  DFFNSRX2TS \destinationAddressbuffer_reg[7][3]  ( .D(n2559), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4743) );
  DFFNSRX2TS \destinationAddressbuffer_reg[7][5]  ( .D(n2557), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4731) );
  DFFNSRX2TS \dataoutbuffer_reg[6][0]  ( .D(n2642), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4716) );
  DFFNSRX2TS \dataoutbuffer_reg[6][2]  ( .D(n2640), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4700) );
  DFFNSRX2TS \dataoutbuffer_reg[6][3]  ( .D(n2639), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4685) );
  DFFNSRX2TS \dataoutbuffer_reg[6][5]  ( .D(n2637), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4669) );
  DFFNSRX2TS \dataoutbuffer_reg[6][7]  ( .D(n2635), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4651) );
  DFFNSRX2TS \dataoutbuffer_reg[6][8]  ( .D(n2634), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4646) );
  DFFNSRX2TS \dataoutbuffer_reg[6][9]  ( .D(n2633), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4635) );
  DFFNSRX2TS \dataoutbuffer_reg[6][11]  ( .D(n2631), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4619) );
  DFFNSRX2TS \dataoutbuffer_reg[6][14]  ( .D(n2628), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4590) );
  DFFNSRX2TS \dataoutbuffer_reg[6][15]  ( .D(n2627), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4583) );
  DFFNSRX2TS \dataoutbuffer_reg[6][16]  ( .D(n2626), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4570) );
  DFFNSRX2TS \dataoutbuffer_reg[6][17]  ( .D(n2625), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4565) );
  DFFNSRX2TS \dataoutbuffer_reg[6][19]  ( .D(n2623), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4543) );
  DFFNSRX2TS \dataoutbuffer_reg[6][22]  ( .D(n2620), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4520) );
  DFFNSRX2TS \dataoutbuffer_reg[6][24]  ( .D(n2618), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4502) );
  DFFNSRX2TS \dataoutbuffer_reg[6][26]  ( .D(n2616), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4482) );
  DFFNSRX2TS \dataoutbuffer_reg[6][27]  ( .D(n2615), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4471) );
  DFFNSRX2TS \dataoutbuffer_reg[6][28]  ( .D(n2614), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4462) );
  DFFNSRX2TS \dataoutbuffer_reg[6][30]  ( .D(n2612), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4446) );
  DFFNSRX2TS \dataoutbuffer_reg[6][31]  ( .D(n2611), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4435) );
  DFFNSRX2TS \destinationAddressbuffer_reg[7][0]  ( .D(n2562), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4775) );
  DFFNSRX2TS \destinationAddressbuffer_reg[7][4]  ( .D(n2558), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4733) );
  DFFNSRX2TS \dataoutbuffer_reg[6][1]  ( .D(n2641), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4704) );
  DFFNSRX2TS \dataoutbuffer_reg[6][6]  ( .D(n2636), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4657) );
  DFFNSRX2TS \dataoutbuffer_reg[6][10]  ( .D(n2632), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4621) );
  DFFNSRX2TS \dataoutbuffer_reg[6][12]  ( .D(n2630), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4609) );
  DFFNSRX2TS \dataoutbuffer_reg[6][13]  ( .D(n2629), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4598) );
  DFFNSRX2TS \dataoutbuffer_reg[6][20]  ( .D(n2622), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4531) );
  DFFNSRX2TS \dataoutbuffer_reg[6][21]  ( .D(n2621), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4524) );
  DFFNSRX2TS \dataoutbuffer_reg[6][23]  ( .D(n2619), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4504) );
  DFFNSRX2TS \dataoutbuffer_reg[6][29]  ( .D(n2613), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4454) );
  DFFNSRX2TS \destinationAddressbuffer_reg[6][5]  ( .D(n2543), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4728) );
  DFFNSRX2TS \requesterAddressbuffer_reg[2][2]  ( .D(n2850), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][2] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[2][3]  ( .D(n2849), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][3] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[2][5]  ( .D(n2847), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][5] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[0][0]  ( .D(n2840), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][0] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[0][1]  ( .D(n2839), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][1] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[0][2]  ( .D(n2838), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][2] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[0][4]  ( .D(n2836), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][4] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[2][0]  ( .D(n2852), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][0] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[2][1]  ( .D(n2851), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][1] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[2][4]  ( .D(n2848), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][4] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[0][3]  ( .D(n2837), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][3] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[0][5]  ( .D(n2835), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][5] ) );
  DFFNSRX2TS \readOutbuffer_reg[3]  ( .D(n2566), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[3]) );
  DFFNSRX2TS \readOutbuffer_reg[6]  ( .D(n2569), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n19) );
  DFFNSRX2TS \writeOutbuffer_reg[7]  ( .D(n2578), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n24) );
  DFFNSRX2TS \readOutbuffer_reg[5]  ( .D(n2568), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n32) );
  DFFNSRX2TS \readOutbuffer_reg[1]  ( .D(n2564), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n25) );
  DFFNSRX2TS \readOutbuffer_reg[0]  ( .D(n2563), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n33) );
  DFFNSRX2TS \requesterAddressbuffer_reg[7][0]  ( .D(n2882), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n31) );
  DFFNSRX2TS \requesterAddressbuffer_reg[7][1]  ( .D(n2881), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n29) );
  DFFNSRX2TS \requesterAddressbuffer_reg[7][3]  ( .D(n2879), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n30) );
  DFFNSRX2TS \requesterAddressbuffer_reg[7][2]  ( .D(n2880), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n28) );
  DFFNSRX2TS \requesterAddressbuffer_reg[7][4]  ( .D(n2878), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n27) );
  DFFNSRX2TS \requesterAddressbuffer_reg[7][5]  ( .D(n2877), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n26) );
  DFFNSRX2TS \writeOutbuffer_reg[1]  ( .D(n2572), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[1]), .QN(n151) );
  DFFNSRX2TS \writeOutbuffer_reg[2]  ( .D(n2573), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[2]), .QN(n154) );
  DFFNSRX2TS \dataoutbuffer_reg[3][7]  ( .D(n2731), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n109), .QN(n4654) );
  DFFNSRX2TS \dataoutbuffer_reg[2][2]  ( .D(n2768), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n146), .QN(n4697) );
  DFFNSRX2TS \dataoutbuffer_reg[2][16]  ( .D(n2754), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n144), .QN(n4573) );
  DFFNSRX2TS \dataoutbuffer_reg[2][22]  ( .D(n2748), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n143), .QN(n4519) );
  DFFNSRX2TS \dataoutbuffer_reg[2][24]  ( .D(n2746), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n142), .QN(n4501) );
  DFFNSRX2TS \dataoutbuffer_reg[2][31]  ( .D(n2739), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n141), .QN(n4438) );
  DFFNSRX2TS \dataoutbuffer_reg[0][0]  ( .D(n2834), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n108), .QN(n4715) );
  DFFNSRX2TS \dataoutbuffer_reg[0][1]  ( .D(n2833), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n107), .QN(n4708) );
  DFFNSRX2TS \dataoutbuffer_reg[0][2]  ( .D(n2832), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n106), .QN(n4699) );
  DFFNSRX2TS \dataoutbuffer_reg[0][5]  ( .D(n2829), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n105), .QN(n4672) );
  DFFNSRX2TS \dataoutbuffer_reg[0][9]  ( .D(n2825), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n104), .QN(n4636) );
  DFFNSRX2TS \dataoutbuffer_reg[0][20]  ( .D(n2814), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n103), .QN(n4537) );
  DFFNSRX2TS \dataoutbuffer_reg[0][23]  ( .D(n2811), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n102), .QN(n4510) );
  DFFNSRX2TS \dataoutbuffer_reg[0][27]  ( .D(n2807), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n101), .QN(n4474) );
  DFFNSRX2TS \dataoutbuffer_reg[0][28]  ( .D(n2806), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n100), .QN(n4465) );
  DFFNSRX2TS \dataoutbuffer_reg[3][2]  ( .D(n2736), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n99), .QN(n4698) );
  DFFNSRX2TS \dataoutbuffer_reg[3][4]  ( .D(n2734), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n98), .QN(n4678) );
  DFFNSRX2TS \dataoutbuffer_reg[3][5]  ( .D(n2733), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n97), .QN(n4671) );
  DFFNSRX2TS \dataoutbuffer_reg[3][13]  ( .D(n2725), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n96), .QN(n4597) );
  DFFNSRX2TS \dataoutbuffer_reg[3][15]  ( .D(n2723), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n95), .QN(n4579) );
  DFFNSRX2TS \dataoutbuffer_reg[3][18]  ( .D(n2720), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n94), .QN(n4554) );
  DFFNSRX2TS \dataoutbuffer_reg[3][20]  ( .D(n2718), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n93), .QN(n4538) );
  DFFNSRX2TS \dataoutbuffer_reg[3][23]  ( .D(n2715), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n92), .QN(n4511) );
  DFFNSRX2TS \dataoutbuffer_reg[3][25]  ( .D(n2713), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n91), .QN(n4487) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][2]  ( .D(n2504), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n90), .QN(n4752) );
  DFFNSRX2TS \destinationAddressbuffer_reg[2][0]  ( .D(n2492), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n137), .QN(n4770) );
  DFFNSRX2TS \destinationAddressbuffer_reg[2][1]  ( .D(n2491), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n136), .QN(n4763) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][0]  ( .D(n2464), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n89), .QN(n4774) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][4]  ( .D(n2460), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n88), .QN(n4736) );
  DFFNSRX2TS \dataoutbuffer_reg[3][0]  ( .D(n2738), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n87), .QN(n4711) );
  DFFNSRX2TS \dataoutbuffer_reg[3][1]  ( .D(n2737), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n86), .QN(n4702) );
  DFFNSRX2TS \dataoutbuffer_reg[3][3]  ( .D(n2735), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n85), .QN(n4688) );
  DFFNSRX2TS \dataoutbuffer_reg[3][6]  ( .D(n2732), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n84), .QN(n4661) );
  DFFNSRX2TS \dataoutbuffer_reg[3][8]  ( .D(n2730), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n83), .QN(n4639) );
  DFFNSRX2TS \dataoutbuffer_reg[3][9]  ( .D(n2729), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n82), .QN(n4632) );
  DFFNSRX2TS \dataoutbuffer_reg[3][10]  ( .D(n2728), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n81), .QN(n4623) );
  DFFNSRX2TS \dataoutbuffer_reg[3][11]  ( .D(n2727), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n80), .QN(n4616) );
  DFFNSRX2TS \dataoutbuffer_reg[3][12]  ( .D(n2726), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n79), .QN(n4605) );
  DFFNSRX2TS \dataoutbuffer_reg[3][14]  ( .D(n2724), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n78), .QN(n4589) );
  DFFNSRX2TS \dataoutbuffer_reg[3][16]  ( .D(n2722), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n77), .QN(n4567) );
  DFFNSRX2TS \dataoutbuffer_reg[3][17]  ( .D(n2721), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n76), .QN(n4558) );
  DFFNSRX2TS \dataoutbuffer_reg[3][19]  ( .D(n2719), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n75), .QN(n4546) );
  DFFNSRX2TS \dataoutbuffer_reg[3][21]  ( .D(n2717), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n74), .QN(n4526) );
  DFFNSRX2TS \dataoutbuffer_reg[3][22]  ( .D(n2716), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n73), .QN(n4515) );
  DFFNSRX2TS \dataoutbuffer_reg[3][24]  ( .D(n2714), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n72), .QN(n4499) );
  DFFNSRX2TS \dataoutbuffer_reg[3][26]  ( .D(n2712), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n71), .QN(n4483) );
  DFFNSRX2TS \dataoutbuffer_reg[3][27]  ( .D(n2711), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n70), .QN(n4472) );
  DFFNSRX2TS \dataoutbuffer_reg[3][28]  ( .D(n2710), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n69), .QN(n4463) );
  DFFNSRX2TS \dataoutbuffer_reg[3][29]  ( .D(n2709), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n68), .QN(n4452) );
  DFFNSRX2TS \dataoutbuffer_reg[3][30]  ( .D(n2708), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n67), .QN(n4447) );
  DFFNSRX2TS \dataoutbuffer_reg[3][31]  ( .D(n2707), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n66), .QN(n4434) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][0]  ( .D(n2506), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n65), .QN(n4773) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][1]  ( .D(n2505), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n64), .QN(n4766) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][3]  ( .D(n2503), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n63), .QN(n4748) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][4]  ( .D(n2502), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n62), .QN(n4735) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][5]  ( .D(n2501), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n61), .QN(n4730) );
  DFFNSRX2TS \dataoutbuffer_reg[2][3]  ( .D(n2767), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n132), .QN(n4684) );
  DFFNSRX2TS \dataoutbuffer_reg[2][4]  ( .D(n2766), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n131), .QN(n4677) );
  DFFNSRX2TS \dataoutbuffer_reg[2][5]  ( .D(n2765), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n130), .QN(n4670) );
  DFFNSRX2TS \dataoutbuffer_reg[2][14]  ( .D(n2756), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n123), .QN(n4585) );
  DFFNSRX2TS \dataoutbuffer_reg[2][15]  ( .D(n2755), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n122), .QN(n4578) );
  DFFNSRX2TS \dataoutbuffer_reg[2][17]  ( .D(n2753), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n121), .QN(n4562) );
  DFFNSRX2TS \dataoutbuffer_reg[2][30]  ( .D(n2740), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n111), .QN(n4443) );
  DFFNSRX2TS \dataoutbuffer_reg[0][3]  ( .D(n2831), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n60), .QN(n4686) );
  DFFNSRX2TS \dataoutbuffer_reg[0][4]  ( .D(n2830), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n59), .QN(n4675) );
  DFFNSRX2TS \dataoutbuffer_reg[0][6]  ( .D(n2828), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n58), .QN(n4659) );
  DFFNSRX2TS \dataoutbuffer_reg[0][7]  ( .D(n2827), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n57), .QN(n4650) );
  DFFNSRX2TS \dataoutbuffer_reg[0][8]  ( .D(n2826), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n56), .QN(n4645) );
  DFFNSRX2TS \dataoutbuffer_reg[0][10]  ( .D(n2824), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n55), .QN(n4625) );
  DFFNSRX2TS \dataoutbuffer_reg[0][11]  ( .D(n2823), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n54), .QN(n4612) );
  DFFNSRX2TS \dataoutbuffer_reg[0][12]  ( .D(n2822), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n53), .QN(n4607) );
  DFFNSRX2TS \dataoutbuffer_reg[0][13]  ( .D(n2821), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n52), .QN(n4600) );
  DFFNSRX2TS \dataoutbuffer_reg[0][14]  ( .D(n2820), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n51), .QN(n4587) );
  DFFNSRX2TS \dataoutbuffer_reg[0][15]  ( .D(n2819), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n50), .QN(n4580) );
  DFFNSRX2TS \dataoutbuffer_reg[0][16]  ( .D(n2818), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n49), .QN(n4569) );
  DFFNSRX2TS \dataoutbuffer_reg[0][17]  ( .D(n2817), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n48), .QN(n4560) );
  DFFNSRX2TS \dataoutbuffer_reg[0][18]  ( .D(n2816), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n47), .QN(n4551) );
  DFFNSRX2TS \dataoutbuffer_reg[0][19]  ( .D(n2815), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n46), .QN(n4542) );
  DFFNSRX2TS \dataoutbuffer_reg[0][21]  ( .D(n2813), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n45), .QN(n4528) );
  DFFNSRX2TS \dataoutbuffer_reg[0][22]  ( .D(n2812), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n44), .QN(n4513) );
  DFFNSRX2TS \dataoutbuffer_reg[0][24]  ( .D(n2810), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n43), .QN(n4497) );
  DFFNSRX2TS \dataoutbuffer_reg[0][25]  ( .D(n2809), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n42), .QN(n4488) );
  DFFNSRX2TS \dataoutbuffer_reg[0][26]  ( .D(n2808), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n41), .QN(n4481) );
  DFFNSRX2TS \dataoutbuffer_reg[0][29]  ( .D(n2805), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n40), .QN(n4456) );
  DFFNSRX2TS \dataoutbuffer_reg[0][30]  ( .D(n2804), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n39), .QN(n4445) );
  DFFNSRX2TS \dataoutbuffer_reg[0][31]  ( .D(n2803), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n38), .QN(n4432) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][1]  ( .D(n2463), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n37), .QN(n4760) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][2]  ( .D(n2462), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n36), .QN(n4755) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][3]  ( .D(n2461), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n35), .QN(n4744) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][5]  ( .D(n2459), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n34), .QN(n4724) );
  DFFNSRX2TS \writeOutbuffer_reg[0]  ( .D(n2571), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[0]), .QN(n156) );
  DFFNSRX2TS \writeOutbuffer_reg[3]  ( .D(n2574), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[3]), .QN(n155) );
  DFFNSRX2TS \writeOutbuffer_reg[6]  ( .D(n2577), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[6]), .QN(n152) );
  DFFNSRX2TS \readOutbuffer_reg[7]  ( .D(n2570), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[7]), .QN(n149) );
  DFFNSRX2TS \readOutbuffer_reg[2]  ( .D(n2565), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[2]), .QN(n150) );
  DFFNSRX2TS \readOutbuffer_reg[4]  ( .D(n2567), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[4]), .QN(n148) );
  DFFNSRX2TS \read_reg_reg[0]  ( .D(n2889), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n9), .QN(n16) );
  DFFNSRX2TS full_reg_reg ( .D(N4718), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        n4844), .QN(n157) );
  DFFNSRX2TS writeOut_reg ( .D(n2449), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        writeOut), .QN(n4841) );
  DFFNSRX2TS \requesterAddressOut_reg[0]  ( .D(n2434), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[0]), .QN(n4845) );
  DFFNSRX2TS \requesterAddressOut_reg[3]  ( .D(n2431), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[3]), .QN(n4846) );
  DFFNSRX2TS readOut_reg ( .D(n2450), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        readOut), .QN(n4843) );
  DFFNSRX2TS \destinationAddressOut_reg[0]  ( .D(n2440), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[0]), .QN(n4768) );
  DFFNSRX2TS \destinationAddressOut_reg[1]  ( .D(n2439), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[1]), .QN(n4759) );
  DFFNSRX2TS \destinationAddressOut_reg[2]  ( .D(n2438), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[2]), .QN(n4750) );
  DFFNSRX2TS \destinationAddressOut_reg[3]  ( .D(n2437), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[3]), .QN(n4741) );
  DFFNSRX2TS \destinationAddressOut_reg[4]  ( .D(n2436), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[4]), .QN(n4732) );
  DFFNSRX2TS \destinationAddressOut_reg[5]  ( .D(n2435), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[5]), .QN(n4723) );
  DFFNSRX2TS \requesterAddressOut_reg[1]  ( .D(n2433), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[1]), .QN(n4722) );
  DFFNSRX2TS \requesterAddressOut_reg[2]  ( .D(n2432), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[2]), .QN(n4721) );
  DFFNSRX2TS \requesterAddressOut_reg[4]  ( .D(n2430), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[4]), .QN(n4720) );
  DFFNSRX2TS \requesterAddressOut_reg[5]  ( .D(n2429), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[5]), .QN(n4719) );
  DFFNSRX2TS \dataOut_reg[0]  ( .D(n2428), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[0]), .QN(n4710) );
  DFFNSRX2TS \dataOut_reg[1]  ( .D(n2427), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[1]), .QN(n4701) );
  DFFNSRX2TS \dataOut_reg[2]  ( .D(n2426), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[2]), .QN(n4692) );
  DFFNSRX2TS \dataOut_reg[3]  ( .D(n2425), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[3]), .QN(n4683) );
  DFFNSRX2TS \dataOut_reg[4]  ( .D(n2424), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[4]), .QN(n4674) );
  DFFNSRX2TS \dataOut_reg[5]  ( .D(n2423), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[5]), .QN(n4665) );
  DFFNSRX2TS \dataOut_reg[6]  ( .D(n2422), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[6]), .QN(n4656) );
  DFFNSRX2TS \dataOut_reg[7]  ( .D(n2421), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[7]), .QN(n4647) );
  DFFNSRX2TS \dataOut_reg[8]  ( .D(n2420), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[8]), .QN(n4638) );
  DFFNSRX2TS \dataOut_reg[9]  ( .D(n2419), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[9]), .QN(n4629) );
  DFFNSRX2TS \dataOut_reg[10]  ( .D(n2418), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[10]), .QN(n4620) );
  DFFNSRX2TS \dataOut_reg[11]  ( .D(n2417), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[11]), .QN(n4611) );
  DFFNSRX2TS \dataOut_reg[12]  ( .D(n2416), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[12]), .QN(n4602) );
  DFFNSRX2TS \dataOut_reg[13]  ( .D(n2415), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[13]), .QN(n4593) );
  DFFNSRX2TS \dataOut_reg[14]  ( .D(n2414), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[14]), .QN(n4584) );
  DFFNSRX2TS \dataOut_reg[15]  ( .D(n2413), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[15]), .QN(n4575) );
  DFFNSRX2TS \dataOut_reg[16]  ( .D(n2412), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[16]), .QN(n4566) );
  DFFNSRX2TS \dataOut_reg[17]  ( .D(n2411), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[17]), .QN(n4557) );
  DFFNSRX2TS \dataOut_reg[18]  ( .D(n2410), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[18]), .QN(n4548) );
  DFFNSRX2TS \dataOut_reg[19]  ( .D(n2409), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[19]), .QN(n4539) );
  DFFNSRX2TS \dataOut_reg[20]  ( .D(n2408), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[20]), .QN(n4530) );
  DFFNSRX2TS \dataOut_reg[21]  ( .D(n2407), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[21]), .QN(n4521) );
  DFFNSRX2TS \dataOut_reg[22]  ( .D(n2406), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[22]), .QN(n4512) );
  DFFNSRX2TS \dataOut_reg[23]  ( .D(n2405), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[23]), .QN(n4503) );
  DFFNSRX2TS \dataOut_reg[24]  ( .D(n2404), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[24]), .QN(n4494) );
  DFFNSRX2TS \dataOut_reg[25]  ( .D(n2403), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[25]), .QN(n4485) );
  DFFNSRX2TS \dataOut_reg[26]  ( .D(n2402), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[26]), .QN(n4476) );
  DFFNSRX2TS \dataOut_reg[27]  ( .D(n2401), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[27]), .QN(n4467) );
  DFFNSRX2TS \dataOut_reg[28]  ( .D(n2400), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[28]), .QN(n4458) );
  DFFNSRX2TS \dataOut_reg[29]  ( .D(n2399), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[29]), .QN(n4449) );
  DFFNSRX2TS \dataOut_reg[30]  ( .D(n2398), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[30]), .QN(n4440) );
  DFFNSRX2TS \dataOut_reg[31]  ( .D(n2397), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[31]), .QN(n4431) );
  DFFNSRX2TS \destinationAddressOut_reg[6]  ( .D(n2448), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[6]) );
  DFFNSRX2TS \destinationAddressOut_reg[7]  ( .D(n2447), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[7]) );
  DFFNSRX2TS \destinationAddressOut_reg[8]  ( .D(n2446), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[8]) );
  DFFNSRX2TS \destinationAddressOut_reg[9]  ( .D(n2445), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[9]) );
  DFFNSRX2TS \destinationAddressOut_reg[10]  ( .D(n2444), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[10]) );
  DFFNSRX2TS \destinationAddressOut_reg[11]  ( .D(n2443), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[11]) );
  DFFNSRX2TS \destinationAddressOut_reg[12]  ( .D(n2442), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[12]) );
  DFFNSRX2TS \destinationAddressOut_reg[13]  ( .D(n2441), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[13]) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][10]  ( .D(n2524), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4808) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][4]  ( .D(n2530), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4738) );
  DFFNSRXLTS \dataoutbuffer_reg[5][0]  ( .D(n2674), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4718) );
  DFFNSRXLTS \dataoutbuffer_reg[5][2]  ( .D(n2672), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4696) );
  DFFNSRXLTS \dataoutbuffer_reg[5][3]  ( .D(n2671), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4691) );
  DFFNSRXLTS \dataoutbuffer_reg[5][4]  ( .D(n2670), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4680) );
  DFFNSRXLTS \dataoutbuffer_reg[5][5]  ( .D(n2669), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4673) );
  DFFNSRXLTS \dataoutbuffer_reg[5][6]  ( .D(n2668), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4660) );
  DFFNSRXLTS \dataoutbuffer_reg[5][7]  ( .D(n2667), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4653) );
  DFFNSRXLTS \dataoutbuffer_reg[5][8]  ( .D(n2666), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4644) );
  DFFNSRXLTS \dataoutbuffer_reg[5][9]  ( .D(n2665), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4633) );
  DFFNSRXLTS \dataoutbuffer_reg[5][10]  ( .D(n2664), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4622) );
  DFFNSRXLTS \dataoutbuffer_reg[5][12]  ( .D(n2662), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4608) );
  DFFNSRXLTS \dataoutbuffer_reg[5][13]  ( .D(n2661), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4599) );
  DFFNSRXLTS \dataoutbuffer_reg[5][14]  ( .D(n2660), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4586) );
  DFFNSRXLTS \dataoutbuffer_reg[5][17]  ( .D(n2657), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4563) );
  DFFNSRXLTS \dataoutbuffer_reg[5][18]  ( .D(n2656), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4552) );
  DFFNSRXLTS \dataoutbuffer_reg[5][19]  ( .D(n2655), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4545) );
  DFFNSRXLTS \dataoutbuffer_reg[5][20]  ( .D(n2654), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4532) );
  DFFNSRXLTS \dataoutbuffer_reg[5][21]  ( .D(n2653), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4525) );
  DFFNSRXLTS \dataoutbuffer_reg[5][22]  ( .D(n2652), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4518) );
  DFFNSRXLTS \dataoutbuffer_reg[5][23]  ( .D(n2651), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4507) );
  DFFNSRXLTS \dataoutbuffer_reg[5][24]  ( .D(n2650), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4500) );
  DFFNSRXLTS \dataoutbuffer_reg[5][25]  ( .D(n2649), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4493) );
  DFFNSRXLTS \dataoutbuffer_reg[5][26]  ( .D(n2648), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4478) );
  DFFNSRXLTS \dataoutbuffer_reg[5][27]  ( .D(n2647), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4469) );
  DFFNSRXLTS \dataoutbuffer_reg[5][28]  ( .D(n2646), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4466) );
  DFFNSRXLTS \dataoutbuffer_reg[5][29]  ( .D(n2645), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4455) );
  DFFNSRXLTS \dataoutbuffer_reg[5][30]  ( .D(n2644), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4444) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][0]  ( .D(n2534), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4772) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][1]  ( .D(n2533), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4765) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][2]  ( .D(n2532), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4756) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][3]  ( .D(n2531), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4747) );
  DFFNSRXLTS \dataoutbuffer_reg[5][1]  ( .D(n2673), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4706) );
  DFFNSRXLTS \dataoutbuffer_reg[5][11]  ( .D(n2663), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4614) );
  DFFNSRXLTS \dataoutbuffer_reg[5][15]  ( .D(n2659), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4576) );
  DFFNSRXLTS \dataoutbuffer_reg[5][16]  ( .D(n2658), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4571) );
  DFFNSRXLTS \dataoutbuffer_reg[5][31]  ( .D(n2643), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4436) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][4]  ( .D(n2474), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4734) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][4]  ( .D(n2516), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4737) );
  DFFNSRXLTS \dataoutbuffer_reg[1][0]  ( .D(n2802), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4717) );
  DFFNSRXLTS \dataoutbuffer_reg[1][1]  ( .D(n2801), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4705) );
  DFFNSRXLTS \dataoutbuffer_reg[1][3]  ( .D(n2799), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4687) );
  DFFNSRXLTS \dataoutbuffer_reg[1][4]  ( .D(n2798), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4682) );
  DFFNSRXLTS \dataoutbuffer_reg[1][6]  ( .D(n2796), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4658) );
  DFFNSRXLTS \dataoutbuffer_reg[1][7]  ( .D(n2795), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4655) );
  DFFNSRXLTS \dataoutbuffer_reg[1][9]  ( .D(n2793), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4631) );
  DFFNSRXLTS \dataoutbuffer_reg[1][11]  ( .D(n2791), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4613) );
  DFFNSRXLTS \dataoutbuffer_reg[1][12]  ( .D(n2790), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4610) );
  DFFNSRXLTS \dataoutbuffer_reg[1][13]  ( .D(n2789), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4601) );
  DFFNSRXLTS \dataoutbuffer_reg[1][14]  ( .D(n2788), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4588) );
  DFFNSRXLTS \dataoutbuffer_reg[1][15]  ( .D(n2787), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4581) );
  DFFNSRXLTS \dataoutbuffer_reg[1][16]  ( .D(n2786), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4574) );
  DFFNSRXLTS \dataoutbuffer_reg[1][17]  ( .D(n2785), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4559) );
  DFFNSRXLTS \dataoutbuffer_reg[1][18]  ( .D(n2784), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4556) );
  DFFNSRXLTS \dataoutbuffer_reg[1][21]  ( .D(n2781), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4523) );
  DFFNSRXLTS \dataoutbuffer_reg[1][23]  ( .D(n2779), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4505) );
  DFFNSRXLTS \dataoutbuffer_reg[1][24]  ( .D(n2778), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4496) );
  DFFNSRXLTS \dataoutbuffer_reg[1][25]  ( .D(n2777), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4491) );
  DFFNSRXLTS \dataoutbuffer_reg[1][26]  ( .D(n2776), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4484) );
  DFFNSRXLTS \dataoutbuffer_reg[1][28]  ( .D(n2774), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4460) );
  DFFNSRXLTS \dataoutbuffer_reg[1][29]  ( .D(n2773), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4453) );
  DFFNSRXLTS \dataoutbuffer_reg[1][30]  ( .D(n2772), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4448) );
  DFFNSRXLTS \dataoutbuffer_reg[1][31]  ( .D(n2771), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4439) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][0]  ( .D(n2478), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4776) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][1]  ( .D(n2477), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4767) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][2]  ( .D(n2476), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4758) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][3]  ( .D(n2475), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4745) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][5]  ( .D(n2473), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4725) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][0]  ( .D(n2548), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4771) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][1]  ( .D(n2547), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4762) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][2]  ( .D(n2546), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4753) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][3]  ( .D(n2545), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4742) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][0]  ( .D(n2520), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4769) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][1]  ( .D(n2519), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4764) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][2]  ( .D(n2518), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4751) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][3]  ( .D(n2517), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4746) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][5]  ( .D(n2515), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4726) );
  DFFNSRXLTS \dataoutbuffer_reg[1][2]  ( .D(n2800), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4693) );
  DFFNSRXLTS \dataoutbuffer_reg[1][5]  ( .D(n2797), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4666) );
  DFFNSRXLTS \dataoutbuffer_reg[1][8]  ( .D(n2794), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4641) );
  DFFNSRXLTS \dataoutbuffer_reg[1][10]  ( .D(n2792), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4627) );
  DFFNSRXLTS \dataoutbuffer_reg[1][19]  ( .D(n2783), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4544) );
  DFFNSRXLTS \dataoutbuffer_reg[1][20]  ( .D(n2782), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4533) );
  DFFNSRXLTS \dataoutbuffer_reg[1][22]  ( .D(n2780), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4517) );
  DFFNSRXLTS \dataoutbuffer_reg[1][27]  ( .D(n2775), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4468) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][4]  ( .D(n2544), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4739) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][0]  ( .D(n2858), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][0] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][1]  ( .D(n2857), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][1] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][2]  ( .D(n2856), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][2] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][3]  ( .D(n2855), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][3] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][5]  ( .D(n2853), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][5] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][4]  ( .D(n2854), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][4] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[6][1]  ( .D(n2875), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][1] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[6][2]  ( .D(n2874), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][2] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[6][3]  ( .D(n2873), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][3] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[6][4]  ( .D(n2872), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][4] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[6][5]  ( .D(n2871), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][5] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[6][0]  ( .D(n2876), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][0] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[5][0]  ( .D(n2870), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6277) );
  DFFNSRXLTS \requesterAddressbuffer_reg[5][1]  ( .D(n2869), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6276) );
  DFFNSRXLTS \requesterAddressbuffer_reg[5][2]  ( .D(n2868), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6275) );
  DFFNSRXLTS \requesterAddressbuffer_reg[5][3]  ( .D(n2867), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6274) );
  DFFNSRXLTS \requesterAddressbuffer_reg[5][4]  ( .D(n2866), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6273) );
  DFFNSRXLTS \requesterAddressbuffer_reg[5][5]  ( .D(n2865), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6272) );
  DFFNSRXLTS \writeOutbuffer_reg[5]  ( .D(n2576), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n6271) );
  DFFNSRXLTS \requesterAddressbuffer_reg[4][4]  ( .D(n2860), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6270) );
  DFFNSRXLTS \requesterAddressbuffer_reg[4][5]  ( .D(n2859), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6269) );
  DFFNSRXLTS \requesterAddressbuffer_reg[4][0]  ( .D(n2864), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6262) );
  DFFNSRXLTS \requesterAddressbuffer_reg[4][1]  ( .D(n2863), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6261) );
  DFFNSRXLTS \requesterAddressbuffer_reg[4][2]  ( .D(n2862), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6260) );
  DFFNSRXLTS \requesterAddressbuffer_reg[4][3]  ( .D(n2861), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6259) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][0]  ( .D(n2846), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6268) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][1]  ( .D(n2845), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6267) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][2]  ( .D(n2844), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6266) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][3]  ( .D(n2843), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6265) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][4]  ( .D(n2842), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6264) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][5]  ( .D(n2841), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6263) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][6]  ( .D(n2528), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4834) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][7]  ( .D(n2527), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4828) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][8]  ( .D(n2526), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4822) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][9]  ( .D(n2525), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4812) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][11]  ( .D(n2523), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4798) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][12]  ( .D(n2522), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4792) );
  DFFNSRX2TS \read_reg_reg[1]  ( .D(n2883), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n10), .QN(n443) );
  DFFNSRX2TS \read_reg_reg[2]  ( .D(n2884), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n8), .QN(n440) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][5]  ( .D(n2529), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4729) );
  DFFNSRXLTS \dataoutbuffer_reg[4][31]  ( .D(n2675), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4433) );
  DFFNSRXLTS \dataoutbuffer_reg[4][30]  ( .D(n2676), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4441) );
  DFFNSRXLTS \dataoutbuffer_reg[4][29]  ( .D(n2677), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4457) );
  DFFNSRXLTS \dataoutbuffer_reg[4][28]  ( .D(n2678), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4459) );
  DFFNSRXLTS \dataoutbuffer_reg[4][27]  ( .D(n2679), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4470) );
  DFFNSRXLTS \dataoutbuffer_reg[4][26]  ( .D(n2680), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4477) );
  DFFNSRXLTS \dataoutbuffer_reg[4][25]  ( .D(n2681), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4490) );
  DFFNSRXLTS \dataoutbuffer_reg[4][24]  ( .D(n2682), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4495) );
  DFFNSRXLTS \dataoutbuffer_reg[4][23]  ( .D(n2683), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4506) );
  DFFNSRXLTS \dataoutbuffer_reg[4][22]  ( .D(n2684), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4516) );
  DFFNSRXLTS \dataoutbuffer_reg[4][21]  ( .D(n2685), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4527) );
  DFFNSRXLTS \dataoutbuffer_reg[4][20]  ( .D(n2686), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4536) );
  DFFNSRXLTS \dataoutbuffer_reg[4][19]  ( .D(n2687), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4541) );
  DFFNSRXLTS \dataoutbuffer_reg[4][18]  ( .D(n2688), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4549) );
  DFFNSRXLTS \dataoutbuffer_reg[4][17]  ( .D(n2689), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4564) );
  DFFNSRXLTS \dataoutbuffer_reg[4][16]  ( .D(n2690), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4568) );
  DFFNSRXLTS \dataoutbuffer_reg[4][15]  ( .D(n2691), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4582) );
  DFFNSRXLTS \dataoutbuffer_reg[4][14]  ( .D(n2692), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4591) );
  DFFNSRXLTS \dataoutbuffer_reg[4][13]  ( .D(n2693), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4594) );
  DFFNSRXLTS \dataoutbuffer_reg[4][12]  ( .D(n2694), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4606) );
  DFFNSRXLTS \dataoutbuffer_reg[4][11]  ( .D(n2695), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4617) );
  DFFNSRXLTS \dataoutbuffer_reg[4][10]  ( .D(n2696), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4624) );
  DFFNSRXLTS \dataoutbuffer_reg[4][9]  ( .D(n2697), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4634) );
  DFFNSRXLTS \dataoutbuffer_reg[4][8]  ( .D(n2698), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4640) );
  DFFNSRXLTS \dataoutbuffer_reg[4][7]  ( .D(n2699), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4652) );
  DFFNSRXLTS \dataoutbuffer_reg[4][6]  ( .D(n2700), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4662) );
  DFFNSRXLTS \dataoutbuffer_reg[4][5]  ( .D(n2701), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4668) );
  DFFNSRXLTS \dataoutbuffer_reg[4][4]  ( .D(n2702), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4679) );
  DFFNSRXLTS \dataoutbuffer_reg[4][3]  ( .D(n2703), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4690) );
  DFFNSRXLTS \dataoutbuffer_reg[4][2]  ( .D(n2704), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4695) );
  DFFNSRXLTS \dataoutbuffer_reg[4][1]  ( .D(n2705), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4703) );
  DFFNSRXLTS \dataoutbuffer_reg[4][0]  ( .D(n2706), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4714) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][13]  ( .D(n2521), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4782) );
  DFFNSRXLTS empty_reg_reg ( .D(n2885), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        n6257), .QN(n4842) );
  DFFNSRXLTS \write_reg_reg[0]  ( .D(n2888), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n18), .QN(n5327) );
  DFFNSRXLTS \write_reg_reg[1]  ( .D(n2887), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n14), .QN(n5323) );
  DFFNSRXLTS \write_reg_reg[2]  ( .D(n2886), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n15), .QN(n5326) );
  DFFNSRX1TS \dataoutbuffer_reg[2][1]  ( .D(n2769), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n140), .QN(n4709) );
  DFFNSRX1TS \dataoutbuffer_reg[2][0]  ( .D(n2770), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n147), .QN(n4713) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][2]  ( .D(n2490), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n110), .QN(n4757) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][5]  ( .D(n2487), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n133), .QN(n4727) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][4]  ( .D(n2488), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n134), .QN(n4740) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][3]  ( .D(n2489), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n135), .QN(n4749) );
  DFFNSRX1TS \dataoutbuffer_reg[2][29]  ( .D(n2741), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n112), .QN(n4450) );
  DFFNSRX1TS \dataoutbuffer_reg[2][28]  ( .D(n2742), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n113), .QN(n4461) );
  DFFNSRX1TS \dataoutbuffer_reg[2][26]  ( .D(n2744), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n114), .QN(n4479) );
  DFFNSRX1TS \dataoutbuffer_reg[2][25]  ( .D(n2745), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n115), .QN(n4486) );
  DFFNSRX1TS \dataoutbuffer_reg[2][23]  ( .D(n2747), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n116), .QN(n4508) );
  DFFNSRX1TS \dataoutbuffer_reg[2][21]  ( .D(n2749), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n117), .QN(n4522) );
  DFFNSRX1TS \dataoutbuffer_reg[2][20]  ( .D(n2750), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n118), .QN(n4535) );
  DFFNSRX1TS \dataoutbuffer_reg[2][19]  ( .D(n2751), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n119), .QN(n4540) );
  DFFNSRX1TS \dataoutbuffer_reg[2][18]  ( .D(n2752), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n120), .QN(n4553) );
  DFFNSRX1TS \dataoutbuffer_reg[2][13]  ( .D(n2757), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n124), .QN(n4596) );
  DFFNSRX1TS \dataoutbuffer_reg[2][12]  ( .D(n2758), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n125), .QN(n4603) );
  DFFNSRX1TS \dataoutbuffer_reg[2][11]  ( .D(n2759), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n126), .QN(n4618) );
  DFFNSRX1TS \dataoutbuffer_reg[2][9]  ( .D(n2761), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n127), .QN(n4630) );
  DFFNSRX1TS \dataoutbuffer_reg[2][8]  ( .D(n2762), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n128), .QN(n4643) );
  DFFNSRX1TS \dataoutbuffer_reg[2][7]  ( .D(n2763), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n129), .QN(n4648) );
  DFFNSRX1TS \dataoutbuffer_reg[2][27]  ( .D(n2743), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n138), .QN(n4475) );
  DFFNSRX1TS \dataoutbuffer_reg[2][10]  ( .D(n2760), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n139), .QN(n4626) );
  DFFNSRX1TS \dataoutbuffer_reg[2][6]  ( .D(n2764), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n145), .QN(n4663) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][8]  ( .D(n2512), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4821) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][7]  ( .D(n2513), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4825) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][6]  ( .D(n2514), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4837) );
  DFFNSRX1TS \writeOutbuffer_reg[4]  ( .D(n2575), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[4]), .QN(n153) );
  NOR2XLTS U2 ( .A(n5521), .B(n6310), .Y(n6114) );
  INVX2TS U3 ( .A(n5333), .Y(n6310) );
  OAI22X2TS U4 ( .A0(n5534), .A1(n352), .B0(n283), .B1(n231), .Y(n5580) );
  OAI211XLTS U5 ( .A0(n4729), .A1(n3401), .B0(n5460), .C0(n5459), .Y(n2529) );
  OAI221X4TS U6 ( .A0(readIn_SOUTH), .A1(n6289), .B0(n3828), .B1(n5567), .C0(
        n5566), .Y(n5571) );
  NOR3X2TS U7 ( .A(n6288), .B(n569), .C(n5325), .Y(n5567) );
  AND3X2TS U8 ( .A(n223), .B(n237), .C(n5426), .Y(n6175) );
  NAND3X1TS U9 ( .A(n5472), .B(n5447), .C(n6296), .Y(n5426) );
  OAI22X2TS U10 ( .A0(n5520), .A1(n350), .B0(n282), .B1(n6283), .Y(n5575) );
  OA21X2TS U11 ( .A0(n5539), .A1(n5425), .B0(n5523), .Y(n5520) );
  AOI221X2TS U12 ( .A0(n263), .A1(n5355), .B0(n6287), .B1(n289), .C0(n261), 
        .Y(n5539) );
  INVX2TS U13 ( .A(n5355), .Y(n6287) );
  INVXLTS U14 ( .A(n5573), .Y(n1) );
  CLKINVX2TS U15 ( .A(n1), .Y(n2) );
  BUFX4TS U16 ( .A(n3325), .Y(n3324) );
  INVXLTS U17 ( .A(n5447), .Y(n6295) );
  INVX4TS U18 ( .A(n5447), .Y(n276) );
  XOR2X4TS U19 ( .A(n5332), .B(n15), .Y(n5447) );
  BUFX3TS U20 ( .A(n3457), .Y(n3455) );
  AO21X1TS U21 ( .A0(n230), .A1(n5458), .B0(n565), .Y(n12) );
  AOI21X1TS U22 ( .A0(n229), .A1(n5402), .B0(n6306), .Y(n5537) );
  AOI21X1TS U23 ( .A0(n447), .A1(n234), .B0(n561), .Y(n5558) );
  INVX2TS U24 ( .A(n5400), .Y(n6296) );
  OAI21X1TS U25 ( .A0(n5328), .A1(n5539), .B0(n6289), .Y(n5449) );
  NAND2X1TS U26 ( .A(n6290), .B(selectBit_EAST), .Y(n5495) );
  INVX2TS U27 ( .A(n5400), .Y(n444) );
  AOI21X1TS U28 ( .A0(n447), .A1(n5365), .B0(n564), .Y(n5530) );
  AOI21X1TS U29 ( .A0(n5497), .A1(n5506), .B0(n562), .Y(n5572) );
  CLKBUFX2TS U30 ( .A(n3763), .Y(n3757) );
  CLKBUFX2TS U31 ( .A(n3763), .Y(n3759) );
  CLKBUFX2TS U32 ( .A(n3762), .Y(n3761) );
  AND3X2TS U33 ( .A(n226), .B(n5554), .C(n5558), .Y(n6191) );
  OAI21X1TS U34 ( .A0(n5495), .A1(n5546), .B0(n5426), .Y(n5547) );
  CLKBUFX2TS U35 ( .A(n3762), .Y(n3760) );
  CLKBUFX2TS U36 ( .A(n3763), .Y(n3758) );
  CLKBUFX2TS U37 ( .A(n3762), .Y(n3756) );
  OA21XLTS U38 ( .A0(n6290), .A1(n5448), .B0(n5527), .Y(n5526) );
  CLKBUFX2TS U39 ( .A(n5558), .Y(n222) );
  OA21XLTS U40 ( .A0(n5449), .A1(n5448), .B0(n5554), .Y(n5553) );
  NOR3X1TS U41 ( .A(n5561), .B(n5562), .C(n5559), .Y(n5560) );
  INVX2TS U42 ( .A(n5539), .Y(n6288) );
  CLKBUFX2TS U43 ( .A(n3429), .Y(n3419) );
  AOI222XLTS U44 ( .A0(\requesterAddressbuffer[6][5] ), .A1(n699), .B0(n3455), 
        .B1(n4253), .C0(n365), .C1(n4411), .Y(n6194) );
  AOI222XLTS U45 ( .A0(n379), .A1(n130), .B0(n4158), .B1(n1728), .C0(n4315), 
        .C1(n3765), .Y(n5962) );
  AOI222XLTS U46 ( .A0(n3918), .A1(n3706), .B0(n455), .B1(n3439), .C0(n4074), 
        .C1(n6204), .Y(n5658) );
  AOI222XLTS U47 ( .A0(n3900), .A1(n3704), .B0(n467), .B1(n3438), .C0(n4056), 
        .C1(n3427), .Y(n5670) );
  AOI222XLTS U48 ( .A0(n3894), .A1(n3704), .B0(n471), .B1(n3445), .C0(n4050), 
        .C1(n3426), .Y(n5674) );
  AOI222XLTS U49 ( .A0(n3891), .A1(n3703), .B0(n473), .B1(n3445), .C0(n4047), 
        .C1(n3427), .Y(n5676) );
  AOI222XLTS U50 ( .A0(n3870), .A1(n3702), .B0(n487), .B1(n3437), .C0(n4026), 
        .C1(n3423), .Y(n5690) );
  AOI222XLTS U51 ( .A0(n3867), .A1(n3701), .B0(n489), .B1(n3437), .C0(n4023), 
        .C1(n3422), .Y(n5692) );
  AOI222XLTS U52 ( .A0(n3861), .A1(n3701), .B0(n493), .B1(n3437), .C0(n4017), 
        .C1(n3422), .Y(n5696) );
  AOI222XLTS U53 ( .A0(n3849), .A1(n3700), .B0(n508), .B1(n3436), .C0(n4005), 
        .C1(n3423), .Y(n5704) );
  AOI222XLTS U54 ( .A0(n3834), .A1(n3699), .B0(n536), .B1(n3434), .C0(n3990), 
        .C1(n3420), .Y(n5714) );
  AOI222XLTS U55 ( .A0(n3924), .A1(n3706), .B0(n451), .B1(n3440), .C0(n4080), 
        .C1(n3430), .Y(n5654) );
  AOI222XLTS U56 ( .A0(n3921), .A1(n3706), .B0(n453), .B1(n3440), .C0(n4077), 
        .C1(n3430), .Y(n5656) );
  AOI222XLTS U57 ( .A0(n3915), .A1(n3706), .B0(n457), .B1(n3439), .C0(n4071), 
        .C1(n3426), .Y(n5660) );
  AOI222XLTS U58 ( .A0(n3912), .A1(n3705), .B0(n459), .B1(n3439), .C0(n4068), 
        .C1(n3424), .Y(n5662) );
  AOI222XLTS U59 ( .A0(n3909), .A1(n3705), .B0(n461), .B1(n3439), .C0(n4065), 
        .C1(n3424), .Y(n5664) );
  AOI222XLTS U60 ( .A0(n3903), .A1(n3705), .B0(n465), .B1(n3438), .C0(n4059), 
        .C1(n3424), .Y(n5668) );
  AOI222XLTS U61 ( .A0(n3897), .A1(n3704), .B0(n469), .B1(n3438), .C0(n4053), 
        .C1(n3431), .Y(n5672) );
  AOI222XLTS U62 ( .A0(n3888), .A1(n3703), .B0(n475), .B1(n3445), .C0(n4044), 
        .C1(n3428), .Y(n5678) );
  AOI222XLTS U63 ( .A0(n3882), .A1(n3703), .B0(n479), .B1(n3443), .C0(n4038), 
        .C1(n3426), .Y(n5682) );
  AOI222XLTS U64 ( .A0(n3879), .A1(n3702), .B0(n481), .B1(n3443), .C0(n4035), 
        .C1(n3426), .Y(n5684) );
  AOI222XLTS U65 ( .A0(n3876), .A1(n3702), .B0(n483), .B1(n3443), .C0(n4032), 
        .C1(n3423), .Y(n5686) );
  AOI222XLTS U66 ( .A0(n3873), .A1(n3702), .B0(n485), .B1(n3446), .C0(n4029), 
        .C1(n3423), .Y(n5688) );
  AOI222XLTS U67 ( .A0(n3864), .A1(n3701), .B0(n491), .B1(n3437), .C0(n4020), 
        .C1(n3422), .Y(n5694) );
  AOI222XLTS U68 ( .A0(n3858), .A1(n3701), .B0(n495), .B1(n3436), .C0(n4014), 
        .C1(n3422), .Y(n5698) );
  AOI222XLTS U69 ( .A0(n3855), .A1(n3700), .B0(n501), .B1(n3436), .C0(n4011), 
        .C1(n3421), .Y(n5700) );
  AOI222XLTS U70 ( .A0(n3852), .A1(n3700), .B0(n505), .B1(n3436), .C0(n4008), 
        .C1(n3421), .Y(n5702) );
  AOI222XLTS U71 ( .A0(n3846), .A1(n3700), .B0(n510), .B1(n3435), .C0(n4002), 
        .C1(n3421), .Y(n5706) );
  AOI222XLTS U72 ( .A0(n3840), .A1(n3699), .B0(n515), .B1(n3435), .C0(n3996), 
        .C1(n3420), .Y(n5710) );
  AOI222XLTS U73 ( .A0(n3837), .A1(n3699), .B0(n526), .B1(n3435), .C0(n3993), 
        .C1(n3420), .Y(n5712) );
  AOI222XLTS U74 ( .A0(n3831), .A1(n3704), .B0(n541), .B1(n3434), .C0(n3987), 
        .C1(n3420), .Y(n5716) );
  AOI222XLTS U75 ( .A0(n3906), .A1(n3705), .B0(n464), .B1(n3438), .C0(n4062), 
        .C1(n3424), .Y(n5666) );
  AOI222XLTS U76 ( .A0(n3885), .A1(n3703), .B0(n478), .B1(n3443), .C0(n4041), 
        .C1(n3429), .Y(n5680) );
  AOI222XLTS U77 ( .A0(n3843), .A1(n3699), .B0(n514), .B1(n3435), .C0(n3999), 
        .C1(n3421), .Y(n5708) );
  AOI222XLTS U78 ( .A0(n4293), .A1(n3455), .B0(n4138), .B1(n3417), .C0(n3982), 
        .C1(n3712), .Y(n5474) );
  AOI222XLTS U79 ( .A0(n4287), .A1(n3455), .B0(n4132), .B1(n3417), .C0(n3976), 
        .C1(n3710), .Y(n5476) );
  AOI222XLTS U80 ( .A0(n4290), .A1(n3455), .B0(n4135), .B1(n3418), .C0(n3979), 
        .C1(n3710), .Y(n5475) );
  NOR2BX1TS U81 ( .AN(n5354), .B(n6240), .Y(n5494) );
  OA22X2TS U82 ( .A0(n6254), .A1(n6243), .B0(n4880), .B1(n279), .Y(n3) );
  NOR2BX1TS U83 ( .AN(n222), .B(n281), .Y(n6189) );
  CLKBUFX2TS U84 ( .A(n557), .Y(n3265) );
  OA22X1TS U85 ( .A0(n5566), .A1(n6303), .B0(n262), .B1(n5496), .Y(n562) );
  CLKBUFX2TS U86 ( .A(n6130), .Y(n834) );
  CLKBUFX2TS U87 ( .A(n6127), .Y(n786) );
  NOR2BX1TS U88 ( .AN(n5530), .B(n280), .Y(n6128) );
  OA22X1TS U89 ( .A0(n5549), .A1(n352), .B0(n282), .B1(n233), .Y(n565) );
  OA22X1TS U90 ( .A0(n5526), .A1(n351), .B0(n5496), .B1(n6283), .Y(n564) );
  CLKBUFX2TS U91 ( .A(n3480), .Y(n3474) );
  OR2X2TS U92 ( .A(n6230), .B(n257), .Y(n4) );
  AND3X2TS U93 ( .A(n5558), .B(n281), .C(n5553), .Y(n5) );
  INVX2TS U94 ( .A(n7), .Y(n366) );
  INVX1TS U95 ( .A(n367), .Y(n268) );
  INVX2TS U96 ( .A(n268), .Y(n270) );
  CLKBUFX2TS U97 ( .A(n6172), .Y(n3283) );
  INVX2TS U98 ( .A(n196), .Y(n352) );
  INVX2TS U99 ( .A(n3), .Y(n216) );
  INVX2TS U100 ( .A(selectBit_NORTH), .Y(n6254) );
  AOI32X1TS U101 ( .A0(n6241), .A1(n556), .A2(n163), .B0(n4847), .B1(
        selectBit_SOUTH), .Y(n4848) );
  OAI21X1TS U102 ( .A0(n5403), .A1(n351), .B0(n558), .Y(n557) );
  INVX2TS U103 ( .A(n244), .Y(n245) );
  INVX2TS U104 ( .A(n244), .Y(n359) );
  INVX2TS U105 ( .A(n244), .Y(n357) );
  INVX2TS U106 ( .A(n246), .Y(n248) );
  NAND2XLTS U107 ( .A(n5549), .B(n224), .Y(n5585) );
  AOI21XLTS U108 ( .A0(n556), .A1(n5324), .B0(n227), .Y(n5399) );
  OR2XLTS U109 ( .A(n556), .B(n5324), .Y(n21) );
  NAND2X1TS U110 ( .A(n5324), .B(selectBit_SOUTH), .Y(n5325) );
  CLKINVX2TS U111 ( .A(n5325), .Y(n6) );
  XNOR2X1TS U112 ( .A(selectBit_NORTH), .B(selectBit_EAST), .Y(n4847) );
  NOR2X2TS U113 ( .A(n253), .B(n205), .Y(n5331) );
  CLKBUFX2TS U114 ( .A(n6188), .Y(n3365) );
  CLKBUFX2TS U115 ( .A(n5530), .Y(n221) );
  INVX2TS U116 ( .A(n5581), .Y(n6307) );
  OA22X1TS U117 ( .A0(n5560), .A1(n350), .B0(n262), .B1(n283), .Y(n563) );
  NAND2X1TS U118 ( .A(n557), .B(n5404), .Y(n442) );
  INVX2TS U119 ( .A(n5580), .Y(n6306) );
  CLKBUFX2TS U120 ( .A(n5), .Y(n3722) );
  AOI21X1TS U121 ( .A0(n263), .A1(n230), .B0(n563), .Y(n5565) );
  NOR2X1TS U122 ( .A(n279), .B(n6290), .Y(n5401) );
  CLKBUFX2TS U123 ( .A(n3330), .Y(n3325) );
  CLKBUFX2TS U124 ( .A(n6223), .Y(n3523) );
  CLKBUFX2TS U125 ( .A(n563), .Y(n703) );
  AOI21X1TS U126 ( .A0(n229), .A1(n261), .B0(n6309), .Y(n5333) );
  CLKBUFX2TS U127 ( .A(n736), .Y(n716) );
  NAND2X1TS U128 ( .A(n5534), .B(n218), .Y(n5581) );
  CLKBUFX2TS U129 ( .A(n3391), .Y(n3390) );
  AOI2BB1X1TS U130 ( .A0N(n6288), .A1N(n5425), .B0(n5547), .Y(n5549) );
  INVX2TS U131 ( .A(n5567), .Y(n6289) );
  CLKBUFX2TS U132 ( .A(n5565), .Y(n158) );
  NAND2X1TS U133 ( .A(n557), .B(n5404), .Y(n5538) );
  AOI21X1TS U134 ( .A0(n5543), .A1(n5401), .B0(n6298), .Y(n5541) );
  CLKBUFX2TS U135 ( .A(n3430), .Y(n3417) );
  CLKBUFX2TS U136 ( .A(n3713), .Y(n3708) );
  CLKBUFX2TS U137 ( .A(n828), .Y(n827) );
  CLKBUFX2TS U138 ( .A(n785), .Y(n777) );
  CLKBUFX2TS U139 ( .A(n801), .Y(n787) );
  CLKBUFX2TS U140 ( .A(n3525), .Y(n3522) );
  CLKBUFX2TS U141 ( .A(n3282), .Y(n3275) );
  CLKBUFX2TS U142 ( .A(n3429), .Y(n3418) );
  AOI222XLTS U143 ( .A0(n3984), .A1(n3359), .B0(n4297), .B1(n204), .C0(n4140), 
        .C1(n3395), .Y(n5450) );
  AOI222XLTS U144 ( .A0(n3986), .A1(n3328), .B0(n541), .B1(n3309), .C0(n3831), 
        .C1(n3286), .Y(n5844) );
  AOI222XLTS U145 ( .A0(n3989), .A1(n3329), .B0(n537), .B1(n3305), .C0(n3834), 
        .C1(n3286), .Y(n5842) );
  AOI222XLTS U146 ( .A0(n3992), .A1(n3315), .B0(n531), .B1(n3305), .C0(n3837), 
        .C1(n3286), .Y(n5840) );
  AOI222XLTS U147 ( .A0(n3995), .A1(n3315), .B0(n516), .B1(n3304), .C0(n3840), 
        .C1(n3286), .Y(n5838) );
  AOI222XLTS U148 ( .A0(n3998), .A1(n3315), .B0(n512), .B1(n3305), .C0(n3843), 
        .C1(n3296), .Y(n5836) );
  AOI222XLTS U149 ( .A0(n4001), .A1(n3315), .B0(n511), .B1(n3305), .C0(n3846), 
        .C1(n3297), .Y(n5834) );
  AOI222XLTS U150 ( .A0(n4004), .A1(n3316), .B0(n509), .B1(n3303), .C0(n3849), 
        .C1(n3288), .Y(n5832) );
  AOI222XLTS U151 ( .A0(n4007), .A1(n3316), .B0(n505), .B1(n3303), .C0(n3852), 
        .C1(n3296), .Y(n5830) );
  AOI222XLTS U152 ( .A0(n4010), .A1(n3316), .B0(n503), .B1(n3304), .C0(n3855), 
        .C1(n3297), .Y(n5828) );
  AOI222XLTS U153 ( .A0(n4013), .A1(n3319), .B0(n495), .B1(n3303), .C0(n3858), 
        .C1(n3287), .Y(n5826) );
  AOI222XLTS U154 ( .A0(n4016), .A1(n3316), .B0(n494), .B1(n3304), .C0(n3861), 
        .C1(n3287), .Y(n5824) );
  AOI222XLTS U155 ( .A0(n4019), .A1(n3317), .B0(n492), .B1(n3304), .C0(n3864), 
        .C1(n3287), .Y(n5822) );
  AOI222XLTS U156 ( .A0(n4022), .A1(n3317), .B0(n490), .B1(n3309), .C0(n3867), 
        .C1(n3287), .Y(n5820) );
  AOI222XLTS U157 ( .A0(n4025), .A1(n3317), .B0(n487), .B1(n3303), .C0(n3870), 
        .C1(n3288), .Y(n5818) );
  AOI222XLTS U158 ( .A0(n4028), .A1(n3317), .B0(n486), .B1(n3312), .C0(n3873), 
        .C1(n3288), .Y(n5816) );
  AOI222XLTS U159 ( .A0(n4031), .A1(n3318), .B0(n484), .B1(n3302), .C0(n3876), 
        .C1(n3288), .Y(n5814) );
  AOI222XLTS U160 ( .A0(n4034), .A1(n3318), .B0(n482), .B1(n3301), .C0(n3879), 
        .C1(n3289), .Y(n5812) );
  AOI222XLTS U161 ( .A0(n4037), .A1(n3318), .B0(n480), .B1(n3313), .C0(n3882), 
        .C1(n3289), .Y(n5810) );
  AOI222XLTS U162 ( .A0(n4040), .A1(n3318), .B0(n477), .B1(n3312), .C0(n3885), 
        .C1(n3289), .Y(n5808) );
  AOI222XLTS U163 ( .A0(n4043), .A1(n3319), .B0(n476), .B1(n3313), .C0(n3888), 
        .C1(n3289), .Y(n5806) );
  AOI222XLTS U164 ( .A0(n4046), .A1(n3319), .B0(n474), .B1(n3302), .C0(n3891), 
        .C1(n3290), .Y(n5804) );
  AOI222XLTS U165 ( .A0(n4049), .A1(n3319), .B0(n472), .B1(n3312), .C0(n3894), 
        .C1(n3290), .Y(n5802) );
  AOI222XLTS U166 ( .A0(n4052), .A1(n3320), .B0(n470), .B1(n3302), .C0(n3897), 
        .C1(n3290), .Y(n5800) );
  AOI222XLTS U167 ( .A0(n4055), .A1(n3320), .B0(n467), .B1(n3302), .C0(n3900), 
        .C1(n3290), .Y(n5798) );
  AOI222XLTS U168 ( .A0(n4058), .A1(n3320), .B0(n465), .B1(n3310), .C0(n3903), 
        .C1(n3291), .Y(n5796) );
  AOI222XLTS U169 ( .A0(n4061), .A1(n3320), .B0(n463), .B1(n3313), .C0(n3906), 
        .C1(n3291), .Y(n5794) );
  AOI222XLTS U170 ( .A0(n4064), .A1(n3321), .B0(n461), .B1(n6174), .C0(n3909), 
        .C1(n3291), .Y(n5792) );
  AOI222XLTS U171 ( .A0(n4067), .A1(n3321), .B0(n460), .B1(n3301), .C0(n3912), 
        .C1(n3291), .Y(n5790) );
  AOI222XLTS U172 ( .A0(n4070), .A1(n3321), .B0(n457), .B1(n3301), .C0(n3915), 
        .C1(n3292), .Y(n5788) );
  AOI222XLTS U173 ( .A0(n4073), .A1(n3321), .B0(n456), .B1(n3311), .C0(n3918), 
        .C1(n3292), .Y(n5786) );
  AOI222XLTS U174 ( .A0(n4076), .A1(n3322), .B0(n453), .B1(n3301), .C0(n3921), 
        .C1(n3292), .Y(n5784) );
  AOI222XLTS U175 ( .A0(n4079), .A1(n3322), .B0(n452), .B1(n3314), .C0(n3924), 
        .C1(n3292), .Y(n5782) );
  AOI222XLTS U176 ( .A0(n4115), .A1(n3393), .B0(n3373), .B1(n192), .C0(n4272), 
        .C1(n213), .Y(n5459) );
  AOI222XLTS U177 ( .A0(n3911), .A1(n835), .B0(n459), .B1(n804), .C0(n4224), 
        .C1(n794), .Y(n5982) );
  AOI222XLTS U178 ( .A0(n3896), .A1(n826), .B0(n469), .B1(n807), .C0(n4209), 
        .C1(n793), .Y(n5992) );
  AOI222XLTS U179 ( .A0(n3890), .A1(n824), .B0(n473), .B1(n807), .C0(n4203), 
        .C1(n793), .Y(n5996) );
  AOI222XLTS U180 ( .A0(n3887), .A1(n824), .B0(n475), .B1(n808), .C0(n4200), 
        .C1(n792), .Y(n5998) );
  AOI222XLTS U181 ( .A0(n3860), .A1(n821), .B0(n493), .B1(n810), .C0(n4173), 
        .C1(n790), .Y(n6016) );
  AOI222XLTS U182 ( .A0(n3854), .A1(n821), .B0(n501), .B1(n810), .C0(n4167), 
        .C1(n789), .Y(n6020) );
  AOI222XLTS U183 ( .A0(n3845), .A1(n820), .B0(n510), .B1(n811), .C0(n4158), 
        .C1(n789), .Y(n6026) );
  AOI222XLTS U184 ( .A0(n3836), .A1(n820), .B0(n526), .B1(n811), .C0(n4149), 
        .C1(n788), .Y(n6032) );
  AOI222XLTS U185 ( .A0(n3923), .A1(n834), .B0(n451), .B1(n805), .C0(n4236), 
        .C1(n795), .Y(n5974) );
  AOI222XLTS U186 ( .A0(n3920), .A1(n830), .B0(n454), .B1(n804), .C0(n4233), 
        .C1(n795), .Y(n5976) );
  AOI222XLTS U187 ( .A0(n3917), .A1(n835), .B0(n455), .B1(n805), .C0(n4230), 
        .C1(n795), .Y(n5978) );
  AOI222XLTS U188 ( .A0(n3914), .A1(n828), .B0(n458), .B1(n804), .C0(n4227), 
        .C1(n795), .Y(n5980) );
  AOI222XLTS U189 ( .A0(n3908), .A1(n829), .B0(n462), .B1(n806), .C0(n4221), 
        .C1(n794), .Y(n5984) );
  AOI222XLTS U190 ( .A0(n3905), .A1(n826), .B0(n464), .B1(n806), .C0(n4218), 
        .C1(n794), .Y(n5986) );
  AOI222XLTS U191 ( .A0(n3902), .A1(n826), .B0(n466), .B1(n805), .C0(n4215), 
        .C1(n794), .Y(n5988) );
  AOI222XLTS U192 ( .A0(n3899), .A1(n826), .B0(n468), .B1(n807), .C0(n4212), 
        .C1(n793), .Y(n5990) );
  AOI222XLTS U193 ( .A0(n3893), .A1(n824), .B0(n471), .B1(n805), .C0(n4206), 
        .C1(n793), .Y(n5994) );
  AOI222XLTS U194 ( .A0(n3884), .A1(n823), .B0(n478), .B1(n806), .C0(n4197), 
        .C1(n792), .Y(n6000) );
  AOI222XLTS U195 ( .A0(n3881), .A1(n823), .B0(n479), .B1(n808), .C0(n4194), 
        .C1(n792), .Y(n6002) );
  AOI222XLTS U196 ( .A0(n3878), .A1(n823), .B0(n481), .B1(n804), .C0(n4191), 
        .C1(n792), .Y(n6004) );
  AOI222XLTS U197 ( .A0(n3875), .A1(n823), .B0(n483), .B1(n807), .C0(n4188), 
        .C1(n791), .Y(n6006) );
  AOI222XLTS U198 ( .A0(n3872), .A1(n822), .B0(n485), .B1(n806), .C0(n4185), 
        .C1(n791), .Y(n6008) );
  AOI222XLTS U199 ( .A0(n3869), .A1(n822), .B0(n488), .B1(n809), .C0(n4182), 
        .C1(n791), .Y(n6010) );
  AOI222XLTS U200 ( .A0(n3866), .A1(n822), .B0(n489), .B1(n808), .C0(n4179), 
        .C1(n790), .Y(n6012) );
  AOI222XLTS U201 ( .A0(n3863), .A1(n822), .B0(n491), .B1(n810), .C0(n4176), 
        .C1(n790), .Y(n6014) );
  AOI222XLTS U202 ( .A0(n3857), .A1(n824), .B0(n496), .B1(n809), .C0(n4170), 
        .C1(n790), .Y(n6018) );
  AOI222XLTS U203 ( .A0(n3851), .A1(n821), .B0(n507), .B1(n809), .C0(n4164), 
        .C1(n789), .Y(n6022) );
  AOI222XLTS U204 ( .A0(n3848), .A1(n821), .B0(n508), .B1(n809), .C0(n4161), 
        .C1(n791), .Y(n6024) );
  AOI222XLTS U205 ( .A0(n3842), .A1(n820), .B0(n514), .B1(n811), .C0(n4155), 
        .C1(n789), .Y(n6028) );
  AOI222XLTS U206 ( .A0(n3839), .A1(n820), .B0(n515), .B1(n810), .C0(n4152), 
        .C1(n788), .Y(n6030) );
  AOI222XLTS U207 ( .A0(n3833), .A1(n819), .B0(n536), .B1(n811), .C0(n4146), 
        .C1(n788), .Y(n6034) );
  AOI222XLTS U208 ( .A0(n3830), .A1(n819), .B0(n543), .B1(n808), .C0(n4143), 
        .C1(n788), .Y(n6036) );
  AOI222XLTS U209 ( .A0(n3817), .A1(n779), .B0(n3825), .B1(n800), .C0(n3812), 
        .C1(n834), .Y(n5577) );
  AOI222XLTS U210 ( .A0(n4080), .A1(n3519), .B0(n452), .B1(n3498), .C0(n4236), 
        .C1(n3489), .Y(n5590) );
  AOI222XLTS U211 ( .A0(n4077), .A1(n3519), .B0(n454), .B1(n3498), .C0(n4233), 
        .C1(n3489), .Y(n5592) );
  AOI222XLTS U212 ( .A0(n4074), .A1(n3518), .B0(n456), .B1(n3509), .C0(n4230), 
        .C1(n3489), .Y(n5594) );
  AOI222XLTS U213 ( .A0(n4071), .A1(n3518), .B0(n458), .B1(n3509), .C0(n4227), 
        .C1(n3489), .Y(n5596) );
  AOI222XLTS U214 ( .A0(n4068), .A1(n3518), .B0(n460), .B1(n6222), .C0(n4224), 
        .C1(n3488), .Y(n5598) );
  AOI222XLTS U215 ( .A0(n4065), .A1(n3518), .B0(n462), .B1(n3507), .C0(n4221), 
        .C1(n3488), .Y(n5600) );
  AOI222XLTS U216 ( .A0(n4062), .A1(n3525), .B0(n463), .B1(n3508), .C0(n4218), 
        .C1(n3488), .Y(n5602) );
  AOI222XLTS U217 ( .A0(n4059), .A1(n3523), .B0(n466), .B1(n3508), .C0(n4215), 
        .C1(n3488), .Y(n5604) );
  AOI222XLTS U218 ( .A0(n4056), .A1(n3527), .B0(n468), .B1(n3508), .C0(n4212), 
        .C1(n3491), .Y(n5606) );
  AOI222XLTS U219 ( .A0(n4053), .A1(n3528), .B0(n470), .B1(n6222), .C0(n4209), 
        .C1(n3491), .Y(n5608) );
  AOI222XLTS U220 ( .A0(n4050), .A1(n3526), .B0(n472), .B1(n3511), .C0(n4206), 
        .C1(n3490), .Y(n5610) );
  AOI222XLTS U221 ( .A0(n4047), .A1(n3525), .B0(n474), .B1(n3507), .C0(n4203), 
        .C1(n3494), .Y(n5612) );
  AOI222XLTS U222 ( .A0(n4044), .A1(n3525), .B0(n476), .B1(n3506), .C0(n4200), 
        .C1(n3493), .Y(n5614) );
  AOI222XLTS U223 ( .A0(n4041), .A1(n3517), .B0(n477), .B1(n3505), .C0(n4197), 
        .C1(n3491), .Y(n5616) );
  AOI222XLTS U224 ( .A0(n4038), .A1(n3517), .B0(n480), .B1(n3499), .C0(n4194), 
        .C1(n3494), .Y(n5618) );
  AOI222XLTS U225 ( .A0(n4035), .A1(n3517), .B0(n482), .B1(n3499), .C0(n4191), 
        .C1(n3493), .Y(n5620) );
  AOI222XLTS U226 ( .A0(n4032), .A1(n3517), .B0(n484), .B1(n3499), .C0(n4188), 
        .C1(n3495), .Y(n5622) );
  AOI222XLTS U227 ( .A0(n4029), .A1(n3516), .B0(n486), .B1(n3499), .C0(n4185), 
        .C1(n3492), .Y(n5624) );
  AOI222XLTS U228 ( .A0(n4026), .A1(n3516), .B0(n488), .B1(n3500), .C0(n4182), 
        .C1(n3495), .Y(n5626) );
  AOI222XLTS U229 ( .A0(n4023), .A1(n3516), .B0(n490), .B1(n3500), .C0(n4179), 
        .C1(n3487), .Y(n5628) );
  AOI222XLTS U230 ( .A0(n4020), .A1(n3516), .B0(n492), .B1(n3500), .C0(n4176), 
        .C1(n3487), .Y(n5630) );
  AOI222XLTS U231 ( .A0(n4017), .A1(n3515), .B0(n494), .B1(n3500), .C0(n4173), 
        .C1(n3487), .Y(n5632) );
  AOI222XLTS U232 ( .A0(n4014), .A1(n3515), .B0(n496), .B1(n3501), .C0(n4170), 
        .C1(n3487), .Y(n5634) );
  AOI222XLTS U233 ( .A0(n4011), .A1(n3515), .B0(n503), .B1(n3501), .C0(n4167), 
        .C1(n3486), .Y(n5636) );
  AOI222XLTS U234 ( .A0(n4008), .A1(n3515), .B0(n507), .B1(n3501), .C0(n4164), 
        .C1(n3486), .Y(n5638) );
  AOI222XLTS U235 ( .A0(n4005), .A1(n3514), .B0(n509), .B1(n3501), .C0(n4161), 
        .C1(n3486), .Y(n5640) );
  AOI222XLTS U236 ( .A0(n4002), .A1(n3514), .B0(n511), .B1(n3502), .C0(n4158), 
        .C1(n3486), .Y(n5642) );
  AOI222XLTS U237 ( .A0(n3999), .A1(n3514), .B0(n512), .B1(n3502), .C0(n4155), 
        .C1(n3485), .Y(n5644) );
  AOI222XLTS U238 ( .A0(n3996), .A1(n3514), .B0(n516), .B1(n3502), .C0(n4152), 
        .C1(n3485), .Y(n5646) );
  AOI222XLTS U239 ( .A0(n3993), .A1(n3513), .B0(n531), .B1(n3502), .C0(n4149), 
        .C1(n3485), .Y(n5648) );
  AOI222XLTS U240 ( .A0(n3990), .A1(n3513), .B0(n537), .B1(n3503), .C0(n4146), 
        .C1(n3485), .Y(n5650) );
  AOI222XLTS U241 ( .A0(n3987), .A1(n3513), .B0(n543), .B1(n3503), .C0(n4143), 
        .C1(n3484), .Y(n5652) );
  AOI222XLTS U242 ( .A0(n4140), .A1(n781), .B0(destinationAddressIn_SOUTH[13]), 
        .B1(n6128), .C0(n3985), .C1(n829), .Y(n5356) );
  AOI222XLTS U243 ( .A0(n4296), .A1(n3278), .B0(n3985), .B1(n3284), .C0(n4141), 
        .C1(n3328), .Y(n5427) );
  AND2X2TS U244 ( .A(n5560), .B(n5565), .Y(n7) );
  CLKBUFX2TS U245 ( .A(n3722), .Y(n3720) );
  CLKINVX2TS U246 ( .A(n5537), .Y(n217) );
  CLKBUFX2TS U247 ( .A(n3723), .Y(n3718) );
  CLKBUFX2TS U248 ( .A(n5), .Y(n3723) );
  CLKBUFX2TS U249 ( .A(n3722), .Y(n3719) );
  CLKBUFX2TS U250 ( .A(n3720), .Y(n3717) );
  CLKBUFX2TS U251 ( .A(n3722), .Y(n3721) );
  CLKBUFX2TS U252 ( .A(n3720), .Y(n3716) );
  CLKINVX2TS U253 ( .A(n3752), .Y(n377) );
  CLKBUFX2TS U254 ( .A(n6309), .Y(n3782) );
  INVX2TS U255 ( .A(n217), .Y(n218) );
  INVX2TS U256 ( .A(n5575), .Y(n6309) );
  INVX1TS U257 ( .A(n376), .Y(n271) );
  BUFX3TS U258 ( .A(n6189), .Y(n200) );
  NAND3XLTS U259 ( .A(n221), .B(n280), .C(n5526), .Y(n5578) );
  AND2X2TS U260 ( .A(n205), .B(n5364), .Y(n11) );
  CLKBUFX2TS U261 ( .A(n6112), .Y(n736) );
  CLKBUFX2TS U262 ( .A(n6143), .Y(n870) );
  OR3X1TS U263 ( .A(n6299), .B(n214), .C(n5538), .Y(n13) );
  OR3X1TS U264 ( .A(n349), .B(n257), .C(n443), .Y(n17) );
  XOR2X1TS U265 ( .A(n5355), .B(n14), .Y(n20) );
  AND2X2TS U266 ( .A(n6), .B(n568), .Y(n22) );
  NAND2BX1TS U267 ( .AN(n5378), .B(n5399), .Y(n5546) );
  INVX2TS U268 ( .A(n13), .Y(n376) );
  CLKINVX2TS U269 ( .A(n376), .Y(n274) );
  CLKINVX2TS U270 ( .A(n332), .Y(n333) );
  OR2X2TS U271 ( .A(n6239), .B(n18), .Y(n23) );
  INVXLTS U272 ( .A(n189), .Y(n159) );
  CLKBUFX2TS U273 ( .A(readReady), .Y(n160) );
  CLKBUFX2TS U274 ( .A(selectBit_WEST), .Y(n161) );
  INVXLTS U275 ( .A(n6243), .Y(n162) );
  CLKBUFX2TS U276 ( .A(selectBit_NORTH), .Y(n163) );
  INVXLTS U277 ( .A(readRequesterAddress[0]), .Y(n164) );
  INVXLTS U278 ( .A(n164), .Y(n165) );
  INVXLTS U279 ( .A(n164), .Y(n166) );
  INVXLTS U280 ( .A(n164), .Y(n167) );
  INVXLTS U281 ( .A(n164), .Y(n168) );
  INVXLTS U282 ( .A(readRequesterAddress[1]), .Y(n169) );
  INVXLTS U283 ( .A(n169), .Y(n170) );
  INVXLTS U284 ( .A(n169), .Y(n171) );
  INVXLTS U285 ( .A(n169), .Y(n172) );
  INVXLTS U286 ( .A(n169), .Y(n173) );
  INVXLTS U287 ( .A(readRequesterAddress[2]), .Y(n174) );
  INVXLTS U288 ( .A(n174), .Y(n175) );
  INVXLTS U289 ( .A(n174), .Y(n176) );
  INVXLTS U290 ( .A(n174), .Y(n177) );
  INVXLTS U291 ( .A(n174), .Y(n178) );
  INVXLTS U292 ( .A(readRequesterAddress[3]), .Y(n179) );
  INVXLTS U293 ( .A(n179), .Y(n180) );
  INVXLTS U294 ( .A(n179), .Y(n181) );
  INVXLTS U295 ( .A(n179), .Y(n182) );
  INVXLTS U296 ( .A(n179), .Y(n183) );
  INVXLTS U297 ( .A(readRequesterAddress[4]), .Y(n184) );
  INVXLTS U298 ( .A(n184), .Y(n185) );
  INVXLTS U299 ( .A(n184), .Y(n186) );
  INVXLTS U300 ( .A(n184), .Y(n187) );
  INVXLTS U301 ( .A(n184), .Y(n188) );
  INVXLTS U302 ( .A(readRequesterAddress[5]), .Y(n189) );
  INVXLTS U303 ( .A(n189), .Y(n190) );
  INVXLTS U304 ( .A(n189), .Y(n191) );
  INVXLTS U305 ( .A(n189), .Y(n192) );
  INVXLTS U306 ( .A(n8), .Y(n193) );
  INVXLTS U307 ( .A(n10), .Y(n194) );
  INVXLTS U308 ( .A(n6287), .Y(n195) );
  INVXLTS U309 ( .A(n6303), .Y(n196) );
  CLKBUFX2TS U310 ( .A(n6189), .Y(n436) );
  INVX2TS U311 ( .A(n200), .Y(n197) );
  INVXLTS U312 ( .A(n202), .Y(n198) );
  INVX2TS U313 ( .A(n197), .Y(n199) );
  CLKBUFX2TS U314 ( .A(n199), .Y(n201) );
  CLKBUFX2TS U315 ( .A(n199), .Y(n213) );
  CLKINVX2TS U316 ( .A(n200), .Y(n202) );
  INVXLTS U317 ( .A(n202), .Y(n203) );
  INVXLTS U318 ( .A(n202), .Y(n204) );
  INVXLTS U319 ( .A(n18), .Y(n205) );
  CLKBUFX2TS U320 ( .A(n199), .Y(n206) );
  CLKBUFX2TS U321 ( .A(n6189), .Y(n207) );
  CLKBUFX2TS U322 ( .A(n199), .Y(n212) );
  INVXLTS U323 ( .A(n197), .Y(n208) );
  INVXLTS U324 ( .A(n197), .Y(n209) );
  INVXLTS U325 ( .A(n197), .Y(n210) );
  INVXLTS U326 ( .A(n202), .Y(n211) );
  AOI222XLTS U327 ( .A0(n3959), .A1(n3708), .B0(n3441), .B1(n190), .C0(n4116), 
        .C1(n3419), .Y(n5482) );
  CLKBUFX2TS U328 ( .A(n5539), .Y(n214) );
  INVXLTS U329 ( .A(n3), .Y(n215) );
  CLKBUFX2TS U330 ( .A(n5572), .Y(n219) );
  CLKBUFX2TS U331 ( .A(n5520), .Y(n220) );
  INVX2TS U332 ( .A(n12), .Y(n223) );
  INVX1TS U333 ( .A(n12), .Y(n224) );
  INVX2TS U334 ( .A(n5555), .Y(n225) );
  INVXLTS U335 ( .A(n225), .Y(n226) );
  INVXLTS U336 ( .A(n21), .Y(n227) );
  INVXLTS U337 ( .A(n21), .Y(n228) );
  INVXLTS U338 ( .A(n23), .Y(n229) );
  INVXLTS U339 ( .A(n23), .Y(n230) );
  INVXLTS U340 ( .A(n5402), .Y(n231) );
  INVXLTS U341 ( .A(n231), .Y(n232) );
  INVXLTS U342 ( .A(n5458), .Y(n233) );
  INVXLTS U343 ( .A(n233), .Y(n234) );
  INVXLTS U344 ( .A(n20), .Y(n235) );
  INVXLTS U345 ( .A(n20), .Y(n236) );
  INVX2TS U346 ( .A(n5546), .Y(n237) );
  CLKINVX1TS U347 ( .A(n237), .Y(n238) );
  INVXLTS U348 ( .A(n17), .Y(n239) );
  INVXLTS U349 ( .A(n17), .Y(n240) );
  INVXLTS U350 ( .A(n4), .Y(n241) );
  INVXLTS U351 ( .A(n353), .Y(n242) );
  INVXLTS U352 ( .A(n246), .Y(n243) );
  CLKINVX2TS U353 ( .A(n6159), .Y(n244) );
  CLKINVX2TS U354 ( .A(n6159), .Y(n246) );
  INVXLTS U355 ( .A(n246), .Y(n247) );
  INVXLTS U356 ( .A(n3715), .Y(n249) );
  INVXLTS U357 ( .A(n249), .Y(n250) );
  INVXLTS U358 ( .A(n271), .Y(n374) );
  INVXLTS U359 ( .A(n3752), .Y(n251) );
  INVXLTS U360 ( .A(n6309), .Y(n252) );
  CLKINVX2TS U361 ( .A(n4851), .Y(n253) );
  CLKINVX1TS U362 ( .A(n4851), .Y(n6252) );
  INVXLTS U363 ( .A(n425), .Y(n254) );
  INVX2TS U364 ( .A(n434), .Y(n435) );
  INVXLTS U365 ( .A(n6242), .Y(n255) );
  INVXLTS U366 ( .A(n255), .Y(n256) );
  INVXLTS U367 ( .A(n440), .Y(n257) );
  INVXLTS U368 ( .A(n443), .Y(n258) );
  INVXLTS U369 ( .A(n433), .Y(n259) );
  INVXLTS U370 ( .A(n5365), .Y(n260) );
  INVXLTS U371 ( .A(n260), .Y(n261) );
  INVXLTS U372 ( .A(n5506), .Y(n262) );
  INVXLTS U373 ( .A(n262), .Y(n263) );
  INVX1TS U374 ( .A(n4880), .Y(n264) );
  INVXLTS U375 ( .A(n264), .Y(n265) );
  INVXLTS U376 ( .A(n7), .Y(n266) );
  INVXLTS U377 ( .A(n266), .Y(n267) );
  INVXLTS U378 ( .A(n268), .Y(n269) );
  INVXLTS U379 ( .A(n271), .Y(n272) );
  INVXLTS U380 ( .A(n271), .Y(n273) );
  INVXLTS U381 ( .A(n274), .Y(n275) );
  NAND3X1TS U382 ( .A(n6296), .B(n5472), .C(n276), .Y(n5521) );
  INVXLTS U383 ( .A(n5323), .Y(n277) );
  INVX2TS U384 ( .A(n6241), .Y(n278) );
  INVX1TS U385 ( .A(n278), .Y(n279) );
  INVX2TS U386 ( .A(n22), .Y(n280) );
  INVXLTS U387 ( .A(n22), .Y(n281) );
  INVXLTS U388 ( .A(n11), .Y(n282) );
  INVXLTS U389 ( .A(n11), .Y(n283) );
  INVXLTS U390 ( .A(n295), .Y(n284) );
  INVXLTS U391 ( .A(n284), .Y(n285) );
  INVXLTS U392 ( .A(n284), .Y(n286) );
  INVXLTS U393 ( .A(n5295), .Y(n287) );
  INVXLTS U394 ( .A(n287), .Y(n288) );
  INVXLTS U395 ( .A(n15), .Y(n289) );
  INVXLTS U396 ( .A(n3752), .Y(n290) );
  INVXLTS U397 ( .A(n290), .Y(n291) );
  INVXLTS U398 ( .A(n290), .Y(n292) );
  INVXLTS U399 ( .A(n4), .Y(n293) );
  INVXLTS U400 ( .A(n274), .Y(n294) );
  INVXLTS U401 ( .A(n13), .Y(n295) );
  INVXLTS U402 ( .A(n251), .Y(n296) );
  INVXLTS U403 ( .A(n378), .Y(n297) );
  INVXLTS U404 ( .A(n297), .Y(n298) );
  INVXLTS U405 ( .A(n252), .Y(n299) );
  INVXLTS U406 ( .A(n6244), .Y(n300) );
  INVXLTS U407 ( .A(n300), .Y(n301) );
  INVXLTS U408 ( .A(n300), .Y(n302) );
  INVXLTS U409 ( .A(destinationAddressIn_NORTH[6]), .Y(n303) );
  INVXLTS U410 ( .A(destinationAddressIn_NORTH[6]), .Y(n304) );
  INVXLTS U411 ( .A(destinationAddressIn_NORTH[6]), .Y(n305) );
  INVXLTS U412 ( .A(n6245), .Y(n306) );
  INVXLTS U413 ( .A(n306), .Y(n307) );
  INVXLTS U414 ( .A(n306), .Y(n308) );
  INVXLTS U415 ( .A(n6250), .Y(n309) );
  INVXLTS U416 ( .A(n309), .Y(n310) );
  INVXLTS U417 ( .A(n309), .Y(n311) );
  INVXLTS U418 ( .A(n6248), .Y(n312) );
  INVXLTS U419 ( .A(n312), .Y(n313) );
  INVXLTS U420 ( .A(n312), .Y(n314) );
  INVXLTS U421 ( .A(n6247), .Y(n315) );
  INVXLTS U422 ( .A(n315), .Y(n316) );
  INVXLTS U423 ( .A(n315), .Y(n317) );
  INVXLTS U424 ( .A(n6251), .Y(n318) );
  INVXLTS U425 ( .A(n318), .Y(n319) );
  INVXLTS U426 ( .A(n318), .Y(n320) );
  INVXLTS U427 ( .A(n6249), .Y(n321) );
  INVXLTS U428 ( .A(n321), .Y(n322) );
  INVXLTS U429 ( .A(n321), .Y(n323) );
  INVXLTS U430 ( .A(n6246), .Y(n324) );
  INVXLTS U431 ( .A(n324), .Y(n325) );
  INVXLTS U432 ( .A(n324), .Y(n326) );
  INVXLTS U433 ( .A(n5589), .Y(n327) );
  INVXLTS U434 ( .A(n327), .Y(n328) );
  INVXLTS U435 ( .A(n327), .Y(n329) );
  INVXLTS U436 ( .A(n3778), .Y(n330) );
  INVXLTS U437 ( .A(n3778), .Y(n331) );
  INVX1TS U438 ( .A(n5576), .Y(n332) );
  INVXLTS U439 ( .A(n332), .Y(n334) );
  INVXLTS U440 ( .A(n5585), .Y(n335) );
  INVXLTS U441 ( .A(n335), .Y(n336) );
  INVXLTS U442 ( .A(n335), .Y(n337) );
  CLKBUFX2TS U443 ( .A(n5581), .Y(n338) );
  CLKBUFX2TS U444 ( .A(n5581), .Y(n339) );
  INVXLTS U445 ( .A(n377), .Y(n340) );
  INVXLTS U446 ( .A(n377), .Y(n341) );
  INVXLTS U447 ( .A(n383), .Y(n342) );
  INVXLTS U448 ( .A(n342), .Y(n343) );
  INVXLTS U449 ( .A(n342), .Y(n344) );
  INVXLTS U450 ( .A(n342), .Y(n345) );
  INVXLTS U451 ( .A(n5575), .Y(n346) );
  INVXLTS U452 ( .A(n342), .Y(n347) );
  INVXLTS U453 ( .A(n16), .Y(n348) );
  INVXLTS U454 ( .A(n16), .Y(n349) );
  INVXLTS U455 ( .A(n5364), .Y(n350) );
  INVXLTS U456 ( .A(n5364), .Y(n351) );
  INVX2TS U457 ( .A(n6159), .Y(n353) );
  INVXLTS U458 ( .A(n353), .Y(n354) );
  INVXLTS U459 ( .A(n353), .Y(n355) );
  INVXLTS U460 ( .A(n353), .Y(n356) );
  INVXLTS U461 ( .A(n386), .Y(n358) );
  INVXLTS U462 ( .A(n386), .Y(n360) );
  INVXLTS U463 ( .A(n386), .Y(n361) );
  INVXLTS U464 ( .A(n246), .Y(n362) );
  INVXLTS U465 ( .A(n437), .Y(n363) );
  INVXLTS U466 ( .A(n266), .Y(n364) );
  INVXLTS U467 ( .A(n266), .Y(n365) );
  INVXLTS U468 ( .A(n366), .Y(n367) );
  INVXLTS U469 ( .A(n366), .Y(n368) );
  INVXLTS U470 ( .A(n366), .Y(n369) );
  INVXLTS U471 ( .A(n13), .Y(n370) );
  INVXLTS U472 ( .A(n274), .Y(n371) );
  INVXLTS U473 ( .A(n284), .Y(n372) );
  INVXLTS U474 ( .A(n284), .Y(n373) );
  INVXLTS U475 ( .A(n271), .Y(n375) );
  INVXLTS U476 ( .A(n251), .Y(n378) );
  INVXLTS U477 ( .A(n377), .Y(n379) );
  INVXLTS U478 ( .A(n251), .Y(n380) );
  INVXLTS U479 ( .A(n251), .Y(n381) );
  INVXLTS U480 ( .A(n252), .Y(n382) );
  INVXLTS U481 ( .A(n5575), .Y(n383) );
  INVXLTS U482 ( .A(n252), .Y(n384) );
  INVXLTS U483 ( .A(n252), .Y(n385) );
  INVX2TS U484 ( .A(n6159), .Y(n386) );
  INVX2TS U523 ( .A(selectBit_SOUTH), .Y(n6243) );
  CLKAND2X2TS U524 ( .A(n5558), .B(n6297), .Y(n6188) );
  NOR2BX1TS U525 ( .AN(n235), .B(n5399), .Y(n5555) );
  XOR2X1TS U526 ( .A(n4873), .B(n216), .Y(n4865) );
  NAND3X1TS U527 ( .A(n5494), .B(n5400), .C(n276), .Y(n5542) );
  INVXLTS U528 ( .A(n5527), .Y(n6300) );
  CLKAND2X2TS U529 ( .A(n5530), .B(n6300), .Y(n6130) );
  AND3XLTS U530 ( .A(n226), .B(n5527), .C(n5530), .Y(n6127) );
  OAI2BB1XLTS U531 ( .A0N(n4851), .A1N(n4879), .B0(n4850), .Y(n4862) );
  OAI2BB1X1TS U532 ( .A0N(n4880), .A1N(selectBit_EAST), .B0(n4848), .Y(n4851)
         );
  XOR2X1TS U533 ( .A(n205), .B(n6252), .Y(n5354) );
  XOR2X4TS U534 ( .A(n5329), .B(n216), .Y(n5400) );
  NOR3BX1TS U535 ( .AN(n5472), .B(n276), .C(n444), .Y(n5559) );
  NAND2X1TS U536 ( .A(n5559), .B(n5565), .Y(n6209) );
  INVXLTS U537 ( .A(n5554), .Y(n6297) );
  NAND3X1TS U538 ( .A(n5572), .B(n6289), .C(n5566), .Y(n5589) );
  NOR2X1TS U539 ( .A(n5568), .B(n5569), .Y(n5566) );
  NOR2X2TS U540 ( .A(n6254), .B(n570), .Y(n5355) );
  CLKINVX2TS U541 ( .A(n5), .Y(n425) );
  INVX2TS U542 ( .A(n425), .Y(n426) );
  CLKINVX2TS U543 ( .A(n3721), .Y(n427) );
  INVX2TS U544 ( .A(n427), .Y(n428) );
  CLKINVX2TS U545 ( .A(n3718), .Y(n429) );
  INVX2TS U546 ( .A(n429), .Y(n430) );
  CLKINVX2TS U547 ( .A(n3719), .Y(n431) );
  INVX2TS U548 ( .A(n431), .Y(n432) );
  XNOR2X4TS U549 ( .A(n555), .B(n5331), .Y(n5329) );
  OAI22XLTS U550 ( .A0(n5534), .A1(n350), .B0(n282), .B1(n231), .Y(n433) );
  CLKINVX2TS U551 ( .A(n5532), .Y(n434) );
  NOR3BX1TS U552 ( .AN(n224), .B(n5547), .C(n6291), .Y(n6172) );
  AND3XLTS U553 ( .A(n5523), .B(n228), .C(n5333), .Y(n6112) );
  INVXLTS U554 ( .A(n227), .Y(n6291) );
  CLKINVX2TS U555 ( .A(n3714), .Y(n437) );
  CLKBUFX2TS U556 ( .A(n7), .Y(n3715) );
  OAI22XLTS U557 ( .A0(n220), .A1(n350), .B0(n282), .B1(n6283), .Y(n438) );
  OAI22XLTS U558 ( .A0(n5520), .A1(n351), .B0(n283), .B1(n6283), .Y(n439) );
  CLKBUFX2TS U559 ( .A(n6309), .Y(n3781) );
  CLKBUFX2TS U560 ( .A(n6237), .Y(n441) );
  NOR3XLTS U561 ( .A(n6293), .B(n6298), .C(n442), .Y(n5582) );
  NOR2XLTS U562 ( .A(n5542), .B(n5538), .Y(n6159) );
  NOR3BXLTS U563 ( .AN(n5494), .B(n276), .C(n444), .Y(n5568) );
  OR2X2TS U564 ( .A(n5313), .B(n6256), .Y(n5291) );
  INVX2TS U565 ( .A(n5291), .Y(n445) );
  INVX2TS U566 ( .A(n5291), .Y(n446) );
  CLKBUFX2TS U567 ( .A(n5497), .Y(n447) );
  OAI31XLTS U568 ( .A0(n5497), .A1(n6), .A2(n195), .B0(n196), .Y(n5496) );
  INVX2TS U569 ( .A(n3709), .Y(n448) );
  INVX1TS U570 ( .A(n6209), .Y(n6304) );
  INVX2TS U571 ( .A(n5303), .Y(n449) );
  OAI32XLTS U572 ( .A0(n4877), .A1(n6237), .A2(n4876), .B0(n449), .B1(n157), 
        .Y(N4718) );
  INVX2TS U573 ( .A(n3669), .Y(n450) );
  CLKBUFX2TS U574 ( .A(cacheDataOut[31]), .Y(n451) );
  CLKBUFX2TS U575 ( .A(cacheDataOut[31]), .Y(n452) );
  CLKBUFX2TS U576 ( .A(cacheDataOut[30]), .Y(n453) );
  CLKBUFX2TS U577 ( .A(cacheDataOut[30]), .Y(n454) );
  CLKBUFX2TS U578 ( .A(cacheDataOut[29]), .Y(n455) );
  CLKBUFX2TS U579 ( .A(cacheDataOut[29]), .Y(n456) );
  CLKBUFX2TS U580 ( .A(cacheDataOut[28]), .Y(n457) );
  CLKBUFX2TS U581 ( .A(cacheDataOut[28]), .Y(n458) );
  CLKBUFX2TS U582 ( .A(cacheDataOut[27]), .Y(n459) );
  CLKBUFX2TS U583 ( .A(cacheDataOut[27]), .Y(n460) );
  CLKBUFX2TS U584 ( .A(cacheDataOut[26]), .Y(n461) );
  CLKBUFX2TS U585 ( .A(cacheDataOut[26]), .Y(n462) );
  CLKBUFX2TS U586 ( .A(cacheDataOut[25]), .Y(n463) );
  CLKBUFX2TS U587 ( .A(cacheDataOut[25]), .Y(n464) );
  CLKBUFX2TS U588 ( .A(cacheDataOut[24]), .Y(n465) );
  CLKBUFX2TS U589 ( .A(cacheDataOut[24]), .Y(n466) );
  CLKBUFX2TS U590 ( .A(cacheDataOut[23]), .Y(n467) );
  CLKBUFX2TS U591 ( .A(cacheDataOut[23]), .Y(n468) );
  CLKBUFX2TS U592 ( .A(cacheDataOut[22]), .Y(n469) );
  CLKBUFX2TS U593 ( .A(cacheDataOut[22]), .Y(n470) );
  CLKBUFX2TS U594 ( .A(cacheDataOut[21]), .Y(n471) );
  CLKBUFX2TS U595 ( .A(cacheDataOut[21]), .Y(n472) );
  CLKBUFX2TS U596 ( .A(cacheDataOut[20]), .Y(n473) );
  CLKBUFX2TS U597 ( .A(cacheDataOut[20]), .Y(n474) );
  CLKBUFX2TS U598 ( .A(cacheDataOut[19]), .Y(n475) );
  CLKBUFX2TS U599 ( .A(cacheDataOut[19]), .Y(n476) );
  CLKBUFX2TS U600 ( .A(cacheDataOut[18]), .Y(n477) );
  CLKBUFX2TS U601 ( .A(cacheDataOut[18]), .Y(n478) );
  CLKBUFX2TS U602 ( .A(cacheDataOut[17]), .Y(n479) );
  CLKBUFX2TS U603 ( .A(cacheDataOut[17]), .Y(n480) );
  CLKBUFX2TS U604 ( .A(cacheDataOut[16]), .Y(n481) );
  CLKBUFX2TS U605 ( .A(cacheDataOut[16]), .Y(n482) );
  CLKBUFX2TS U606 ( .A(cacheDataOut[15]), .Y(n483) );
  CLKBUFX2TS U607 ( .A(cacheDataOut[15]), .Y(n484) );
  CLKBUFX2TS U608 ( .A(cacheDataOut[14]), .Y(n485) );
  CLKBUFX2TS U609 ( .A(cacheDataOut[14]), .Y(n486) );
  CLKBUFX2TS U610 ( .A(cacheDataOut[13]), .Y(n487) );
  CLKBUFX2TS U611 ( .A(cacheDataOut[13]), .Y(n488) );
  CLKBUFX2TS U612 ( .A(cacheDataOut[12]), .Y(n489) );
  CLKBUFX2TS U613 ( .A(cacheDataOut[12]), .Y(n490) );
  CLKBUFX2TS U614 ( .A(cacheDataOut[11]), .Y(n491) );
  CLKBUFX2TS U615 ( .A(cacheDataOut[11]), .Y(n492) );
  CLKBUFX2TS U616 ( .A(cacheDataOut[10]), .Y(n493) );
  CLKBUFX2TS U617 ( .A(cacheDataOut[10]), .Y(n494) );
  CLKBUFX2TS U618 ( .A(cacheDataOut[9]), .Y(n495) );
  CLKBUFX2TS U619 ( .A(cacheDataOut[9]), .Y(n496) );
  CLKBUFX2TS U620 ( .A(cacheDataOut[8]), .Y(n501) );
  CLKBUFX2TS U621 ( .A(cacheDataOut[8]), .Y(n503) );
  CLKBUFX2TS U622 ( .A(cacheDataOut[7]), .Y(n505) );
  CLKBUFX2TS U623 ( .A(cacheDataOut[7]), .Y(n507) );
  CLKBUFX2TS U624 ( .A(cacheDataOut[6]), .Y(n508) );
  CLKBUFX2TS U625 ( .A(cacheDataOut[6]), .Y(n509) );
  CLKBUFX2TS U626 ( .A(cacheDataOut[5]), .Y(n510) );
  CLKBUFX2TS U627 ( .A(cacheDataOut[5]), .Y(n511) );
  CLKBUFX2TS U628 ( .A(cacheDataOut[4]), .Y(n512) );
  CLKBUFX2TS U629 ( .A(cacheDataOut[4]), .Y(n514) );
  CLKBUFX2TS U630 ( .A(cacheDataOut[3]), .Y(n515) );
  CLKBUFX2TS U631 ( .A(cacheDataOut[3]), .Y(n516) );
  CLKBUFX2TS U632 ( .A(cacheDataOut[2]), .Y(n526) );
  CLKBUFX2TS U633 ( .A(cacheDataOut[2]), .Y(n531) );
  CLKBUFX2TS U634 ( .A(cacheDataOut[1]), .Y(n536) );
  CLKBUFX2TS U635 ( .A(cacheDataOut[1]), .Y(n537) );
  CLKBUFX2TS U636 ( .A(cacheDataOut[0]), .Y(n541) );
  CLKBUFX2TS U637 ( .A(cacheDataOut[0]), .Y(n543) );
  CLKBUFX2TS U638 ( .A(n6226), .Y(n544) );
  CLKBUFX2TS U639 ( .A(n6226), .Y(n545) );
  CLKBUFX2TS U640 ( .A(n5582), .Y(n546) );
  CLKBUFX2TS U641 ( .A(n5582), .Y(n548) );
  CLKBUFX2TS U642 ( .A(n2), .Y(n551) );
  CLKBUFX2TS U643 ( .A(n2), .Y(n554) );
  INVXLTS U644 ( .A(n2), .Y(n6311) );
  NOR3XLTS U645 ( .A(n238), .B(n6302), .C(n6310), .Y(n5573) );
  CLKBUFX2TS U646 ( .A(n5323), .Y(n555) );
  CLKAND2X2TS U647 ( .A(n5537), .B(n5471), .Y(n6145) );
  CLKBUFX2TS U648 ( .A(n6243), .Y(n556) );
  NOR3X1TS U649 ( .A(n6286), .B(n5327), .C(n6253), .Y(n4869) );
  INVX1TS U650 ( .A(n5582), .Y(n6305) );
  CLKBUFX2TS U651 ( .A(n6311), .Y(n3796) );
  NAND2X1TS U652 ( .A(n5520), .B(n5333), .Y(n5576) );
  CLKINVX2TS U653 ( .A(n5543), .Y(n6293) );
  AND2XLTS U654 ( .A(n5568), .B(n219), .Y(n6220) );
  INVX2TS U655 ( .A(n3224), .Y(n558) );
  AND2XLTS U656 ( .A(n5569), .B(n5572), .Y(n6223) );
  NOR2X1TS U657 ( .A(n5531), .B(n5495), .Y(n5562) );
  INVXLTS U658 ( .A(n3214), .Y(n3209) );
  INVXLTS U659 ( .A(n3213), .Y(n3210) );
  INVXLTS U660 ( .A(n3212), .Y(n3211) );
  CLKBUFX2TS U661 ( .A(n853), .Y(n850) );
  CLKBUFX2TS U662 ( .A(n3546), .Y(n3543) );
  CLKBUFX2TS U663 ( .A(n702), .Y(n699) );
  CLKBUFX2TS U664 ( .A(n702), .Y(n698) );
  CLKBUFX2TS U665 ( .A(n853), .Y(n851) );
  CLKBUFX2TS U666 ( .A(n3415), .Y(n3412) );
  CLKBUFX2TS U667 ( .A(n3349), .Y(n3346) );
  CLKBUFX2TS U668 ( .A(n3415), .Y(n3413) );
  CLKBUFX2TS U669 ( .A(n3349), .Y(n3347) );
  AND2XLTS U670 ( .A(n435), .B(n5537), .Y(n560) );
  NOR2XLTS U671 ( .A(n6291), .B(n236), .Y(n5471) );
  INVX1TS U672 ( .A(n5578), .Y(n6308) );
  OR2XLTS U673 ( .A(n442), .B(n6288), .Y(n559) );
  CLKBUFX2TS U674 ( .A(n685), .Y(n680) );
  AND3XLTS U675 ( .A(n5472), .B(n5400), .C(n6295), .Y(n5532) );
  NAND3XLTS U676 ( .A(n5494), .B(n5447), .C(n6296), .Y(n5554) );
  NAND3XLTS U677 ( .A(n444), .B(n5494), .C(n6295), .Y(n5527) );
  NAND2XLTS U678 ( .A(n5399), .B(n5378), .Y(n5531) );
  NAND2XLTS U679 ( .A(n228), .B(n235), .Y(n5425) );
  AND2XLTS U680 ( .A(n5562), .B(n5565), .Y(n6204) );
  AND2XLTS U681 ( .A(n5561), .B(n158), .Y(n6206) );
  AND2XLTS U682 ( .A(n5572), .B(n5567), .Y(n6221) );
  NOR2X1TS U683 ( .A(n277), .B(n15), .Y(n5365) );
  AOI221X2TS U684 ( .A0(n6294), .A1(n5401), .B0(n289), .B1(n5471), .C0(n5532), 
        .Y(n5534) );
  INVX1TS U685 ( .A(n5531), .Y(n6294) );
  NOR2X1TS U686 ( .A(n5354), .B(n6240), .Y(n5472) );
  AOI32XLTS U687 ( .A0(n222), .A1(n5557), .A2(n5556), .B0(n3414), .B1(n32), 
        .Y(n2568) );
  AOI32XLTS U688 ( .A0(n226), .A1(n5554), .A2(n3820), .B0(n5553), .B1(n5552), 
        .Y(n5556) );
  AOI32XLTS U689 ( .A0(n221), .A1(n5529), .A2(n5528), .B0(n850), .B1(n25), .Y(
        n2564) );
  AOI32XLTS U690 ( .A0(n226), .A1(n5527), .A2(n3821), .B0(n5526), .B1(n5552), 
        .Y(n5528) );
  INVX2TS U691 ( .A(n5364), .Y(n6303) );
  AND2XLTS U692 ( .A(n265), .B(n4878), .Y(n5322) );
  AND2XLTS U693 ( .A(n4879), .B(n6241), .Y(n4878) );
  NOR2X1TS U694 ( .A(n6239), .B(n5327), .Y(n5497) );
  OAI32XLTS U695 ( .A0(n3822), .A1(n435), .A2(n5531), .B0(n6292), .B1(n256), 
        .Y(n5533) );
  NOR2X1TS U696 ( .A(n289), .B(n568), .Y(n5506) );
  NOR2X1TS U697 ( .A(n15), .B(n569), .Y(n5402) );
  NOR2X1TS U698 ( .A(n277), .B(n289), .Y(n5458) );
  NOR2X1TS U699 ( .A(n348), .B(n5327), .Y(n4853) );
  NOR3X1TS U700 ( .A(n440), .B(n9), .C(n194), .Y(n5294) );
  OAI211XLTS U701 ( .A0(n3210), .A1(n3835), .B0(n5971), .C0(n5970), .Y(n2769)
         );
  OAI211XLTS U702 ( .A0(n3210), .A1(n3832), .B0(n5973), .C0(n5972), .Y(n2770)
         );
  OAI211XLTS U703 ( .A0(n3201), .A1(n3952), .B0(n5394), .C0(n5393), .Y(n2490)
         );
  OAI211XLTS U704 ( .A0(n3202), .A1(n3922), .B0(n5913), .C0(n5912), .Y(n2740)
         );
  OAI211XLTS U705 ( .A0(n3203), .A1(n3919), .B0(n5915), .C0(n5914), .Y(n2741)
         );
  OAI211XLTS U706 ( .A0(n3203), .A1(n3916), .B0(n5917), .C0(n5916), .Y(n2742)
         );
  OAI211XLTS U707 ( .A0(n3203), .A1(n3910), .B0(n5921), .C0(n5920), .Y(n2744)
         );
  OAI211XLTS U708 ( .A0(n3204), .A1(n3907), .B0(n5923), .C0(n5922), .Y(n2745)
         );
  OAI211XLTS U709 ( .A0(n3204), .A1(n3901), .B0(n5927), .C0(n5926), .Y(n2747)
         );
  OAI211XLTS U710 ( .A0(n3205), .A1(n3895), .B0(n5931), .C0(n5930), .Y(n2749)
         );
  OAI211XLTS U711 ( .A0(n3205), .A1(n3892), .B0(n5933), .C0(n5932), .Y(n2750)
         );
  OAI211XLTS U712 ( .A0(n3205), .A1(n3889), .B0(n5935), .C0(n5934), .Y(n2751)
         );
  OAI211XLTS U713 ( .A0(n3205), .A1(n3886), .B0(n5937), .C0(n5936), .Y(n2752)
         );
  OAI211XLTS U714 ( .A0(n3206), .A1(n3883), .B0(n5939), .C0(n5938), .Y(n2753)
         );
  OAI211XLTS U715 ( .A0(n3206), .A1(n3877), .B0(n5943), .C0(n5942), .Y(n2755)
         );
  OAI211XLTS U716 ( .A0(n3206), .A1(n3874), .B0(n5945), .C0(n5944), .Y(n2756)
         );
  OAI211XLTS U717 ( .A0(n3207), .A1(n3871), .B0(n5947), .C0(n5946), .Y(n2757)
         );
  OAI211XLTS U718 ( .A0(n3207), .A1(n3868), .B0(n5949), .C0(n5948), .Y(n2758)
         );
  OAI211XLTS U719 ( .A0(n3207), .A1(n3865), .B0(n5951), .C0(n5950), .Y(n2759)
         );
  OAI211XLTS U720 ( .A0(n3208), .A1(n3859), .B0(n5955), .C0(n5954), .Y(n2761)
         );
  OAI211XLTS U721 ( .A0(n3208), .A1(n3856), .B0(n5957), .C0(n5956), .Y(n2762)
         );
  OAI211XLTS U722 ( .A0(n3208), .A1(n3853), .B0(n5959), .C0(n5958), .Y(n2763)
         );
  OAI211XLTS U723 ( .A0(n3209), .A1(n3847), .B0(n5963), .C0(n5962), .Y(n2765)
         );
  OAI211XLTS U724 ( .A0(n3209), .A1(n3844), .B0(n5965), .C0(n5964), .Y(n2766)
         );
  OAI211XLTS U725 ( .A0(n3209), .A1(n3841), .B0(n5967), .C0(n5966), .Y(n2767)
         );
  OAI211XLTS U726 ( .A0(n3201), .A1(n3961), .B0(n5388), .C0(n5387), .Y(n2487)
         );
  OAI211XLTS U727 ( .A0(n3201), .A1(n3958), .B0(n5390), .C0(n5389), .Y(n2488)
         );
  OAI211XLTS U728 ( .A0(n3201), .A1(n3955), .B0(n5392), .C0(n5391), .Y(n2489)
         );
  OAI211XLTS U729 ( .A0(n3202), .A1(n3949), .B0(n5396), .C0(n5395), .Y(n2491)
         );
  OAI211XLTS U730 ( .A0(n3202), .A1(n3946), .B0(n5398), .C0(n5397), .Y(n2492)
         );
  OAI211XLTS U731 ( .A0(n3203), .A1(n3913), .B0(n5919), .C0(n5918), .Y(n2743)
         );
  OAI211XLTS U732 ( .A0(n3207), .A1(n3862), .B0(n5953), .C0(n5952), .Y(n2760)
         );
  OAI211XLTS U733 ( .A0(n3202), .A1(n3925), .B0(n5911), .C0(n5910), .Y(n2739)
         );
  OAI211XLTS U734 ( .A0(n3204), .A1(n3904), .B0(n5925), .C0(n5924), .Y(n2746)
         );
  OAI211XLTS U735 ( .A0(n3204), .A1(n3898), .B0(n5929), .C0(n5928), .Y(n2748)
         );
  OAI211XLTS U736 ( .A0(n3206), .A1(n3880), .B0(n5941), .C0(n5940), .Y(n2754)
         );
  OAI211XLTS U737 ( .A0(n3208), .A1(n3850), .B0(n5961), .C0(n5960), .Y(n2764)
         );
  OAI211XLTS U738 ( .A0(n3209), .A1(n3838), .B0(n5969), .C0(n5968), .Y(n2768)
         );
  OAI211XLTS U739 ( .A0(n4099), .A1(n3789), .B0(n6103), .C0(n6102), .Y(n2835)
         );
  OAI211XLTS U740 ( .A0(n4096), .A1(n3789), .B0(n6105), .C0(n6104), .Y(n2836)
         );
  OAI211XLTS U741 ( .A0(n4093), .A1(n3790), .B0(n6107), .C0(n6106), .Y(n2837)
         );
  OAI211XLTS U742 ( .A0(n4090), .A1(n3790), .B0(n6109), .C0(n6108), .Y(n2838)
         );
  OAI211XLTS U743 ( .A0(n4087), .A1(n3790), .B0(n6111), .C0(n6110), .Y(n2839)
         );
  OAI211XLTS U744 ( .A0(n4084), .A1(n3790), .B0(n6116), .C0(n6115), .Y(n2840)
         );
  OAI211XLTS U745 ( .A0(n3940), .A1(n3210), .B0(n6136), .C0(n6135), .Y(n2848)
         );
  OAI211XLTS U746 ( .A0(n3943), .A1(n3210), .B0(n6134), .C0(n6133), .Y(n2847)
         );
  OAI211XLTS U747 ( .A0(n3931), .A1(n3211), .B0(n6142), .C0(n6141), .Y(n2851)
         );
  OAI211XLTS U748 ( .A0(n3928), .A1(n3211), .B0(n6147), .C0(n6146), .Y(n2852)
         );
  OAI211XLTS U749 ( .A0(n3937), .A1(n3211), .B0(n6138), .C0(n6137), .Y(n2849)
         );
  OAI211XLTS U750 ( .A0(n3934), .A1(n3211), .B0(n6140), .C0(n6139), .Y(n2850)
         );
  OAI211XLTS U751 ( .A0(n3789), .A1(n3991), .B0(n6099), .C0(n6098), .Y(n2833)
         );
  OAI211XLTS U752 ( .A0(n3789), .A1(n3988), .B0(n6101), .C0(n6100), .Y(n2834)
         );
  OAI211XLTS U753 ( .A0(n3783), .A1(n4117), .B0(n5343), .C0(n5342), .Y(n2459)
         );
  OAI211XLTS U754 ( .A0(n3783), .A1(n4111), .B0(n5347), .C0(n5346), .Y(n2461)
         );
  OAI211XLTS U755 ( .A0(n3783), .A1(n4108), .B0(n5349), .C0(n5348), .Y(n2462)
         );
  OAI211XLTS U756 ( .A0(n3784), .A1(n4105), .B0(n5351), .C0(n5350), .Y(n2463)
         );
  OAI211XLTS U757 ( .A0(n3784), .A1(n4081), .B0(n6039), .C0(n6038), .Y(n2803)
         );
  OAI211XLTS U758 ( .A0(n3784), .A1(n4078), .B0(n6041), .C0(n6040), .Y(n2804)
         );
  OAI211XLTS U759 ( .A0(n3785), .A1(n4075), .B0(n6043), .C0(n6042), .Y(n2805)
         );
  OAI211XLTS U760 ( .A0(n3785), .A1(n4066), .B0(n6049), .C0(n6048), .Y(n2808)
         );
  OAI211XLTS U761 ( .A0(n3786), .A1(n4063), .B0(n6051), .C0(n6050), .Y(n2809)
         );
  OAI211XLTS U762 ( .A0(n3786), .A1(n4060), .B0(n6053), .C0(n6052), .Y(n2810)
         );
  OAI211XLTS U763 ( .A0(n3786), .A1(n4054), .B0(n6057), .C0(n6056), .Y(n2812)
         );
  OAI211XLTS U764 ( .A0(n3787), .A1(n4051), .B0(n6059), .C0(n6058), .Y(n2813)
         );
  OAI211XLTS U765 ( .A0(n3787), .A1(n4045), .B0(n6063), .C0(n6062), .Y(n2815)
         );
  OAI211XLTS U766 ( .A0(n3787), .A1(n4042), .B0(n6065), .C0(n6064), .Y(n2816)
         );
  OAI211XLTS U767 ( .A0(n3793), .A1(n4039), .B0(n6067), .C0(n6066), .Y(n2817)
         );
  OAI211XLTS U768 ( .A0(n3794), .A1(n4036), .B0(n6069), .C0(n6068), .Y(n2818)
         );
  OAI211XLTS U769 ( .A0(n3796), .A1(n4033), .B0(n6071), .C0(n6070), .Y(n2819)
         );
  OAI211XLTS U770 ( .A0(n3791), .A1(n4030), .B0(n6073), .C0(n6072), .Y(n2820)
         );
  OAI211XLTS U771 ( .A0(n3792), .A1(n4027), .B0(n6075), .C0(n6074), .Y(n2821)
         );
  OAI211XLTS U772 ( .A0(n3795), .A1(n4024), .B0(n6077), .C0(n6076), .Y(n2822)
         );
  OAI211XLTS U773 ( .A0(n3792), .A1(n4021), .B0(n6079), .C0(n6078), .Y(n2823)
         );
  OAI211XLTS U774 ( .A0(n3796), .A1(n4018), .B0(n6081), .C0(n6080), .Y(n2824)
         );
  OAI211XLTS U775 ( .A0(n3796), .A1(n4012), .B0(n6085), .C0(n6084), .Y(n2826)
         );
  OAI211XLTS U776 ( .A0(n3794), .A1(n4009), .B0(n6087), .C0(n6086), .Y(n2827)
         );
  OAI211XLTS U777 ( .A0(n3793), .A1(n4006), .B0(n6089), .C0(n6088), .Y(n2828)
         );
  OAI211XLTS U778 ( .A0(n3788), .A1(n4000), .B0(n6093), .C0(n6092), .Y(n2830)
         );
  OAI211XLTS U779 ( .A0(n3788), .A1(n3997), .B0(n6095), .C0(n6094), .Y(n2831)
         );
  OAI211XLTS U780 ( .A0(n3783), .A1(n4114), .B0(n5345), .C0(n5344), .Y(n2460)
         );
  OAI211XLTS U781 ( .A0(n3784), .A1(n4102), .B0(n5353), .C0(n5352), .Y(n2464)
         );
  OAI211XLTS U782 ( .A0(n3785), .A1(n4072), .B0(n6045), .C0(n6044), .Y(n2806)
         );
  OAI211XLTS U783 ( .A0(n3785), .A1(n4069), .B0(n6047), .C0(n6046), .Y(n2807)
         );
  OAI211XLTS U784 ( .A0(n3786), .A1(n4057), .B0(n6055), .C0(n6054), .Y(n2811)
         );
  OAI211XLTS U785 ( .A0(n3787), .A1(n4048), .B0(n6061), .C0(n6060), .Y(n2814)
         );
  OAI211XLTS U786 ( .A0(n3794), .A1(n4015), .B0(n6083), .C0(n6082), .Y(n2825)
         );
  OAI211XLTS U787 ( .A0(n3788), .A1(n4003), .B0(n6091), .C0(n6090), .Y(n2829)
         );
  OAI211XLTS U788 ( .A0(n3788), .A1(n3994), .B0(n6097), .C0(n6096), .Y(n2832)
         );
  OAI32XLTS U789 ( .A0(n3822), .A1(n6302), .A2(n238), .B0(n5521), .B1(n3816), 
        .Y(n5522) );
  AOI22XLTS U790 ( .A0(n5525), .A1(n5524), .B0(n3781), .B1(n33), .Y(n2563) );
  AOI31XLTS U791 ( .A0(n5523), .A1(n228), .A2(readIn_SOUTH), .B0(n5522), .Y(
        n5524) );
  OAI22XLTS U792 ( .A0(n214), .A1(n256), .B0(n6288), .B1(n3829), .Y(n5540) );
  NOR2X1TS U793 ( .A(n4844), .B(n5322), .Y(n5364) );
  NAND2XLTS U794 ( .A(n3815), .B(n435), .Y(n5536) );
  AOI21XLTS U795 ( .A0(n3827), .A1(n5549), .B0(n5548), .Y(n5550) );
  AOI2BB2XLTS U796 ( .B0(readReady), .B1(selectBit_WEST), .A0N(n4879), .A1N(
        n6252), .Y(n4873) );
  OAI211XLTS U797 ( .A0(n3943), .A1(n6209), .B0(n6195), .C0(n6194), .Y(n2871)
         );
  AOI22XLTS U798 ( .A0(n3434), .A1(n159), .B0(n3417), .B1(n4097), .Y(n6195) );
  OAI211XLTS U799 ( .A0(n3940), .A1(n6209), .B0(n6197), .C0(n6196), .Y(n2872)
         );
  OAI211XLTS U800 ( .A0(n3937), .A1(n448), .B0(n6199), .C0(n6198), .Y(n2873)
         );
  OAI211XLTS U801 ( .A0(n3934), .A1(n448), .B0(n6201), .C0(n6200), .Y(n2874)
         );
  OAI211XLTS U802 ( .A0(n3931), .A1(n448), .B0(n6203), .C0(n6202), .Y(n2875)
         );
  OAI211XLTS U803 ( .A0(n3928), .A1(n448), .B0(n6208), .C0(n6207), .Y(n2876)
         );
  AOI22XLTS U804 ( .A0(n3433), .A1(n166), .B0(n3417), .B1(n4082), .Y(n6208) );
  OAI211XLTS U805 ( .A0(n3530), .A1(n30), .B0(n6215), .C0(n6214), .Y(n2879) );
  OAI211XLTS U806 ( .A0(n3529), .A1(n29), .B0(n6219), .C0(n6218), .Y(n2881) );
  OAI211XLTS U807 ( .A0(n3530), .A1(n26), .B0(n6211), .C0(n6210), .Y(n2877) );
  OAI211XLTS U808 ( .A0(n3529), .A1(n27), .B0(n6213), .C0(n6212), .Y(n2878) );
  OAI211XLTS U809 ( .A0(n3529), .A1(n28), .B0(n6217), .C0(n6216), .Y(n2880) );
  OAI211XLTS U810 ( .A0(n3530), .A1(n31), .B0(n6225), .C0(n6224), .Y(n2882) );
  OAI211XLTS U811 ( .A0(n3399), .A1(n6274), .B0(n6183), .C0(n6182), .Y(n2867)
         );
  OAI211XLTS U812 ( .A0(n3398), .A1(n6275), .B0(n6185), .C0(n6184), .Y(n2868)
         );
  OAI211XLTS U813 ( .A0(n3398), .A1(n6276), .B0(n6187), .C0(n6186), .Y(n2869)
         );
  OAI211XLTS U814 ( .A0(n3399), .A1(n6272), .B0(n6179), .C0(n6178), .Y(n2865)
         );
  OAI211XLTS U815 ( .A0(n3398), .A1(n6273), .B0(n6181), .C0(n6180), .Y(n2866)
         );
  OAI211XLTS U816 ( .A0(n3399), .A1(n6277), .B0(n6193), .C0(n6192), .Y(n2870)
         );
  OAI211XLTS U817 ( .A0(n3333), .A1(n6259), .B0(n6167), .C0(n6166), .Y(n2861)
         );
  OAI211XLTS U818 ( .A0(n3332), .A1(n6260), .B0(n6169), .C0(n6168), .Y(n2862)
         );
  OAI211XLTS U819 ( .A0(n3332), .A1(n6261), .B0(n6171), .C0(n6170), .Y(n2863)
         );
  OAI211XLTS U820 ( .A0(n3333), .A1(n6262), .B0(n6177), .C0(n6176), .Y(n2864)
         );
  OAI211XLTS U821 ( .A0(n3333), .A1(n6269), .B0(n6163), .C0(n6162), .Y(n2859)
         );
  OAI211XLTS U822 ( .A0(n3332), .A1(n6270), .B0(n6165), .C0(n6164), .Y(n2860)
         );
  OAI211XLTS U823 ( .A0(n837), .A1(n6265), .B0(n6122), .C0(n6121), .Y(n2843)
         );
  OAI211XLTS U824 ( .A0(n836), .A1(n6266), .B0(n6124), .C0(n6123), .Y(n2844)
         );
  OAI211XLTS U825 ( .A0(n836), .A1(n6267), .B0(n6126), .C0(n6125), .Y(n2845)
         );
  OAI211XLTS U826 ( .A0(n837), .A1(n6263), .B0(n6118), .C0(n6117), .Y(n2841)
         );
  OAI211XLTS U827 ( .A0(n836), .A1(n6264), .B0(n6120), .C0(n6119), .Y(n2842)
         );
  OAI211XLTS U828 ( .A0(n837), .A1(n6268), .B0(n6132), .C0(n6131), .Y(n2846)
         );
  OAI211XLTS U829 ( .A0(n4099), .A1(n3744), .B0(n6149), .C0(n6148), .Y(n2853)
         );
  OAI211XLTS U830 ( .A0(n4093), .A1(n3745), .B0(n6153), .C0(n6152), .Y(n2855)
         );
  OAI211XLTS U831 ( .A0(n4090), .A1(n3745), .B0(n6155), .C0(n6154), .Y(n2856)
         );
  OAI211XLTS U832 ( .A0(n4087), .A1(n3745), .B0(n6157), .C0(n6156), .Y(n2857)
         );
  OAI211XLTS U833 ( .A0(n4084), .A1(n3745), .B0(n6161), .C0(n6160), .Y(n2858)
         );
  OAI211XLTS U834 ( .A0(n4096), .A1(n3744), .B0(n6151), .C0(n6150), .Y(n2854)
         );
  OAI211XLTS U835 ( .A0(n4733), .A1(n3542), .B0(n5511), .C0(n5510), .Y(n2558)
         );
  INVXLTS U836 ( .A(n3544), .Y(n3542) );
  OAI211XLTS U837 ( .A0(n4454), .A1(n695), .B0(n5659), .C0(n5658), .Y(n2613)
         );
  OAI211XLTS U838 ( .A0(n4504), .A1(n694), .B0(n5671), .C0(n5670), .Y(n2619)
         );
  OAI211XLTS U839 ( .A0(n4524), .A1(n693), .B0(n5675), .C0(n5674), .Y(n2621)
         );
  OAI211XLTS U840 ( .A0(n4531), .A1(n693), .B0(n5677), .C0(n5676), .Y(n2622)
         );
  OAI211XLTS U841 ( .A0(n4598), .A1(n691), .B0(n5691), .C0(n5690), .Y(n2629)
         );
  OAI211XLTS U842 ( .A0(n4609), .A1(n691), .B0(n5693), .C0(n5692), .Y(n2630)
         );
  OAI211XLTS U843 ( .A0(n4621), .A1(n690), .B0(n5697), .C0(n5696), .Y(n2632)
         );
  OAI211XLTS U844 ( .A0(n4657), .A1(n689), .B0(n5705), .C0(n5704), .Y(n2636)
         );
  OAI211XLTS U845 ( .A0(n4704), .A1(n688), .B0(n5715), .C0(n5714), .Y(n2641)
         );
  AOI22XLTS U846 ( .A0(n4145), .A1(n3447), .B0(n4302), .B1(n367), .Y(n5715) );
  OAI211XLTS U847 ( .A0(n4435), .A1(n696), .B0(n5655), .C0(n5654), .Y(n2611)
         );
  OAI211XLTS U848 ( .A0(n4446), .A1(n696), .B0(n5657), .C0(n5656), .Y(n2612)
         );
  OAI211XLTS U849 ( .A0(n4462), .A1(n695), .B0(n5661), .C0(n5660), .Y(n2614)
         );
  OAI211XLTS U850 ( .A0(n4471), .A1(n695), .B0(n5663), .C0(n5662), .Y(n2615)
         );
  OAI211XLTS U851 ( .A0(n4482), .A1(n695), .B0(n5665), .C0(n5664), .Y(n2616)
         );
  OAI211XLTS U852 ( .A0(n4502), .A1(n694), .B0(n5669), .C0(n5668), .Y(n2618)
         );
  OAI211XLTS U853 ( .A0(n4520), .A1(n694), .B0(n5673), .C0(n5672), .Y(n2620)
         );
  OAI211XLTS U854 ( .A0(n4543), .A1(n693), .B0(n5679), .C0(n5678), .Y(n2623)
         );
  OAI211XLTS U855 ( .A0(n4565), .A1(n692), .B0(n5683), .C0(n5682), .Y(n2625)
         );
  OAI211XLTS U856 ( .A0(n4570), .A1(n692), .B0(n5685), .C0(n5684), .Y(n2626)
         );
  OAI211XLTS U857 ( .A0(n4583), .A1(n692), .B0(n5687), .C0(n5686), .Y(n2627)
         );
  OAI211XLTS U858 ( .A0(n4590), .A1(n691), .B0(n5689), .C0(n5688), .Y(n2628)
         );
  OAI211XLTS U859 ( .A0(n4619), .A1(n691), .B0(n5695), .C0(n5694), .Y(n2631)
         );
  OAI211XLTS U860 ( .A0(n4635), .A1(n690), .B0(n5699), .C0(n5698), .Y(n2633)
         );
  OAI211XLTS U861 ( .A0(n4646), .A1(n690), .B0(n5701), .C0(n5700), .Y(n2634)
         );
  OAI211XLTS U862 ( .A0(n4651), .A1(n690), .B0(n5703), .C0(n5702), .Y(n2635)
         );
  OAI211XLTS U863 ( .A0(n4669), .A1(n689), .B0(n5707), .C0(n5706), .Y(n2637)
         );
  OAI211XLTS U864 ( .A0(n4685), .A1(n689), .B0(n5711), .C0(n5710), .Y(n2639)
         );
  OAI211XLTS U865 ( .A0(n4700), .A1(n688), .B0(n5713), .C0(n5712), .Y(n2640)
         );
  OAI211XLTS U866 ( .A0(n4716), .A1(n693), .B0(n5717), .C0(n5716), .Y(n2642)
         );
  AOI22XLTS U867 ( .A0(n4142), .A1(n3447), .B0(n4299), .B1(n267), .Y(n5717) );
  OAI211XLTS U868 ( .A0(n4492), .A1(n694), .B0(n5667), .C0(n5666), .Y(n2617)
         );
  OAI211XLTS U869 ( .A0(n4555), .A1(n692), .B0(n5681), .C0(n5680), .Y(n2624)
         );
  OAI211XLTS U870 ( .A0(n4681), .A1(n689), .B0(n5709), .C0(n5708), .Y(n2638)
         );
  OAI211XLTS U871 ( .A0(n4728), .A1(n688), .B0(n5483), .C0(n5482), .Y(n2543)
         );
  OAI211XLTS U872 ( .A0(n4731), .A1(n3532), .B0(n5509), .C0(n5508), .Y(n2557)
         );
  OAI211XLTS U873 ( .A0(n4437), .A1(n3540), .B0(n5591), .C0(n5590), .Y(n2579)
         );
  OAI211XLTS U874 ( .A0(n4442), .A1(n3540), .B0(n5593), .C0(n5592), .Y(n2580)
         );
  OAI211XLTS U875 ( .A0(n4451), .A1(n3540), .B0(n5595), .C0(n5594), .Y(n2581)
         );
  OAI211XLTS U876 ( .A0(n4464), .A1(n3540), .B0(n5597), .C0(n5596), .Y(n2582)
         );
  OAI211XLTS U877 ( .A0(n4473), .A1(n3539), .B0(n5599), .C0(n5598), .Y(n2583)
         );
  OAI211XLTS U878 ( .A0(n4480), .A1(n3539), .B0(n5601), .C0(n5600), .Y(n2584)
         );
  OAI211XLTS U879 ( .A0(n4489), .A1(n3539), .B0(n5603), .C0(n5602), .Y(n2585)
         );
  OAI211XLTS U880 ( .A0(n4498), .A1(n3539), .B0(n5605), .C0(n5604), .Y(n2586)
         );
  OAI211XLTS U881 ( .A0(n4509), .A1(n3538), .B0(n5607), .C0(n5606), .Y(n2587)
         );
  OAI211XLTS U882 ( .A0(n4514), .A1(n3538), .B0(n5609), .C0(n5608), .Y(n2588)
         );
  OAI211XLTS U883 ( .A0(n4529), .A1(n3538), .B0(n5611), .C0(n5610), .Y(n2589)
         );
  OAI211XLTS U884 ( .A0(n4534), .A1(n3538), .B0(n5613), .C0(n5612), .Y(n2590)
         );
  OAI211XLTS U885 ( .A0(n4547), .A1(n3537), .B0(n5615), .C0(n5614), .Y(n2591)
         );
  OAI211XLTS U886 ( .A0(n4550), .A1(n3537), .B0(n5617), .C0(n5616), .Y(n2592)
         );
  OAI211XLTS U887 ( .A0(n4561), .A1(n3537), .B0(n5619), .C0(n5618), .Y(n2593)
         );
  OAI211XLTS U888 ( .A0(n4572), .A1(n3537), .B0(n5621), .C0(n5620), .Y(n2594)
         );
  OAI211XLTS U889 ( .A0(n4577), .A1(n3536), .B0(n5623), .C0(n5622), .Y(n2595)
         );
  OAI211XLTS U890 ( .A0(n4592), .A1(n3536), .B0(n5625), .C0(n5624), .Y(n2596)
         );
  OAI211XLTS U891 ( .A0(n4595), .A1(n3536), .B0(n5627), .C0(n5626), .Y(n2597)
         );
  OAI211XLTS U892 ( .A0(n4604), .A1(n3535), .B0(n5629), .C0(n5628), .Y(n2598)
         );
  OAI211XLTS U893 ( .A0(n4615), .A1(n3535), .B0(n5631), .C0(n5630), .Y(n2599)
         );
  OAI211XLTS U894 ( .A0(n4628), .A1(n3535), .B0(n5633), .C0(n5632), .Y(n2600)
         );
  OAI211XLTS U895 ( .A0(n4637), .A1(n3535), .B0(n5635), .C0(n5634), .Y(n2601)
         );
  OAI211XLTS U896 ( .A0(n4642), .A1(n3534), .B0(n5637), .C0(n5636), .Y(n2602)
         );
  OAI211XLTS U897 ( .A0(n4649), .A1(n3534), .B0(n5639), .C0(n5638), .Y(n2603)
         );
  OAI211XLTS U898 ( .A0(n4664), .A1(n3536), .B0(n5641), .C0(n5640), .Y(n2604)
         );
  OAI211XLTS U899 ( .A0(n4667), .A1(n3534), .B0(n5643), .C0(n5642), .Y(n2605)
         );
  OAI211XLTS U900 ( .A0(n4676), .A1(n3534), .B0(n5645), .C0(n5644), .Y(n2606)
         );
  OAI211XLTS U901 ( .A0(n4689), .A1(n3533), .B0(n5647), .C0(n5646), .Y(n2607)
         );
  OAI211XLTS U902 ( .A0(n4694), .A1(n3533), .B0(n5649), .C0(n5648), .Y(n2608)
         );
  OAI211XLTS U903 ( .A0(n4707), .A1(n3533), .B0(n5651), .C0(n5650), .Y(n2609)
         );
  OAI211XLTS U904 ( .A0(n4712), .A1(n3533), .B0(n5653), .C0(n5652), .Y(n2610)
         );
  OAI211XLTS U905 ( .A0(n4775), .A1(n3541), .B0(n5519), .C0(n5518), .Y(n2562)
         );
  OAI211XLTS U906 ( .A0(n4743), .A1(n3541), .B0(n5513), .C0(n5512), .Y(n2559)
         );
  OAI211XLTS U907 ( .A0(n4754), .A1(n3541), .B0(n5515), .C0(n5514), .Y(n2560)
         );
  OAI211XLTS U908 ( .A0(n4761), .A1(n3541), .B0(n5517), .C0(n5516), .Y(n2561)
         );
  OAI211XLTS U909 ( .A0(n4436), .A1(n3409), .B0(n5719), .C0(n5718), .Y(n2643)
         );
  OAI211XLTS U910 ( .A0(n4571), .A1(n3406), .B0(n5749), .C0(n5748), .Y(n2658)
         );
  OAI211XLTS U911 ( .A0(n4576), .A1(n3405), .B0(n5751), .C0(n5750), .Y(n2659)
         );
  OAI211XLTS U912 ( .A0(n4614), .A1(n3404), .B0(n5759), .C0(n5758), .Y(n2663)
         );
  OAI211XLTS U913 ( .A0(n4706), .A1(n3402), .B0(n5779), .C0(n5778), .Y(n2673)
         );
  OAI211XLTS U914 ( .A0(n4444), .A1(n3409), .B0(n5721), .C0(n5720), .Y(n2644)
         );
  OAI211XLTS U915 ( .A0(n4455), .A1(n3409), .B0(n5723), .C0(n5722), .Y(n2645)
         );
  OAI211XLTS U916 ( .A0(n4466), .A1(n3409), .B0(n5725), .C0(n5724), .Y(n2646)
         );
  OAI211XLTS U917 ( .A0(n4469), .A1(n3408), .B0(n5727), .C0(n5726), .Y(n2647)
         );
  OAI211XLTS U918 ( .A0(n4478), .A1(n3408), .B0(n5729), .C0(n5728), .Y(n2648)
         );
  OAI211XLTS U919 ( .A0(n4493), .A1(n3408), .B0(n5731), .C0(n5730), .Y(n2649)
         );
  OAI211XLTS U920 ( .A0(n4500), .A1(n3408), .B0(n5733), .C0(n5732), .Y(n2650)
         );
  OAI211XLTS U921 ( .A0(n4507), .A1(n3407), .B0(n5735), .C0(n5734), .Y(n2651)
         );
  OAI211XLTS U922 ( .A0(n4518), .A1(n3407), .B0(n5737), .C0(n5736), .Y(n2652)
         );
  OAI211XLTS U923 ( .A0(n4525), .A1(n3407), .B0(n5739), .C0(n5738), .Y(n2653)
         );
  OAI211XLTS U924 ( .A0(n4532), .A1(n3407), .B0(n5741), .C0(n5740), .Y(n2654)
         );
  OAI211XLTS U925 ( .A0(n4545), .A1(n3406), .B0(n5743), .C0(n5742), .Y(n2655)
         );
  OAI211XLTS U926 ( .A0(n4552), .A1(n3406), .B0(n5745), .C0(n5744), .Y(n2656)
         );
  OAI211XLTS U927 ( .A0(n4563), .A1(n3406), .B0(n5747), .C0(n5746), .Y(n2657)
         );
  OAI211XLTS U928 ( .A0(n4586), .A1(n3405), .B0(n5753), .C0(n5752), .Y(n2660)
         );
  OAI211XLTS U929 ( .A0(n4599), .A1(n3405), .B0(n5755), .C0(n5754), .Y(n2661)
         );
  OAI211XLTS U930 ( .A0(n4608), .A1(n3404), .B0(n5757), .C0(n5756), .Y(n2662)
         );
  OAI211XLTS U931 ( .A0(n4622), .A1(n3404), .B0(n5761), .C0(n5760), .Y(n2664)
         );
  OAI211XLTS U932 ( .A0(n4633), .A1(n3404), .B0(n5763), .C0(n5762), .Y(n2665)
         );
  OAI211XLTS U933 ( .A0(n4644), .A1(n3403), .B0(n5765), .C0(n5764), .Y(n2666)
         );
  OAI211XLTS U934 ( .A0(n4653), .A1(n3403), .B0(n5767), .C0(n5766), .Y(n2667)
         );
  OAI211XLTS U935 ( .A0(n4660), .A1(n3405), .B0(n5769), .C0(n5768), .Y(n2668)
         );
  OAI211XLTS U936 ( .A0(n4673), .A1(n3403), .B0(n5771), .C0(n5770), .Y(n2669)
         );
  OAI211XLTS U937 ( .A0(n4680), .A1(n3403), .B0(n5773), .C0(n5772), .Y(n2670)
         );
  OAI211XLTS U938 ( .A0(n4691), .A1(n3402), .B0(n5775), .C0(n5774), .Y(n2671)
         );
  OAI211XLTS U939 ( .A0(n4696), .A1(n3402), .B0(n5777), .C0(n5776), .Y(n2672)
         );
  OAI211XLTS U940 ( .A0(n4718), .A1(n3402), .B0(n5781), .C0(n5780), .Y(n2674)
         );
  OAI211XLTS U941 ( .A0(n4747), .A1(n3410), .B0(n5464), .C0(n5463), .Y(n2531)
         );
  OAI211XLTS U942 ( .A0(n4756), .A1(n3410), .B0(n5466), .C0(n5465), .Y(n2532)
         );
  OAI211XLTS U943 ( .A0(n4765), .A1(n3410), .B0(n5468), .C0(n5467), .Y(n2533)
         );
  OAI211XLTS U944 ( .A0(n4772), .A1(n3410), .B0(n5470), .C0(n5469), .Y(n2534)
         );
  OAI211XLTS U945 ( .A0(n4726), .A1(n3335), .B0(n5436), .C0(n5435), .Y(n2515)
         );
  OAI211XLTS U946 ( .A0(n4441), .A1(n3343), .B0(n5785), .C0(n5784), .Y(n2676)
         );
  OAI211XLTS U947 ( .A0(n4459), .A1(n3343), .B0(n5789), .C0(n5788), .Y(n2678)
         );
  OAI211XLTS U948 ( .A0(n4470), .A1(n3342), .B0(n5791), .C0(n5790), .Y(n2679)
         );
  OAI211XLTS U949 ( .A0(n4477), .A1(n3342), .B0(n5793), .C0(n5792), .Y(n2680)
         );
  OAI211XLTS U950 ( .A0(n4490), .A1(n3342), .B0(n5795), .C0(n5794), .Y(n2681)
         );
  OAI211XLTS U951 ( .A0(n4495), .A1(n3342), .B0(n5797), .C0(n5796), .Y(n2682)
         );
  OAI211XLTS U952 ( .A0(n4506), .A1(n3341), .B0(n5799), .C0(n5798), .Y(n2683)
         );
  OAI211XLTS U953 ( .A0(n4549), .A1(n3340), .B0(n5809), .C0(n5808), .Y(n2688)
         );
  OAI211XLTS U954 ( .A0(n4594), .A1(n3339), .B0(n5819), .C0(n5818), .Y(n2693)
         );
  OAI211XLTS U955 ( .A0(n4634), .A1(n3338), .B0(n5827), .C0(n5826), .Y(n2697)
         );
  OAI211XLTS U956 ( .A0(n4652), .A1(n3337), .B0(n5831), .C0(n5830), .Y(n2699)
         );
  OAI211XLTS U957 ( .A0(n4668), .A1(n3337), .B0(n5835), .C0(n5834), .Y(n2701)
         );
  OAI211XLTS U958 ( .A0(n4679), .A1(n3337), .B0(n5837), .C0(n5836), .Y(n2702)
         );
  OAI211XLTS U959 ( .A0(n4695), .A1(n3336), .B0(n5841), .C0(n5840), .Y(n2704)
         );
  OAI211XLTS U960 ( .A0(n4433), .A1(n3343), .B0(n5783), .C0(n5782), .Y(n2675)
         );
  OAI211XLTS U961 ( .A0(n4457), .A1(n3343), .B0(n5787), .C0(n5786), .Y(n2677)
         );
  OAI211XLTS U962 ( .A0(n4516), .A1(n3341), .B0(n5801), .C0(n5800), .Y(n2684)
         );
  OAI211XLTS U963 ( .A0(n4527), .A1(n3341), .B0(n5803), .C0(n5802), .Y(n2685)
         );
  OAI211XLTS U964 ( .A0(n4536), .A1(n3341), .B0(n5805), .C0(n5804), .Y(n2686)
         );
  OAI211XLTS U965 ( .A0(n4541), .A1(n3340), .B0(n5807), .C0(n5806), .Y(n2687)
         );
  OAI211XLTS U966 ( .A0(n4568), .A1(n3340), .B0(n5813), .C0(n5812), .Y(n2690)
         );
  OAI211XLTS U967 ( .A0(n4606), .A1(n3338), .B0(n5821), .C0(n5820), .Y(n2694)
         );
  OAI211XLTS U968 ( .A0(n4617), .A1(n3338), .B0(n5823), .C0(n5822), .Y(n2695)
         );
  OAI211XLTS U969 ( .A0(n4624), .A1(n3338), .B0(n5825), .C0(n5824), .Y(n2696)
         );
  OAI211XLTS U970 ( .A0(n4640), .A1(n3337), .B0(n5829), .C0(n5828), .Y(n2698)
         );
  OAI211XLTS U971 ( .A0(n4662), .A1(n3339), .B0(n5833), .C0(n5832), .Y(n2700)
         );
  OAI211XLTS U972 ( .A0(n4703), .A1(n3336), .B0(n5843), .C0(n5842), .Y(n2705)
         );
  OAI211XLTS U973 ( .A0(n4714), .A1(n3336), .B0(n5845), .C0(n5844), .Y(n2706)
         );
  OAI211XLTS U974 ( .A0(n4564), .A1(n3340), .B0(n5811), .C0(n5810), .Y(n2689)
         );
  OAI211XLTS U975 ( .A0(n4582), .A1(n3339), .B0(n5815), .C0(n5814), .Y(n2691)
         );
  OAI211XLTS U976 ( .A0(n4591), .A1(n3339), .B0(n5817), .C0(n5816), .Y(n2692)
         );
  OAI211XLTS U977 ( .A0(n4690), .A1(n3336), .B0(n5839), .C0(n5838), .Y(n2703)
         );
  OAI211XLTS U978 ( .A0(n4742), .A1(n697), .B0(n5487), .C0(n5486), .Y(n2545)
         );
  OAI211XLTS U979 ( .A0(n4753), .A1(n697), .B0(n5489), .C0(n5488), .Y(n2546)
         );
  OAI211XLTS U980 ( .A0(n4762), .A1(n696), .B0(n5491), .C0(n5490), .Y(n2547)
         );
  OAI211XLTS U981 ( .A0(n4771), .A1(n696), .B0(n5493), .C0(n5492), .Y(n2548)
         );
  OAI211XLTS U982 ( .A0(n4746), .A1(n3344), .B0(n5440), .C0(n5439), .Y(n2517)
         );
  OAI211XLTS U983 ( .A0(n4751), .A1(n3344), .B0(n5442), .C0(n5441), .Y(n2518)
         );
  OAI211XLTS U984 ( .A0(n4764), .A1(n3344), .B0(n5444), .C0(n5443), .Y(n2519)
         );
  OAI211XLTS U985 ( .A0(n4769), .A1(n3344), .B0(n5446), .C0(n5445), .Y(n2520)
         );
  OAI211XLTS U986 ( .A0(n4739), .A1(n697), .B0(n5485), .C0(n5484), .Y(n2544)
         );
  OAI211XLTS U987 ( .A0(n4738), .A1(n3411), .B0(n5462), .C0(n5461), .Y(n2530)
         );
  INVXLTS U988 ( .A(n3412), .Y(n3411) );
  OAI211XLTS U989 ( .A0(n4725), .A1(n839), .B0(n5367), .C0(n5366), .Y(n2473)
         );
  OAI211XLTS U990 ( .A0(n4468), .A1(n846), .B0(n5983), .C0(n5982), .Y(n2775)
         );
  OAI211XLTS U991 ( .A0(n4517), .A1(n845), .B0(n5993), .C0(n5992), .Y(n2780)
         );
  OAI211XLTS U992 ( .A0(n4533), .A1(n845), .B0(n5997), .C0(n5996), .Y(n2782)
         );
  OAI211XLTS U993 ( .A0(n4544), .A1(n844), .B0(n5999), .C0(n5998), .Y(n2783)
         );
  OAI211XLTS U994 ( .A0(n4627), .A1(n842), .B0(n6017), .C0(n6016), .Y(n2792)
         );
  OAI211XLTS U995 ( .A0(n4641), .A1(n841), .B0(n6021), .C0(n6020), .Y(n2794)
         );
  OAI211XLTS U996 ( .A0(n4666), .A1(n841), .B0(n6027), .C0(n6026), .Y(n2797)
         );
  OAI211XLTS U997 ( .A0(n4693), .A1(n840), .B0(n6033), .C0(n6032), .Y(n2800)
         );
  OAI211XLTS U998 ( .A0(n4439), .A1(n847), .B0(n5975), .C0(n5974), .Y(n2771)
         );
  OAI211XLTS U999 ( .A0(n4448), .A1(n847), .B0(n5977), .C0(n5976), .Y(n2772)
         );
  OAI211XLTS U1000 ( .A0(n4453), .A1(n847), .B0(n5979), .C0(n5978), .Y(n2773)
         );
  OAI211XLTS U1001 ( .A0(n4460), .A1(n847), .B0(n5981), .C0(n5980), .Y(n2774)
         );
  OAI211XLTS U1002 ( .A0(n4484), .A1(n846), .B0(n5985), .C0(n5984), .Y(n2776)
         );
  OAI211XLTS U1003 ( .A0(n4491), .A1(n846), .B0(n5987), .C0(n5986), .Y(n2777)
         );
  OAI211XLTS U1004 ( .A0(n4496), .A1(n846), .B0(n5989), .C0(n5988), .Y(n2778)
         );
  OAI211XLTS U1005 ( .A0(n4505), .A1(n845), .B0(n5991), .C0(n5990), .Y(n2779)
         );
  OAI211XLTS U1006 ( .A0(n4523), .A1(n845), .B0(n5995), .C0(n5994), .Y(n2781)
         );
  OAI211XLTS U1007 ( .A0(n4556), .A1(n844), .B0(n6001), .C0(n6000), .Y(n2784)
         );
  OAI211XLTS U1008 ( .A0(n4559), .A1(n844), .B0(n6003), .C0(n6002), .Y(n2785)
         );
  OAI211XLTS U1009 ( .A0(n4574), .A1(n844), .B0(n6005), .C0(n6004), .Y(n2786)
         );
  OAI211XLTS U1010 ( .A0(n4581), .A1(n843), .B0(n6007), .C0(n6006), .Y(n2787)
         );
  OAI211XLTS U1011 ( .A0(n4588), .A1(n843), .B0(n6009), .C0(n6008), .Y(n2788)
         );
  OAI211XLTS U1012 ( .A0(n4601), .A1(n843), .B0(n6011), .C0(n6010), .Y(n2789)
         );
  OAI211XLTS U1013 ( .A0(n4610), .A1(n842), .B0(n6013), .C0(n6012), .Y(n2790)
         );
  OAI211XLTS U1014 ( .A0(n4613), .A1(n842), .B0(n6015), .C0(n6014), .Y(n2791)
         );
  OAI211XLTS U1015 ( .A0(n4631), .A1(n842), .B0(n6019), .C0(n6018), .Y(n2793)
         );
  OAI211XLTS U1016 ( .A0(n4655), .A1(n841), .B0(n6023), .C0(n6022), .Y(n2795)
         );
  OAI211XLTS U1017 ( .A0(n4658), .A1(n843), .B0(n6025), .C0(n6024), .Y(n2796)
         );
  OAI211XLTS U1018 ( .A0(n4682), .A1(n841), .B0(n6029), .C0(n6028), .Y(n2798)
         );
  OAI211XLTS U1019 ( .A0(n4687), .A1(n840), .B0(n6031), .C0(n6030), .Y(n2799)
         );
  OAI211XLTS U1020 ( .A0(n4705), .A1(n840), .B0(n6035), .C0(n6034), .Y(n2801)
         );
  OAI211XLTS U1021 ( .A0(n4717), .A1(n840), .B0(n6037), .C0(n6036), .Y(n2802)
         );
  OAI211XLTS U1022 ( .A0(n4737), .A1(n3345), .B0(n5438), .C0(n5437), .Y(n2516)
         );
  INVXLTS U1023 ( .A(n3346), .Y(n3345) );
  OAI211XLTS U1024 ( .A0(n4745), .A1(n848), .B0(n5371), .C0(n5370), .Y(n2475)
         );
  OAI211XLTS U1025 ( .A0(n4758), .A1(n848), .B0(n5373), .C0(n5372), .Y(n2476)
         );
  OAI211XLTS U1026 ( .A0(n4767), .A1(n848), .B0(n5375), .C0(n5374), .Y(n2477)
         );
  OAI211XLTS U1027 ( .A0(n4776), .A1(n848), .B0(n5377), .C0(n5376), .Y(n2478)
         );
  OAI211XLTS U1028 ( .A0(n4734), .A1(n849), .B0(n5369), .C0(n5368), .Y(n2474)
         );
  INVXLTS U1029 ( .A(n851), .Y(n849) );
  OAI211XLTS U1030 ( .A0(n3738), .A1(n4114), .B0(n5416), .C0(n5415), .Y(n2502)
         );
  OAI211XLTS U1031 ( .A0(n3738), .A1(n4111), .B0(n5418), .C0(n5417), .Y(n2503)
         );
  OAI211XLTS U1032 ( .A0(n3738), .A1(n4108), .B0(n5420), .C0(n5419), .Y(n2504)
         );
  OAI211XLTS U1033 ( .A0(n3738), .A1(n4117), .B0(n5414), .C0(n5413), .Y(n2501)
         );
  OAI211XLTS U1034 ( .A0(n3744), .A1(n3991), .B0(n5907), .C0(n5906), .Y(n2737)
         );
  OAI211XLTS U1035 ( .A0(n3744), .A1(n3988), .B0(n5909), .C0(n5908), .Y(n2738)
         );
  OAI211XLTS U1036 ( .A0(n3747), .A1(n4105), .B0(n5422), .C0(n5421), .Y(n2505)
         );
  OAI211XLTS U1037 ( .A0(n3751), .A1(n4102), .B0(n5424), .C0(n5423), .Y(n2506)
         );
  OAI211XLTS U1038 ( .A0(n3746), .A1(n4081), .B0(n5847), .C0(n5846), .Y(n2707)
         );
  OAI211XLTS U1039 ( .A0(n3748), .A1(n4078), .B0(n5849), .C0(n5848), .Y(n2708)
         );
  OAI211XLTS U1040 ( .A0(n3750), .A1(n4075), .B0(n5851), .C0(n5850), .Y(n2709)
         );
  OAI211XLTS U1041 ( .A0(n3746), .A1(n4072), .B0(n5853), .C0(n5852), .Y(n2710)
         );
  OAI211XLTS U1042 ( .A0(n3749), .A1(n4069), .B0(n5855), .C0(n5854), .Y(n2711)
         );
  OAI211XLTS U1043 ( .A0(n3750), .A1(n4066), .B0(n5857), .C0(n5856), .Y(n2712)
         );
  OAI211XLTS U1044 ( .A0(n3748), .A1(n4060), .B0(n5861), .C0(n5860), .Y(n2714)
         );
  OAI211XLTS U1045 ( .A0(n3749), .A1(n4054), .B0(n5865), .C0(n5864), .Y(n2716)
         );
  OAI211XLTS U1046 ( .A0(n3739), .A1(n4051), .B0(n5867), .C0(n5866), .Y(n2717)
         );
  OAI211XLTS U1047 ( .A0(n3739), .A1(n4045), .B0(n5871), .C0(n5870), .Y(n2719)
         );
  OAI211XLTS U1048 ( .A0(n3740), .A1(n4039), .B0(n5875), .C0(n5874), .Y(n2721)
         );
  OAI211XLTS U1049 ( .A0(n3740), .A1(n4036), .B0(n5877), .C0(n5876), .Y(n2722)
         );
  OAI211XLTS U1050 ( .A0(n3740), .A1(n4030), .B0(n5881), .C0(n5880), .Y(n2724)
         );
  OAI211XLTS U1051 ( .A0(n3741), .A1(n4024), .B0(n5885), .C0(n5884), .Y(n2726)
         );
  OAI211XLTS U1052 ( .A0(n3741), .A1(n4021), .B0(n5887), .C0(n5886), .Y(n2727)
         );
  OAI211XLTS U1053 ( .A0(n3741), .A1(n4018), .B0(n5889), .C0(n5888), .Y(n2728)
         );
  OAI211XLTS U1054 ( .A0(n3742), .A1(n4015), .B0(n5891), .C0(n5890), .Y(n2729)
         );
  OAI211XLTS U1055 ( .A0(n3742), .A1(n4012), .B0(n5893), .C0(n5892), .Y(n2730)
         );
  OAI211XLTS U1056 ( .A0(n3742), .A1(n4006), .B0(n5897), .C0(n5896), .Y(n2732)
         );
  OAI211XLTS U1057 ( .A0(n3743), .A1(n3997), .B0(n5903), .C0(n5902), .Y(n2735)
         );
  OAI211XLTS U1058 ( .A0(n3747), .A1(n4063), .B0(n5859), .C0(n5858), .Y(n2713)
         );
  OAI211XLTS U1059 ( .A0(n3749), .A1(n4057), .B0(n5863), .C0(n5862), .Y(n2715)
         );
  OAI211XLTS U1060 ( .A0(n3739), .A1(n4048), .B0(n5869), .C0(n5868), .Y(n2718)
         );
  OAI211XLTS U1061 ( .A0(n3739), .A1(n4042), .B0(n5873), .C0(n5872), .Y(n2720)
         );
  OAI211XLTS U1062 ( .A0(n3740), .A1(n4033), .B0(n5879), .C0(n5878), .Y(n2723)
         );
  OAI211XLTS U1063 ( .A0(n3741), .A1(n4027), .B0(n5883), .C0(n5882), .Y(n2725)
         );
  OAI211XLTS U1064 ( .A0(n3743), .A1(n4003), .B0(n5899), .C0(n5898), .Y(n2733)
         );
  OAI211XLTS U1065 ( .A0(n3743), .A1(n4000), .B0(n5901), .C0(n5900), .Y(n2734)
         );
  OAI211XLTS U1066 ( .A0(n3743), .A1(n3994), .B0(n5905), .C0(n5904), .Y(n2736)
         );
  OAI211XLTS U1067 ( .A0(n3742), .A1(n4009), .B0(n5895), .C0(n5894), .Y(n2731)
         );
  XNOR2XLTS U1068 ( .A(n6239), .B(n6252), .Y(n4849) );
  AOI32XLTS U1069 ( .A0(n160), .A1(n6240), .A2(n6252), .B0(n161), .B1(n4849), 
        .Y(n4850) );
  AOI32XLTS U1070 ( .A0(n219), .A1(n5571), .A2(n5570), .B0(n3543), .B1(n149), 
        .Y(n2570) );
  AOI32XLTS U1071 ( .A0(n158), .A1(n5564), .A2(n5563), .B0(n700), .B1(n19), 
        .Y(n2569) );
  NAND2XLTS U1072 ( .A(n3814), .B(n5559), .Y(n5564) );
  NAND2XLTS U1073 ( .A(n5555), .B(n278), .Y(n5448) );
  NAND3XLTS U1074 ( .A(n4878), .B(n6254), .C(n162), .Y(n5313) );
  NAND3XLTS U1075 ( .A(n265), .B(n4879), .C(n278), .Y(n5314) );
  NAND3XLTS U1076 ( .A(n4878), .B(n556), .C(n163), .Y(n5312) );
  NAND4XLTS U1077 ( .A(n161), .B(n265), .C(n6239), .D(n279), .Y(n5315) );
  NAND4XLTS U1078 ( .A(n160), .B(n265), .C(n279), .D(n6240), .Y(n5311) );
  CLKBUFX2TS U1079 ( .A(n5323), .Y(n569) );
  CLKBUFX2TS U1080 ( .A(n5327), .Y(n570) );
  NOR3X1TS U1081 ( .A(n258), .B(n8), .C(n349), .Y(n5295) );
  OAI2BB2XLTS U1082 ( .B0(n6263), .B1(n3577), .A0N(
        \requesterAddressbuffer[2][5] ), .A1N(n240), .Y(n5138) );
  OAI2BB2XLTS U1083 ( .B0(n6264), .B1(n3577), .A0N(
        \requesterAddressbuffer[2][4] ), .A1N(n240), .Y(n5146) );
  OAI2BB2XLTS U1084 ( .B0(n6266), .B1(n3576), .A0N(
        \requesterAddressbuffer[2][2] ), .A1N(n239), .Y(n5162) );
  OAI2BB2XLTS U1085 ( .B0(n6267), .B1(n3576), .A0N(
        \requesterAddressbuffer[2][1] ), .A1N(n239), .Y(n5170) );
  OAI2BB2XLTS U1086 ( .B0(n6265), .B1(n3576), .A0N(
        \requesterAddressbuffer[2][3] ), .A1N(n240), .Y(n5154) );
  OAI2BB2XLTS U1087 ( .B0(n6268), .B1(n3576), .A0N(
        \requesterAddressbuffer[2][0] ), .A1N(n240), .Y(n5178) );
  NAND2X1TS U1088 ( .A(n10), .B(n348), .Y(n6230) );
  CLKBUFX2TS U1089 ( .A(n3750), .Y(n3739) );
  CLKBUFX2TS U1090 ( .A(n3748), .Y(n3740) );
  CLKBUFX2TS U1091 ( .A(n3748), .Y(n3741) );
  CLKBUFX2TS U1092 ( .A(n3747), .Y(n3743) );
  CLKBUFX2TS U1093 ( .A(n3747), .Y(n3742) );
  CLKBUFX2TS U1094 ( .A(n3746), .Y(n3744) );
  CLKBUFX2TS U1095 ( .A(n3746), .Y(n3745) );
  CLKBUFX2TS U1096 ( .A(n3751), .Y(n3746) );
  CLKBUFX2TS U1097 ( .A(n3751), .Y(n3748) );
  CLKBUFX2TS U1098 ( .A(n3751), .Y(n3747) );
  CLKBUFX2TS U1099 ( .A(n3734), .Y(n3725) );
  CLKBUFX2TS U1100 ( .A(n3732), .Y(n3731) );
  CLKBUFX2TS U1101 ( .A(n3732), .Y(n3730) );
  CLKBUFX2TS U1102 ( .A(n3733), .Y(n3728) );
  CLKBUFX2TS U1103 ( .A(n3733), .Y(n3727) );
  CLKBUFX2TS U1104 ( .A(n3697), .Y(n3685) );
  CLKBUFX2TS U1105 ( .A(n3696), .Y(n3686) );
  CLKBUFX2TS U1106 ( .A(n3696), .Y(n3687) );
  CLKBUFX2TS U1107 ( .A(n3695), .Y(n3688) );
  CLKBUFX2TS U1108 ( .A(n3694), .Y(n3689) );
  CLKBUFX2TS U1109 ( .A(n3694), .Y(n3690) );
  CLKBUFX2TS U1110 ( .A(n3693), .Y(n3691) );
  CLKBUFX2TS U1111 ( .A(n3693), .Y(n3692) );
  CLKBUFX2TS U1112 ( .A(n3737), .Y(n3729) );
  CLKBUFX2TS U1113 ( .A(n3734), .Y(n3726) );
  CLKBUFX2TS U1114 ( .A(n3709), .Y(n3707) );
  CLKBUFX2TS U1115 ( .A(n3709), .Y(n3706) );
  CLKBUFX2TS U1116 ( .A(n3711), .Y(n3702) );
  CLKBUFX2TS U1117 ( .A(n3711), .Y(n3701) );
  CLKBUFX2TS U1118 ( .A(n3712), .Y(n3700) );
  CLKBUFX2TS U1119 ( .A(n3710), .Y(n3704) );
  CLKBUFX2TS U1120 ( .A(n3709), .Y(n3705) );
  CLKBUFX2TS U1121 ( .A(n3710), .Y(n3703) );
  CLKBUFX2TS U1122 ( .A(n3712), .Y(n3699) );
  CLKBUFX2TS U1123 ( .A(n3806), .Y(n3798) );
  CLKBUFX2TS U1124 ( .A(n3804), .Y(n3803) );
  CLKBUFX2TS U1125 ( .A(n3804), .Y(n3802) );
  CLKBUFX2TS U1126 ( .A(n3805), .Y(n3801) );
  CLKBUFX2TS U1127 ( .A(n3805), .Y(n3800) );
  CLKBUFX2TS U1128 ( .A(n3806), .Y(n3799) );
  CLKBUFX2TS U1129 ( .A(n3793), .Y(n3784) );
  CLKBUFX2TS U1130 ( .A(n3793), .Y(n3785) );
  CLKBUFX2TS U1131 ( .A(n3792), .Y(n3786) );
  CLKBUFX2TS U1132 ( .A(n3792), .Y(n3787) );
  CLKBUFX2TS U1133 ( .A(n3791), .Y(n3788) );
  CLKBUFX2TS U1134 ( .A(n3749), .Y(n3738) );
  CLKBUFX2TS U1135 ( .A(n3750), .Y(n3749) );
  CLKBUFX2TS U1136 ( .A(n3791), .Y(n3789) );
  CLKBUFX2TS U1137 ( .A(n3791), .Y(n3790) );
  CLKBUFX2TS U1138 ( .A(n3809), .Y(n3807) );
  CLKBUFX2TS U1139 ( .A(n3810), .Y(n3804) );
  CLKBUFX2TS U1140 ( .A(n3810), .Y(n3805) );
  CLKBUFX2TS U1141 ( .A(n3810), .Y(n3806) );
  CLKBUFX2TS U1142 ( .A(n3737), .Y(n3732) );
  CLKBUFX2TS U1143 ( .A(n3736), .Y(n3733) );
  CLKBUFX2TS U1144 ( .A(n3713), .Y(n3711) );
  CLKBUFX2TS U1145 ( .A(n3698), .Y(n3696) );
  CLKBUFX2TS U1146 ( .A(n3698), .Y(n3695) );
  CLKBUFX2TS U1147 ( .A(n3698), .Y(n3694) );
  CLKBUFX2TS U1148 ( .A(n3698), .Y(n3693) );
  CLKBUFX2TS U1149 ( .A(n3736), .Y(n3734) );
  CLKBUFX2TS U1150 ( .A(n6304), .Y(n3709) );
  CLKBUFX2TS U1151 ( .A(n3713), .Y(n3710) );
  CLKBUFX2TS U1152 ( .A(n3713), .Y(n3712) );
  CLKBUFX2TS U1153 ( .A(n3795), .Y(n3793) );
  CLKBUFX2TS U1154 ( .A(n3795), .Y(n3792) );
  CLKBUFX2TS U1155 ( .A(n3796), .Y(n3791) );
  CLKBUFX2TS U1156 ( .A(n6305), .Y(n3750) );
  CLKBUFX2TS U1157 ( .A(n6305), .Y(n3751) );
  CLKBUFX2TS U1158 ( .A(n784), .Y(n769) );
  CLKBUFX2TS U1159 ( .A(n784), .Y(n770) );
  CLKBUFX2TS U1160 ( .A(n781), .Y(n776) );
  CLKBUFX2TS U1161 ( .A(n782), .Y(n774) );
  CLKBUFX2TS U1162 ( .A(n782), .Y(n773) );
  CLKBUFX2TS U1163 ( .A(n781), .Y(n775) );
  CLKBUFX2TS U1164 ( .A(n783), .Y(n772) );
  CLKBUFX2TS U1165 ( .A(n783), .Y(n771) );
  CLKBUFX2TS U1166 ( .A(n3474), .Y(n3472) );
  CLKBUFX2TS U1167 ( .A(n3475), .Y(n3471) );
  CLKBUFX2TS U1168 ( .A(n3476), .Y(n3469) );
  CLKBUFX2TS U1169 ( .A(n3476), .Y(n3468) );
  CLKBUFX2TS U1170 ( .A(n3477), .Y(n3467) );
  CLKBUFX2TS U1171 ( .A(n3477), .Y(n3466) );
  CLKBUFX2TS U1172 ( .A(n3478), .Y(n3465) );
  CLKBUFX2TS U1173 ( .A(n3478), .Y(n3464) );
  CLKBUFX2TS U1174 ( .A(n3475), .Y(n3470) );
  CLKBUFX2TS U1175 ( .A(n868), .Y(n854) );
  CLKBUFX2TS U1176 ( .A(n3735), .Y(n3724) );
  CLKBUFX2TS U1177 ( .A(n3736), .Y(n3735) );
  CLKBUFX2TS U1178 ( .A(n868), .Y(n855) );
  CLKBUFX2TS U1179 ( .A(n3777), .Y(n3768) );
  CLKBUFX2TS U1180 ( .A(n866), .Y(n858) );
  CLKBUFX2TS U1181 ( .A(n865), .Y(n860) );
  CLKBUFX2TS U1182 ( .A(n864), .Y(n862) );
  CLKBUFX2TS U1183 ( .A(n865), .Y(n861) );
  CLKBUFX2TS U1184 ( .A(n866), .Y(n859) );
  CLKBUFX2TS U1185 ( .A(n867), .Y(n857) );
  CLKBUFX2TS U1186 ( .A(n867), .Y(n856) );
  CLKBUFX2TS U1187 ( .A(n3775), .Y(n3774) );
  CLKBUFX2TS U1188 ( .A(n3775), .Y(n3773) );
  CLKBUFX2TS U1189 ( .A(n3780), .Y(n3772) );
  CLKBUFX2TS U1190 ( .A(n3776), .Y(n3771) );
  CLKBUFX2TS U1191 ( .A(n3776), .Y(n3770) );
  CLKBUFX2TS U1192 ( .A(n3777), .Y(n3769) );
  CLKBUFX2TS U1193 ( .A(n327), .Y(n3697) );
  CLKBUFX2TS U1194 ( .A(n832), .Y(n818) );
  CLKBUFX2TS U1195 ( .A(n3395), .Y(n3381) );
  CLKBUFX2TS U1196 ( .A(n3395), .Y(n3382) );
  CLKBUFX2TS U1197 ( .A(n832), .Y(n819) );
  CLKBUFX2TS U1198 ( .A(n3474), .Y(n3473) );
  CLKBUFX2TS U1199 ( .A(n3325), .Y(n3323) );
  CLKBUFX2TS U1200 ( .A(n829), .Y(n826) );
  CLKBUFX2TS U1201 ( .A(n830), .Y(n823) );
  CLKBUFX2TS U1202 ( .A(n830), .Y(n822) );
  CLKBUFX2TS U1203 ( .A(n829), .Y(n824) );
  CLKBUFX2TS U1204 ( .A(n831), .Y(n821) );
  CLKBUFX2TS U1205 ( .A(n831), .Y(n820) );
  CLKBUFX2TS U1206 ( .A(n3326), .Y(n3322) );
  CLKBUFX2TS U1207 ( .A(n3326), .Y(n3321) );
  CLKBUFX2TS U1208 ( .A(n3327), .Y(n3320) );
  CLKBUFX2TS U1209 ( .A(n3327), .Y(n3319) );
  CLKBUFX2TS U1210 ( .A(n3329), .Y(n3316) );
  CLKBUFX2TS U1211 ( .A(n3391), .Y(n3389) );
  CLKBUFX2TS U1212 ( .A(n3392), .Y(n3388) );
  CLKBUFX2TS U1213 ( .A(n3393), .Y(n3386) );
  CLKBUFX2TS U1214 ( .A(n3393), .Y(n3385) );
  CLKBUFX2TS U1215 ( .A(n3392), .Y(n3387) );
  CLKBUFX2TS U1216 ( .A(n3394), .Y(n3384) );
  CLKBUFX2TS U1217 ( .A(n3394), .Y(n3383) );
  CLKBUFX2TS U1218 ( .A(n766), .Y(n752) );
  CLKBUFX2TS U1219 ( .A(n766), .Y(n753) );
  CLKBUFX2TS U1220 ( .A(n3197), .Y(n1602) );
  CLKBUFX2TS U1221 ( .A(n3197), .Y(n1653) );
  CLKBUFX2TS U1222 ( .A(n3328), .Y(n3318) );
  CLKBUFX2TS U1223 ( .A(n3328), .Y(n3317) );
  CLKBUFX2TS U1224 ( .A(n3329), .Y(n3315) );
  CLKBUFX2TS U1225 ( .A(n765), .Y(n754) );
  CLKBUFX2TS U1226 ( .A(n3196), .Y(n1654) );
  CLKBUFX2TS U1227 ( .A(n763), .Y(n758) );
  CLKBUFX2TS U1228 ( .A(n764), .Y(n757) );
  CLKBUFX2TS U1229 ( .A(n3195), .Y(n1817) );
  CLKBUFX2TS U1230 ( .A(n3195), .Y(n1797) );
  CLKBUFX2TS U1231 ( .A(n762), .Y(n761) );
  CLKBUFX2TS U1232 ( .A(n762), .Y(n760) );
  CLKBUFX2TS U1233 ( .A(n763), .Y(n759) );
  CLKBUFX2TS U1234 ( .A(n764), .Y(n756) );
  CLKBUFX2TS U1235 ( .A(n765), .Y(n755) );
  CLKBUFX2TS U1236 ( .A(n3194), .Y(n1822) );
  CLKBUFX2TS U1237 ( .A(n3194), .Y(n1894) );
  CLKBUFX2TS U1238 ( .A(n3196), .Y(n1728) );
  CLKBUFX2TS U1239 ( .A(n3298), .Y(n3284) );
  CLKBUFX2TS U1240 ( .A(n3298), .Y(n3285) );
  CLKBUFX2TS U1241 ( .A(n3764), .Y(n3755) );
  CLKBUFX2TS U1242 ( .A(n3764), .Y(n3754) );
  CLKBUFX2TS U1243 ( .A(n3293), .Y(n3291) );
  CLKBUFX2TS U1244 ( .A(n3293), .Y(n3292) );
  CLKBUFX2TS U1245 ( .A(n3294), .Y(n3290) );
  CLKBUFX2TS U1246 ( .A(n3295), .Y(n3287) );
  CLKBUFX2TS U1247 ( .A(n3294), .Y(n3289) );
  CLKBUFX2TS U1248 ( .A(n3295), .Y(n3288) );
  CLKBUFX2TS U1249 ( .A(n3296), .Y(n3286) );
  CLKBUFX2TS U1250 ( .A(n3808), .Y(n3797) );
  CLKBUFX2TS U1251 ( .A(n3809), .Y(n3808) );
  CLKBUFX2TS U1252 ( .A(n3794), .Y(n3783) );
  CLKBUFX2TS U1253 ( .A(n3795), .Y(n3794) );
  INVX2TS U1254 ( .A(n3244), .Y(n3241) );
  INVX2TS U1255 ( .A(n3248), .Y(n3240) );
  INVX2TS U1256 ( .A(n3243), .Y(n3242) );
  CLKBUFX2TS U1257 ( .A(n3363), .Y(n3350) );
  CLKBUFX2TS U1258 ( .A(n3363), .Y(n3351) );
  CLKBUFX2TS U1259 ( .A(n3361), .Y(n3355) );
  CLKBUFX2TS U1260 ( .A(n3361), .Y(n3354) );
  CLKBUFX2TS U1261 ( .A(n3360), .Y(n3356) );
  CLKBUFX2TS U1262 ( .A(n3362), .Y(n3353) );
  CLKBUFX2TS U1263 ( .A(n3362), .Y(n3352) );
  CLKBUFX2TS U1264 ( .A(n749), .Y(n737) );
  CLKBUFX2TS U1265 ( .A(n747), .Y(n739) );
  CLKBUFX2TS U1266 ( .A(n746), .Y(n740) );
  CLKBUFX2TS U1267 ( .A(n747), .Y(n738) );
  CLKBUFX2TS U1268 ( .A(n746), .Y(n741) );
  CLKBUFX2TS U1269 ( .A(n745), .Y(n742) );
  CLKBUFX2TS U1270 ( .A(n745), .Y(n743) );
  CLKBUFX2TS U1271 ( .A(n332), .Y(n3809) );
  CLKBUFX2TS U1272 ( .A(n3248), .Y(n3243) );
  CLKBUFX2TS U1273 ( .A(n3248), .Y(n3244) );
  CLKBUFX2TS U1274 ( .A(n3217), .Y(n3212) );
  CLKBUFX2TS U1275 ( .A(n3217), .Y(n3214) );
  CLKBUFX2TS U1276 ( .A(n3217), .Y(n3213) );
  CLKBUFX2TS U1277 ( .A(n870), .Y(n863) );
  CLKBUFX2TS U1278 ( .A(n870), .Y(n864) );
  CLKBUFX2TS U1279 ( .A(n870), .Y(n865) );
  CLKBUFX2TS U1280 ( .A(n869), .Y(n866) );
  CLKBUFX2TS U1281 ( .A(n869), .Y(n867) );
  CLKBUFX2TS U1282 ( .A(n869), .Y(n868) );
  CLKBUFX2TS U1283 ( .A(n3330), .Y(n3328) );
  CLKBUFX2TS U1284 ( .A(n3331), .Y(n3329) );
  CLKBUFX2TS U1285 ( .A(n3198), .Y(n3195) );
  CLKBUFX2TS U1286 ( .A(n6114), .Y(n762) );
  CLKBUFX2TS U1287 ( .A(n767), .Y(n763) );
  CLKBUFX2TS U1288 ( .A(n767), .Y(n764) );
  CLKBUFX2TS U1289 ( .A(n767), .Y(n765) );
  CLKBUFX2TS U1290 ( .A(n6307), .Y(n3762) );
  CLKBUFX2TS U1291 ( .A(n3199), .Y(n3193) );
  CLKBUFX2TS U1292 ( .A(n6307), .Y(n3763) );
  CLKBUFX2TS U1293 ( .A(n3766), .Y(n3764) );
  CLKBUFX2TS U1294 ( .A(n3199), .Y(n3194) );
  CLKBUFX2TS U1295 ( .A(n3766), .Y(n3765) );
  CLKBUFX2TS U1296 ( .A(n3198), .Y(n3196) );
  CLKBUFX2TS U1297 ( .A(n3299), .Y(n3298) );
  CLKBUFX2TS U1298 ( .A(n3299), .Y(n3297) );
  CLKBUFX2TS U1299 ( .A(n786), .Y(n779) );
  CLKBUFX2TS U1300 ( .A(n3780), .Y(n3775) );
  CLKBUFX2TS U1301 ( .A(n786), .Y(n780) );
  CLKBUFX2TS U1302 ( .A(n833), .Y(n830) );
  CLKBUFX2TS U1303 ( .A(n785), .Y(n782) );
  CLKBUFX2TS U1304 ( .A(n834), .Y(n829) );
  CLKBUFX2TS U1305 ( .A(n786), .Y(n781) );
  CLKBUFX2TS U1306 ( .A(n3779), .Y(n3776) );
  CLKBUFX2TS U1307 ( .A(n833), .Y(n831) );
  CLKBUFX2TS U1308 ( .A(n785), .Y(n783) );
  CLKBUFX2TS U1309 ( .A(n3300), .Y(n3293) );
  CLKBUFX2TS U1310 ( .A(n3396), .Y(n3393) );
  CLKBUFX2TS U1311 ( .A(n6191), .Y(n3392) );
  CLKBUFX2TS U1312 ( .A(n3396), .Y(n3394) );
  CLKBUFX2TS U1313 ( .A(n3396), .Y(n3395) );
  CLKBUFX2TS U1314 ( .A(n3479), .Y(n3476) );
  CLKBUFX2TS U1315 ( .A(n3479), .Y(n3477) );
  CLKBUFX2TS U1316 ( .A(n3479), .Y(n3478) );
  CLKBUFX2TS U1317 ( .A(n3480), .Y(n3475) );
  CLKBUFX2TS U1318 ( .A(n767), .Y(n766) );
  CLKBUFX2TS U1319 ( .A(n833), .Y(n832) );
  CLKBUFX2TS U1320 ( .A(n3779), .Y(n3777) );
  CLKBUFX2TS U1321 ( .A(n785), .Y(n784) );
  CLKBUFX2TS U1322 ( .A(n3198), .Y(n3197) );
  CLKBUFX2TS U1323 ( .A(n3300), .Y(n3294) );
  CLKBUFX2TS U1324 ( .A(n3300), .Y(n3295) );
  CLKBUFX2TS U1325 ( .A(n3299), .Y(n3296) );
  CLKBUFX2TS U1326 ( .A(n3330), .Y(n3326) );
  CLKBUFX2TS U1327 ( .A(n3330), .Y(n3327) );
  CLKBUFX2TS U1328 ( .A(n335), .Y(n3737) );
  CLKBUFX2TS U1329 ( .A(n335), .Y(n3736) );
  CLKBUFX2TS U1330 ( .A(n6311), .Y(n3795) );
  CLKBUFX2TS U1331 ( .A(n332), .Y(n3810) );
  CLKBUFX2TS U1332 ( .A(n7), .Y(n3714) );
  CLKBUFX2TS U1333 ( .A(n6304), .Y(n3713) );
  CLKBUFX2TS U1334 ( .A(n327), .Y(n3698) );
  CLKBUFX2TS U1335 ( .A(n3281), .Y(n3267) );
  CLKBUFX2TS U1336 ( .A(n3281), .Y(n3268) );
  CLKBUFX2TS U1337 ( .A(n3278), .Y(n3274) );
  CLKBUFX2TS U1338 ( .A(n3278), .Y(n3273) );
  CLKBUFX2TS U1339 ( .A(n3280), .Y(n3270) );
  CLKBUFX2TS U1340 ( .A(n3458), .Y(n3454) );
  CLKBUFX2TS U1341 ( .A(n3459), .Y(n3452) );
  CLKBUFX2TS U1342 ( .A(n3460), .Y(n3450) );
  CLKBUFX2TS U1343 ( .A(n3460), .Y(n3449) );
  CLKBUFX2TS U1344 ( .A(n3461), .Y(n3447) );
  CLKBUFX2TS U1345 ( .A(n3279), .Y(n3272) );
  CLKBUFX2TS U1346 ( .A(n3279), .Y(n3271) );
  CLKBUFX2TS U1347 ( .A(n3280), .Y(n3269) );
  CLKBUFX2TS U1348 ( .A(n3458), .Y(n3453) );
  CLKBUFX2TS U1349 ( .A(n3459), .Y(n3451) );
  CLKBUFX2TS U1350 ( .A(n3461), .Y(n3448) );
  CLKBUFX2TS U1351 ( .A(n3430), .Y(n3416) );
  CLKBUFX2TS U1352 ( .A(n734), .Y(n704) );
  CLKBUFX2TS U1353 ( .A(n3778), .Y(n3767) );
  CLKBUFX2TS U1354 ( .A(n3779), .Y(n3778) );
  CLKBUFX2TS U1355 ( .A(n734), .Y(n705) );
  CLKBUFX2TS U1356 ( .A(n732), .Y(n711) );
  CLKBUFX2TS U1357 ( .A(n732), .Y(n708) );
  CLKBUFX2TS U1358 ( .A(n733), .Y(n707) );
  CLKBUFX2TS U1359 ( .A(n716), .Y(n714) );
  CLKBUFX2TS U1360 ( .A(n729), .Y(n712) );
  CLKBUFX2TS U1361 ( .A(n733), .Y(n706) );
  CLKBUFX2TS U1362 ( .A(n3358), .Y(n3357) );
  CLKBUFX2TS U1363 ( .A(n3523), .Y(n3520) );
  CLKBUFX2TS U1364 ( .A(n3524), .Y(n3519) );
  CLKBUFX2TS U1365 ( .A(n3524), .Y(n3518) );
  CLKBUFX2TS U1366 ( .A(n3526), .Y(n3517) );
  CLKBUFX2TS U1367 ( .A(n3526), .Y(n3516) );
  CLKBUFX2TS U1368 ( .A(n3527), .Y(n3515) );
  CLKBUFX2TS U1369 ( .A(n3527), .Y(n3514) );
  CLKBUFX2TS U1370 ( .A(n3528), .Y(n3513) );
  CLKBUFX2TS U1371 ( .A(n3528), .Y(n3512) );
  CLKBUFX2TS U1372 ( .A(n3495), .Y(n3481) );
  CLKBUFX2TS U1373 ( .A(n3495), .Y(n3482) );
  CLKBUFX2TS U1374 ( .A(n3494), .Y(n3483) );
  CLKBUFX2TS U1375 ( .A(n3427), .Y(n3423) );
  CLKBUFX2TS U1376 ( .A(n3427), .Y(n3422) );
  CLKBUFX2TS U1377 ( .A(n3428), .Y(n3420) );
  CLKBUFX2TS U1378 ( .A(n3490), .Y(n3489) );
  CLKBUFX2TS U1379 ( .A(n3490), .Y(n3488) );
  CLKBUFX2TS U1380 ( .A(n3492), .Y(n3487) );
  CLKBUFX2TS U1381 ( .A(n3493), .Y(n3486) );
  CLKBUFX2TS U1382 ( .A(n3493), .Y(n3485) );
  CLKBUFX2TS U1383 ( .A(n3494), .Y(n3484) );
  CLKBUFX2TS U1384 ( .A(n3432), .Y(n3424) );
  CLKBUFX2TS U1385 ( .A(n3428), .Y(n3421) );
  CLKBUFX2TS U1386 ( .A(n3523), .Y(n3521) );
  CLKBUFX2TS U1387 ( .A(n796), .Y(n795) );
  CLKBUFX2TS U1388 ( .A(n796), .Y(n794) );
  CLKBUFX2TS U1389 ( .A(n797), .Y(n793) );
  CLKBUFX2TS U1390 ( .A(n797), .Y(n792) );
  CLKBUFX2TS U1391 ( .A(n798), .Y(n790) );
  CLKBUFX2TS U1392 ( .A(n798), .Y(n791) );
  CLKBUFX2TS U1393 ( .A(n799), .Y(n789) );
  CLKBUFX2TS U1394 ( .A(n799), .Y(n788) );
  CLKBUFX2TS U1395 ( .A(n3763), .Y(n3753) );
  INVX2TS U1396 ( .A(n3543), .Y(n3539) );
  INVX2TS U1397 ( .A(n3543), .Y(n3538) );
  INVX2TS U1398 ( .A(n3543), .Y(n3537) );
  INVX2TS U1399 ( .A(n3545), .Y(n3531) );
  INVX2TS U1400 ( .A(n3545), .Y(n3532) );
  INVX2TS U1401 ( .A(n3546), .Y(n3535) );
  INVX2TS U1402 ( .A(n3545), .Y(n3536) );
  INVX2TS U1403 ( .A(n3546), .Y(n3534) );
  INVX2TS U1404 ( .A(n562), .Y(n3533) );
  INVX2TS U1405 ( .A(n3246), .Y(n3232) );
  INVX2TS U1406 ( .A(n3247), .Y(n3233) );
  INVX2TS U1407 ( .A(n3245), .Y(n3239) );
  CLKBUFX2TS U1408 ( .A(n3247), .Y(n3245) );
  INVX2TS U1409 ( .A(n3246), .Y(n3238) );
  CLKBUFX2TS U1410 ( .A(n3247), .Y(n3246) );
  INVX2TS U1411 ( .A(n3247), .Y(n3237) );
  INVX2TS U1412 ( .A(n3246), .Y(n3236) );
  INVX2TS U1413 ( .A(n3248), .Y(n3234) );
  INVX2TS U1414 ( .A(n3245), .Y(n3235) );
  INVX2TS U1415 ( .A(n3216), .Y(n3205) );
  INVX2TS U1416 ( .A(n3215), .Y(n3201) );
  INVX2TS U1417 ( .A(n3215), .Y(n3203) );
  INVX2TS U1418 ( .A(n3215), .Y(n3207) );
  INVX2TS U1419 ( .A(n3216), .Y(n3202) );
  INVX2TS U1420 ( .A(n3215), .Y(n3204) );
  INVX2TS U1421 ( .A(n3216), .Y(n3206) );
  INVX2TS U1422 ( .A(n3216), .Y(n3208) );
  INVX2TS U1423 ( .A(n3544), .Y(n3529) );
  INVX2TS U1424 ( .A(n3544), .Y(n3530) );
  CLKBUFX2TS U1425 ( .A(n3365), .Y(n3359) );
  CLKBUFX2TS U1426 ( .A(n3364), .Y(n3361) );
  CLKBUFX2TS U1427 ( .A(n3365), .Y(n3360) );
  CLKBUFX2TS U1428 ( .A(n3364), .Y(n3362) );
  CLKBUFX2TS U1429 ( .A(n3364), .Y(n3363) );
  INVX2TS U1430 ( .A(n3260), .Y(n3250) );
  INVX2TS U1431 ( .A(n3260), .Y(n3249) );
  INVX2TS U1432 ( .A(n3261), .Y(n3251) );
  INVX2TS U1433 ( .A(n3261), .Y(n3252) );
  INVX2TS U1434 ( .A(n3262), .Y(n3253) );
  INVX2TS U1435 ( .A(n3263), .Y(n3254) );
  INVX2TS U1436 ( .A(n3263), .Y(n3255) );
  INVX2TS U1437 ( .A(n3264), .Y(n3257) );
  INVX2TS U1438 ( .A(n3264), .Y(n3256) );
  INVX2TS U1439 ( .A(n3262), .Y(n3259) );
  INVX2TS U1440 ( .A(n701), .Y(n696) );
  INVX2TS U1441 ( .A(n701), .Y(n695) );
  INVX2TS U1442 ( .A(n698), .Y(n691) );
  INVX2TS U1443 ( .A(n698), .Y(n690) );
  INVX2TS U1444 ( .A(n699), .Y(n693) );
  INVX2TS U1445 ( .A(n702), .Y(n694) );
  INVX2TS U1446 ( .A(n699), .Y(n692) );
  INVX2TS U1447 ( .A(n698), .Y(n689) );
  INVX2TS U1448 ( .A(n850), .Y(n846) );
  INVX2TS U1449 ( .A(n850), .Y(n845) );
  INVX2TS U1450 ( .A(n850), .Y(n844) );
  INVX2TS U1451 ( .A(n3413), .Y(n3408) );
  INVX2TS U1452 ( .A(n3414), .Y(n3407) );
  INVX2TS U1453 ( .A(n3415), .Y(n3406) );
  INVX2TS U1454 ( .A(n3347), .Y(n3342) );
  INVX2TS U1455 ( .A(n3348), .Y(n3341) );
  INVX2TS U1456 ( .A(n3349), .Y(n3340) );
  INVX2TS U1457 ( .A(n853), .Y(n838) );
  INVX2TS U1458 ( .A(n3413), .Y(n3400) );
  INVX2TS U1459 ( .A(n3347), .Y(n3334) );
  INVX2TS U1460 ( .A(n564), .Y(n839) );
  INVX2TS U1461 ( .A(n3413), .Y(n3401) );
  INVX2TS U1462 ( .A(n3347), .Y(n3335) );
  INVX2TS U1463 ( .A(n851), .Y(n842) );
  INVX2TS U1464 ( .A(n851), .Y(n843) );
  INVX2TS U1465 ( .A(n851), .Y(n841) );
  INVX2TS U1466 ( .A(n3346), .Y(n3338) );
  INVX2TS U1467 ( .A(n3346), .Y(n3337) );
  INVX2TS U1468 ( .A(n3412), .Y(n3404) );
  INVX2TS U1469 ( .A(n3412), .Y(n3405) );
  INVX2TS U1470 ( .A(n3412), .Y(n3403) );
  INVX2TS U1471 ( .A(n3413), .Y(n3402) );
  INVX2TS U1472 ( .A(n564), .Y(n840) );
  INVX2TS U1473 ( .A(n3346), .Y(n3339) );
  INVX2TS U1474 ( .A(n3347), .Y(n3336) );
  INVX2TS U1475 ( .A(n3265), .Y(n3258) );
  INVX2TS U1476 ( .A(n699), .Y(n697) );
  INVX2TS U1477 ( .A(n852), .Y(n836) );
  INVX2TS U1478 ( .A(n3414), .Y(n3398) );
  INVX2TS U1479 ( .A(n3348), .Y(n3332) );
  INVX2TS U1480 ( .A(n852), .Y(n837) );
  INVX2TS U1481 ( .A(n3348), .Y(n3333) );
  INVX2TS U1482 ( .A(n3414), .Y(n3399) );
  CLKBUFX2TS U1483 ( .A(n750), .Y(n749) );
  CLKBUFX2TS U1484 ( .A(n750), .Y(n748) );
  CLKBUFX2TS U1485 ( .A(n751), .Y(n747) );
  CLKBUFX2TS U1486 ( .A(n751), .Y(n746) );
  CLKBUFX2TS U1487 ( .A(n751), .Y(n745) );
  CLKBUFX2TS U1488 ( .A(n3229), .Y(n3218) );
  CLKBUFX2TS U1489 ( .A(n3228), .Y(n3220) );
  CLKBUFX2TS U1490 ( .A(n1598), .Y(n886) );
  CLKBUFX2TS U1491 ( .A(n1598), .Y(n871) );
  CLKBUFX2TS U1492 ( .A(n3229), .Y(n3219) );
  CLKBUFX2TS U1493 ( .A(n1571), .Y(n919) );
  CLKBUFX2TS U1494 ( .A(n1535), .Y(n955) );
  CLKBUFX2TS U1495 ( .A(n1535), .Y(n959) );
  CLKBUFX2TS U1496 ( .A(n1598), .Y(n970) );
  CLKBUFX2TS U1497 ( .A(n3227), .Y(n3223) );
  CLKBUFX2TS U1498 ( .A(n3228), .Y(n3221) );
  CLKBUFX2TS U1499 ( .A(n1571), .Y(n936) );
  CLKBUFX2TS U1500 ( .A(n1535), .Y(n957) );
  CLKBUFX2TS U1501 ( .A(n1533), .Y(n986) );
  CLKBUFX2TS U1502 ( .A(n1533), .Y(n1402) );
  CLKBUFX2TS U1503 ( .A(n3227), .Y(n3222) );
  CLKBUFX2TS U1504 ( .A(n3444), .Y(n3434) );
  CLKBUFX2TS U1505 ( .A(n816), .Y(n805) );
  CLKBUFX2TS U1506 ( .A(n815), .Y(n807) );
  CLKBUFX2TS U1507 ( .A(n816), .Y(n806) );
  CLKBUFX2TS U1508 ( .A(n814), .Y(n809) );
  CLKBUFX2TS U1509 ( .A(n814), .Y(n810) );
  CLKBUFX2TS U1510 ( .A(n813), .Y(n811) );
  CLKBUFX2TS U1511 ( .A(n3311), .Y(n3303) );
  CLKBUFX2TS U1512 ( .A(n3310), .Y(n3305) );
  CLKBUFX2TS U1513 ( .A(n3379), .Y(n3367) );
  CLKBUFX2TS U1514 ( .A(n3378), .Y(n3369) );
  CLKBUFX2TS U1515 ( .A(n6190), .Y(n3368) );
  CLKBUFX2TS U1516 ( .A(n3377), .Y(n3371) );
  CLKBUFX2TS U1517 ( .A(n3377), .Y(n3372) );
  CLKBUFX2TS U1518 ( .A(n3378), .Y(n3370) );
  CLKBUFX2TS U1519 ( .A(n3442), .Y(n3439) );
  CLKBUFX2TS U1520 ( .A(n3442), .Y(n3437) );
  CLKBUFX2TS U1521 ( .A(n3442), .Y(n3436) );
  CLKBUFX2TS U1522 ( .A(n3509), .Y(n3498) );
  CLKBUFX2TS U1523 ( .A(n3507), .Y(n3499) );
  CLKBUFX2TS U1524 ( .A(n3507), .Y(n3500) );
  CLKBUFX2TS U1525 ( .A(n3506), .Y(n3501) );
  CLKBUFX2TS U1526 ( .A(n3506), .Y(n3502) );
  CLKBUFX2TS U1527 ( .A(n3505), .Y(n3503) );
  CLKBUFX2TS U1528 ( .A(n3505), .Y(n3504) );
  CLKBUFX2TS U1529 ( .A(n815), .Y(n808) );
  CLKBUFX2TS U1530 ( .A(n3312), .Y(n3302) );
  CLKBUFX2TS U1531 ( .A(n3311), .Y(n3304) );
  CLKBUFX2TS U1532 ( .A(n3442), .Y(n3438) );
  CLKBUFX2TS U1533 ( .A(n3444), .Y(n3435) );
  CLKBUFX2TS U1534 ( .A(n6205), .Y(n3440) );
  CLKBUFX2TS U1535 ( .A(n3309), .Y(n3308) );
  CLKBUFX2TS U1536 ( .A(n3310), .Y(n3306) );
  CLKBUFX2TS U1537 ( .A(n813), .Y(n812) );
  CLKBUFX2TS U1538 ( .A(n3309), .Y(n3307) );
  CLKBUFX2TS U1539 ( .A(n3376), .Y(n3375) );
  CLKBUFX2TS U1540 ( .A(n3377), .Y(n3373) );
  CLKBUFX2TS U1541 ( .A(n3376), .Y(n3374) );
  CLKBUFX2TS U1542 ( .A(n6205), .Y(n3441) );
  CLKBUFX2TS U1543 ( .A(n3573), .Y(n3561) );
  CLKBUFX2TS U1544 ( .A(n3573), .Y(n3569) );
  CLKBUFX2TS U1545 ( .A(n3570), .Y(n3568) );
  CLKBUFX2TS U1546 ( .A(n3570), .Y(n3567) );
  CLKBUFX2TS U1547 ( .A(n3571), .Y(n3566) );
  CLKBUFX2TS U1548 ( .A(n3571), .Y(n3565) );
  CLKBUFX2TS U1549 ( .A(n3572), .Y(n3564) );
  CLKBUFX2TS U1550 ( .A(n3573), .Y(n3562) );
  CLKBUFX2TS U1551 ( .A(n3572), .Y(n3563) );
  CLKBUFX2TS U1552 ( .A(n3559), .Y(n3548) );
  CLKBUFX2TS U1553 ( .A(n3557), .Y(n3549) );
  CLKBUFX2TS U1554 ( .A(n3557), .Y(n3550) );
  CLKBUFX2TS U1555 ( .A(n3556), .Y(n3551) );
  CLKBUFX2TS U1556 ( .A(n3555), .Y(n3554) );
  CLKBUFX2TS U1557 ( .A(n3556), .Y(n3552) );
  CLKBUFX2TS U1558 ( .A(n3555), .Y(n3553) );
  CLKBUFX2TS U1559 ( .A(n3667), .Y(n3655) );
  CLKBUFX2TS U1560 ( .A(n3634), .Y(n3632) );
  CLKBUFX2TS U1561 ( .A(n3667), .Y(n3656) );
  CLKBUFX2TS U1562 ( .A(n6281), .Y(n3631) );
  CLKBUFX2TS U1563 ( .A(n6281), .Y(n3630) );
  CLKBUFX2TS U1564 ( .A(n3668), .Y(n3657) );
  CLKBUFX2TS U1565 ( .A(n3666), .Y(n3658) );
  CLKBUFX2TS U1566 ( .A(n3635), .Y(n3628) );
  CLKBUFX2TS U1567 ( .A(n3666), .Y(n3659) );
  CLKBUFX2TS U1568 ( .A(n3636), .Y(n3627) );
  CLKBUFX2TS U1569 ( .A(n3665), .Y(n3660) );
  CLKBUFX2TS U1570 ( .A(n3637), .Y(n3624) );
  CLKBUFX2TS U1571 ( .A(n3636), .Y(n3626) );
  CLKBUFX2TS U1572 ( .A(n3637), .Y(n3625) );
  CLKBUFX2TS U1573 ( .A(n3635), .Y(n3629) );
  CLKBUFX2TS U1574 ( .A(n3665), .Y(n3661) );
  CLKBUFX2TS U1575 ( .A(n3664), .Y(n3662) );
  CLKBUFX2TS U1576 ( .A(n3664), .Y(n3663) );
  CLKBUFX2TS U1577 ( .A(n6143), .Y(n869) );
  CLKBUFX2TS U1578 ( .A(n3545), .Y(n3544) );
  CLKBUFX2TS U1579 ( .A(n6306), .Y(n3752) );
  CLKBUFX2TS U1580 ( .A(n802), .Y(n801) );
  CLKBUFX2TS U1581 ( .A(n3432), .Y(n3427) );
  CLKBUFX2TS U1582 ( .A(n3496), .Y(n3495) );
  CLKBUFX2TS U1583 ( .A(n3497), .Y(n3490) );
  CLKBUFX2TS U1584 ( .A(n3497), .Y(n3491) );
  CLKBUFX2TS U1585 ( .A(n3496), .Y(n3493) );
  CLKBUFX2TS U1586 ( .A(n3497), .Y(n3492) );
  CLKBUFX2TS U1587 ( .A(n3431), .Y(n3429) );
  CLKBUFX2TS U1588 ( .A(n3432), .Y(n3426) );
  CLKBUFX2TS U1589 ( .A(n3431), .Y(n3428) );
  CLKBUFX2TS U1590 ( .A(n3496), .Y(n3494) );
  CLKBUFX2TS U1591 ( .A(n3431), .Y(n3430) );
  CLKBUFX2TS U1592 ( .A(n802), .Y(n800) );
  CLKBUFX2TS U1593 ( .A(n3283), .Y(n3276) );
  CLKBUFX2TS U1594 ( .A(n3231), .Y(n3224) );
  CLKBUFX2TS U1595 ( .A(n803), .Y(n796) );
  CLKBUFX2TS U1596 ( .A(n803), .Y(n797) );
  CLKBUFX2TS U1597 ( .A(n803), .Y(n798) );
  CLKBUFX2TS U1598 ( .A(n3283), .Y(n3277) );
  CLKBUFX2TS U1599 ( .A(n3283), .Y(n3278) );
  CLKBUFX2TS U1600 ( .A(n3282), .Y(n3281) );
  CLKBUFX2TS U1601 ( .A(n3462), .Y(n3460) );
  CLKBUFX2TS U1602 ( .A(n6223), .Y(n3524) );
  CLKBUFX2TS U1603 ( .A(n6223), .Y(n3526) );
  CLKBUFX2TS U1604 ( .A(n3524), .Y(n3527) );
  CLKBUFX2TS U1605 ( .A(n3523), .Y(n3528) );
  CLKBUFX2TS U1606 ( .A(n6223), .Y(n3525) );
  CLKBUFX2TS U1607 ( .A(n802), .Y(n799) );
  CLKBUFX2TS U1608 ( .A(n3282), .Y(n3279) );
  CLKBUFX2TS U1609 ( .A(n3282), .Y(n3280) );
  CLKBUFX2TS U1610 ( .A(n3463), .Y(n3457) );
  CLKBUFX2TS U1611 ( .A(n3463), .Y(n3458) );
  CLKBUFX2TS U1612 ( .A(n3462), .Y(n3459) );
  CLKBUFX2TS U1613 ( .A(n3462), .Y(n3461) );
  CLKBUFX2TS U1614 ( .A(n6114), .Y(n768) );
  CLKBUFX2TS U1615 ( .A(n835), .Y(n828) );
  CLKBUFX2TS U1616 ( .A(n6130), .Y(n835) );
  CLKBUFX2TS U1617 ( .A(n3200), .Y(n3192) );
  CLKBUFX2TS U1618 ( .A(n6145), .Y(n3200) );
  CLKBUFX2TS U1619 ( .A(n6175), .Y(n3331) );
  CLKBUFX2TS U1620 ( .A(n735), .Y(n732) );
  CLKBUFX2TS U1621 ( .A(n3397), .Y(n3391) );
  CLKBUFX2TS U1622 ( .A(n6191), .Y(n3397) );
  CLKBUFX2TS U1623 ( .A(n3366), .Y(n3358) );
  CLKBUFX2TS U1624 ( .A(n6188), .Y(n3366) );
  CLKBUFX2TS U1625 ( .A(n736), .Y(n728) );
  CLKBUFX2TS U1626 ( .A(n736), .Y(n729) );
  CLKBUFX2TS U1627 ( .A(n735), .Y(n733) );
  CLKBUFX2TS U1628 ( .A(n735), .Y(n734) );
  CLKBUFX2TS U1629 ( .A(n6145), .Y(n3199) );
  CLKBUFX2TS U1630 ( .A(n6145), .Y(n3198) );
  CLKBUFX2TS U1631 ( .A(n6173), .Y(n3299) );
  CLKBUFX2TS U1632 ( .A(n6173), .Y(n3300) );
  CLKBUFX2TS U1633 ( .A(n6220), .Y(n3480) );
  CLKBUFX2TS U1634 ( .A(n6191), .Y(n3396) );
  CLKBUFX2TS U1635 ( .A(n6220), .Y(n3479) );
  CLKBUFX2TS U1636 ( .A(n6130), .Y(n833) );
  CLKBUFX2TS U1637 ( .A(n6127), .Y(n785) );
  CLKBUFX2TS U1638 ( .A(n6114), .Y(n767) );
  CLKBUFX2TS U1639 ( .A(n6307), .Y(n3766) );
  CLKBUFX2TS U1640 ( .A(n6308), .Y(n3780) );
  CLKBUFX2TS U1641 ( .A(n6308), .Y(n3779) );
  CLKBUFX2TS U1642 ( .A(n6175), .Y(n3330) );
  CLKBUFX2TS U1643 ( .A(n560), .Y(n3215) );
  CLKBUFX2TS U1644 ( .A(n560), .Y(n3216) );
  CLKBUFX2TS U1645 ( .A(n559), .Y(n3247) );
  CLKBUFX2TS U1646 ( .A(n559), .Y(n3248) );
  CLKBUFX2TS U1647 ( .A(n560), .Y(n3217) );
  CLKBUFX2TS U1648 ( .A(n701), .Y(n700) );
  CLKBUFX2TS U1649 ( .A(n736), .Y(n715) );
  CLKBUFX2TS U1650 ( .A(n3462), .Y(n3456) );
  CLKBUFX2TS U1651 ( .A(n3428), .Y(n3425) );
  INVX2TS U1652 ( .A(n3546), .Y(n3541) );
  INVX2TS U1653 ( .A(n3544), .Y(n3540) );
  CLKBUFX2TS U1654 ( .A(n3266), .Y(n3260) );
  CLKBUFX2TS U1655 ( .A(n3265), .Y(n3264) );
  CLKBUFX2TS U1656 ( .A(n3266), .Y(n3261) );
  CLKBUFX2TS U1657 ( .A(n3266), .Y(n3262) );
  CLKBUFX2TS U1658 ( .A(n3265), .Y(n3263) );
  CLKBUFX2TS U1659 ( .A(n853), .Y(n852) );
  CLKBUFX2TS U1660 ( .A(n3415), .Y(n3414) );
  CLKBUFX2TS U1661 ( .A(n3349), .Y(n3348) );
  CLKBUFX2TS U1662 ( .A(n6188), .Y(n3364) );
  INVX2TS U1663 ( .A(n5471), .Y(n6292) );
  INVX2TS U1664 ( .A(n703), .Y(n686) );
  INVX2TS U1665 ( .A(n703), .Y(n687) );
  INVX2TS U1666 ( .A(n703), .Y(n688) );
  INVX2TS U1667 ( .A(n565), .Y(n3344) );
  INVX2TS U1668 ( .A(n852), .Y(n848) );
  INVX2TS U1669 ( .A(n852), .Y(n847) );
  INVX2TS U1670 ( .A(n565), .Y(n3343) );
  INVX2TS U1671 ( .A(n561), .Y(n3410) );
  INVX2TS U1672 ( .A(n561), .Y(n3409) );
  CLKBUFX2TS U1673 ( .A(n6129), .Y(n816) );
  CLKBUFX2TS U1674 ( .A(n6129), .Y(n814) );
  CLKBUFX2TS U1675 ( .A(n6129), .Y(n813) );
  CLKBUFX2TS U1676 ( .A(n6144), .Y(n1598) );
  CLKBUFX2TS U1677 ( .A(n3230), .Y(n3229) );
  CLKBUFX2TS U1678 ( .A(n3231), .Y(n3225) );
  CLKBUFX2TS U1679 ( .A(n3231), .Y(n3226) );
  CLKBUFX2TS U1680 ( .A(n3230), .Y(n3228) );
  CLKBUFX2TS U1681 ( .A(n3314), .Y(n3310) );
  CLKBUFX2TS U1682 ( .A(n3314), .Y(n3309) );
  CLKBUFX2TS U1683 ( .A(n6190), .Y(n3378) );
  CLKBUFX2TS U1684 ( .A(n3380), .Y(n3377) );
  CLKBUFX2TS U1685 ( .A(n3380), .Y(n3376) );
  CLKBUFX2TS U1686 ( .A(n3510), .Y(n3509) );
  CLKBUFX2TS U1687 ( .A(n3510), .Y(n3508) );
  CLKBUFX2TS U1688 ( .A(n3511), .Y(n3507) );
  CLKBUFX2TS U1689 ( .A(n3511), .Y(n3506) );
  CLKBUFX2TS U1690 ( .A(n3511), .Y(n3505) );
  CLKBUFX2TS U1691 ( .A(n814), .Y(n815) );
  CLKBUFX2TS U1692 ( .A(n6144), .Y(n1571) );
  CLKBUFX2TS U1693 ( .A(n6144), .Y(n1535) );
  CLKBUFX2TS U1694 ( .A(n1571), .Y(n1533) );
  CLKBUFX2TS U1695 ( .A(n3230), .Y(n3227) );
  CLKBUFX2TS U1696 ( .A(n6174), .Y(n3312) );
  CLKBUFX2TS U1697 ( .A(n3314), .Y(n3311) );
  CLKBUFX2TS U1698 ( .A(n6205), .Y(n3442) );
  CLKBUFX2TS U1699 ( .A(n3446), .Y(n3443) );
  CLKBUFX2TS U1700 ( .A(n3446), .Y(n3444) );
  CLKBUFX2TS U1701 ( .A(n6113), .Y(n750) );
  CLKBUFX2TS U1702 ( .A(n6113), .Y(n751) );
  INVX2TS U1703 ( .A(n684), .Y(n669) );
  INVX2TS U1704 ( .A(n685), .Y(n670) );
  INVX2TS U1705 ( .A(n683), .Y(n679) );
  INVX2TS U1706 ( .A(n683), .Y(n678) );
  INVX2TS U1707 ( .A(n680), .Y(n677) );
  INVX2TS U1708 ( .A(n680), .Y(n676) );
  INVX2TS U1709 ( .A(n680), .Y(n675) );
  INVX2TS U1710 ( .A(n684), .Y(n673) );
  INVX2TS U1711 ( .A(n684), .Y(n672) );
  INVX2TS U1712 ( .A(n684), .Y(n674) );
  INVX2TS U1713 ( .A(n680), .Y(n671) );
  CLKBUFX2TS U1714 ( .A(n3445), .Y(n3433) );
  CLKBUFX2TS U1715 ( .A(n3446), .Y(n3445) );
  CLKBUFX2TS U1716 ( .A(n817), .Y(n804) );
  CLKBUFX2TS U1717 ( .A(n813), .Y(n817) );
  CLKBUFX2TS U1718 ( .A(n3313), .Y(n3301) );
  CLKBUFX2TS U1719 ( .A(n6174), .Y(n3313) );
  CLKBUFX2TS U1720 ( .A(n6190), .Y(n3379) );
  CLKBUFX2TS U1721 ( .A(n649), .Y(n637) );
  CLKBUFX2TS U1722 ( .A(n647), .Y(n645) );
  CLKBUFX2TS U1723 ( .A(n646), .Y(n644) );
  CLKBUFX2TS U1724 ( .A(n646), .Y(n643) );
  CLKBUFX2TS U1725 ( .A(n647), .Y(n642) );
  CLKBUFX2TS U1726 ( .A(n647), .Y(n641) );
  CLKBUFX2TS U1727 ( .A(n649), .Y(n638) );
  CLKBUFX2TS U1728 ( .A(n648), .Y(n640) );
  CLKBUFX2TS U1729 ( .A(n648), .Y(n639) );
  INVX2TS U1730 ( .A(n605), .Y(n604) );
  INVX2TS U1731 ( .A(n606), .Y(n603) );
  INVX2TS U1732 ( .A(n607), .Y(n602) );
  CLKBUFX2TS U1733 ( .A(n3575), .Y(n3570) );
  CLKBUFX2TS U1734 ( .A(n3574), .Y(n3571) );
  CLKBUFX2TS U1735 ( .A(n3574), .Y(n3573) );
  CLKBUFX2TS U1736 ( .A(n3574), .Y(n3572) );
  CLKBUFX2TS U1737 ( .A(n3560), .Y(n3557) );
  CLKBUFX2TS U1738 ( .A(n3560), .Y(n3556) );
  CLKBUFX2TS U1739 ( .A(n3560), .Y(n3555) );
  CLKBUFX2TS U1740 ( .A(n583), .Y(n571) );
  CLKBUFX2TS U1741 ( .A(n583), .Y(n572) );
  CLKBUFX2TS U1742 ( .A(n582), .Y(n573) );
  CLKBUFX2TS U1743 ( .A(n584), .Y(n574) );
  CLKBUFX2TS U1744 ( .A(n582), .Y(n575) );
  CLKBUFX2TS U1745 ( .A(n581), .Y(n576) );
  CLKBUFX2TS U1746 ( .A(n580), .Y(n579) );
  CLKBUFX2TS U1747 ( .A(n581), .Y(n577) );
  CLKBUFX2TS U1748 ( .A(n580), .Y(n578) );
  CLKBUFX2TS U1749 ( .A(n632), .Y(n611) );
  CLKBUFX2TS U1750 ( .A(n626), .Y(n612) );
  CLKBUFX2TS U1751 ( .A(n627), .Y(n613) );
  CLKBUFX2TS U1752 ( .A(n627), .Y(n614) );
  CLKBUFX2TS U1753 ( .A(n626), .Y(n621) );
  CLKBUFX2TS U1754 ( .A(n625), .Y(n624) );
  CLKBUFX2TS U1755 ( .A(n626), .Y(n622) );
  CLKBUFX2TS U1756 ( .A(n625), .Y(n623) );
  CLKBUFX2TS U1757 ( .A(n3558), .Y(n3547) );
  CLKBUFX2TS U1758 ( .A(n3559), .Y(n3558) );
  INVX2TS U1759 ( .A(reset), .Y(n4430) );
  CLKBUFX2TS U1760 ( .A(n3605), .Y(n3593) );
  CLKBUFX2TS U1761 ( .A(n3650), .Y(n3648) );
  CLKBUFX2TS U1762 ( .A(n3605), .Y(n3594) );
  CLKBUFX2TS U1763 ( .A(n3651), .Y(n3647) );
  CLKBUFX2TS U1764 ( .A(n3651), .Y(n3646) );
  CLKBUFX2TS U1765 ( .A(n3683), .Y(n3670) );
  CLKBUFX2TS U1766 ( .A(n3653), .Y(n3645) );
  CLKBUFX2TS U1767 ( .A(n3652), .Y(n3644) );
  CLKBUFX2TS U1768 ( .A(n3679), .Y(n3671) );
  CLKBUFX2TS U1769 ( .A(n3606), .Y(n3595) );
  CLKBUFX2TS U1770 ( .A(n3652), .Y(n3643) );
  CLKBUFX2TS U1771 ( .A(n3680), .Y(n3672) );
  CLKBUFX2TS U1772 ( .A(n3604), .Y(n3596) );
  CLKBUFX2TS U1773 ( .A(n3652), .Y(n3642) );
  CLKBUFX2TS U1774 ( .A(n3680), .Y(n3673) );
  CLKBUFX2TS U1775 ( .A(n3604), .Y(n3597) );
  CLKBUFX2TS U1776 ( .A(n3653), .Y(n3641) );
  CLKBUFX2TS U1777 ( .A(n3679), .Y(n3674) );
  CLKBUFX2TS U1778 ( .A(n3603), .Y(n3598) );
  CLKBUFX2TS U1779 ( .A(n3653), .Y(n3640) );
  CLKBUFX2TS U1780 ( .A(n3591), .Y(n3576) );
  CLKBUFX2TS U1781 ( .A(n3591), .Y(n3577) );
  CLKBUFX2TS U1782 ( .A(n3619), .Y(n3609) );
  CLKBUFX2TS U1783 ( .A(n3587), .Y(n3583) );
  CLKBUFX2TS U1784 ( .A(n3588), .Y(n3582) );
  CLKBUFX2TS U1785 ( .A(n3617), .Y(n3613) );
  CLKBUFX2TS U1786 ( .A(n3589), .Y(n3581) );
  CLKBUFX2TS U1787 ( .A(n3617), .Y(n3612) );
  CLKBUFX2TS U1788 ( .A(n3589), .Y(n3580) );
  CLKBUFX2TS U1789 ( .A(n3618), .Y(n3611) );
  CLKBUFX2TS U1790 ( .A(n3590), .Y(n3579) );
  CLKBUFX2TS U1791 ( .A(n3618), .Y(n3610) );
  CLKBUFX2TS U1792 ( .A(n3590), .Y(n3578) );
  CLKBUFX2TS U1793 ( .A(n3651), .Y(n3649) );
  CLKBUFX2TS U1794 ( .A(n3603), .Y(n3599) );
  CLKBUFX2TS U1795 ( .A(n3679), .Y(n3675) );
  CLKBUFX2TS U1796 ( .A(n3602), .Y(n3601) );
  CLKBUFX2TS U1797 ( .A(n3639), .Y(n3634) );
  CLKBUFX2TS U1798 ( .A(n3668), .Y(n3667) );
  CLKBUFX2TS U1799 ( .A(n3669), .Y(n3666) );
  CLKBUFX2TS U1800 ( .A(n3669), .Y(n3665) );
  CLKBUFX2TS U1801 ( .A(n3638), .Y(n3636) );
  CLKBUFX2TS U1802 ( .A(n3638), .Y(n3637) );
  CLKBUFX2TS U1803 ( .A(n3638), .Y(n3635) );
  CLKBUFX2TS U1804 ( .A(n3669), .Y(n3664) );
  CLKBUFX2TS U1805 ( .A(n3587), .Y(n3584) );
  CLKBUFX2TS U1806 ( .A(n3639), .Y(n3633) );
  CLKBUFX2TS U1807 ( .A(n3602), .Y(n3600) );
  CLKBUFX2TS U1808 ( .A(n3678), .Y(n3676) );
  CLKBUFX2TS U1809 ( .A(n3678), .Y(n3677) );
  AND2X2TS U1810 ( .A(n223), .B(n6301), .Y(n6173) );
  INVX2TS U1811 ( .A(n5521), .Y(n6302) );
  CLKBUFX2TS U1812 ( .A(n562), .Y(n3546) );
  CLKBUFX2TS U1813 ( .A(n563), .Y(n701) );
  CLKBUFX2TS U1814 ( .A(n563), .Y(n702) );
  CLKBUFX2TS U1815 ( .A(n562), .Y(n3545) );
  CLKBUFX2TS U1816 ( .A(n6172), .Y(n3282) );
  CLKBUFX2TS U1817 ( .A(n6128), .Y(n802) );
  CLKBUFX2TS U1818 ( .A(n6128), .Y(n803) );
  CLKBUFX2TS U1819 ( .A(n6221), .Y(n3497) );
  CLKBUFX2TS U1820 ( .A(n6204), .Y(n3432) );
  CLKBUFX2TS U1821 ( .A(n6221), .Y(n3496) );
  CLKBUFX2TS U1822 ( .A(n6204), .Y(n3431) );
  CLKBUFX2TS U1823 ( .A(n6206), .Y(n3463) );
  CLKBUFX2TS U1824 ( .A(n6206), .Y(n3462) );
  CLKBUFX2TS U1825 ( .A(n6158), .Y(n3231) );
  CLKBUFX2TS U1826 ( .A(n6112), .Y(n735) );
  INVX2TS U1827 ( .A(n5542), .Y(n6298) );
  INVX2TS U1828 ( .A(n5541), .Y(n6299) );
  CLKBUFX2TS U1829 ( .A(n561), .Y(n3415) );
  CLKBUFX2TS U1830 ( .A(n564), .Y(n853) );
  CLKBUFX2TS U1831 ( .A(n565), .Y(n3349) );
  CLKBUFX2TS U1832 ( .A(n557), .Y(n3266) );
  INVX2TS U1833 ( .A(n5426), .Y(n6301) );
  CLKBUFX2TS U1834 ( .A(n609), .Y(n605) );
  CLKBUFX2TS U1835 ( .A(n609), .Y(n606) );
  CLKBUFX2TS U1836 ( .A(n609), .Y(n607) );
  AND2X2TS U1837 ( .A(n5481), .B(n5365), .Y(n6113) );
  CLKBUFX2TS U1838 ( .A(n649), .Y(n646) );
  CLKBUFX2TS U1839 ( .A(n650), .Y(n647) );
  CLKBUFX2TS U1840 ( .A(n651), .Y(n649) );
  CLKBUFX2TS U1841 ( .A(n651), .Y(n648) );
  CLKBUFX2TS U1842 ( .A(n6190), .Y(n3380) );
  CLKBUFX2TS U1843 ( .A(n6222), .Y(n3510) );
  CLKBUFX2TS U1844 ( .A(n6222), .Y(n3511) );
  CLKBUFX2TS U1845 ( .A(n6158), .Y(n3230) );
  CLKBUFX2TS U1846 ( .A(n6174), .Y(n3314) );
  CLKBUFX2TS U1847 ( .A(n6205), .Y(n3446) );
  CLKBUFX2TS U1848 ( .A(n683), .Y(n681) );
  CLKBUFX2TS U1849 ( .A(n683), .Y(n682) );
  CLKBUFX2TS U1850 ( .A(n650), .Y(n636) );
  CLKBUFX2TS U1851 ( .A(n651), .Y(n650) );
  INVX2TS U1852 ( .A(n566), .Y(n585) );
  INVX2TS U1853 ( .A(n566), .Y(n586) );
  INVX2TS U1854 ( .A(n608), .Y(n587) );
  INVX2TS U1855 ( .A(n608), .Y(n597) );
  INVX2TS U1856 ( .A(n608), .Y(n598) );
  INVX2TS U1857 ( .A(n607), .Y(n599) );
  INVX2TS U1858 ( .A(n608), .Y(n600) );
  INVX2TS U1859 ( .A(n609), .Y(n601) );
  CLKBUFX2TS U1860 ( .A(n634), .Y(n632) );
  CLKBUFX2TS U1861 ( .A(n584), .Y(n583) );
  CLKBUFX2TS U1862 ( .A(n5226), .Y(n582) );
  CLKBUFX2TS U1863 ( .A(n635), .Y(n627) );
  CLKBUFX2TS U1864 ( .A(n635), .Y(n626) );
  CLKBUFX2TS U1865 ( .A(n584), .Y(n581) );
  CLKBUFX2TS U1866 ( .A(n635), .Y(n625) );
  CLKBUFX2TS U1867 ( .A(n584), .Y(n580) );
  CLKBUFX2TS U1868 ( .A(n6258), .Y(n3575) );
  CLKBUFX2TS U1869 ( .A(n6258), .Y(n3574) );
  CLKBUFX2TS U1870 ( .A(n5291), .Y(n3559) );
  CLKBUFX2TS U1871 ( .A(n5291), .Y(n3560) );
  CLKBUFX2TS U1872 ( .A(n633), .Y(n610) );
  CLKBUFX2TS U1873 ( .A(n634), .Y(n633) );
  CLKBUFX2TS U1874 ( .A(n4274), .Y(n4275) );
  CLKBUFX2TS U1875 ( .A(n4277), .Y(n4278) );
  CLKBUFX2TS U1876 ( .A(n4274), .Y(n4276) );
  CLKBUFX2TS U1877 ( .A(n4277), .Y(n4279) );
  INVX2TS U1878 ( .A(n3823), .Y(n3820) );
  CLKBUFX2TS U1879 ( .A(n3592), .Y(n3587) );
  CLKBUFX2TS U1880 ( .A(n3683), .Y(n3682) );
  CLKBUFX2TS U1881 ( .A(n3606), .Y(n3605) );
  CLKBUFX2TS U1882 ( .A(n6279), .Y(n3588) );
  CLKBUFX2TS U1883 ( .A(n3683), .Y(n3681) );
  CLKBUFX2TS U1884 ( .A(n4), .Y(n3651) );
  CLKBUFX2TS U1885 ( .A(n3622), .Y(n3617) );
  CLKBUFX2TS U1886 ( .A(n3588), .Y(n3589) );
  CLKBUFX2TS U1887 ( .A(n3654), .Y(n3652) );
  CLKBUFX2TS U1888 ( .A(n3684), .Y(n3680) );
  CLKBUFX2TS U1889 ( .A(n3607), .Y(n3604) );
  CLKBUFX2TS U1890 ( .A(n3621), .Y(n3618) );
  CLKBUFX2TS U1891 ( .A(n3684), .Y(n3679) );
  CLKBUFX2TS U1892 ( .A(n3607), .Y(n3603) );
  CLKBUFX2TS U1893 ( .A(n6279), .Y(n3590) );
  CLKBUFX2TS U1894 ( .A(n3654), .Y(n3653) );
  CLKBUFX2TS U1895 ( .A(n3621), .Y(n3619) );
  CLKBUFX2TS U1896 ( .A(n3588), .Y(n3591) );
  CLKBUFX2TS U1897 ( .A(n3607), .Y(n3602) );
  CLKBUFX2TS U1898 ( .A(n663), .Y(n657) );
  CLKBUFX2TS U1899 ( .A(n663), .Y(n656) );
  CLKBUFX2TS U1900 ( .A(n664), .Y(n655) );
  CLKBUFX2TS U1901 ( .A(n664), .Y(n654) );
  CLKBUFX2TS U1902 ( .A(n665), .Y(n653) );
  CLKBUFX2TS U1903 ( .A(n665), .Y(n652) );
  CLKBUFX2TS U1904 ( .A(n3620), .Y(n3608) );
  CLKBUFX2TS U1905 ( .A(n3621), .Y(n3620) );
  INVX2TS U1906 ( .A(n5365), .Y(n6283) );
  CLKBUFX2TS U1907 ( .A(n3654), .Y(n3650) );
  CLKBUFX2TS U1908 ( .A(n3684), .Y(n3678) );
  CLKBUFX2TS U1909 ( .A(n6282), .Y(n3668) );
  CLKBUFX2TS U1910 ( .A(n6282), .Y(n3669) );
  CLKBUFX2TS U1911 ( .A(n6281), .Y(n3639) );
  CLKBUFX2TS U1912 ( .A(n6281), .Y(n3638) );
  CLKBUFX2TS U1913 ( .A(n3616), .Y(n3614) );
  CLKBUFX2TS U1914 ( .A(n3616), .Y(n3615) );
  CLKBUFX2TS U1915 ( .A(n3586), .Y(n3585) );
  OA22X1TS U1916 ( .A0(n5553), .A1(n352), .B0(n5496), .B1(n233), .Y(n561) );
  XNOR2X1TS U1917 ( .A(n6278), .B(n6238), .Y(n4868) );
  OAI21X1TS U1918 ( .A0(n6), .A1(n235), .B0(n280), .Y(n5378) );
  OAI2BB1X1TS U1919 ( .A0N(n215), .A1N(n5331), .B0(n5330), .Y(n5332) );
  OAI21X1TS U1920 ( .A0(n5331), .A1(n215), .B0(n277), .Y(n5330) );
  NOR2X1TS U1921 ( .A(n236), .B(n5399), .Y(n5543) );
  NOR2X1TS U1922 ( .A(n4865), .B(n6286), .Y(n4870) );
  AOI21X2TS U1923 ( .A0(n237), .A1(n5401), .B0(n6302), .Y(n5523) );
  NOR2X1TS U1924 ( .A(n5404), .B(n6303), .Y(n6158) );
  INVX2TS U1925 ( .A(n4864), .Y(n6286) );
  INVX2TS U1926 ( .A(n5449), .Y(n6290) );
  OR2X2TS U1927 ( .A(n4870), .B(n4869), .Y(n4871) );
  AOI21X1TS U1928 ( .A0(n232), .A1(n6290), .B0(n6299), .Y(n5403) );
  NAND2X1TS U1929 ( .A(n232), .B(n5497), .Y(n5404) );
  INVX2TS U1930 ( .A(n216), .Y(n6255) );
  NOR2BX1TS U1931 ( .AN(n229), .B(n351), .Y(n5481) );
  AND2X2TS U1932 ( .A(n5481), .B(n232), .Y(n6144) );
  AND2X2TS U1933 ( .A(n5507), .B(n263), .Y(n6222) );
  AND2X2TS U1934 ( .A(n5507), .B(n261), .Y(n6129) );
  AND2X2TS U1935 ( .A(n5481), .B(n5506), .Y(n6205) );
  AND2X2TS U1936 ( .A(n5507), .B(n5458), .Y(n6190) );
  AND2X2TS U1937 ( .A(n5481), .B(n234), .Y(n6174) );
  CLKBUFX2TS U1938 ( .A(n685), .Y(n684) );
  CLKBUFX2TS U1939 ( .A(n685), .Y(n683) );
  CLKBUFX2TS U1940 ( .A(n5290), .Y(n651) );
  CLKBUFX2TS U1941 ( .A(n566), .Y(n608) );
  CLKBUFX2TS U1942 ( .A(n566), .Y(n609) );
  NAND2X1TS U1943 ( .A(n352), .B(n4430), .Y(n6236) );
  CLKBUFX2TS U1944 ( .A(destinationAddressIn_SOUTH[6]), .Y(n4274) );
  CLKBUFX2TS U1945 ( .A(destinationAddressIn_SOUTH[7]), .Y(n4277) );
  CLKBUFX2TS U1946 ( .A(n5289), .Y(n634) );
  CLKBUFX2TS U1947 ( .A(n5289), .Y(n635) );
  CLKBUFX2TS U1948 ( .A(n5226), .Y(n584) );
  CLKBUFX2TS U1949 ( .A(n4301), .Y(n4302) );
  CLKBUFX2TS U1950 ( .A(n4412), .Y(n4413) );
  CLKBUFX2TS U1951 ( .A(n4385), .Y(n4386) );
  CLKBUFX2TS U1952 ( .A(n4367), .Y(n4368) );
  CLKBUFX2TS U1953 ( .A(n4361), .Y(n4362) );
  CLKBUFX2TS U1954 ( .A(n4358), .Y(n4359) );
  CLKBUFX2TS U1955 ( .A(n4337), .Y(n4338) );
  CLKBUFX2TS U1956 ( .A(n4334), .Y(n4335) );
  CLKBUFX2TS U1957 ( .A(n4328), .Y(n4329) );
  CLKBUFX2TS U1958 ( .A(n4316), .Y(n4317) );
  CLKBUFX2TS U1959 ( .A(n4391), .Y(n4392) );
  CLKBUFX2TS U1960 ( .A(n4388), .Y(n4389) );
  CLKBUFX2TS U1961 ( .A(n4382), .Y(n4383) );
  CLKBUFX2TS U1962 ( .A(n4379), .Y(n4380) );
  CLKBUFX2TS U1963 ( .A(n4376), .Y(n4377) );
  CLKBUFX2TS U1964 ( .A(n4370), .Y(n4371) );
  CLKBUFX2TS U1965 ( .A(n4364), .Y(n4365) );
  CLKBUFX2TS U1966 ( .A(n4355), .Y(n4356) );
  CLKBUFX2TS U1967 ( .A(n4346), .Y(n4347) );
  CLKBUFX2TS U1968 ( .A(n4331), .Y(n4332) );
  CLKBUFX2TS U1969 ( .A(n4325), .Y(n4326) );
  CLKBUFX2TS U1970 ( .A(n4322), .Y(n4323) );
  CLKBUFX2TS U1971 ( .A(n4319), .Y(n4320) );
  CLKBUFX2TS U1972 ( .A(n4313), .Y(n4314) );
  CLKBUFX2TS U1973 ( .A(n4304), .Y(n4305) );
  CLKBUFX2TS U1974 ( .A(n4427), .Y(n4428) );
  CLKBUFX2TS U1975 ( .A(n4421), .Y(n4422) );
  CLKBUFX2TS U1976 ( .A(n4418), .Y(n4419) );
  CLKBUFX2TS U1977 ( .A(n4415), .Y(n4416) );
  CLKBUFX2TS U1978 ( .A(n4298), .Y(n4299) );
  CLKBUFX2TS U1979 ( .A(n4349), .Y(n4350) );
  CLKBUFX2TS U1980 ( .A(n4343), .Y(n4344) );
  CLKBUFX2TS U1981 ( .A(n4340), .Y(n4341) );
  CLKBUFX2TS U1982 ( .A(n4307), .Y(n4308) );
  CLKBUFX2TS U1983 ( .A(n4424), .Y(n4425) );
  CLKBUFX2TS U1984 ( .A(n4373), .Y(n4374) );
  CLKBUFX2TS U1985 ( .A(n4352), .Y(n4353) );
  CLKBUFX2TS U1986 ( .A(n4310), .Y(n4311) );
  CLKBUFX2TS U1987 ( .A(n4409), .Y(n4410) );
  CLKBUFX2TS U1988 ( .A(n4406), .Y(n4407) );
  CLKBUFX2TS U1989 ( .A(n4400), .Y(n4401) );
  CLKBUFX2TS U1990 ( .A(n4403), .Y(n4404) );
  CLKBUFX2TS U1991 ( .A(n4397), .Y(n4398) );
  CLKBUFX2TS U1992 ( .A(n4394), .Y(n4395) );
  INVX2TS U1993 ( .A(n3925), .Y(n3923) );
  INVX2TS U1994 ( .A(n3922), .Y(n3920) );
  INVX2TS U1995 ( .A(n3919), .Y(n3917) );
  INVX2TS U1996 ( .A(n3916), .Y(n3914) );
  INVX2TS U1997 ( .A(n3913), .Y(n3911) );
  INVX2TS U1998 ( .A(n3910), .Y(n3908) );
  INVX2TS U1999 ( .A(n3907), .Y(n3905) );
  INVX2TS U2000 ( .A(n3904), .Y(n3902) );
  INVX2TS U2001 ( .A(n3901), .Y(n3899) );
  INVX2TS U2002 ( .A(n3898), .Y(n3896) );
  INVX2TS U2003 ( .A(n3895), .Y(n3893) );
  INVX2TS U2004 ( .A(n3892), .Y(n3890) );
  INVX2TS U2005 ( .A(n3889), .Y(n3887) );
  INVX2TS U2006 ( .A(n3886), .Y(n3884) );
  INVX2TS U2007 ( .A(n3883), .Y(n3881) );
  INVX2TS U2008 ( .A(n3880), .Y(n3878) );
  INVX2TS U2009 ( .A(n3877), .Y(n3875) );
  INVX2TS U2010 ( .A(n3874), .Y(n3872) );
  INVX2TS U2011 ( .A(n3871), .Y(n3869) );
  INVX2TS U2012 ( .A(n3868), .Y(n3866) );
  INVX2TS U2013 ( .A(n3865), .Y(n3863) );
  INVX2TS U2014 ( .A(n3862), .Y(n3860) );
  INVX2TS U2015 ( .A(n3859), .Y(n3857) );
  INVX2TS U2016 ( .A(n3856), .Y(n3854) );
  INVX2TS U2017 ( .A(n3853), .Y(n3851) );
  INVX2TS U2018 ( .A(n3850), .Y(n3848) );
  INVX2TS U2019 ( .A(n3847), .Y(n3845) );
  INVX2TS U2020 ( .A(n3844), .Y(n3842) );
  INVX2TS U2021 ( .A(n3841), .Y(n3839) );
  INVX2TS U2022 ( .A(n3838), .Y(n3836) );
  INVX2TS U2023 ( .A(n3835), .Y(n3833) );
  INVX2TS U2024 ( .A(n3832), .Y(n3830) );
  INVX2TS U2025 ( .A(n3946), .Y(n3944) );
  INVX2TS U2026 ( .A(n3961), .Y(n3959) );
  INVX2TS U2027 ( .A(n3955), .Y(n3953) );
  INVX2TS U2028 ( .A(n3952), .Y(n3950) );
  INVX2TS U2029 ( .A(n3949), .Y(n3947) );
  INVX2TS U2030 ( .A(n3958), .Y(n3956) );
  INVX2TS U2031 ( .A(n3943), .Y(n3941) );
  INVX2TS U2032 ( .A(n3940), .Y(n3938) );
  INVX2TS U2033 ( .A(n3934), .Y(n3932) );
  INVX2TS U2034 ( .A(n3937), .Y(n3935) );
  INVX2TS U2035 ( .A(n3931), .Y(n3929) );
  INVX2TS U2036 ( .A(n3928), .Y(n3926) );
  INVX2TS U2037 ( .A(n6226), .Y(n6258) );
  INVX2TS U2038 ( .A(n4096), .Y(n4094) );
  INVX2TS U2039 ( .A(n4099), .Y(n4097) );
  INVX2TS U2040 ( .A(n4090), .Y(n4088) );
  INVX2TS U2041 ( .A(n4093), .Y(n4091) );
  INVX2TS U2042 ( .A(n4087), .Y(n4085) );
  INVX2TS U2043 ( .A(n4084), .Y(n4082) );
  INVX2TS U2044 ( .A(n4249), .Y(n4247) );
  INVX2TS U2045 ( .A(n4246), .Y(n4244) );
  INVX2TS U2046 ( .A(n4243), .Y(n4241) );
  INVX2TS U2047 ( .A(n4240), .Y(n4238) );
  INVX2TS U2048 ( .A(n4255), .Y(n4253) );
  INVX2TS U2049 ( .A(n4252), .Y(n4250) );
  INVX2TS U2050 ( .A(n3816), .Y(n3815) );
  CLKBUFX2TS U2051 ( .A(n4427), .Y(n4429) );
  CLKBUFX2TS U2052 ( .A(n4424), .Y(n4426) );
  CLKBUFX2TS U2053 ( .A(n4421), .Y(n4423) );
  CLKBUFX2TS U2054 ( .A(n4415), .Y(n4417) );
  CLKBUFX2TS U2055 ( .A(n4412), .Y(n4414) );
  CLKBUFX2TS U2056 ( .A(n4418), .Y(n4420) );
  CLKBUFX2TS U2057 ( .A(n4388), .Y(n4390) );
  CLKBUFX2TS U2058 ( .A(n4385), .Y(n4387) );
  CLKBUFX2TS U2059 ( .A(n4376), .Y(n4378) );
  CLKBUFX2TS U2060 ( .A(n4373), .Y(n4375) );
  CLKBUFX2TS U2061 ( .A(n4361), .Y(n4363) );
  CLKBUFX2TS U2062 ( .A(n4355), .Y(n4357) );
  CLKBUFX2TS U2063 ( .A(n4352), .Y(n4354) );
  CLKBUFX2TS U2064 ( .A(n4349), .Y(n4351) );
  CLKBUFX2TS U2065 ( .A(n4343), .Y(n4345) );
  CLKBUFX2TS U2066 ( .A(n4340), .Y(n4342) );
  CLKBUFX2TS U2067 ( .A(n4337), .Y(n4339) );
  CLKBUFX2TS U2068 ( .A(n4334), .Y(n4336) );
  CLKBUFX2TS U2069 ( .A(n4331), .Y(n4333) );
  CLKBUFX2TS U2070 ( .A(n4328), .Y(n4330) );
  CLKBUFX2TS U2071 ( .A(n4322), .Y(n4324) );
  CLKBUFX2TS U2072 ( .A(n4310), .Y(n4312) );
  CLKBUFX2TS U2073 ( .A(n4307), .Y(n4309) );
  CLKBUFX2TS U2074 ( .A(n4382), .Y(n4384) );
  CLKBUFX2TS U2075 ( .A(n4379), .Y(n4381) );
  CLKBUFX2TS U2076 ( .A(n4367), .Y(n4369) );
  CLKBUFX2TS U2077 ( .A(n4358), .Y(n4360) );
  CLKBUFX2TS U2078 ( .A(n4325), .Y(n4327) );
  CLKBUFX2TS U2079 ( .A(n4313), .Y(n4315) );
  CLKBUFX2TS U2080 ( .A(n4301), .Y(n4303) );
  CLKBUFX2TS U2081 ( .A(n4391), .Y(n4393) );
  CLKBUFX2TS U2082 ( .A(n4370), .Y(n4372) );
  CLKBUFX2TS U2083 ( .A(n4364), .Y(n4366) );
  CLKBUFX2TS U2084 ( .A(n4346), .Y(n4348) );
  CLKBUFX2TS U2085 ( .A(n4316), .Y(n4318) );
  CLKBUFX2TS U2086 ( .A(n4304), .Y(n4306) );
  CLKBUFX2TS U2087 ( .A(n4298), .Y(n4300) );
  CLKBUFX2TS U2088 ( .A(n4319), .Y(n4321) );
  INVX2TS U2089 ( .A(n4021), .Y(n4019) );
  INVX2TS U2090 ( .A(n3991), .Y(n3989) );
  INVX2TS U2091 ( .A(n4078), .Y(n4076) );
  INVX2TS U2092 ( .A(n4075), .Y(n4073) );
  INVX2TS U2093 ( .A(n4072), .Y(n4070) );
  INVX2TS U2094 ( .A(n4069), .Y(n4067) );
  INVX2TS U2095 ( .A(n4066), .Y(n4064) );
  INVX2TS U2096 ( .A(n4063), .Y(n4061) );
  INVX2TS U2097 ( .A(n4057), .Y(n4055) );
  INVX2TS U2098 ( .A(n4051), .Y(n4049) );
  INVX2TS U2099 ( .A(n4048), .Y(n4046) );
  INVX2TS U2100 ( .A(n4045), .Y(n4043) );
  INVX2TS U2101 ( .A(n4042), .Y(n4040) );
  INVX2TS U2102 ( .A(n4027), .Y(n4025) );
  INVX2TS U2103 ( .A(n4024), .Y(n4022) );
  INVX2TS U2104 ( .A(n4018), .Y(n4016) );
  INVX2TS U2105 ( .A(n4015), .Y(n4013) );
  INVX2TS U2106 ( .A(n4012), .Y(n4010) );
  INVX2TS U2107 ( .A(n4009), .Y(n4007) );
  INVX2TS U2108 ( .A(n4003), .Y(n4001) );
  INVX2TS U2109 ( .A(n4000), .Y(n3998) );
  INVX2TS U2110 ( .A(n4081), .Y(n4079) );
  INVX2TS U2111 ( .A(n4060), .Y(n4058) );
  INVX2TS U2112 ( .A(n4054), .Y(n4052) );
  INVX2TS U2113 ( .A(n4036), .Y(n4034) );
  INVX2TS U2114 ( .A(n4006), .Y(n4004) );
  INVX2TS U2115 ( .A(n3994), .Y(n3992) );
  INVX2TS U2116 ( .A(n3988), .Y(n3986) );
  INVX2TS U2117 ( .A(n4039), .Y(n4037) );
  INVX2TS U2118 ( .A(n4033), .Y(n4031) );
  INVX2TS U2119 ( .A(n4030), .Y(n4028) );
  INVX2TS U2120 ( .A(n3997), .Y(n3995) );
  INVX2TS U2121 ( .A(n4117), .Y(n4115) );
  INVX2TS U2122 ( .A(n4114), .Y(n4112) );
  INVX2TS U2123 ( .A(n4111), .Y(n4109) );
  INVX2TS U2124 ( .A(n4108), .Y(n4106) );
  INVX2TS U2125 ( .A(n4105), .Y(n4103) );
  INVX2TS U2126 ( .A(n4102), .Y(n4100) );
  CLKBUFX2TS U2127 ( .A(n3980), .Y(n3981) );
  CLKBUFX2TS U2128 ( .A(n3968), .Y(n3969) );
  CLKBUFX2TS U2129 ( .A(n3962), .Y(n3963) );
  CLKBUFX2TS U2130 ( .A(n3977), .Y(n3978) );
  CLKBUFX2TS U2131 ( .A(n3971), .Y(n3972) );
  CLKBUFX2TS U2132 ( .A(n3983), .Y(n3984) );
  CLKBUFX2TS U2133 ( .A(n3974), .Y(n3975) );
  CLKBUFX2TS U2134 ( .A(n3965), .Y(n3966) );
  CLKBUFX2TS U2135 ( .A(n4292), .Y(n4293) );
  CLKBUFX2TS U2136 ( .A(n4286), .Y(n4287) );
  CLKBUFX2TS U2137 ( .A(n4283), .Y(n4284) );
  CLKBUFX2TS U2138 ( .A(n4295), .Y(n4296) );
  CLKBUFX2TS U2139 ( .A(n4289), .Y(n4290) );
  CLKBUFX2TS U2140 ( .A(n4280), .Y(n4281) );
  CLKBUFX2TS U2141 ( .A(n4139), .Y(n4140) );
  CLKBUFX2TS U2142 ( .A(n4136), .Y(n4137) );
  CLKBUFX2TS U2143 ( .A(n4130), .Y(n4131) );
  CLKBUFX2TS U2144 ( .A(n4124), .Y(n4125) );
  CLKBUFX2TS U2145 ( .A(n4118), .Y(n4119) );
  CLKBUFX2TS U2146 ( .A(n4133), .Y(n4134) );
  CLKBUFX2TS U2147 ( .A(n4127), .Y(n4128) );
  CLKBUFX2TS U2148 ( .A(n4121), .Y(n4122) );
  CLKBUFX2TS U2149 ( .A(n4136), .Y(n4138) );
  CLKBUFX2TS U2150 ( .A(n4118), .Y(n4120) );
  CLKBUFX2TS U2151 ( .A(n3980), .Y(n3982) );
  CLKBUFX2TS U2152 ( .A(n3974), .Y(n3976) );
  CLKBUFX2TS U2153 ( .A(n3962), .Y(n3964) );
  CLKBUFX2TS U2154 ( .A(n4130), .Y(n4132) );
  CLKBUFX2TS U2155 ( .A(n4127), .Y(n4129) );
  CLKBUFX2TS U2156 ( .A(n3971), .Y(n3973) );
  CLKBUFX2TS U2157 ( .A(n3983), .Y(n3985) );
  CLKBUFX2TS U2158 ( .A(n4139), .Y(n4141) );
  CLKBUFX2TS U2159 ( .A(n3977), .Y(n3979) );
  CLKBUFX2TS U2160 ( .A(n4133), .Y(n4135) );
  CLKBUFX2TS U2161 ( .A(n3968), .Y(n3970) );
  CLKBUFX2TS U2162 ( .A(n4124), .Y(n4126) );
  CLKBUFX2TS U2163 ( .A(n3965), .Y(n3967) );
  CLKBUFX2TS U2164 ( .A(n4121), .Y(n4123) );
  CLKBUFX2TS U2165 ( .A(n4292), .Y(n4294) );
  CLKBUFX2TS U2166 ( .A(n4280), .Y(n4282) );
  CLKBUFX2TS U2167 ( .A(n4289), .Y(n4291) );
  CLKBUFX2TS U2168 ( .A(n4283), .Y(n4285) );
  CLKBUFX2TS U2169 ( .A(n4295), .Y(n4297) );
  CLKBUFX2TS U2170 ( .A(n4286), .Y(n4288) );
  CLKBUFX2TS U2171 ( .A(n4406), .Y(n4408) );
  CLKBUFX2TS U2172 ( .A(n4397), .Y(n4399) );
  CLKBUFX2TS U2173 ( .A(n4394), .Y(n4396) );
  CLKBUFX2TS U2174 ( .A(n4409), .Y(n4411) );
  CLKBUFX2TS U2175 ( .A(n4403), .Y(n4405) );
  CLKBUFX2TS U2176 ( .A(n4400), .Y(n4402) );
  CLKBUFX2TS U2177 ( .A(n3823), .Y(n3822) );
  INVX2TS U2178 ( .A(n3829), .Y(n3827) );
  INVX2TS U2179 ( .A(n3813), .Y(n3811) );
  INVX2TS U2180 ( .A(n3826), .Y(n3824) );
  INVX2TS U2181 ( .A(n3819), .Y(n3817) );
  INVX2TS U2182 ( .A(n3871), .Y(n3870) );
  INVX2TS U2183 ( .A(n3919), .Y(n3918) );
  INVX2TS U2184 ( .A(n3895), .Y(n3894) );
  INVX2TS U2185 ( .A(n3868), .Y(n3867) );
  INVX2TS U2186 ( .A(n3862), .Y(n3861) );
  INVX2TS U2187 ( .A(n3850), .Y(n3849) );
  INVX2TS U2188 ( .A(n3925), .Y(n3924) );
  INVX2TS U2189 ( .A(n3922), .Y(n3921) );
  INVX2TS U2190 ( .A(n3910), .Y(n3909) );
  INVX2TS U2191 ( .A(n3904), .Y(n3903) );
  INVX2TS U2192 ( .A(n3898), .Y(n3897) );
  INVX2TS U2193 ( .A(n3889), .Y(n3888) );
  INVX2TS U2194 ( .A(n3880), .Y(n3879) );
  INVX2TS U2195 ( .A(n3865), .Y(n3864) );
  INVX2TS U2196 ( .A(n3856), .Y(n3855) );
  INVX2TS U2197 ( .A(n3916), .Y(n3915) );
  INVX2TS U2198 ( .A(n3913), .Y(n3912) );
  INVX2TS U2199 ( .A(n3901), .Y(n3900) );
  INVX2TS U2200 ( .A(n3892), .Y(n3891) );
  INVX2TS U2201 ( .A(n3859), .Y(n3858) );
  INVX2TS U2202 ( .A(n3847), .Y(n3846) );
  INVX2TS U2203 ( .A(n3838), .Y(n3837) );
  INVX2TS U2204 ( .A(n3835), .Y(n3834) );
  INVX2TS U2205 ( .A(n3832), .Y(n3831) );
  INVX2TS U2206 ( .A(n3853), .Y(n3852) );
  INVX2TS U2207 ( .A(n3883), .Y(n3882) );
  INVX2TS U2208 ( .A(n3877), .Y(n3876) );
  INVX2TS U2209 ( .A(n3874), .Y(n3873) );
  INVX2TS U2210 ( .A(n3841), .Y(n3840) );
  INVX2TS U2211 ( .A(n3907), .Y(n3906) );
  INVX2TS U2212 ( .A(n3886), .Y(n3885) );
  INVX2TS U2213 ( .A(n3844), .Y(n3843) );
  INVX2TS U2214 ( .A(n3961), .Y(n3960) );
  INVX2TS U2215 ( .A(n3958), .Y(n3957) );
  INVX2TS U2216 ( .A(n3955), .Y(n3954) );
  INVX2TS U2217 ( .A(n3949), .Y(n3948) );
  INVX2TS U2218 ( .A(n3946), .Y(n3945) );
  INVX2TS U2219 ( .A(n3952), .Y(n3951) );
  INVX2TS U2220 ( .A(n3813), .Y(n3812) );
  INVX2TS U2221 ( .A(n4270), .Y(n4269) );
  INVX2TS U2222 ( .A(n4258), .Y(n4257) );
  INVX2TS U2223 ( .A(n4273), .Y(n4272) );
  INVX2TS U2224 ( .A(n4267), .Y(n4266) );
  INVX2TS U2225 ( .A(n4264), .Y(n4263) );
  INVX2TS U2226 ( .A(n4261), .Y(n4260) );
  INVX2TS U2227 ( .A(n4234), .Y(n4233) );
  INVX2TS U2228 ( .A(n4231), .Y(n4230) );
  INVX2TS U2229 ( .A(n4228), .Y(n4227) );
  INVX2TS U2230 ( .A(n4225), .Y(n4224) );
  INVX2TS U2231 ( .A(n4222), .Y(n4221) );
  INVX2TS U2232 ( .A(n4219), .Y(n4218) );
  INVX2TS U2233 ( .A(n4213), .Y(n4212) );
  INVX2TS U2234 ( .A(n4207), .Y(n4206) );
  INVX2TS U2235 ( .A(n4204), .Y(n4203) );
  INVX2TS U2236 ( .A(n4201), .Y(n4200) );
  INVX2TS U2237 ( .A(n4198), .Y(n4197) );
  INVX2TS U2238 ( .A(n4195), .Y(n4194) );
  INVX2TS U2239 ( .A(n4189), .Y(n4188) );
  INVX2TS U2240 ( .A(n4186), .Y(n4185) );
  INVX2TS U2241 ( .A(n4183), .Y(n4182) );
  INVX2TS U2242 ( .A(n4180), .Y(n4179) );
  INVX2TS U2243 ( .A(n4177), .Y(n4176) );
  INVX2TS U2244 ( .A(n4174), .Y(n4173) );
  INVX2TS U2245 ( .A(n4171), .Y(n4170) );
  INVX2TS U2246 ( .A(n4168), .Y(n4167) );
  INVX2TS U2247 ( .A(n4165), .Y(n4164) );
  INVX2TS U2248 ( .A(n4159), .Y(n4158) );
  INVX2TS U2249 ( .A(n4156), .Y(n4155) );
  INVX2TS U2250 ( .A(n4153), .Y(n4152) );
  INVX2TS U2251 ( .A(n4147), .Y(n4146) );
  INVX2TS U2252 ( .A(n4237), .Y(n4236) );
  INVX2TS U2253 ( .A(n4216), .Y(n4215) );
  INVX2TS U2254 ( .A(n4210), .Y(n4209) );
  INVX2TS U2255 ( .A(n4192), .Y(n4191) );
  INVX2TS U2256 ( .A(n4162), .Y(n4161) );
  INVX2TS U2257 ( .A(n4150), .Y(n4149) );
  INVX2TS U2258 ( .A(n4144), .Y(n4143) );
  INVX2TS U2259 ( .A(n3826), .Y(n3825) );
  INVX2TS U2260 ( .A(n4255), .Y(n4254) );
  INVX2TS U2261 ( .A(n4252), .Y(n4251) );
  INVX2TS U2262 ( .A(n4246), .Y(n4245) );
  INVX2TS U2263 ( .A(n4249), .Y(n4248) );
  INVX2TS U2264 ( .A(n4243), .Y(n4242) );
  INVX2TS U2265 ( .A(n4240), .Y(n4239) );
  INVX2TS U2266 ( .A(n3819), .Y(n3818) );
  INVX2TS U2267 ( .A(n4081), .Y(n4080) );
  INVX2TS U2268 ( .A(n4078), .Y(n4077) );
  INVX2TS U2269 ( .A(n4075), .Y(n4074) );
  INVX2TS U2270 ( .A(n4072), .Y(n4071) );
  INVX2TS U2271 ( .A(n4069), .Y(n4068) );
  INVX2TS U2272 ( .A(n4066), .Y(n4065) );
  INVX2TS U2273 ( .A(n4060), .Y(n4059) );
  INVX2TS U2274 ( .A(n4057), .Y(n4056) );
  INVX2TS U2275 ( .A(n4054), .Y(n4053) );
  INVX2TS U2276 ( .A(n4051), .Y(n4050) );
  INVX2TS U2277 ( .A(n4048), .Y(n4047) );
  INVX2TS U2278 ( .A(n4045), .Y(n4044) );
  INVX2TS U2279 ( .A(n4039), .Y(n4038) );
  INVX2TS U2280 ( .A(n4036), .Y(n4035) );
  INVX2TS U2281 ( .A(n4033), .Y(n4032) );
  INVX2TS U2282 ( .A(n4030), .Y(n4029) );
  INVX2TS U2283 ( .A(n4027), .Y(n4026) );
  INVX2TS U2284 ( .A(n4024), .Y(n4023) );
  INVX2TS U2285 ( .A(n4021), .Y(n4020) );
  INVX2TS U2286 ( .A(n4018), .Y(n4017) );
  INVX2TS U2287 ( .A(n4015), .Y(n4014) );
  INVX2TS U2288 ( .A(n4012), .Y(n4011) );
  INVX2TS U2289 ( .A(n4009), .Y(n4008) );
  INVX2TS U2290 ( .A(n4006), .Y(n4005) );
  INVX2TS U2291 ( .A(n4003), .Y(n4002) );
  INVX2TS U2292 ( .A(n3997), .Y(n3996) );
  INVX2TS U2293 ( .A(n3994), .Y(n3993) );
  INVX2TS U2294 ( .A(n3991), .Y(n3990) );
  INVX2TS U2295 ( .A(n3988), .Y(n3987) );
  INVX2TS U2296 ( .A(n4063), .Y(n4062) );
  INVX2TS U2297 ( .A(n4042), .Y(n4041) );
  INVX2TS U2298 ( .A(n4000), .Y(n3999) );
  INVX2TS U2299 ( .A(n4102), .Y(n4101) );
  INVX2TS U2300 ( .A(n4117), .Y(n4116) );
  INVX2TS U2301 ( .A(n4111), .Y(n4110) );
  INVX2TS U2302 ( .A(n4108), .Y(n4107) );
  INVX2TS U2303 ( .A(n4105), .Y(n4104) );
  INVX2TS U2304 ( .A(n4114), .Y(n4113) );
  INVX2TS U2305 ( .A(n4099), .Y(n4098) );
  INVX2TS U2306 ( .A(n4096), .Y(n4095) );
  INVX2TS U2307 ( .A(n4093), .Y(n4092) );
  INVX2TS U2308 ( .A(n4090), .Y(n4089) );
  INVX2TS U2309 ( .A(n4087), .Y(n4086) );
  INVX2TS U2310 ( .A(n4084), .Y(n4083) );
  INVX2TS U2311 ( .A(n3937), .Y(n3936) );
  INVX2TS U2312 ( .A(n3934), .Y(n3933) );
  INVX2TS U2313 ( .A(n3931), .Y(n3930) );
  INVX2TS U2314 ( .A(n3928), .Y(n3927) );
  INVX2TS U2315 ( .A(n3943), .Y(n3942) );
  INVX2TS U2316 ( .A(n3940), .Y(n3939) );
  INVX2TS U2317 ( .A(n3829), .Y(n3828) );
  INVX2TS U2318 ( .A(n3816), .Y(n3814) );
  INVX2TS U2319 ( .A(n4273), .Y(n4271) );
  INVX2TS U2320 ( .A(n4267), .Y(n4265) );
  INVX2TS U2321 ( .A(n4261), .Y(n4259) );
  INVX2TS U2322 ( .A(n4258), .Y(n4256) );
  INVX2TS U2323 ( .A(n4264), .Y(n4262) );
  INVX2TS U2324 ( .A(n4183), .Y(n4181) );
  INVX2TS U2325 ( .A(n4231), .Y(n4229) );
  INVX2TS U2326 ( .A(n4207), .Y(n4205) );
  INVX2TS U2327 ( .A(n4180), .Y(n4178) );
  INVX2TS U2328 ( .A(n4174), .Y(n4172) );
  INVX2TS U2329 ( .A(n4162), .Y(n4160) );
  INVX2TS U2330 ( .A(n4237), .Y(n4235) );
  INVX2TS U2331 ( .A(n4234), .Y(n4232) );
  INVX2TS U2332 ( .A(n4222), .Y(n4220) );
  INVX2TS U2333 ( .A(n4216), .Y(n4214) );
  INVX2TS U2334 ( .A(n4210), .Y(n4208) );
  INVX2TS U2335 ( .A(n4201), .Y(n4199) );
  INVX2TS U2336 ( .A(n4192), .Y(n4190) );
  INVX2TS U2337 ( .A(n4177), .Y(n4175) );
  INVX2TS U2338 ( .A(n4168), .Y(n4166) );
  INVX2TS U2339 ( .A(n4228), .Y(n4226) );
  INVX2TS U2340 ( .A(n4225), .Y(n4223) );
  INVX2TS U2341 ( .A(n4213), .Y(n4211) );
  INVX2TS U2342 ( .A(n4204), .Y(n4202) );
  INVX2TS U2343 ( .A(n4171), .Y(n4169) );
  INVX2TS U2344 ( .A(n4159), .Y(n4157) );
  INVX2TS U2345 ( .A(n4150), .Y(n4148) );
  INVX2TS U2346 ( .A(n4147), .Y(n4145) );
  INVX2TS U2347 ( .A(n4144), .Y(n4142) );
  INVX2TS U2348 ( .A(n4165), .Y(n4163) );
  INVX2TS U2349 ( .A(n4195), .Y(n4193) );
  INVX2TS U2350 ( .A(n4189), .Y(n4187) );
  INVX2TS U2351 ( .A(n4186), .Y(n4184) );
  INVX2TS U2352 ( .A(n4153), .Y(n4151) );
  INVX2TS U2353 ( .A(n4270), .Y(n4268) );
  INVX2TS U2354 ( .A(n4219), .Y(n4217) );
  INVX2TS U2355 ( .A(n4198), .Y(n4196) );
  INVX2TS U2356 ( .A(n4156), .Y(n4154) );
  INVX2TS U2357 ( .A(n4856), .Y(n6285) );
  INVX2TS U2358 ( .A(n4853), .Y(n6284) );
  CLKBUFX2TS U2359 ( .A(n667), .Y(n661) );
  CLKBUFX2TS U2360 ( .A(n667), .Y(n662) );
  CLKBUFX2TS U2361 ( .A(n666), .Y(n663) );
  CLKBUFX2TS U2362 ( .A(n666), .Y(n664) );
  CLKBUFX2TS U2363 ( .A(n666), .Y(n665) );
  CLKBUFX2TS U2364 ( .A(n17), .Y(n3683) );
  CLKBUFX2TS U2365 ( .A(n287), .Y(n3606) );
  CLKBUFX2TS U2366 ( .A(n287), .Y(n3607) );
  CLKBUFX2TS U2367 ( .A(n6280), .Y(n3622) );
  CLKBUFX2TS U2368 ( .A(n17), .Y(n3684) );
  CLKBUFX2TS U2369 ( .A(n4), .Y(n3654) );
  CLKBUFX2TS U2370 ( .A(n6280), .Y(n3621) );
  INVX2TS U2371 ( .A(n5294), .Y(n6282) );
  CLKBUFX2TS U2372 ( .A(n3623), .Y(n3616) );
  CLKBUFX2TS U2373 ( .A(n6280), .Y(n3623) );
  CLKBUFX2TS U2374 ( .A(n3592), .Y(n3586) );
  CLKBUFX2TS U2375 ( .A(n6279), .Y(n3592) );
  INVX2TS U2376 ( .A(n5306), .Y(n6281) );
  CLKBUFX2TS U2377 ( .A(n660), .Y(n658) );
  CLKBUFX2TS U2378 ( .A(n660), .Y(n659) );
  NOR2X1TS U2379 ( .A(n6293), .B(n5495), .Y(n5569) );
  AOI21X1TS U2380 ( .A0(n6254), .A1(n570), .B0(n5355), .Y(n5324) );
  XNOR2X1TS U2381 ( .A(n4866), .B(n4870), .Y(n6235) );
  XNOR2X1TS U2382 ( .A(n4869), .B(n569), .Y(n4866) );
  XNOR2X1TS U2383 ( .A(n194), .B(n6235), .Y(n4867) );
  NOR2X1TS U2384 ( .A(n555), .B(n5325), .Y(n5328) );
  OAI211X1TS U2385 ( .A0(n4861), .A1(n4860), .B0(n4859), .C0(n4858), .Y(n4864)
         );
  NAND3BX1TS U2386 ( .AN(n6231), .B(n6229), .C(n4856), .Y(n4859) );
  OAI21X1TS U2387 ( .A0(n6255), .A1(n4873), .B0(n4857), .Y(n4858) );
  OAI32X1TS U2388 ( .A0(n4857), .A1(n6255), .A2(n4873), .B0(n6231), .B1(n4865), 
        .Y(n4860) );
  INVX2TS U2389 ( .A(n4862), .Y(n6253) );
  XOR2X1TS U2390 ( .A(n4875), .B(n4874), .Y(n6234) );
  NOR3X1TS U2391 ( .A(n4873), .B(n6286), .C(n6255), .Y(n4874) );
  XNOR2X1TS U2392 ( .A(n5326), .B(n4872), .Y(n4875) );
  AOI22X1TS U2393 ( .A0(n4871), .A1(n14), .B0(n4870), .B1(n4869), .Y(n4872) );
  XOR2X1TS U2394 ( .A(n4863), .B(n18), .Y(n6238) );
  NAND2X1TS U2395 ( .A(n4862), .B(n4864), .Y(n4863) );
  OAI221XLTS U2396 ( .A0(n328), .A1(n302), .B0(n3529), .B1(n24), .C0(n5588), 
        .Y(n2578) );
  AOI222XLTS U2397 ( .A0(n3811), .A1(n3473), .B0(n3825), .B1(n3483), .C0(n3818), .C1(n3521), .Y(n5588) );
  OAI221XLTS U2398 ( .A0(n431), .A1(n6244), .B0(n3398), .B1(n6271), .C0(n5586), 
        .Y(n2576) );
  AOI222XLTS U2399 ( .A0(n3811), .A1(n3365), .B0(n3825), .B1(n204), .C0(n3817), 
        .C1(n3397), .Y(n5586) );
  AOI211X1TS U2400 ( .A0(n6231), .A1(n4865), .B0(n6285), .C0(n6253), .Y(n4861)
         );
  NOR2X1TS U2401 ( .A(n6292), .B(n5326), .Y(n5561) );
  OAI33XLTS U2402 ( .A0(n6242), .A1(n6291), .A2(n5547), .B0(n3822), .B1(n6301), 
        .B2(n238), .Y(n5548) );
  NAND2X1TS U2403 ( .A(n3814), .B(n6300), .Y(n5529) );
  INVX2TS U2404 ( .A(n3822), .Y(n3821) );
  NAND2X1TS U2405 ( .A(n3814), .B(n6297), .Y(n5557) );
  NOR2X1TS U2406 ( .A(n5314), .B(n6256), .Y(n5290) );
  NOR2X1TS U2407 ( .A(n5315), .B(n6256), .Y(n5289) );
  OAI2BB2XLTS U2408 ( .B0(n281), .B1(n6242), .A0N(n281), .A1N(n3827), .Y(n5552) );
  INVX2TS U2409 ( .A(n5321), .Y(n685) );
  NAND4X1TS U2410 ( .A(n5315), .B(n5313), .C(n5311), .D(n4881), .Y(n5321) );
  AND3X2TS U2411 ( .A(n5303), .B(n5314), .C(n5312), .Y(n4881) );
  AND2X2TS U2412 ( .A(n447), .B(n196), .Y(n5507) );
  OAI222X1TS U2413 ( .A0(n3816), .A1(n5315), .B0(n3823), .B1(n5314), .C0(n256), 
        .C1(n5313), .Y(n5316) );
  OR2X2TS U2414 ( .A(n5312), .B(n6256), .Y(n566) );
  OAI211X1TS U2415 ( .A0(n3829), .A1(n5312), .B0(n5311), .C0(n6257), .Y(n5317)
         );
  INVX2TS U2416 ( .A(n5303), .Y(n6256) );
  NOR2X1TS U2417 ( .A(n6257), .B(reset), .Y(n6226) );
  NAND2X1TS U2418 ( .A(n196), .B(n4430), .Y(n6237) );
  NOR2X1TS U2419 ( .A(n5311), .B(n449), .Y(n5226) );
  INVX2TS U2420 ( .A(readIn_NORTH), .Y(n3829) );
  INVX2TS U2421 ( .A(writeIn_SOUTH), .Y(n3826) );
  INVX2TS U2422 ( .A(writeIn_WEST), .Y(n3813) );
  OAI221XLTS U2423 ( .A0(n301), .A1(n5312), .B0(n3819), .B1(n5314), .C0(n6257), 
        .Y(n5302) );
  INVX2TS U2424 ( .A(readIn_WEST), .Y(n3816) );
  INVX2TS U2425 ( .A(requesterAddressIn_EAST[5]), .Y(n4099) );
  INVX2TS U2426 ( .A(requesterAddressIn_EAST[3]), .Y(n4093) );
  INVX2TS U2427 ( .A(requesterAddressIn_EAST[4]), .Y(n4096) );
  INVX2TS U2428 ( .A(requesterAddressIn_EAST[2]), .Y(n4090) );
  INVX2TS U2429 ( .A(requesterAddressIn_EAST[1]), .Y(n4087) );
  INVX2TS U2430 ( .A(requesterAddressIn_EAST[0]), .Y(n4084) );
  INVX2TS U2431 ( .A(requesterAddressIn_WEST[4]), .Y(n3940) );
  INVX2TS U2432 ( .A(requesterAddressIn_WEST[1]), .Y(n3931) );
  INVX2TS U2433 ( .A(requesterAddressIn_WEST[0]), .Y(n3928) );
  INVX2TS U2434 ( .A(requesterAddressIn_WEST[5]), .Y(n3943) );
  INVX2TS U2435 ( .A(requesterAddressIn_WEST[3]), .Y(n3937) );
  INVX2TS U2436 ( .A(requesterAddressIn_WEST[2]), .Y(n3934) );
  INVX2TS U2437 ( .A(dataIn_EAST[31]), .Y(n4081) );
  INVX2TS U2438 ( .A(dataIn_EAST[30]), .Y(n4078) );
  INVX2TS U2439 ( .A(dataIn_EAST[29]), .Y(n4075) );
  INVX2TS U2440 ( .A(dataIn_EAST[26]), .Y(n4066) );
  INVX2TS U2441 ( .A(dataIn_EAST[24]), .Y(n4060) );
  INVX2TS U2442 ( .A(dataIn_EAST[22]), .Y(n4054) );
  INVX2TS U2443 ( .A(dataIn_EAST[21]), .Y(n4051) );
  INVX2TS U2444 ( .A(dataIn_EAST[19]), .Y(n4045) );
  INVX2TS U2445 ( .A(dataIn_EAST[17]), .Y(n4039) );
  INVX2TS U2446 ( .A(dataIn_EAST[16]), .Y(n4036) );
  INVX2TS U2447 ( .A(dataIn_EAST[14]), .Y(n4030) );
  INVX2TS U2448 ( .A(dataIn_EAST[12]), .Y(n4024) );
  INVX2TS U2449 ( .A(dataIn_EAST[11]), .Y(n4021) );
  INVX2TS U2450 ( .A(dataIn_EAST[10]), .Y(n4018) );
  INVX2TS U2451 ( .A(dataIn_EAST[8]), .Y(n4012) );
  INVX2TS U2452 ( .A(dataIn_EAST[6]), .Y(n4006) );
  INVX2TS U2453 ( .A(dataIn_EAST[3]), .Y(n3997) );
  INVX2TS U2454 ( .A(dataIn_EAST[25]), .Y(n4063) );
  INVX2TS U2455 ( .A(dataIn_EAST[18]), .Y(n4042) );
  INVX2TS U2456 ( .A(dataIn_EAST[15]), .Y(n4033) );
  INVX2TS U2457 ( .A(dataIn_EAST[13]), .Y(n4027) );
  INVX2TS U2458 ( .A(dataIn_EAST[4]), .Y(n4000) );
  INVX2TS U2459 ( .A(dataIn_EAST[28]), .Y(n4072) );
  INVX2TS U2460 ( .A(dataIn_EAST[27]), .Y(n4069) );
  INVX2TS U2461 ( .A(dataIn_EAST[23]), .Y(n4057) );
  INVX2TS U2462 ( .A(dataIn_EAST[20]), .Y(n4048) );
  INVX2TS U2463 ( .A(dataIn_EAST[9]), .Y(n4015) );
  INVX2TS U2464 ( .A(dataIn_EAST[5]), .Y(n4003) );
  INVX2TS U2465 ( .A(dataIn_EAST[2]), .Y(n3994) );
  INVX2TS U2466 ( .A(dataIn_EAST[1]), .Y(n3991) );
  INVX2TS U2467 ( .A(dataIn_EAST[0]), .Y(n3988) );
  INVX2TS U2468 ( .A(dataIn_EAST[7]), .Y(n4009) );
  INVX2TS U2469 ( .A(destinationAddressIn_EAST[5]), .Y(n4117) );
  INVX2TS U2470 ( .A(destinationAddressIn_EAST[3]), .Y(n4111) );
  INVX2TS U2471 ( .A(destinationAddressIn_EAST[1]), .Y(n4105) );
  INVX2TS U2472 ( .A(destinationAddressIn_EAST[4]), .Y(n4114) );
  INVX2TS U2473 ( .A(destinationAddressIn_EAST[0]), .Y(n4102) );
  INVX2TS U2474 ( .A(destinationAddressIn_EAST[2]), .Y(n4108) );
  INVX2TS U2475 ( .A(writeIn_EAST), .Y(n3819) );
  INVX2TS U2476 ( .A(destinationAddressIn_SOUTH[0]), .Y(n4258) );
  INVX2TS U2477 ( .A(requesterAddressIn_SOUTH[5]), .Y(n4255) );
  INVX2TS U2478 ( .A(requesterAddressIn_SOUTH[4]), .Y(n4252) );
  INVX2TS U2479 ( .A(requesterAddressIn_SOUTH[2]), .Y(n4246) );
  INVX2TS U2480 ( .A(destinationAddressIn_SOUTH[5]), .Y(n4273) );
  INVX2TS U2481 ( .A(destinationAddressIn_SOUTH[3]), .Y(n4267) );
  INVX2TS U2482 ( .A(destinationAddressIn_SOUTH[2]), .Y(n4264) );
  INVX2TS U2483 ( .A(destinationAddressIn_SOUTH[1]), .Y(n4261) );
  INVX2TS U2484 ( .A(dataIn_SOUTH[30]), .Y(n4234) );
  INVX2TS U2485 ( .A(dataIn_SOUTH[29]), .Y(n4231) );
  INVX2TS U2486 ( .A(dataIn_SOUTH[26]), .Y(n4222) );
  INVX2TS U2487 ( .A(dataIn_SOUTH[21]), .Y(n4207) );
  INVX2TS U2488 ( .A(dataIn_SOUTH[19]), .Y(n4201) );
  INVX2TS U2489 ( .A(dataIn_SOUTH[13]), .Y(n4183) );
  INVX2TS U2490 ( .A(dataIn_SOUTH[12]), .Y(n4180) );
  INVX2TS U2491 ( .A(dataIn_SOUTH[11]), .Y(n4177) );
  INVX2TS U2492 ( .A(dataIn_SOUTH[10]), .Y(n4174) );
  INVX2TS U2493 ( .A(dataIn_SOUTH[8]), .Y(n4168) );
  INVX2TS U2494 ( .A(requesterAddressIn_SOUTH[3]), .Y(n4249) );
  INVX2TS U2495 ( .A(requesterAddressIn_SOUTH[1]), .Y(n4243) );
  INVX2TS U2496 ( .A(requesterAddressIn_SOUTH[0]), .Y(n4240) );
  INVX2TS U2497 ( .A(dataIn_SOUTH[28]), .Y(n4228) );
  INVX2TS U2498 ( .A(dataIn_SOUTH[27]), .Y(n4225) );
  INVX2TS U2499 ( .A(dataIn_SOUTH[23]), .Y(n4213) );
  INVX2TS U2500 ( .A(dataIn_SOUTH[20]), .Y(n4204) );
  INVX2TS U2501 ( .A(dataIn_SOUTH[9]), .Y(n4171) );
  INVX2TS U2502 ( .A(dataIn_SOUTH[5]), .Y(n4159) );
  INVX2TS U2503 ( .A(dataIn_SOUTH[1]), .Y(n4147) );
  INVX2TS U2504 ( .A(dataIn_SOUTH[31]), .Y(n4237) );
  INVX2TS U2505 ( .A(dataIn_SOUTH[24]), .Y(n4216) );
  INVX2TS U2506 ( .A(dataIn_SOUTH[22]), .Y(n4210) );
  INVX2TS U2507 ( .A(dataIn_SOUTH[16]), .Y(n4192) );
  INVX2TS U2508 ( .A(dataIn_SOUTH[6]), .Y(n4162) );
  INVX2TS U2509 ( .A(dataIn_SOUTH[2]), .Y(n4150) );
  INVX2TS U2510 ( .A(dataIn_SOUTH[0]), .Y(n4144) );
  INVX2TS U2511 ( .A(dataIn_SOUTH[7]), .Y(n4165) );
  INVX2TS U2512 ( .A(dataIn_SOUTH[17]), .Y(n4195) );
  INVX2TS U2513 ( .A(dataIn_SOUTH[15]), .Y(n4189) );
  INVX2TS U2514 ( .A(dataIn_SOUTH[14]), .Y(n4186) );
  INVX2TS U2515 ( .A(dataIn_SOUTH[3]), .Y(n4153) );
  INVX2TS U2516 ( .A(destinationAddressIn_SOUTH[4]), .Y(n4270) );
  INVX2TS U2517 ( .A(dataIn_SOUTH[25]), .Y(n4219) );
  INVX2TS U2518 ( .A(dataIn_SOUTH[18]), .Y(n4198) );
  INVX2TS U2519 ( .A(dataIn_SOUTH[4]), .Y(n4156) );
  INVX2TS U2520 ( .A(dataIn_WEST[31]), .Y(n3925) );
  INVX2TS U2521 ( .A(dataIn_WEST[30]), .Y(n3922) );
  INVX2TS U2522 ( .A(dataIn_WEST[29]), .Y(n3919) );
  INVX2TS U2523 ( .A(dataIn_WEST[26]), .Y(n3910) );
  INVX2TS U2524 ( .A(dataIn_WEST[24]), .Y(n3904) );
  INVX2TS U2525 ( .A(dataIn_WEST[22]), .Y(n3898) );
  INVX2TS U2526 ( .A(dataIn_WEST[21]), .Y(n3895) );
  INVX2TS U2527 ( .A(dataIn_WEST[19]), .Y(n3889) );
  INVX2TS U2528 ( .A(dataIn_WEST[16]), .Y(n3880) );
  INVX2TS U2529 ( .A(dataIn_WEST[13]), .Y(n3871) );
  INVX2TS U2530 ( .A(dataIn_WEST[12]), .Y(n3868) );
  INVX2TS U2531 ( .A(dataIn_WEST[11]), .Y(n3865) );
  INVX2TS U2532 ( .A(dataIn_WEST[10]), .Y(n3862) );
  INVX2TS U2533 ( .A(dataIn_WEST[8]), .Y(n3856) );
  INVX2TS U2534 ( .A(dataIn_WEST[6]), .Y(n3850) );
  INVX2TS U2535 ( .A(dataIn_WEST[28]), .Y(n3916) );
  INVX2TS U2536 ( .A(dataIn_WEST[27]), .Y(n3913) );
  INVX2TS U2537 ( .A(dataIn_WEST[23]), .Y(n3901) );
  INVX2TS U2538 ( .A(dataIn_WEST[20]), .Y(n3892) );
  INVX2TS U2539 ( .A(dataIn_WEST[9]), .Y(n3859) );
  INVX2TS U2540 ( .A(dataIn_WEST[5]), .Y(n3847) );
  INVX2TS U2541 ( .A(dataIn_WEST[2]), .Y(n3838) );
  INVX2TS U2542 ( .A(dataIn_WEST[1]), .Y(n3835) );
  INVX2TS U2543 ( .A(dataIn_WEST[0]), .Y(n3832) );
  INVX2TS U2544 ( .A(dataIn_WEST[7]), .Y(n3853) );
  INVX2TS U2545 ( .A(dataIn_WEST[17]), .Y(n3883) );
  INVX2TS U2546 ( .A(dataIn_WEST[15]), .Y(n3877) );
  INVX2TS U2547 ( .A(dataIn_WEST[14]), .Y(n3874) );
  INVX2TS U2548 ( .A(dataIn_WEST[3]), .Y(n3841) );
  INVX2TS U2549 ( .A(dataIn_WEST[25]), .Y(n3907) );
  INVX2TS U2550 ( .A(dataIn_WEST[18]), .Y(n3886) );
  INVX2TS U2551 ( .A(dataIn_WEST[4]), .Y(n3844) );
  INVX2TS U2552 ( .A(destinationAddressIn_WEST[0]), .Y(n3946) );
  INVX2TS U2553 ( .A(destinationAddressIn_WEST[5]), .Y(n3961) );
  INVX2TS U2554 ( .A(destinationAddressIn_WEST[3]), .Y(n3955) );
  INVX2TS U2555 ( .A(destinationAddressIn_WEST[2]), .Y(n3952) );
  INVX2TS U2556 ( .A(destinationAddressIn_WEST[1]), .Y(n3949) );
  INVX2TS U2557 ( .A(destinationAddressIn_WEST[4]), .Y(n3958) );
  NOR2BX1TS U2558 ( .AN(n6237), .B(n6233), .Y(n2885) );
  AOI31X1TS U2559 ( .A0(n6232), .A1(n6285), .A2(n6231), .B0(n3574), .Y(n6233)
         );
  XNOR2X1TS U2560 ( .A(n6230), .B(n6229), .Y(n6232) );
  CLKBUFX2TS U2561 ( .A(destinationAddressIn_EAST[12]), .Y(n4136) );
  CLKBUFX2TS U2562 ( .A(destinationAddressIn_EAST[6]), .Y(n4118) );
  CLKBUFX2TS U2563 ( .A(destinationAddressIn_WEST[12]), .Y(n3980) );
  CLKBUFX2TS U2564 ( .A(destinationAddressIn_SOUTH[12]), .Y(n4292) );
  CLKBUFX2TS U2565 ( .A(destinationAddressIn_WEST[6]), .Y(n3962) );
  CLKBUFX2TS U2566 ( .A(destinationAddressIn_EAST[10]), .Y(n4130) );
  CLKBUFX2TS U2567 ( .A(destinationAddressIn_SOUTH[10]), .Y(n4286) );
  CLKBUFX2TS U2568 ( .A(destinationAddressIn_WEST[10]), .Y(n3974) );
  CLKBUFX2TS U2569 ( .A(destinationAddressIn_EAST[9]), .Y(n4127) );
  CLKBUFX2TS U2570 ( .A(destinationAddressIn_WEST[9]), .Y(n3971) );
  CLKBUFX2TS U2571 ( .A(destinationAddressIn_SOUTH[9]), .Y(n4283) );
  CLKBUFX2TS U2572 ( .A(destinationAddressIn_WEST[13]), .Y(n3983) );
  CLKBUFX2TS U2573 ( .A(destinationAddressIn_EAST[13]), .Y(n4139) );
  CLKBUFX2TS U2574 ( .A(destinationAddressIn_SOUTH[13]), .Y(n4295) );
  CLKBUFX2TS U2575 ( .A(destinationAddressIn_WEST[11]), .Y(n3977) );
  CLKBUFX2TS U2576 ( .A(destinationAddressIn_EAST[11]), .Y(n4133) );
  CLKBUFX2TS U2577 ( .A(destinationAddressIn_SOUTH[11]), .Y(n4289) );
  CLKBUFX2TS U2578 ( .A(destinationAddressIn_WEST[8]), .Y(n3968) );
  CLKBUFX2TS U2579 ( .A(destinationAddressIn_EAST[8]), .Y(n4124) );
  CLKBUFX2TS U2580 ( .A(destinationAddressIn_SOUTH[8]), .Y(n4280) );
  CLKBUFX2TS U2581 ( .A(destinationAddressIn_WEST[7]), .Y(n3965) );
  CLKBUFX2TS U2582 ( .A(destinationAddressIn_EAST[7]), .Y(n4121) );
  CLKBUFX2TS U2583 ( .A(destinationAddressIn_NORTH[0]), .Y(n4412) );
  CLKBUFX2TS U2584 ( .A(requesterAddressIn_NORTH[5]), .Y(n4409) );
  CLKBUFX2TS U2585 ( .A(requesterAddressIn_NORTH[4]), .Y(n4406) );
  CLKBUFX2TS U2586 ( .A(requesterAddressIn_NORTH[2]), .Y(n4400) );
  CLKBUFX2TS U2587 ( .A(destinationAddressIn_NORTH[5]), .Y(n4427) );
  CLKBUFX2TS U2588 ( .A(destinationAddressIn_NORTH[3]), .Y(n4421) );
  CLKBUFX2TS U2589 ( .A(destinationAddressIn_NORTH[2]), .Y(n4418) );
  CLKBUFX2TS U2590 ( .A(destinationAddressIn_NORTH[1]), .Y(n4415) );
  CLKBUFX2TS U2591 ( .A(dataIn_NORTH[30]), .Y(n4388) );
  CLKBUFX2TS U2592 ( .A(dataIn_NORTH[29]), .Y(n4385) );
  CLKBUFX2TS U2593 ( .A(dataIn_NORTH[26]), .Y(n4376) );
  CLKBUFX2TS U2594 ( .A(dataIn_NORTH[21]), .Y(n4361) );
  CLKBUFX2TS U2595 ( .A(dataIn_NORTH[19]), .Y(n4355) );
  CLKBUFX2TS U2596 ( .A(dataIn_NORTH[13]), .Y(n4337) );
  CLKBUFX2TS U2597 ( .A(dataIn_NORTH[12]), .Y(n4334) );
  CLKBUFX2TS U2598 ( .A(dataIn_NORTH[11]), .Y(n4331) );
  CLKBUFX2TS U2599 ( .A(dataIn_NORTH[10]), .Y(n4328) );
  CLKBUFX2TS U2600 ( .A(dataIn_NORTH[8]), .Y(n4322) );
  CLKBUFX2TS U2601 ( .A(requesterAddressIn_NORTH[3]), .Y(n4403) );
  CLKBUFX2TS U2602 ( .A(requesterAddressIn_NORTH[1]), .Y(n4397) );
  CLKBUFX2TS U2603 ( .A(requesterAddressIn_NORTH[0]), .Y(n4394) );
  CLKBUFX2TS U2604 ( .A(dataIn_NORTH[28]), .Y(n4382) );
  CLKBUFX2TS U2605 ( .A(dataIn_NORTH[27]), .Y(n4379) );
  CLKBUFX2TS U2606 ( .A(dataIn_NORTH[23]), .Y(n4367) );
  CLKBUFX2TS U2607 ( .A(dataIn_NORTH[20]), .Y(n4358) );
  CLKBUFX2TS U2608 ( .A(dataIn_NORTH[9]), .Y(n4325) );
  CLKBUFX2TS U2609 ( .A(dataIn_NORTH[5]), .Y(n4313) );
  CLKBUFX2TS U2610 ( .A(dataIn_NORTH[1]), .Y(n4301) );
  CLKBUFX2TS U2611 ( .A(dataIn_NORTH[31]), .Y(n4391) );
  CLKBUFX2TS U2612 ( .A(dataIn_NORTH[24]), .Y(n4370) );
  CLKBUFX2TS U2613 ( .A(dataIn_NORTH[22]), .Y(n4364) );
  CLKBUFX2TS U2614 ( .A(dataIn_NORTH[16]), .Y(n4346) );
  CLKBUFX2TS U2615 ( .A(dataIn_NORTH[6]), .Y(n4316) );
  CLKBUFX2TS U2616 ( .A(dataIn_NORTH[2]), .Y(n4304) );
  CLKBUFX2TS U2617 ( .A(dataIn_NORTH[0]), .Y(n4298) );
  CLKBUFX2TS U2618 ( .A(dataIn_NORTH[7]), .Y(n4319) );
  CLKBUFX2TS U2619 ( .A(dataIn_NORTH[17]), .Y(n4349) );
  CLKBUFX2TS U2620 ( .A(dataIn_NORTH[15]), .Y(n4343) );
  CLKBUFX2TS U2621 ( .A(dataIn_NORTH[14]), .Y(n4340) );
  CLKBUFX2TS U2622 ( .A(dataIn_NORTH[3]), .Y(n4307) );
  CLKBUFX2TS U2623 ( .A(dataIn_NORTH[25]), .Y(n4373) );
  CLKBUFX2TS U2624 ( .A(dataIn_NORTH[18]), .Y(n4352) );
  CLKBUFX2TS U2625 ( .A(dataIn_NORTH[4]), .Y(n4310) );
  CLKBUFX2TS U2626 ( .A(destinationAddressIn_NORTH[4]), .Y(n4424) );
  INVX2TS U2627 ( .A(readIn_EAST), .Y(n3823) );
  OAI21X1TS U2628 ( .A0(n6257), .A1(n6230), .B0(n4430), .Y(n6228) );
  OAI22X1TS U2629 ( .A0(n3561), .A1(n3644), .B0(n193), .B1(n6228), .Y(n2884)
         );
  XNOR2X1TS U2630 ( .A(n5326), .B(n193), .Y(n6229) );
  AOI21X1TS U2631 ( .A0(n9), .A1(n205), .B0(n4853), .Y(n4856) );
  XNOR2X1TS U2632 ( .A(n6229), .B(n4855), .Y(n4857) );
  AOI21X1TS U2633 ( .A0(n555), .A1(n6284), .B0(n4854), .Y(n4855) );
  AOI21X1TS U2634 ( .A0(n4853), .A1(n14), .B0(n194), .Y(n4854) );
  OAI22X1TS U2635 ( .A0(n6272), .A1(n655), .B0(n26), .B1(n3627), .Y(n5139) );
  OAI22X1TS U2636 ( .A0(n6273), .A1(n654), .B0(n27), .B1(n3626), .Y(n5147) );
  OAI22X1TS U2637 ( .A0(n6275), .A1(n654), .B0(n28), .B1(n3626), .Y(n5163) );
  OAI22X1TS U2638 ( .A0(n6276), .A1(n654), .B0(n29), .B1(n3626), .Y(n5171) );
  OAI22X1TS U2639 ( .A0(n6274), .A1(n654), .B0(n30), .B1(n3626), .Y(n5155) );
  OAI22X1TS U2640 ( .A0(n6277), .A1(n653), .B0(n31), .B1(n3625), .Y(n5179) );
  CLKBUFX2TS U2641 ( .A(n5309), .Y(n667) );
  CLKBUFX2TS U2642 ( .A(n5309), .Y(n666) );
  INVX2TS U2643 ( .A(n5307), .Y(n6280) );
  INVX2TS U2644 ( .A(n5297), .Y(n6279) );
  NOR2X1TS U2645 ( .A(n6230), .B(n193), .Y(n5306) );
  INVX2TS U2646 ( .A(n348), .Y(n6278) );
  CLKBUFX2TS U2647 ( .A(n668), .Y(n660) );
  CLKBUFX2TS U2648 ( .A(n5309), .Y(n668) );
  AOI222XLTS U2649 ( .A0(n4296), .A1(n1602), .B0(destinationAddressIn_EAST[13]), .B1(n869), .C0(n3985), .C1(n3212), .Y(n5379) );
  AOI222XLTS U2650 ( .A0(n3811), .A1(n754), .B0(n3824), .B1(n716), .C0(n3817), 
        .C1(n2), .Y(n5574) );
  AOI222XLTS U2651 ( .A0(n4290), .A1(n1602), .B0(destinationAddressIn_EAST[11]), .B1(n864), .C0(n3979), .C1(n3212), .Y(n5381) );
  AOI222XLTS U2652 ( .A0(n4284), .A1(n1653), .B0(destinationAddressIn_EAST[9]), 
        .B1(n867), .C0(n3973), .C1(n3213), .Y(n5383) );
  AOI222XLTS U2653 ( .A0(n4278), .A1(n1653), .B0(destinationAddressIn_EAST[7]), 
        .B1(n863), .C0(n3967), .C1(n3214), .Y(n5385) );
  AOI222XLTS U2654 ( .A0(n3824), .A1(n1654), .B0(n3818), .B1(n863), .C0(n3812), 
        .C1(n3214), .Y(n5579) );
  AOI222XLTS U2655 ( .A0(n4293), .A1(n1602), .B0(destinationAddressIn_EAST[12]), .B1(n864), .C0(n3982), .C1(n3212), .Y(n5380) );
  AOI222XLTS U2656 ( .A0(n4287), .A1(n1602), .B0(destinationAddressIn_EAST[10]), .B1(n864), .C0(n3976), .C1(n3213), .Y(n5382) );
  AOI222XLTS U2657 ( .A0(n4281), .A1(n1653), .B0(destinationAddressIn_EAST[8]), 
        .B1(n863), .C0(n3970), .C1(n3213), .Y(n5384) );
  AOI222XLTS U2658 ( .A0(n4275), .A1(n1653), .B0(destinationAddressIn_EAST[6]), 
        .B1(n863), .C0(n3964), .C1(n3214), .Y(n5386) );
  AOI222XLTS U2659 ( .A0(n3981), .A1(n752), .B0(n4294), .B1(n715), .C0(n4137), 
        .C1(n554), .Y(n5335) );
  AOI222XLTS U2660 ( .A0(n3969), .A1(n753), .B0(n4282), .B1(n716), .C0(n4125), 
        .C1(n551), .Y(n5339) );
  AOI222XLTS U2661 ( .A0(n3984), .A1(n752), .B0(n4297), .B1(n735), .C0(n4140), 
        .C1(n551), .Y(n5334) );
  AOI222XLTS U2662 ( .A0(n3975), .A1(n752), .B0(n4288), .B1(n715), .C0(n4131), 
        .C1(n554), .Y(n5337) );
  AOI222XLTS U2663 ( .A0(n3963), .A1(n753), .B0(n4276), .B1(n716), .C0(n4119), 
        .C1(n551), .Y(n5341) );
  AOI222XLTS U2664 ( .A0(n3978), .A1(n752), .B0(n4291), .B1(n715), .C0(n4134), 
        .C1(n554), .Y(n5336) );
  AOI222XLTS U2665 ( .A0(n3972), .A1(n753), .B0(n4285), .B1(n715), .C0(n4128), 
        .C1(n551), .Y(n5338) );
  AOI222XLTS U2666 ( .A0(n3966), .A1(n753), .B0(n4279), .B1(n729), .C0(n4122), 
        .C1(n554), .Y(n5340) );
  NOR2X1TS U2667 ( .A(selectBit_SOUTH), .B(selectBit_NORTH), .Y(n4880) );
  INVX2TS U2668 ( .A(selectBit_EAST), .Y(n6241) );
  OAI22X1TS U2669 ( .A0(n6234), .A1(n6237), .B0(n5326), .B1(n6236), .Y(n2886)
         );
  INVX2TS U2670 ( .A(readReady), .Y(n6239) );
  NOR2X1TS U2671 ( .A(selectBit_WEST), .B(readReady), .Y(n4879) );
  INVX2TS U2672 ( .A(selectBit_WEST), .Y(n6240) );
  NAND2X1TS U2673 ( .A(n4868), .B(n4867), .Y(n4877) );
  XNOR2X1TS U2674 ( .A(n257), .B(n6234), .Y(n4876) );
  OAI221XLTS U2675 ( .A0(n268), .A1(n6250), .B0(n4789), .B1(n686), .C0(n5474), 
        .Y(n2536) );
  OAI221XLTS U2676 ( .A0(n268), .A1(n6248), .B0(n4801), .B1(n687), .C0(n5476), 
        .Y(n2538) );
  OAI221XLTS U2677 ( .A0(n366), .A1(n6247), .B0(n4809), .B1(n687), .C0(n5477), 
        .Y(n2539) );
  AOI222XLTS U2678 ( .A0(n4284), .A1(n3463), .B0(n4129), .B1(n3418), .C0(n3973), .C1(n3712), .Y(n5477) );
  OAI221XLTS U2679 ( .A0(n437), .A1(n303), .B0(n4833), .B1(n688), .C0(n5480), 
        .Y(n2542) );
  AOI222XLTS U2680 ( .A0(n4275), .A1(n3463), .B0(n4120), .B1(n3418), .C0(n3964), .C1(n3708), .Y(n5480) );
  OAI221XLTS U2681 ( .A0(n5578), .A1(n6251), .B0(n4778), .B1(n838), .C0(n5356), 
        .Y(n2465) );
  OAI221XLTS U2682 ( .A0(n331), .A1(n310), .B0(n4786), .B1(n837), .C0(n5357), 
        .Y(n2466) );
  AOI222XLTS U2683 ( .A0(n4137), .A1(n777), .B0(destinationAddressIn_SOUTH[12]), .B1(n801), .C0(n3982), .C1(n827), .Y(n5357) );
  OAI221XLTS U2684 ( .A0(n330), .A1(n6249), .B0(n4796), .B1(n838), .C0(n5358), 
        .Y(n2467) );
  AOI222XLTS U2685 ( .A0(n4134), .A1(n777), .B0(destinationAddressIn_SOUTH[11]), .B1(n797), .C0(n3979), .C1(n827), .Y(n5358) );
  OAI221XLTS U2686 ( .A0(n331), .A1(n313), .B0(n4802), .B1(n838), .C0(n5359), 
        .Y(n2468) );
  AOI222XLTS U2687 ( .A0(n4131), .A1(n777), .B0(destinationAddressIn_SOUTH[10]), .B1(n802), .C0(n3976), .C1(n827), .Y(n5359) );
  OAI221XLTS U2688 ( .A0(n330), .A1(n316), .B0(n4814), .B1(n839), .C0(n5360), 
        .Y(n2469) );
  AOI222XLTS U2689 ( .A0(n4128), .A1(n777), .B0(destinationAddressIn_SOUTH[9]), 
        .B1(n787), .C0(n3973), .C1(n827), .Y(n5360) );
  OAI221XLTS U2690 ( .A0(n331), .A1(n6246), .B0(n4818), .B1(n839), .C0(n5361), 
        .Y(n2470) );
  AOI222XLTS U2691 ( .A0(n4125), .A1(n779), .B0(destinationAddressIn_SOUTH[8]), 
        .B1(n787), .C0(n3970), .C1(n834), .Y(n5361) );
  OAI221XLTS U2692 ( .A0(n330), .A1(n6245), .B0(n4826), .B1(n839), .C0(n5362), 
        .Y(n2471) );
  AOI222XLTS U2693 ( .A0(n4122), .A1(n779), .B0(n4277), .B1(n787), .C0(n3967), 
        .C1(n6130), .Y(n5362) );
  OAI221XLTS U2694 ( .A0(n331), .A1(n304), .B0(n4838), .B1(n838), .C0(n5363), 
        .Y(n2472) );
  AOI222XLTS U2695 ( .A0(n4119), .A1(n779), .B0(n4274), .B1(n787), .C0(n3964), 
        .C1(n835), .Y(n5363) );
  OAI221XLTS U2696 ( .A0(n330), .A1(n302), .B0(n836), .B1(n151), .C0(n5577), 
        .Y(n2572) );
  OAI221XLTS U2697 ( .A0(n249), .A1(n322), .B0(n4799), .B1(n686), .C0(n5475), 
        .Y(n2537) );
  OAI221XLTS U2698 ( .A0(n249), .A1(n325), .B0(n4823), .B1(n687), .C0(n5478), 
        .Y(n2540) );
  AOI222XLTS U2699 ( .A0(n4281), .A1(n3457), .B0(n4126), .B1(n3419), .C0(n3970), .C1(n3711), .Y(n5478) );
  OAI221XLTS U2700 ( .A0(n437), .A1(n307), .B0(n4829), .B1(n687), .C0(n5479), 
        .Y(n2541) );
  AOI222XLTS U2701 ( .A0(n4278), .A1(n3457), .B0(n4123), .B1(n3419), .C0(n3967), .C1(n6304), .Y(n5479) );
  OAI221XLTS U2702 ( .A0(n249), .A1(n319), .B0(n4779), .B1(n686), .C0(n5473), 
        .Y(n2535) );
  AOI222XLTS U2703 ( .A0(n4296), .A1(n3461), .B0(n4141), .B1(n3418), .C0(n3985), .C1(n3711), .Y(n5473) );
  OAI221XLTS U2704 ( .A0(n437), .A1(n302), .B0(n686), .B1(n152), .C0(n5587), 
        .Y(n2577) );
  AOI222XLTS U2705 ( .A0(n3824), .A1(n3461), .B0(n3818), .B1(n3419), .C0(n3812), .C1(n3708), .Y(n5587) );
  OAI221XLTS U2706 ( .A0(n3245), .A1(n301), .B0(n3260), .B1(n155), .C0(n5583), 
        .Y(n2574) );
  AOI222XLTS U2707 ( .A0(n3811), .A1(n361), .B0(n3825), .B1(n294), .C0(n3818), 
        .C1(n546), .Y(n5583) );
  OAI221XLTS U2708 ( .A0(n336), .A1(n302), .B0(n3332), .B1(n153), .C0(n5584), 
        .Y(n2575) );
  AOI222XLTS U2709 ( .A0(n3824), .A1(n3276), .B0(n3812), .B1(n3297), .C0(n3817), .C1(n3324), .Y(n5584) );
  OAI221XLTS U2710 ( .A0(n3243), .A1(n323), .B0(n4795), .B1(n3264), .C0(n5407), 
        .Y(n2495) );
  AOI222XLTS U2711 ( .A0(n3978), .A1(n362), .B0(n4291), .B1(n295), .C0(n4135), 
        .C1(n546), .Y(n5407) );
  OAI221XLTS U2712 ( .A0(n3245), .A1(n305), .B0(n4835), .B1(n3264), .C0(n5412), 
        .Y(n2500) );
  AOI222XLTS U2713 ( .A0(n3963), .A1(n248), .B0(n4276), .B1(n295), .C0(n4120), 
        .C1(n546), .Y(n5412) );
  OAI221XLTS U2714 ( .A0(n337), .A1(n311), .B0(n4787), .B1(n3333), .C0(n5428), 
        .Y(n2508) );
  AOI222XLTS U2715 ( .A0(n4293), .A1(n3275), .B0(n3982), .B1(n3284), .C0(n4138), .C1(n3331), .Y(n5428) );
  OAI221XLTS U2716 ( .A0(n337), .A1(n322), .B0(n4793), .B1(n3334), .C0(n5429), 
        .Y(n2509) );
  AOI222XLTS U2717 ( .A0(n4290), .A1(n3275), .B0(n3979), .B1(n3284), .C0(n4135), .C1(n3331), .Y(n5429) );
  OAI221XLTS U2718 ( .A0(n336), .A1(n314), .B0(n4803), .B1(n3334), .C0(n5430), 
        .Y(n2510) );
  AOI222XLTS U2719 ( .A0(n4287), .A1(n3275), .B0(n3976), .B1(n3284), .C0(n4132), .C1(n3325), .Y(n5430) );
  OAI221XLTS U2720 ( .A0(n337), .A1(n326), .B0(n4821), .B1(n3335), .C0(n5432), 
        .Y(n2512) );
  AOI222XLTS U2721 ( .A0(n4281), .A1(n3276), .B0(n3970), .B1(n3285), .C0(n4126), .C1(n3324), .Y(n5432) );
  OAI221XLTS U2722 ( .A0(n5585), .A1(n308), .B0(n4825), .B1(n3335), .C0(n5433), 
        .Y(n2513) );
  AOI222XLTS U2723 ( .A0(n4278), .A1(n3276), .B0(n3967), .B1(n3285), .C0(n4123), .C1(n3324), .Y(n5433) );
  OAI221XLTS U2724 ( .A0(n336), .A1(n303), .B0(n4837), .B1(n3334), .C0(n5434), 
        .Y(n2514) );
  AOI222XLTS U2725 ( .A0(n4275), .A1(n3276), .B0(n3964), .B1(n3285), .C0(n4120), .C1(n3324), .Y(n5434) );
  OAI221XLTS U2726 ( .A0(n329), .A1(n317), .B0(n4813), .B1(n3532), .C0(n5502), 
        .Y(n2553) );
  AOI222XLTS U2727 ( .A0(n3972), .A1(n3474), .B0(n4285), .B1(n3482), .C0(n4129), .C1(n3522), .Y(n5502) );
  OAI221XLTS U2728 ( .A0(n3243), .A1(n310), .B0(n4788), .B1(n3261), .C0(n5406), 
        .Y(n2494) );
  AOI222XLTS U2729 ( .A0(n3981), .A1(n354), .B0(n4294), .B1(n376), .C0(n4138), 
        .C1(n546), .Y(n5406) );
  OAI221XLTS U2730 ( .A0(n3244), .A1(n316), .B0(n4810), .B1(n3262), .C0(n5409), 
        .Y(n2497) );
  AOI222XLTS U2731 ( .A0(n3972), .A1(n354), .B0(n4285), .B1(n275), .C0(n4129), 
        .C1(n5582), .Y(n5409) );
  OAI221XLTS U2732 ( .A0(n3244), .A1(n325), .B0(n4824), .B1(n3263), .C0(n5410), 
        .Y(n2498) );
  AOI222XLTS U2733 ( .A0(n3969), .A1(n356), .B0(n4282), .B1(n294), .C0(n4126), 
        .C1(n548), .Y(n5410) );
  OAI221XLTS U2734 ( .A0(n5589), .A1(n320), .B0(n4780), .B1(n3531), .C0(n5498), 
        .Y(n2549) );
  AOI222XLTS U2735 ( .A0(n3984), .A1(n3479), .B0(n4297), .B1(n3481), .C0(n4141), .C1(n3526), .Y(n5498) );
  OAI221XLTS U2736 ( .A0(n328), .A1(n310), .B0(n4790), .B1(n3530), .C0(n5499), 
        .Y(n2550) );
  AOI222XLTS U2737 ( .A0(n3981), .A1(n3475), .B0(n4294), .B1(n3481), .C0(n4138), .C1(n3522), .Y(n5499) );
  OAI221XLTS U2738 ( .A0(n329), .A1(n322), .B0(n4794), .B1(n3531), .C0(n5500), 
        .Y(n2551) );
  AOI222XLTS U2739 ( .A0(n3978), .A1(n3476), .B0(n4291), .B1(n3481), .C0(n4135), .C1(n3522), .Y(n5500) );
  OAI221XLTS U2740 ( .A0(n329), .A1(n313), .B0(n4804), .B1(n3531), .C0(n5501), 
        .Y(n2552) );
  AOI222XLTS U2741 ( .A0(n3975), .A1(n3477), .B0(n4288), .B1(n3481), .C0(n4132), .C1(n3522), .Y(n5501) );
  OAI221XLTS U2742 ( .A0(n328), .A1(n325), .B0(n4820), .B1(n3532), .C0(n5503), 
        .Y(n2554) );
  AOI222XLTS U2743 ( .A0(n3969), .A1(n3473), .B0(n4282), .B1(n3482), .C0(n4126), .C1(n3521), .Y(n5503) );
  OAI221XLTS U2744 ( .A0(n329), .A1(n307), .B0(n4830), .B1(n3532), .C0(n5504), 
        .Y(n2555) );
  AOI222XLTS U2745 ( .A0(n3966), .A1(n3473), .B0(n4279), .B1(n3482), .C0(n4123), .C1(n3521), .Y(n5504) );
  OAI221XLTS U2746 ( .A0(n5589), .A1(n304), .B0(n4836), .B1(n3531), .C0(n5505), 
        .Y(n2556) );
  AOI222XLTS U2747 ( .A0(n3963), .A1(n3473), .B0(n4276), .B1(n3482), .C0(n4120), .C1(n3521), .Y(n5505) );
  OAI221XLTS U2748 ( .A0(n3243), .A1(n319), .B0(n4781), .B1(n3261), .C0(n5405), 
        .Y(n2493) );
  AOI222XLTS U2749 ( .A0(n3984), .A1(n360), .B0(n4297), .B1(n295), .C0(n4141), 
        .C1(n548), .Y(n5405) );
  OAI221XLTS U2750 ( .A0(n3244), .A1(n313), .B0(n4807), .B1(n3262), .C0(n5408), 
        .Y(n2496) );
  AOI222XLTS U2751 ( .A0(n3975), .A1(n355), .B0(n4288), .B1(n294), .C0(n4132), 
        .C1(n548), .Y(n5408) );
  OAI221XLTS U2752 ( .A0(n3246), .A1(n307), .B0(n4831), .B1(n3263), .C0(n5411), 
        .Y(n2499) );
  AOI222XLTS U2753 ( .A0(n3966), .A1(n355), .B0(n4279), .B1(n294), .C0(n4123), 
        .C1(n548), .Y(n5411) );
  OAI221XLTS U2754 ( .A0(n337), .A1(n319), .B0(n4783), .B1(n3334), .C0(n5427), 
        .Y(n2507) );
  OAI221XLTS U2755 ( .A0(n5585), .A1(n316), .B0(n4815), .B1(n3335), .C0(n5431), 
        .Y(n2511) );
  AOI222XLTS U2756 ( .A0(n4284), .A1(n3275), .B0(n3973), .B1(n3285), .C0(n4129), .C1(n6175), .Y(n5431) );
  OAI221XLTS U2757 ( .A0(n427), .A1(n319), .B0(n4782), .B1(n3400), .C0(n5450), 
        .Y(n2521) );
  OAI221XLTS U2758 ( .A0(n431), .A1(n310), .B0(n4792), .B1(n3399), .C0(n5451), 
        .Y(n2522) );
  AOI222XLTS U2759 ( .A0(n3981), .A1(n3357), .B0(n4294), .B1(n212), .C0(n4137), 
        .C1(n3390), .Y(n5451) );
  OAI221XLTS U2760 ( .A0(n425), .A1(n322), .B0(n4798), .B1(n3400), .C0(n5452), 
        .Y(n2523) );
  AOI222XLTS U2761 ( .A0(n3978), .A1(n3357), .B0(n4291), .B1(n198), .C0(n4134), 
        .C1(n3390), .Y(n5452) );
  OAI221XLTS U2762 ( .A0(n429), .A1(n313), .B0(n4808), .B1(n3400), .C0(n5453), 
        .Y(n2524) );
  AOI222XLTS U2763 ( .A0(n3975), .A1(n3357), .B0(n4288), .B1(n201), .C0(n4131), 
        .C1(n3390), .Y(n5453) );
  OAI221XLTS U2764 ( .A0(n427), .A1(n316), .B0(n4812), .B1(n3401), .C0(n5454), 
        .Y(n2525) );
  AOI222XLTS U2765 ( .A0(n3972), .A1(n3357), .B0(n4285), .B1(n204), .C0(n4128), 
        .C1(n3390), .Y(n5454) );
  OAI221XLTS U2766 ( .A0(n427), .A1(n325), .B0(n4822), .B1(n3401), .C0(n5455), 
        .Y(n2526) );
  AOI222XLTS U2767 ( .A0(n3969), .A1(n3365), .B0(n4282), .B1(n201), .C0(n4125), 
        .C1(n3397), .Y(n5455) );
  OAI221XLTS U2768 ( .A0(n425), .A1(n307), .B0(n4828), .B1(n3401), .C0(n5456), 
        .Y(n2527) );
  AOI222XLTS U2769 ( .A0(n3966), .A1(n3366), .B0(n4279), .B1(n207), .C0(n4122), 
        .C1(n3393), .Y(n5456) );
  OAI221XLTS U2770 ( .A0(n431), .A1(n304), .B0(n4834), .B1(n3400), .C0(n5457), 
        .Y(n2528) );
  AOI222XLTS U2771 ( .A0(n3963), .A1(n3358), .B0(n4276), .B1(n213), .C0(n4119), 
        .C1(n3394), .Y(n5457) );
  AOI22X1TS U2772 ( .A0(n3267), .A1(n4247), .B0(n3724), .B1(n4404), .Y(n6167)
         );
  AOI222XLTS U2773 ( .A0(n3326), .A1(n4092), .B0(n3306), .B1(n182), .C0(n3293), 
        .C1(n3936), .Y(n6166) );
  AOI22X1TS U2774 ( .A0(n3267), .A1(n4244), .B0(n3724), .B1(n4401), .Y(n6169)
         );
  AOI222XLTS U2775 ( .A0(n3331), .A1(n4089), .B0(n3306), .B1(n177), .C0(n3294), 
        .C1(n3933), .Y(n6168) );
  AOI22X1TS U2776 ( .A0(n3267), .A1(n4241), .B0(n3724), .B1(n4398), .Y(n6171)
         );
  AOI222XLTS U2777 ( .A0(n3327), .A1(n4086), .B0(n3306), .B1(n172), .C0(n3295), 
        .C1(n3930), .Y(n6170) );
  AOI22X1TS U2778 ( .A0(n3268), .A1(n4238), .B0(n3724), .B1(n4395), .Y(n6177)
         );
  AOI222XLTS U2779 ( .A0(n3326), .A1(n4083), .B0(n3307), .B1(n167), .C0(n6173), 
        .C1(n3927), .Y(n6176) );
  AOI22X1TS U2780 ( .A0(n3268), .A1(n4253), .B0(n3725), .B1(n4410), .Y(n6163)
         );
  AOI222XLTS U2781 ( .A0(n3329), .A1(n4098), .B0(n3307), .B1(n159), .C0(n3298), 
        .C1(n3942), .Y(n6162) );
  AOI22X1TS U2782 ( .A0(n3267), .A1(n4250), .B0(n3725), .B1(n4407), .Y(n6165)
         );
  AOI222XLTS U2783 ( .A0(n3327), .A1(n4095), .B0(n3307), .B1(n186), .C0(n6173), 
        .C1(n3939), .Y(n6164) );
  AOI22X1TS U2784 ( .A0(n3220), .A1(n191), .B0(n273), .B1(n4253), .Y(n6149) );
  AOI222XLTS U2785 ( .A0(\requesterAddressbuffer[3][5] ), .A1(n3258), .B0(n360), .B1(n3942), .C0(n3233), .C1(n4411), .Y(n6148) );
  AOI22X1TS U2786 ( .A0(n3220), .A1(n185), .B0(n272), .B1(n4250), .Y(n6151) );
  AOI222XLTS U2787 ( .A0(\requesterAddressbuffer[3][4] ), .A1(n3258), .B0(n355), .B1(n3939), .C0(n3233), .C1(n4408), .Y(n6150) );
  AOI22X1TS U2788 ( .A0(n3220), .A1(n180), .B0(n370), .B1(n4247), .Y(n6153) );
  AOI222XLTS U2789 ( .A0(\requesterAddressbuffer[3][3] ), .A1(n3259), .B0(n248), .B1(n3936), .C0(n3232), .C1(n4405), .Y(n6152) );
  AOI22X1TS U2790 ( .A0(n3219), .A1(n175), .B0(n371), .B1(n4244), .Y(n6155) );
  AOI222XLTS U2791 ( .A0(\requesterAddressbuffer[3][2] ), .A1(n3259), .B0(n356), .B1(n3933), .C0(n3232), .C1(n4402), .Y(n6154) );
  AOI22X1TS U2792 ( .A0(n3218), .A1(n170), .B0(n286), .B1(n4241), .Y(n6157) );
  AOI222XLTS U2793 ( .A0(\requesterAddressbuffer[3][1] ), .A1(n3259), .B0(n362), .B1(n3930), .C0(n3232), .C1(n4399), .Y(n6156) );
  AOI22X1TS U2794 ( .A0(n3220), .A1(n166), .B0(n285), .B1(n4238), .Y(n6161) );
  AOI222XLTS U2795 ( .A0(\requesterAddressbuffer[3][0] ), .A1(n3259), .B0(n354), .B1(n3927), .C0(n3232), .C1(n4396), .Y(n6160) );
  AOI22X1TS U2796 ( .A0(n770), .A1(n4097), .B0(n3768), .B1(n4410), .Y(n6118)
         );
  AOI222XLTS U2797 ( .A0(n819), .A1(n3941), .B0(n816), .B1(n190), .C0(n798), 
        .C1(n4254), .Y(n6117) );
  AOI22X1TS U2798 ( .A0(n769), .A1(n4094), .B0(n3768), .B1(n4407), .Y(n6120)
         );
  AOI222XLTS U2799 ( .A0(n818), .A1(n3938), .B0(n815), .B1(n187), .C0(n800), 
        .C1(n4251), .Y(n6119) );
  AOI22X1TS U2800 ( .A0(n769), .A1(n4091), .B0(n3767), .B1(n4404), .Y(n6122)
         );
  AOI222XLTS U2801 ( .A0(n818), .A1(n3935), .B0(n812), .B1(n183), .C0(n800), 
        .C1(n4248), .Y(n6121) );
  AOI22X1TS U2802 ( .A0(n769), .A1(n4088), .B0(n3767), .B1(n4401), .Y(n6124)
         );
  AOI222XLTS U2803 ( .A0(n818), .A1(n3932), .B0(n812), .B1(n178), .C0(n801), 
        .C1(n4245), .Y(n6123) );
  AOI22X1TS U2804 ( .A0(n769), .A1(n4085), .B0(n3767), .B1(n4398), .Y(n6126)
         );
  AOI222XLTS U2805 ( .A0(n818), .A1(n3929), .B0(n812), .B1(n173), .C0(n796), 
        .C1(n4242), .Y(n6125) );
  AOI22X1TS U2806 ( .A0(n770), .A1(n4082), .B0(n3767), .B1(n4395), .Y(n6132)
         );
  AOI222XLTS U2807 ( .A0(n819), .A1(n3926), .B0(n817), .B1(n168), .C0(n798), 
        .C1(n4239), .Y(n6131) );
  AOI22X1TS U2808 ( .A0(n3351), .A1(n3941), .B0(n426), .B1(n4410), .Y(n6179)
         );
  AOI222XLTS U2809 ( .A0(n3382), .A1(n4098), .B0(n3374), .B1(n191), .C0(n436), 
        .C1(n4254), .Y(n6178) );
  AOI22X1TS U2810 ( .A0(n3350), .A1(n3938), .B0(n3716), .B1(n4407), .Y(n6181)
         );
  AOI222XLTS U2811 ( .A0(n3381), .A1(n4095), .B0(n3374), .B1(n188), .C0(n206), 
        .C1(n4251), .Y(n6180) );
  AOI22X1TS U2812 ( .A0(n3350), .A1(n3935), .B0(n3717), .B1(n4404), .Y(n6183)
         );
  AOI222XLTS U2813 ( .A0(n3381), .A1(n4092), .B0(n3373), .B1(n180), .C0(n211), 
        .C1(n4248), .Y(n6182) );
  AOI22X1TS U2814 ( .A0(n3350), .A1(n3932), .B0(n3716), .B1(n4401), .Y(n6185)
         );
  AOI222XLTS U2815 ( .A0(n3381), .A1(n4089), .B0(n3373), .B1(n175), .C0(n206), 
        .C1(n4245), .Y(n6184) );
  AOI22X1TS U2816 ( .A0(n3350), .A1(n3929), .B0(n428), .B1(n4398), .Y(n6187)
         );
  AOI222XLTS U2817 ( .A0(n3381), .A1(n4086), .B0(n3373), .B1(n170), .C0(n201), 
        .C1(n4242), .Y(n6186) );
  AOI22X1TS U2818 ( .A0(n3351), .A1(n3926), .B0(n3716), .B1(n4395), .Y(n6193)
         );
  AOI222XLTS U2819 ( .A0(n3382), .A1(n4083), .B0(n3374), .B1(n165), .C0(n209), 
        .C1(n4239), .Y(n6192) );
  AOI22X1TS U2820 ( .A0(n3434), .A1(n186), .B0(n3416), .B1(n4094), .Y(n6197)
         );
  AOI222XLTS U2821 ( .A0(\requesterAddressbuffer[6][4] ), .A1(n698), .B0(n3456), .B1(n4250), .C0(n364), .C1(n4408), .Y(n6196) );
  AOI22X1TS U2822 ( .A0(n3433), .A1(n176), .B0(n3416), .B1(n4088), .Y(n6201)
         );
  AOI222XLTS U2823 ( .A0(\requesterAddressbuffer[6][2] ), .A1(n701), .B0(n3456), .B1(n4244), .C0(n3714), .C1(n4402), .Y(n6200) );
  AOI22X1TS U2824 ( .A0(n4271), .A1(n3453), .B0(n4428), .B1(n369), .Y(n5483)
         );
  AOI22X1TS U2825 ( .A0(n4229), .A1(n3454), .B0(n4386), .B1(n367), .Y(n5659)
         );
  AOI22X1TS U2826 ( .A0(n4211), .A1(n3452), .B0(n4368), .B1(n250), .Y(n5671)
         );
  AOI22X1TS U2827 ( .A0(n4205), .A1(n3452), .B0(n4362), .B1(n3714), .Y(n5675)
         );
  AOI22X1TS U2828 ( .A0(n4202), .A1(n3452), .B0(n4359), .B1(n369), .Y(n5677)
         );
  AOI22X1TS U2829 ( .A0(n4181), .A1(n3450), .B0(n4338), .B1(n364), .Y(n5691)
         );
  AOI22X1TS U2830 ( .A0(n4178), .A1(n3450), .B0(n4335), .B1(n365), .Y(n5693)
         );
  AOI22X1TS U2831 ( .A0(n4172), .A1(n3449), .B0(n4329), .B1(n267), .Y(n5697)
         );
  AOI22X1TS U2832 ( .A0(n4160), .A1(n3448), .B0(n4317), .B1(n365), .Y(n5705)
         );
  AOI22X1TS U2833 ( .A0(n3956), .A1(n3472), .B0(n4425), .B1(n3697), .Y(n5511)
         );
  AOI222XLTS U2834 ( .A0(n4113), .A1(n3520), .B0(readRequesterAddress[4]), 
        .B1(n3509), .C0(n4269), .C1(n3490), .Y(n5510) );
  AOI22X1TS U2835 ( .A0(n3944), .A1(n3474), .B0(n4413), .B1(n3685), .Y(n5519)
         );
  AOI222XLTS U2836 ( .A0(n4101), .A1(n3519), .B0(readRequesterAddress[0]), 
        .B1(n3498), .C0(n4257), .C1(n3491), .Y(n5518) );
  AOI22X1TS U2837 ( .A0(n4235), .A1(n3458), .B0(n4392), .B1(n270), .Y(n5655)
         );
  AOI22X1TS U2838 ( .A0(n4232), .A1(n3454), .B0(n4389), .B1(n267), .Y(n5657)
         );
  AOI22X1TS U2839 ( .A0(n4226), .A1(n3454), .B0(n4383), .B1(n369), .Y(n5661)
         );
  AOI22X1TS U2840 ( .A0(n4223), .A1(n3454), .B0(n4380), .B1(n250), .Y(n5663)
         );
  AOI22X1TS U2841 ( .A0(n4220), .A1(n3453), .B0(n4377), .B1(n3714), .Y(n5665)
         );
  AOI22X1TS U2842 ( .A0(n4214), .A1(n3453), .B0(n4371), .B1(n368), .Y(n5669)
         );
  AOI22X1TS U2843 ( .A0(n4208), .A1(n3452), .B0(n4365), .B1(n368), .Y(n5673)
         );
  AOI22X1TS U2844 ( .A0(n4199), .A1(n3451), .B0(n4356), .B1(n270), .Y(n5679)
         );
  AOI22X1TS U2845 ( .A0(n4193), .A1(n3451), .B0(n4350), .B1(n363), .Y(n5683)
         );
  AOI22X1TS U2846 ( .A0(n4190), .A1(n3451), .B0(n4347), .B1(n250), .Y(n5685)
         );
  AOI22X1TS U2847 ( .A0(n4187), .A1(n3450), .B0(n4344), .B1(n363), .Y(n5687)
         );
  AOI22X1TS U2848 ( .A0(n4184), .A1(n3450), .B0(n4341), .B1(n365), .Y(n5689)
         );
  AOI22X1TS U2849 ( .A0(n4175), .A1(n3449), .B0(n4332), .B1(n364), .Y(n5695)
         );
  AOI22X1TS U2850 ( .A0(n4169), .A1(n3449), .B0(n4326), .B1(n269), .Y(n5699)
         );
  AOI22X1TS U2851 ( .A0(n4166), .A1(n3449), .B0(n4323), .B1(n363), .Y(n5701)
         );
  AOI22X1TS U2852 ( .A0(n4163), .A1(n3448), .B0(n4320), .B1(n270), .Y(n5703)
         );
  AOI22X1TS U2853 ( .A0(n4157), .A1(n3448), .B0(n4314), .B1(n368), .Y(n5707)
         );
  AOI22X1TS U2854 ( .A0(n4151), .A1(n3447), .B0(n4308), .B1(n363), .Y(n5711)
         );
  AOI22X1TS U2855 ( .A0(n4148), .A1(n3447), .B0(n4305), .B1(n364), .Y(n5713)
         );
  AOI22X1TS U2856 ( .A0(n3959), .A1(n3472), .B0(n4428), .B1(n3697), .Y(n5509)
         );
  AOI222XLTS U2857 ( .A0(n4116), .A1(n3520), .B0(n192), .B1(n3508), .C0(n4272), 
        .C1(n3483), .Y(n5508) );
  AOI22X1TS U2858 ( .A0(n3953), .A1(n3472), .B0(n4422), .B1(n3697), .Y(n5513)
         );
  AOI222XLTS U2859 ( .A0(n4110), .A1(n3520), .B0(readRequesterAddress[3]), 
        .B1(n3510), .C0(n4266), .C1(n3497), .Y(n5512) );
  AOI22X1TS U2860 ( .A0(n3950), .A1(n3472), .B0(n4419), .B1(n3696), .Y(n5515)
         );
  AOI222XLTS U2861 ( .A0(n4107), .A1(n3520), .B0(readRequesterAddress[2]), 
        .B1(n3510), .C0(n4263), .C1(n3496), .Y(n5514) );
  AOI22X1TS U2862 ( .A0(n3947), .A1(n3476), .B0(n4416), .B1(n3685), .Y(n5517)
         );
  AOI222XLTS U2863 ( .A0(n4104), .A1(n3519), .B0(readRequesterAddress[1]), 
        .B1(n3498), .C0(n4260), .C1(n3492), .Y(n5516) );
  AOI22X1TS U2864 ( .A0(n3923), .A1(n3477), .B0(n4393), .B1(n3685), .Y(n5591)
         );
  AOI22X1TS U2865 ( .A0(n3920), .A1(n3480), .B0(n4390), .B1(n3685), .Y(n5593)
         );
  AOI22X1TS U2866 ( .A0(n3917), .A1(n3478), .B0(n4387), .B1(n3696), .Y(n5595)
         );
  AOI22X1TS U2867 ( .A0(n3914), .A1(n3478), .B0(n4384), .B1(n3694), .Y(n5597)
         );
  AOI22X1TS U2868 ( .A0(n3911), .A1(n6220), .B0(n4381), .B1(n3693), .Y(n5599)
         );
  AOI22X1TS U2869 ( .A0(n3908), .A1(n3475), .B0(n4378), .B1(n3695), .Y(n5601)
         );
  AOI22X1TS U2870 ( .A0(n3905), .A1(n3471), .B0(n4375), .B1(n3686), .Y(n5603)
         );
  AOI22X1TS U2871 ( .A0(n3902), .A1(n3471), .B0(n4372), .B1(n3686), .Y(n5605)
         );
  AOI22X1TS U2872 ( .A0(n3899), .A1(n3471), .B0(n4369), .B1(n3686), .Y(n5607)
         );
  AOI22X1TS U2873 ( .A0(n3896), .A1(n3471), .B0(n4366), .B1(n3686), .Y(n5609)
         );
  AOI22X1TS U2874 ( .A0(n3893), .A1(n3470), .B0(n4363), .B1(n3687), .Y(n5611)
         );
  AOI22X1TS U2875 ( .A0(n3890), .A1(n3470), .B0(n4360), .B1(n3687), .Y(n5613)
         );
  AOI22X1TS U2876 ( .A0(n3887), .A1(n3470), .B0(n4357), .B1(n3687), .Y(n5615)
         );
  AOI22X1TS U2877 ( .A0(n3884), .A1(n3469), .B0(n4354), .B1(n3687), .Y(n5617)
         );
  AOI22X1TS U2878 ( .A0(n3881), .A1(n3469), .B0(n4351), .B1(n3695), .Y(n5619)
         );
  AOI22X1TS U2879 ( .A0(n3878), .A1(n3469), .B0(n4348), .B1(n3694), .Y(n5621)
         );
  AOI22X1TS U2880 ( .A0(n3875), .A1(n3469), .B0(n4345), .B1(n3693), .Y(n5623)
         );
  AOI22X1TS U2881 ( .A0(n3872), .A1(n3468), .B0(n4342), .B1(n3695), .Y(n5625)
         );
  AOI22X1TS U2882 ( .A0(n3869), .A1(n3468), .B0(n4339), .B1(n3688), .Y(n5627)
         );
  AOI22X1TS U2883 ( .A0(n3866), .A1(n3468), .B0(n4336), .B1(n3688), .Y(n5629)
         );
  AOI22X1TS U2884 ( .A0(n3863), .A1(n3468), .B0(n4333), .B1(n3688), .Y(n5631)
         );
  AOI22X1TS U2885 ( .A0(n3860), .A1(n3467), .B0(n4330), .B1(n3688), .Y(n5633)
         );
  AOI22X1TS U2886 ( .A0(n3857), .A1(n3467), .B0(n4327), .B1(n3689), .Y(n5635)
         );
  AOI22X1TS U2887 ( .A0(n3854), .A1(n3467), .B0(n4324), .B1(n3689), .Y(n5637)
         );
  AOI22X1TS U2888 ( .A0(n3851), .A1(n3467), .B0(n4321), .B1(n3689), .Y(n5639)
         );
  AOI22X1TS U2889 ( .A0(n3848), .A1(n3466), .B0(n4318), .B1(n3689), .Y(n5641)
         );
  AOI22X1TS U2890 ( .A0(n3845), .A1(n3466), .B0(n4315), .B1(n3690), .Y(n5643)
         );
  AOI22X1TS U2891 ( .A0(n3842), .A1(n3466), .B0(n4312), .B1(n3690), .Y(n5645)
         );
  AOI22X1TS U2892 ( .A0(n3839), .A1(n3466), .B0(n4309), .B1(n3690), .Y(n5647)
         );
  AOI22X1TS U2893 ( .A0(n3836), .A1(n3465), .B0(n4306), .B1(n3690), .Y(n5649)
         );
  AOI22X1TS U2894 ( .A0(n3833), .A1(n3465), .B0(n4303), .B1(n3691), .Y(n5651)
         );
  AOI22X1TS U2895 ( .A0(n3830), .A1(n3465), .B0(n4300), .B1(n3691), .Y(n5653)
         );
  AOI22X1TS U2896 ( .A0(n4217), .A1(n3453), .B0(n4374), .B1(n269), .Y(n5667)
         );
  AOI22X1TS U2897 ( .A0(n4196), .A1(n3451), .B0(n4353), .B1(n367), .Y(n5681)
         );
  AOI22X1TS U2898 ( .A0(n4154), .A1(n3448), .B0(n4311), .B1(n267), .Y(n5709)
         );
  AOI22X1TS U2899 ( .A0(n4067), .A1(n780), .B0(n4380), .B1(n3775), .Y(n5983)
         );
  AOI22X1TS U2900 ( .A0(n4052), .A1(n776), .B0(n4365), .B1(n6308), .Y(n5993)
         );
  AOI22X1TS U2901 ( .A0(n4046), .A1(n775), .B0(n4359), .B1(n3777), .Y(n5997)
         );
  AOI22X1TS U2902 ( .A0(n4043), .A1(n775), .B0(n4356), .B1(n3778), .Y(n5999)
         );
  AOI22X1TS U2903 ( .A0(n4016), .A1(n772), .B0(n4329), .B1(n3771), .Y(n6017)
         );
  AOI22X1TS U2904 ( .A0(n4010), .A1(n772), .B0(n4323), .B1(n3770), .Y(n6021)
         );
  AOI22X1TS U2905 ( .A0(n4001), .A1(n771), .B0(n4314), .B1(n3769), .Y(n6027)
         );
  AOI22X1TS U2906 ( .A0(n3992), .A1(n771), .B0(n4305), .B1(n3769), .Y(n6033)
         );
  AOI22X1TS U2907 ( .A0(n4271), .A1(n3279), .B0(n4429), .B1(n3731), .Y(n5436)
         );
  AOI222XLTS U2908 ( .A0(n4115), .A1(n3323), .B0(n3306), .B1(n192), .C0(n3960), 
        .C1(n3297), .Y(n5435) );
  AOI22X1TS U2909 ( .A0(n4268), .A1(n3281), .B0(n4426), .B1(n3731), .Y(n5438)
         );
  AOI222XLTS U2910 ( .A0(n4112), .A1(n3323), .B0(n3308), .B1(n187), .C0(n3957), 
        .C1(n3300), .Y(n5437) );
  AOI22X1TS U2911 ( .A0(n4265), .A1(n3278), .B0(n4423), .B1(n3731), .Y(n5440)
         );
  AOI222XLTS U2912 ( .A0(n4109), .A1(n3323), .B0(n3308), .B1(n182), .C0(n3954), 
        .C1(n3294), .Y(n5439) );
  AOI22X1TS U2913 ( .A0(n4262), .A1(n3283), .B0(n4420), .B1(n3731), .Y(n5442)
         );
  AOI222XLTS U2914 ( .A0(n4106), .A1(n3323), .B0(n3308), .B1(n177), .C0(n3951), 
        .C1(n3295), .Y(n5441) );
  AOI22X1TS U2915 ( .A0(n4259), .A1(n3281), .B0(n4417), .B1(n3730), .Y(n5444)
         );
  AOI222XLTS U2916 ( .A0(n4103), .A1(n3322), .B0(n3308), .B1(n172), .C0(n3948), 
        .C1(n3296), .Y(n5443) );
  AOI22X1TS U2917 ( .A0(n4256), .A1(n3280), .B0(n4414), .B1(n3730), .Y(n5446)
         );
  AOI222XLTS U2918 ( .A0(n4100), .A1(n3322), .B0(n3307), .B1(n167), .C0(n3945), 
        .C1(n3293), .Y(n5445) );
  AOI22X1TS U2919 ( .A0(n4232), .A1(n3277), .B0(n4389), .B1(n3730), .Y(n5785)
         );
  AOI22X1TS U2920 ( .A0(n4226), .A1(n3277), .B0(n4383), .B1(n3735), .Y(n5789)
         );
  AOI22X1TS U2921 ( .A0(n4223), .A1(n3277), .B0(n4380), .B1(n3737), .Y(n5791)
         );
  AOI22X1TS U2922 ( .A0(n4220), .A1(n3277), .B0(n4377), .B1(n3733), .Y(n5793)
         );
  AOI22X1TS U2923 ( .A0(n4217), .A1(n3274), .B0(n4374), .B1(n3734), .Y(n5795)
         );
  AOI22X1TS U2924 ( .A0(n4214), .A1(n3274), .B0(n4371), .B1(n3736), .Y(n5797)
         );
  AOI22X1TS U2925 ( .A0(n4211), .A1(n3274), .B0(n4368), .B1(n3734), .Y(n5799)
         );
  AOI22X1TS U2926 ( .A0(n4196), .A1(n3272), .B0(n4353), .B1(n3735), .Y(n5809)
         );
  AOI22X1TS U2927 ( .A0(n4181), .A1(n3271), .B0(n4338), .B1(n3728), .Y(n5819)
         );
  AOI22X1TS U2928 ( .A0(n4169), .A1(n3273), .B0(n4326), .B1(n3727), .Y(n5827)
         );
  AOI22X1TS U2929 ( .A0(n4163), .A1(n3270), .B0(n4320), .B1(n3727), .Y(n5831)
         );
  AOI22X1TS U2930 ( .A0(n4157), .A1(n3269), .B0(n4314), .B1(n3726), .Y(n5835)
         );
  AOI22X1TS U2931 ( .A0(n4154), .A1(n3269), .B0(n4311), .B1(n3726), .Y(n5837)
         );
  AOI22X1TS U2932 ( .A0(n4148), .A1(n3269), .B0(n4305), .B1(n3726), .Y(n5841)
         );
  AOI22X1TS U2933 ( .A0(n3923), .A1(n3359), .B0(n4392), .B1(n254), .Y(n5719)
         );
  AOI222XLTS U2934 ( .A0(n4079), .A1(n3392), .B0(cacheDataOut[31]), .B1(n3367), 
        .C0(n4236), .C1(n211), .Y(n5718) );
  AOI22X1TS U2935 ( .A0(n3878), .A1(n3355), .B0(n4347), .B1(n432), .Y(n5749)
         );
  AOI222XLTS U2936 ( .A0(n4034), .A1(n3386), .B0(cacheDataOut[16]), .B1(n3379), 
        .C0(n4191), .C1(n210), .Y(n5748) );
  AOI22X1TS U2937 ( .A0(n3875), .A1(n3355), .B0(n4344), .B1(n428), .Y(n5751)
         );
  AOI222XLTS U2938 ( .A0(n4031), .A1(n3386), .B0(cacheDataOut[15]), .B1(n3369), 
        .C0(n4188), .C1(n198), .Y(n5750) );
  AOI22X1TS U2939 ( .A0(n3863), .A1(n3354), .B0(n4332), .B1(n428), .Y(n5759)
         );
  AOI222XLTS U2940 ( .A0(n4019), .A1(n3385), .B0(cacheDataOut[11]), .B1(n3371), 
        .C0(n4176), .C1(n210), .Y(n5758) );
  AOI22X1TS U2941 ( .A0(n3833), .A1(n3351), .B0(n4302), .B1(n3717), .Y(n5779)
         );
  AOI222XLTS U2942 ( .A0(n3989), .A1(n3382), .B0(cacheDataOut[1]), .B1(n3372), 
        .C0(n4146), .C1(n203), .Y(n5778) );
  AOI22X1TS U2943 ( .A0(n4265), .A1(n3457), .B0(n4422), .B1(n368), .Y(n5487)
         );
  AOI222XLTS U2944 ( .A0(n3953), .A1(n3707), .B0(n3441), .B1(n183), .C0(n4110), 
        .C1(n3425), .Y(n5486) );
  AOI22X1TS U2945 ( .A0(n4262), .A1(n3459), .B0(n4419), .B1(n250), .Y(n5489)
         );
  AOI222XLTS U2946 ( .A0(n3950), .A1(n3707), .B0(n3441), .B1(n178), .C0(n4107), 
        .C1(n3425), .Y(n5488) );
  AOI22X1TS U2947 ( .A0(n4259), .A1(n3458), .B0(n4416), .B1(n369), .Y(n5491)
         );
  AOI222XLTS U2948 ( .A0(n3947), .A1(n3707), .B0(n3440), .B1(n173), .C0(n4104), 
        .C1(n3425), .Y(n5490) );
  AOI22X1TS U2949 ( .A0(n4256), .A1(n3459), .B0(n4413), .B1(n269), .Y(n5493)
         );
  AOI222XLTS U2950 ( .A0(n3944), .A1(n3707), .B0(n3440), .B1(n168), .C0(n4101), 
        .C1(n3425), .Y(n5492) );
  AOI22X1TS U2951 ( .A0(n4115), .A1(n782), .B0(n4428), .B1(n3774), .Y(n5367)
         );
  AOI222XLTS U2952 ( .A0(n3960), .A1(n832), .B0(n812), .B1(n191), .C0(n4272), 
        .C1(n800), .Y(n5366) );
  AOI22X1TS U2953 ( .A0(n4112), .A1(n784), .B0(n4425), .B1(n3774), .Y(n5369)
         );
  AOI222XLTS U2954 ( .A0(n3957), .A1(n832), .B0(n6129), .B1(n188), .C0(n4269), 
        .C1(n803), .Y(n5368) );
  AOI22X1TS U2955 ( .A0(n4109), .A1(n781), .B0(n4422), .B1(n3774), .Y(n5371)
         );
  AOI222XLTS U2956 ( .A0(n3954), .A1(n830), .B0(n816), .B1(n180), .C0(n4266), 
        .C1(n799), .Y(n5370) );
  AOI22X1TS U2957 ( .A0(n4106), .A1(n786), .B0(n4419), .B1(n3774), .Y(n5373)
         );
  AOI222XLTS U2958 ( .A0(n3951), .A1(n831), .B0(n813), .B1(n175), .C0(n4263), 
        .C1(n799), .Y(n5372) );
  AOI22X1TS U2959 ( .A0(n4103), .A1(n784), .B0(n4416), .B1(n3773), .Y(n5375)
         );
  AOI222XLTS U2960 ( .A0(n3948), .A1(n833), .B0(n814), .B1(n170), .C0(n4260), 
        .C1(n796), .Y(n5374) );
  AOI22X1TS U2961 ( .A0(n4100), .A1(n783), .B0(n4413), .B1(n3773), .Y(n5377)
         );
  AOI222XLTS U2962 ( .A0(n3945), .A1(n831), .B0(n817), .B1(n165), .C0(n4257), 
        .C1(n797), .Y(n5376) );
  AOI22X1TS U2963 ( .A0(n4079), .A1(n780), .B0(n4392), .B1(n3773), .Y(n5975)
         );
  AOI22X1TS U2964 ( .A0(n4076), .A1(n783), .B0(n4389), .B1(n3773), .Y(n5977)
         );
  AOI22X1TS U2965 ( .A0(n4073), .A1(n780), .B0(n4386), .B1(n3780), .Y(n5979)
         );
  AOI22X1TS U2966 ( .A0(n4070), .A1(n780), .B0(n4383), .B1(n3777), .Y(n5981)
         );
  AOI22X1TS U2967 ( .A0(n4064), .A1(n782), .B0(n4377), .B1(n3779), .Y(n5985)
         );
  AOI22X1TS U2968 ( .A0(n4061), .A1(n776), .B0(n4374), .B1(n6308), .Y(n5987)
         );
  AOI22X1TS U2969 ( .A0(n4058), .A1(n776), .B0(n4371), .B1(n3776), .Y(n5989)
         );
  AOI22X1TS U2970 ( .A0(n4055), .A1(n776), .B0(n4368), .B1(n3775), .Y(n5991)
         );
  AOI22X1TS U2971 ( .A0(n4049), .A1(n775), .B0(n4362), .B1(n3780), .Y(n5995)
         );
  AOI22X1TS U2972 ( .A0(n4040), .A1(n774), .B0(n4353), .B1(n3776), .Y(n6001)
         );
  AOI22X1TS U2973 ( .A0(n4037), .A1(n774), .B0(n4350), .B1(n3772), .Y(n6003)
         );
  AOI22X1TS U2974 ( .A0(n4034), .A1(n774), .B0(n4347), .B1(n3772), .Y(n6005)
         );
  AOI22X1TS U2975 ( .A0(n4031), .A1(n774), .B0(n4344), .B1(n3772), .Y(n6007)
         );
  AOI22X1TS U2976 ( .A0(n4028), .A1(n773), .B0(n4341), .B1(n3772), .Y(n6009)
         );
  AOI22X1TS U2977 ( .A0(n4025), .A1(n773), .B0(n4338), .B1(n3771), .Y(n6011)
         );
  AOI22X1TS U2978 ( .A0(n4022), .A1(n773), .B0(n4335), .B1(n3771), .Y(n6013)
         );
  AOI22X1TS U2979 ( .A0(n4019), .A1(n773), .B0(n4332), .B1(n3771), .Y(n6015)
         );
  AOI22X1TS U2980 ( .A0(n4013), .A1(n775), .B0(n4326), .B1(n3770), .Y(n6019)
         );
  AOI22X1TS U2981 ( .A0(n4007), .A1(n772), .B0(n4320), .B1(n3770), .Y(n6023)
         );
  AOI22X1TS U2982 ( .A0(n4004), .A1(n772), .B0(n4317), .B1(n3770), .Y(n6025)
         );
  AOI22X1TS U2983 ( .A0(n3998), .A1(n771), .B0(n4311), .B1(n3769), .Y(n6029)
         );
  AOI22X1TS U2984 ( .A0(n3995), .A1(n771), .B0(n4308), .B1(n3769), .Y(n6031)
         );
  AOI22X1TS U2985 ( .A0(n3989), .A1(n770), .B0(n4302), .B1(n3768), .Y(n6035)
         );
  AOI22X1TS U2986 ( .A0(n4235), .A1(n3280), .B0(n4392), .B1(n3730), .Y(n5783)
         );
  AOI22X1TS U2987 ( .A0(n4229), .A1(n3279), .B0(n4386), .B1(n3732), .Y(n5787)
         );
  AOI22X1TS U2988 ( .A0(n4208), .A1(n3274), .B0(n4365), .B1(n3732), .Y(n5801)
         );
  AOI22X1TS U2989 ( .A0(n4205), .A1(n3273), .B0(n4362), .B1(n3737), .Y(n5803)
         );
  AOI22X1TS U2990 ( .A0(n4202), .A1(n3273), .B0(n4359), .B1(n3735), .Y(n5805)
         );
  AOI22X1TS U2991 ( .A0(n4199), .A1(n3273), .B0(n4356), .B1(n3733), .Y(n5807)
         );
  AOI22X1TS U2992 ( .A0(n4190), .A1(n3272), .B0(n4347), .B1(n3729), .Y(n5813)
         );
  AOI22X1TS U2993 ( .A0(n4178), .A1(n3271), .B0(n4335), .B1(n3728), .Y(n5821)
         );
  AOI22X1TS U2994 ( .A0(n4175), .A1(n3271), .B0(n4332), .B1(n3728), .Y(n5823)
         );
  AOI22X1TS U2995 ( .A0(n4172), .A1(n3270), .B0(n4329), .B1(n3728), .Y(n5825)
         );
  AOI22X1TS U2996 ( .A0(n4166), .A1(n3270), .B0(n4323), .B1(n3727), .Y(n5829)
         );
  AOI22X1TS U2997 ( .A0(n4160), .A1(n3270), .B0(n4317), .B1(n3727), .Y(n5833)
         );
  AOI22X1TS U2998 ( .A0(n4145), .A1(n3268), .B0(n4302), .B1(n3725), .Y(n5843)
         );
  AOI22X1TS U2999 ( .A0(n4142), .A1(n3268), .B0(n4299), .B1(n3725), .Y(n5845)
         );
  AOI22X1TS U3000 ( .A0(n3959), .A1(n3359), .B0(n4428), .B1(n3718), .Y(n5460)
         );
  AOI22X1TS U3001 ( .A0(n3956), .A1(n3366), .B0(n4425), .B1(n3721), .Y(n5462)
         );
  AOI222XLTS U3002 ( .A0(n4112), .A1(n3394), .B0(n3375), .B1(n185), .C0(n4269), 
        .C1(n210), .Y(n5461) );
  AOI22X1TS U3003 ( .A0(n3953), .A1(n3366), .B0(n4422), .B1(n5), .Y(n5464) );
  AOI222XLTS U3004 ( .A0(n4109), .A1(n3396), .B0(n3375), .B1(n181), .C0(n4266), 
        .C1(n198), .Y(n5463) );
  AOI22X1TS U3005 ( .A0(n3950), .A1(n6188), .B0(n4419), .B1(n3719), .Y(n5466)
         );
  AOI222XLTS U3006 ( .A0(n4106), .A1(n3395), .B0(n3375), .B1(n176), .C0(n4263), 
        .C1(n200), .Y(n5465) );
  AOI22X1TS U3007 ( .A0(n3947), .A1(n3363), .B0(n4416), .B1(n3720), .Y(n5468)
         );
  AOI222XLTS U3008 ( .A0(n4103), .A1(n3391), .B0(n3375), .B1(n171), .C0(n4260), 
        .C1(n203), .Y(n5467) );
  AOI22X1TS U3009 ( .A0(n3944), .A1(n3359), .B0(n4413), .B1(n3723), .Y(n5470)
         );
  AOI222XLTS U3010 ( .A0(n4100), .A1(n3392), .B0(n3374), .B1(n166), .C0(n4257), 
        .C1(n212), .Y(n5469) );
  AOI22X1TS U3011 ( .A0(n3920), .A1(n3362), .B0(n4389), .B1(n3716), .Y(n5721)
         );
  AOI222XLTS U3012 ( .A0(n4076), .A1(n6191), .B0(cacheDataOut[30]), .B1(n3379), 
        .C0(n4233), .C1(n203), .Y(n5720) );
  AOI22X1TS U3013 ( .A0(n3917), .A1(n3361), .B0(n4386), .B1(n432), .Y(n5723)
         );
  AOI222XLTS U3014 ( .A0(n4073), .A1(n3389), .B0(cacheDataOut[29]), .B1(n3367), 
        .C0(n4230), .C1(n207), .Y(n5722) );
  AOI22X1TS U3015 ( .A0(n3914), .A1(n3361), .B0(n4383), .B1(n254), .Y(n5725)
         );
  AOI222XLTS U3016 ( .A0(n4070), .A1(n3389), .B0(cacheDataOut[28]), .B1(n3378), 
        .C0(n4227), .C1(n208), .Y(n5724) );
  AOI22X1TS U3017 ( .A0(n3911), .A1(n3362), .B0(n4380), .B1(n3719), .Y(n5727)
         );
  AOI222XLTS U3018 ( .A0(n4067), .A1(n3389), .B0(cacheDataOut[27]), .B1(n3379), 
        .C0(n4224), .C1(n207), .Y(n5726) );
  AOI22X1TS U3019 ( .A0(n3908), .A1(n3363), .B0(n4377), .B1(n430), .Y(n5729)
         );
  AOI222XLTS U3020 ( .A0(n4064), .A1(n3389), .B0(cacheDataOut[26]), .B1(n3368), 
        .C0(n4221), .C1(n206), .Y(n5728) );
  AOI22X1TS U3021 ( .A0(n3905), .A1(n3360), .B0(n4374), .B1(n3718), .Y(n5731)
         );
  AOI222XLTS U3022 ( .A0(n4061), .A1(n3388), .B0(cacheDataOut[25]), .B1(n3368), 
        .C0(n4218), .C1(n436), .Y(n5730) );
  AOI22X1TS U3023 ( .A0(n3902), .A1(n3364), .B0(n4371), .B1(n432), .Y(n5733)
         );
  AOI222XLTS U3024 ( .A0(n4058), .A1(n3388), .B0(cacheDataOut[24]), .B1(n3367), 
        .C0(n4215), .C1(n436), .Y(n5732) );
  AOI22X1TS U3025 ( .A0(n3899), .A1(n3360), .B0(n4368), .B1(n432), .Y(n5735)
         );
  AOI222XLTS U3026 ( .A0(n4055), .A1(n3388), .B0(cacheDataOut[23]), .B1(n3369), 
        .C0(n4212), .C1(n212), .Y(n5734) );
  AOI22X1TS U3027 ( .A0(n3896), .A1(n3360), .B0(n4365), .B1(n254), .Y(n5737)
         );
  AOI222XLTS U3028 ( .A0(n4052), .A1(n3388), .B0(cacheDataOut[22]), .B1(n3369), 
        .C0(n4209), .C1(n436), .Y(n5736) );
  AOI22X1TS U3029 ( .A0(n3893), .A1(n3356), .B0(n4362), .B1(n3723), .Y(n5739)
         );
  AOI222XLTS U3030 ( .A0(n4049), .A1(n3387), .B0(cacheDataOut[21]), .B1(n3367), 
        .C0(n4206), .C1(n203), .Y(n5738) );
  AOI22X1TS U3031 ( .A0(n3890), .A1(n3356), .B0(n4359), .B1(n3721), .Y(n5741)
         );
  AOI222XLTS U3032 ( .A0(n4046), .A1(n3387), .B0(cacheDataOut[20]), .B1(n3369), 
        .C0(n4203), .C1(n208), .Y(n5740) );
  AOI22X1TS U3033 ( .A0(n3887), .A1(n3356), .B0(n4356), .B1(n3719), .Y(n5743)
         );
  AOI222XLTS U3034 ( .A0(n4043), .A1(n3387), .B0(cacheDataOut[19]), .B1(n3370), 
        .C0(n4200), .C1(n211), .Y(n5742) );
  AOI22X1TS U3035 ( .A0(n3884), .A1(n3355), .B0(n4353), .B1(n3717), .Y(n5745)
         );
  AOI222XLTS U3036 ( .A0(n4040), .A1(n3386), .B0(cacheDataOut[18]), .B1(n3368), 
        .C0(n4197), .C1(n208), .Y(n5744) );
  AOI22X1TS U3037 ( .A0(n3881), .A1(n3355), .B0(n4350), .B1(n254), .Y(n5747)
         );
  AOI222XLTS U3038 ( .A0(n4037), .A1(n3386), .B0(cacheDataOut[17]), .B1(n3370), 
        .C0(n4194), .C1(n209), .Y(n5746) );
  AOI22X1TS U3039 ( .A0(n3872), .A1(n3354), .B0(n4341), .B1(n426), .Y(n5753)
         );
  AOI222XLTS U3040 ( .A0(n4028), .A1(n3385), .B0(cacheDataOut[14]), .B1(n3368), 
        .C0(n4185), .C1(n198), .Y(n5752) );
  AOI22X1TS U3041 ( .A0(n3869), .A1(n3354), .B0(n4338), .B1(n426), .Y(n5755)
         );
  AOI222XLTS U3042 ( .A0(n4025), .A1(n3385), .B0(cacheDataOut[13]), .B1(n3378), 
        .C0(n4182), .C1(n213), .Y(n5754) );
  AOI22X1TS U3043 ( .A0(n3866), .A1(n3354), .B0(n4335), .B1(n430), .Y(n5757)
         );
  AOI222XLTS U3044 ( .A0(n4022), .A1(n3385), .B0(cacheDataOut[12]), .B1(n3370), 
        .C0(n4179), .C1(n211), .Y(n5756) );
  AOI22X1TS U3045 ( .A0(n3860), .A1(n3353), .B0(n4329), .B1(n3723), .Y(n5761)
         );
  AOI222XLTS U3046 ( .A0(n4016), .A1(n3384), .B0(cacheDataOut[10]), .B1(n3371), 
        .C0(n4173), .C1(n209), .Y(n5760) );
  AOI22X1TS U3047 ( .A0(n3857), .A1(n3356), .B0(n4326), .B1(n430), .Y(n5763)
         );
  AOI222XLTS U3048 ( .A0(n4013), .A1(n3387), .B0(cacheDataOut[9]), .B1(n3376), 
        .C0(n4170), .C1(n210), .Y(n5762) );
  AOI22X1TS U3049 ( .A0(n3854), .A1(n3353), .B0(n4323), .B1(n430), .Y(n5765)
         );
  AOI222XLTS U3050 ( .A0(n4010), .A1(n3384), .B0(cacheDataOut[8]), .B1(n3371), 
        .C0(n4167), .C1(n213), .Y(n5764) );
  AOI22X1TS U3051 ( .A0(n3851), .A1(n3353), .B0(n4320), .B1(n426), .Y(n5767)
         );
  AOI222XLTS U3052 ( .A0(n4007), .A1(n3384), .B0(cacheDataOut[7]), .B1(n3376), 
        .C0(n4164), .C1(n208), .Y(n5766) );
  AOI22X1TS U3053 ( .A0(n3848), .A1(n3353), .B0(n4317), .B1(n3722), .Y(n5769)
         );
  AOI222XLTS U3054 ( .A0(n4004), .A1(n3384), .B0(cacheDataOut[6]), .B1(n3380), 
        .C0(n4161), .C1(n201), .Y(n5768) );
  AOI22X1TS U3055 ( .A0(n3845), .A1(n3352), .B0(n4314), .B1(n3717), .Y(n5771)
         );
  AOI222XLTS U3056 ( .A0(n4001), .A1(n3383), .B0(cacheDataOut[5]), .B1(n3372), 
        .C0(n4158), .C1(n212), .Y(n5770) );
  AOI22X1TS U3057 ( .A0(n3842), .A1(n3352), .B0(n4311), .B1(n3721), .Y(n5773)
         );
  AOI222XLTS U3058 ( .A0(n3998), .A1(n3383), .B0(cacheDataOut[4]), .B1(n3372), 
        .C0(n4155), .C1(n209), .Y(n5772) );
  AOI22X1TS U3059 ( .A0(n3839), .A1(n3352), .B0(n4308), .B1(n428), .Y(n5775)
         );
  AOI222XLTS U3060 ( .A0(n3995), .A1(n3383), .B0(cacheDataOut[3]), .B1(n3371), 
        .C0(n4152), .C1(n204), .Y(n5774) );
  AOI22X1TS U3061 ( .A0(n3836), .A1(n3352), .B0(n4305), .B1(n3718), .Y(n5777)
         );
  AOI222XLTS U3062 ( .A0(n3992), .A1(n3383), .B0(cacheDataOut[2]), .B1(n3372), 
        .C0(n4149), .C1(n206), .Y(n5776) );
  AOI22X1TS U3063 ( .A0(n3830), .A1(n3351), .B0(n4299), .B1(n3720), .Y(n5781)
         );
  AOI222XLTS U3064 ( .A0(n3986), .A1(n3382), .B0(cacheDataOut[0]), .B1(n3370), 
        .C0(n4143), .C1(n207), .Y(n5780) );
  AOI22X1TS U3065 ( .A0(n3986), .A1(n770), .B0(n4299), .B1(n3768), .Y(n6037)
         );
  AOI22X1TS U3066 ( .A0(n4193), .A1(n3272), .B0(n4350), .B1(n3729), .Y(n5811)
         );
  AOI22X1TS U3067 ( .A0(n4187), .A1(n3272), .B0(n4344), .B1(n3729), .Y(n5815)
         );
  AOI22X1TS U3068 ( .A0(n4184), .A1(n3271), .B0(n4341), .B1(n3729), .Y(n5817)
         );
  AOI22X1TS U3069 ( .A0(n4151), .A1(n3269), .B0(n4308), .B1(n3726), .Y(n5839)
         );
  AOI22X1TS U3070 ( .A0(n4268), .A1(n3460), .B0(n4425), .B1(n270), .Y(n5485)
         );
  AOI222XLTS U3071 ( .A0(n3956), .A1(n3708), .B0(n3441), .B1(n185), .C0(n4113), 
        .C1(n3432), .Y(n5484) );
  AOI22X1TS U3072 ( .A0(n1571), .A1(n173), .B0(n854), .B1(n4085), .Y(n6142) );
  AOI222XLTS U3073 ( .A0(\requesterAddressbuffer[2][1] ), .A1(n379), .B0(n3192), .B1(n4242), .C0(n3753), .C1(n4399), .Y(n6141) );
  AOI22X1TS U3074 ( .A0(n871), .A1(n168), .B0(n855), .B1(n4082), .Y(n6147) );
  AOI222XLTS U3075 ( .A0(\requesterAddressbuffer[2][0] ), .A1(n340), .B0(n3200), .B1(n4239), .C0(n3753), .C1(n4396), .Y(n6146) );
  AOI22X1TS U3076 ( .A0(n6144), .A1(n183), .B0(n854), .B1(n4091), .Y(n6138) );
  AOI222XLTS U3077 ( .A0(\requesterAddressbuffer[2][3] ), .A1(n341), .B0(n3200), .B1(n4248), .C0(n3753), .C1(n4405), .Y(n6137) );
  AOI22X1TS U3078 ( .A0(n1535), .A1(n177), .B0(n854), .B1(n4088), .Y(n6140) );
  AOI222XLTS U3079 ( .A0(\requesterAddressbuffer[2][2] ), .A1(n259), .B0(n3200), .B1(n4245), .C0(n3753), .C1(n4402), .Y(n6139) );
  AOI22X1TS U3080 ( .A0(n871), .A1(n187), .B0(n854), .B1(n4094), .Y(n6136) );
  AOI222XLTS U3081 ( .A0(\requesterAddressbuffer[2][4] ), .A1(n378), .B0(n3192), .B1(n4251), .C0(n6307), .C1(n4408), .Y(n6135) );
  AOI22X1TS U3082 ( .A0(n871), .A1(readRequesterAddress[5]), .B0(n855), .B1(
        n4097), .Y(n6134) );
  AOI222XLTS U3083 ( .A0(\requesterAddressbuffer[2][5] ), .A1(n381), .B0(n3193), .B1(n4254), .C0(n3765), .C1(n4411), .Y(n6133) );
  AOI22X1TS U3084 ( .A0(n3433), .A1(n181), .B0(n3416), .B1(n4091), .Y(n6199)
         );
  AOI222XLTS U3085 ( .A0(\requesterAddressbuffer[6][3] ), .A1(n700), .B0(n3456), .B1(n4247), .C0(n3715), .C1(n4405), .Y(n6198) );
  AOI22X1TS U3086 ( .A0(n3433), .A1(n171), .B0(n3416), .B1(n4085), .Y(n6203)
         );
  AOI222XLTS U3087 ( .A0(\requesterAddressbuffer[6][1] ), .A1(n700), .B0(n3456), .B1(n4241), .C0(n3715), .C1(n4399), .Y(n6202) );
  AOI222XLTS U3088 ( .A0(\requesterAddressbuffer[6][0] ), .A1(n700), .B0(n3460), .B1(n4238), .C0(n3715), .C1(n4396), .Y(n6207) );
  AOI22X1TS U3089 ( .A0(n749), .A1(readRequesterAddress[5]), .B0(n705), .B1(
        n4253), .Y(n6103) );
  AOI222XLTS U3090 ( .A0(\requesterAddressbuffer[0][5] ), .A1(n383), .B0(n766), 
        .B1(n3942), .C0(n3806), .C1(n4411), .Y(n6102) );
  AOI22X1TS U3091 ( .A0(n748), .A1(n182), .B0(n704), .B1(n4247), .Y(n6107) );
  AOI222XLTS U3092 ( .A0(\requesterAddressbuffer[0][3] ), .A1(n384), .B0(n768), 
        .B1(n3936), .C0(n3797), .C1(n4405), .Y(n6106) );
  AOI22X1TS U3093 ( .A0(n745), .A1(n186), .B0(n704), .B1(n4250), .Y(n6105) );
  AOI222XLTS U3094 ( .A0(\requesterAddressbuffer[0][4] ), .A1(n346), .B0(n762), 
        .B1(n3939), .C0(n3804), .C1(n4408), .Y(n6104) );
  AOI22X1TS U3095 ( .A0(n750), .A1(n176), .B0(n704), .B1(n4244), .Y(n6109) );
  AOI222XLTS U3096 ( .A0(\requesterAddressbuffer[0][2] ), .A1(n345), .B0(n768), 
        .B1(n3933), .C0(n3797), .C1(n4402), .Y(n6108) );
  AOI22X1TS U3097 ( .A0(n6113), .A1(n172), .B0(n704), .B1(n4241), .Y(n6111) );
  AOI222XLTS U3098 ( .A0(\requesterAddressbuffer[0][1] ), .A1(n3782), .B0(n768), .B1(n3930), .C0(n3797), .C1(n4399), .Y(n6110) );
  AOI22X1TS U3099 ( .A0(n750), .A1(n165), .B0(n705), .B1(n4238), .Y(n6116) );
  AOI222XLTS U3100 ( .A0(\requesterAddressbuffer[0][0] ), .A1(n343), .B0(n763), 
        .B1(n3927), .C0(n3797), .C1(n4396), .Y(n6115) );
  AOI22X1TS U3101 ( .A0(n749), .A1(n190), .B0(n4271), .B1(n714), .Y(n5343) );
  AOI222XLTS U3102 ( .A0(n385), .A1(n34), .B0(n3960), .B1(n754), .C0(n4429), 
        .C1(n3803), .Y(n5342) );
  AOI22X1TS U3103 ( .A0(n737), .A1(n180), .B0(n4265), .B1(n714), .Y(n5347) );
  AOI222XLTS U3104 ( .A0(n3782), .A1(n35), .B0(n3954), .B1(n768), .C0(n4423), 
        .C1(n3803), .Y(n5346) );
  AOI22X1TS U3105 ( .A0(n737), .A1(n178), .B0(n4262), .B1(n714), .Y(n5349) );
  AOI222XLTS U3106 ( .A0(n299), .A1(n36), .B0(n3951), .B1(n762), .C0(n4420), 
        .C1(n3803), .Y(n5348) );
  AOI22X1TS U3107 ( .A0(n745), .A1(n173), .B0(n4259), .B1(n728), .Y(n5351) );
  AOI222XLTS U3108 ( .A0(n299), .A1(n37), .B0(n3948), .B1(n765), .C0(n4417), 
        .C1(n3802), .Y(n5350) );
  AOI22X1TS U3109 ( .A0(n451), .A1(n743), .B0(n4235), .B1(n728), .Y(n6039) );
  AOI222XLTS U3110 ( .A0(n346), .A1(n38), .B0(n3924), .B1(n765), .C0(n4393), 
        .C1(n3802), .Y(n6038) );
  AOI22X1TS U3111 ( .A0(n453), .A1(n748), .B0(n4232), .B1(n732), .Y(n6041) );
  AOI222XLTS U3112 ( .A0(n344), .A1(n39), .B0(n3921), .B1(n764), .C0(n4390), 
        .C1(n3802), .Y(n6040) );
  AOI22X1TS U3113 ( .A0(n455), .A1(n748), .B0(n4229), .B1(n733), .Y(n6043) );
  AOI222XLTS U3114 ( .A0(n3782), .A1(n40), .B0(n3918), .B1(n761), .C0(n4387), 
        .C1(n3801), .Y(n6042) );
  AOI22X1TS U3115 ( .A0(n461), .A1(n740), .B0(n4220), .B1(n734), .Y(n6049) );
  AOI222XLTS U3116 ( .A0(n347), .A1(n41), .B0(n3909), .B1(n761), .C0(n4378), 
        .C1(n3801), .Y(n6048) );
  AOI22X1TS U3117 ( .A0(n463), .A1(n747), .B0(n4217), .B1(n729), .Y(n6051) );
  AOI222XLTS U3118 ( .A0(n344), .A1(n42), .B0(n3906), .B1(n760), .C0(n4375), 
        .C1(n3800), .Y(n6050) );
  AOI22X1TS U3119 ( .A0(n465), .A1(n751), .B0(n4214), .B1(n729), .Y(n6053) );
  AOI222XLTS U3120 ( .A0(n3781), .A1(n43), .B0(n3903), .B1(n760), .C0(n4372), 
        .C1(n3800), .Y(n6052) );
  AOI22X1TS U3121 ( .A0(n469), .A1(n6113), .B0(n4208), .B1(n728), .Y(n6057) );
  AOI222XLTS U3122 ( .A0(n345), .A1(n44), .B0(n3897), .B1(n760), .C0(n4366), 
        .C1(n3800), .Y(n6056) );
  AOI22X1TS U3123 ( .A0(n471), .A1(n738), .B0(n4205), .B1(n712), .Y(n6059) );
  AOI222XLTS U3124 ( .A0(n343), .A1(n45), .B0(n3894), .B1(n759), .C0(n4363), 
        .C1(n3799), .Y(n6058) );
  AOI22X1TS U3125 ( .A0(n475), .A1(n738), .B0(n4199), .B1(n712), .Y(n6063) );
  AOI222XLTS U3126 ( .A0(n383), .A1(n46), .B0(n3888), .B1(n759), .C0(n4357), 
        .C1(n3799), .Y(n6062) );
  AOI22X1TS U3127 ( .A0(n477), .A1(n739), .B0(n4196), .B1(n711), .Y(n6065) );
  AOI222XLTS U3128 ( .A0(n385), .A1(n47), .B0(n3885), .B1(n758), .C0(n4354), 
        .C1(n3799), .Y(n6064) );
  AOI22X1TS U3129 ( .A0(n479), .A1(n738), .B0(n4193), .B1(n711), .Y(n6067) );
  AOI222XLTS U3130 ( .A0(n345), .A1(n48), .B0(n3882), .B1(n758), .C0(n4351), 
        .C1(n3798), .Y(n6066) );
  AOI22X1TS U3131 ( .A0(n481), .A1(n739), .B0(n4190), .B1(n711), .Y(n6069) );
  AOI222XLTS U3132 ( .A0(n384), .A1(n49), .B0(n3879), .B1(n758), .C0(n4348), 
        .C1(n3798), .Y(n6068) );
  AOI22X1TS U3133 ( .A0(n483), .A1(n740), .B0(n4187), .B1(n711), .Y(n6071) );
  AOI222XLTS U3134 ( .A0(n383), .A1(n50), .B0(n3876), .B1(n758), .C0(n4345), 
        .C1(n3798), .Y(n6070) );
  AOI22X1TS U3135 ( .A0(n485), .A1(n739), .B0(n4184), .B1(n708), .Y(n6073) );
  AOI222XLTS U3136 ( .A0(n346), .A1(n51), .B0(n3873), .B1(n757), .C0(n4342), 
        .C1(n3798), .Y(n6072) );
  AOI22X1TS U3137 ( .A0(n487), .A1(n739), .B0(n4181), .B1(n708), .Y(n6075) );
  AOI222XLTS U3138 ( .A0(n347), .A1(n52), .B0(n3870), .B1(n757), .C0(n4339), 
        .C1(n3807), .Y(n6074) );
  AOI22X1TS U3139 ( .A0(n489), .A1(n740), .B0(n4178), .B1(n708), .Y(n6077) );
  AOI222XLTS U3140 ( .A0(n384), .A1(n53), .B0(n3867), .B1(n757), .C0(n4336), 
        .C1(n3809), .Y(n6076) );
  AOI22X1TS U3141 ( .A0(n491), .A1(n740), .B0(n4175), .B1(n708), .Y(n6079) );
  AOI222XLTS U3142 ( .A0(n347), .A1(n54), .B0(n3864), .B1(n757), .C0(n4333), 
        .C1(n3809), .Y(n6078) );
  AOI22X1TS U3143 ( .A0(n493), .A1(n743), .B0(n4172), .B1(n707), .Y(n6081) );
  AOI222XLTS U3144 ( .A0(n344), .A1(n55), .B0(n3861), .B1(n756), .C0(n4330), 
        .C1(n3810), .Y(n6080) );
  AOI22X1TS U3145 ( .A0(n501), .A1(n741), .B0(n4166), .B1(n707), .Y(n6085) );
  AOI222XLTS U3146 ( .A0(n345), .A1(n56), .B0(n3855), .B1(n756), .C0(n4324), 
        .C1(n3808), .Y(n6084) );
  AOI22X1TS U3147 ( .A0(n505), .A1(n741), .B0(n4163), .B1(n707), .Y(n6087) );
  AOI222XLTS U3148 ( .A0(n3781), .A1(n57), .B0(n3852), .B1(n756), .C0(n4321), 
        .C1(n3808), .Y(n6086) );
  AOI22X1TS U3149 ( .A0(n508), .A1(n742), .B0(n4160), .B1(n707), .Y(n6089) );
  AOI222XLTS U3150 ( .A0(n343), .A1(n58), .B0(n3849), .B1(n759), .C0(n4318), 
        .C1(n3808), .Y(n6088) );
  AOI22X1TS U3151 ( .A0(n512), .A1(n742), .B0(n4154), .B1(n706), .Y(n6093) );
  AOI222XLTS U3152 ( .A0(n343), .A1(n59), .B0(n3843), .B1(n755), .C0(n4312), 
        .C1(n3805), .Y(n6092) );
  AOI22X1TS U3153 ( .A0(n515), .A1(n743), .B0(n4151), .B1(n706), .Y(n6095) );
  AOI222XLTS U3154 ( .A0(n3782), .A1(n60), .B0(n3840), .B1(n755), .C0(n4309), 
        .C1(n3806), .Y(n6094) );
  AOI22X1TS U3155 ( .A0(n3218), .A1(n190), .B0(n4271), .B1(n275), .Y(n5414) );
  AOI222XLTS U3156 ( .A0(n3249), .A1(n61), .B0(n3960), .B1(n248), .C0(n4429), 
        .C1(n3242), .Y(n5413) );
  AOI22X1TS U3157 ( .A0(n3218), .A1(n188), .B0(n4268), .B1(n373), .Y(n5416) );
  AOI222XLTS U3158 ( .A0(n3249), .A1(n62), .B0(n3957), .B1(n357), .C0(n4426), 
        .C1(n3242), .Y(n5415) );
  AOI22X1TS U3159 ( .A0(n3218), .A1(n183), .B0(n4265), .B1(n376), .Y(n5418) );
  AOI222XLTS U3160 ( .A0(n3249), .A1(n63), .B0(n3954), .B1(n359), .C0(n4423), 
        .C1(n3242), .Y(n5417) );
  AOI22X1TS U3161 ( .A0(n3219), .A1(n171), .B0(n4259), .B1(n275), .Y(n5422) );
  AOI222XLTS U3162 ( .A0(n3250), .A1(n64), .B0(n3948), .B1(n359), .C0(n4417), 
        .C1(n3241), .Y(n5421) );
  AOI22X1TS U3163 ( .A0(n3219), .A1(n167), .B0(n4256), .B1(n275), .Y(n5424) );
  AOI222XLTS U3164 ( .A0(n3250), .A1(n65), .B0(n3945), .B1(n245), .C0(n4414), 
        .C1(n3241), .Y(n5423) );
  AOI22X1TS U3165 ( .A0(n452), .A1(n3224), .B0(n4235), .B1(n272), .Y(n5847) );
  AOI222XLTS U3166 ( .A0(n3250), .A1(n66), .B0(n3924), .B1(n242), .C0(n4393), 
        .C1(n3241), .Y(n5846) );
  AOI22X1TS U3167 ( .A0(n454), .A1(n6158), .B0(n4232), .B1(n375), .Y(n5849) );
  AOI222XLTS U3168 ( .A0(n3250), .A1(n67), .B0(n3921), .B1(n362), .C0(n4390), 
        .C1(n3241), .Y(n5848) );
  AOI22X1TS U3169 ( .A0(n456), .A1(n3231), .B0(n4229), .B1(n374), .Y(n5851) );
  AOI222XLTS U3170 ( .A0(n3251), .A1(n68), .B0(n3918), .B1(n242), .C0(n4387), 
        .C1(n3240), .Y(n5850) );
  AOI22X1TS U3171 ( .A0(n457), .A1(n3226), .B0(n4226), .B1(n375), .Y(n5853) );
  AOI222XLTS U3172 ( .A0(n3251), .A1(n69), .B0(n3915), .B1(n242), .C0(n4384), 
        .C1(n3240), .Y(n5852) );
  AOI22X1TS U3173 ( .A0(n459), .A1(n3224), .B0(n4223), .B1(n374), .Y(n5855) );
  AOI222XLTS U3174 ( .A0(n3251), .A1(n70), .B0(n3912), .B1(n245), .C0(n4381), 
        .C1(n3240), .Y(n5854) );
  AOI22X1TS U3175 ( .A0(n462), .A1(n3225), .B0(n4220), .B1(n373), .Y(n5857) );
  AOI222XLTS U3176 ( .A0(n3251), .A1(n71), .B0(n3909), .B1(n359), .C0(n4378), 
        .C1(n3240), .Y(n5856) );
  AOI22X1TS U3177 ( .A0(n466), .A1(n3227), .B0(n4214), .B1(n273), .Y(n5861) );
  AOI222XLTS U3178 ( .A0(n3252), .A1(n72), .B0(n3903), .B1(n358), .C0(n4372), 
        .C1(n3239), .Y(n5860) );
  AOI22X1TS U3179 ( .A0(n470), .A1(n3229), .B0(n4208), .B1(n371), .Y(n5865) );
  AOI222XLTS U3180 ( .A0(n3252), .A1(n73), .B0(n3897), .B1(n358), .C0(n4366), 
        .C1(n3239), .Y(n5864) );
  AOI22X1TS U3181 ( .A0(n472), .A1(n3227), .B0(n4205), .B1(n372), .Y(n5867) );
  AOI222XLTS U3182 ( .A0(n3253), .A1(n74), .B0(n3894), .B1(n361), .C0(n4363), 
        .C1(n3238), .Y(n5866) );
  AOI22X1TS U3183 ( .A0(n476), .A1(n3228), .B0(n4199), .B1(n285), .Y(n5871) );
  AOI222XLTS U3184 ( .A0(n3253), .A1(n75), .B0(n3888), .B1(n243), .C0(n4357), 
        .C1(n3238), .Y(n5870) );
  AOI22X1TS U3185 ( .A0(n480), .A1(n3226), .B0(n4193), .B1(n285), .Y(n5875) );
  AOI222XLTS U3186 ( .A0(n3254), .A1(n76), .B0(n3882), .B1(n354), .C0(n4351), 
        .C1(n3237), .Y(n5874) );
  AOI22X1TS U3187 ( .A0(n482), .A1(n3226), .B0(n4190), .B1(n372), .Y(n5877) );
  AOI222XLTS U3188 ( .A0(n3254), .A1(n77), .B0(n3879), .B1(n362), .C0(n4348), 
        .C1(n3237), .Y(n5876) );
  AOI22X1TS U3189 ( .A0(n486), .A1(n3225), .B0(n4184), .B1(n286), .Y(n5881) );
  AOI222XLTS U3190 ( .A0(n3254), .A1(n78), .B0(n3873), .B1(n245), .C0(n4342), 
        .C1(n3237), .Y(n5880) );
  AOI22X1TS U3191 ( .A0(n490), .A1(n3229), .B0(n4178), .B1(n273), .Y(n5885) );
  AOI222XLTS U3192 ( .A0(n3255), .A1(n79), .B0(n3867), .B1(n243), .C0(n4336), 
        .C1(n3236), .Y(n5884) );
  AOI22X1TS U3193 ( .A0(n492), .A1(n3223), .B0(n4175), .B1(n371), .Y(n5887) );
  AOI222XLTS U3194 ( .A0(n3255), .A1(n80), .B0(n3864), .B1(n361), .C0(n4333), 
        .C1(n3236), .Y(n5886) );
  AOI22X1TS U3195 ( .A0(n494), .A1(n3223), .B0(n4172), .B1(n286), .Y(n5889) );
  AOI222XLTS U3196 ( .A0(n3255), .A1(n81), .B0(n3861), .B1(n242), .C0(n4330), 
        .C1(n3236), .Y(n5888) );
  AOI22X1TS U3197 ( .A0(n495), .A1(n3223), .B0(n4169), .B1(n371), .Y(n5891) );
  AOI222XLTS U3198 ( .A0(n3256), .A1(n82), .B0(n3858), .B1(n360), .C0(n4327), 
        .C1(n3235), .Y(n5890) );
  AOI22X1TS U3199 ( .A0(n503), .A1(n3223), .B0(n4166), .B1(n375), .Y(n5893) );
  AOI222XLTS U3200 ( .A0(n3256), .A1(n83), .B0(n3855), .B1(n357), .C0(n4324), 
        .C1(n3235), .Y(n5892) );
  AOI22X1TS U3201 ( .A0(n509), .A1(n3222), .B0(n4160), .B1(n273), .Y(n5897) );
  AOI222XLTS U3202 ( .A0(n3256), .A1(n84), .B0(n3849), .B1(n360), .C0(n4318), 
        .C1(n3235), .Y(n5896) );
  AOI22X1TS U3203 ( .A0(n516), .A1(n3221), .B0(n4151), .B1(n373), .Y(n5903) );
  AOI222XLTS U3204 ( .A0(n3257), .A1(n85), .B0(n3840), .B1(n361), .C0(n4309), 
        .C1(n3234), .Y(n5902) );
  AOI22X1TS U3205 ( .A0(n536), .A1(n3221), .B0(n4145), .B1(n272), .Y(n5907) );
  AOI222XLTS U3206 ( .A0(n3258), .A1(n86), .B0(n3834), .B1(n358), .C0(n4303), 
        .C1(n3233), .Y(n5906) );
  AOI22X1TS U3207 ( .A0(n541), .A1(n3221), .B0(n4142), .B1(n370), .Y(n5909) );
  AOI222XLTS U3208 ( .A0(n3258), .A1(n87), .B0(n3831), .B1(n359), .C0(n4300), 
        .C1(n3233), .Y(n5908) );
  AOI22X1TS U3209 ( .A0(n737), .A1(n188), .B0(n4268), .B1(n714), .Y(n5345) );
  AOI222XLTS U3210 ( .A0(n347), .A1(n88), .B0(n3957), .B1(n766), .C0(n4426), 
        .C1(n3803), .Y(n5344) );
  AOI22X1TS U3211 ( .A0(n737), .A1(n165), .B0(n4256), .B1(n734), .Y(n5353) );
  AOI222XLTS U3212 ( .A0(n382), .A1(n89), .B0(n3945), .B1(n6114), .C0(n4414), 
        .C1(n3802), .Y(n5352) );
  AOI22X1TS U3213 ( .A0(n3219), .A1(n178), .B0(n4262), .B1(n373), .Y(n5420) );
  AOI222XLTS U3214 ( .A0(n3249), .A1(n90), .B0(n3951), .B1(n243), .C0(n4420), 
        .C1(n3242), .Y(n5419) );
  AOI22X1TS U3215 ( .A0(n464), .A1(n3228), .B0(n4217), .B1(n272), .Y(n5859) );
  AOI222XLTS U3216 ( .A0(n3252), .A1(n91), .B0(n3906), .B1(n243), .C0(n4375), 
        .C1(n3239), .Y(n5858) );
  AOI22X1TS U3217 ( .A0(n467), .A1(n6158), .B0(n4211), .B1(n370), .Y(n5863) );
  AOI222XLTS U3218 ( .A0(n3252), .A1(n92), .B0(n3900), .B1(n358), .C0(n4369), 
        .C1(n3239), .Y(n5862) );
  AOI22X1TS U3219 ( .A0(n473), .A1(n3225), .B0(n4202), .B1(n285), .Y(n5869) );
  AOI222XLTS U3220 ( .A0(n3253), .A1(n93), .B0(n3891), .B1(n357), .C0(n4360), 
        .C1(n3238), .Y(n5868) );
  AOI22X1TS U3221 ( .A0(n478), .A1(n3226), .B0(n4196), .B1(n372), .Y(n5873) );
  AOI222XLTS U3222 ( .A0(n3253), .A1(n94), .B0(n3885), .B1(n355), .C0(n4354), 
        .C1(n3238), .Y(n5872) );
  AOI22X1TS U3223 ( .A0(n484), .A1(n3225), .B0(n4187), .B1(n286), .Y(n5879) );
  AOI222XLTS U3224 ( .A0(n3254), .A1(n95), .B0(n3876), .B1(n247), .C0(n4345), 
        .C1(n3237), .Y(n5878) );
  AOI22X1TS U3225 ( .A0(n488), .A1(n3230), .B0(n4181), .B1(n372), .Y(n5883) );
  AOI222XLTS U3226 ( .A0(n3255), .A1(n96), .B0(n3870), .B1(n247), .C0(n4339), 
        .C1(n3236), .Y(n5882) );
  AOI22X1TS U3227 ( .A0(n510), .A1(n3222), .B0(n4157), .B1(n374), .Y(n5899) );
  AOI222XLTS U3228 ( .A0(n3257), .A1(n97), .B0(n3846), .B1(n356), .C0(n4315), 
        .C1(n3234), .Y(n5898) );
  AOI22X1TS U3229 ( .A0(n514), .A1(n3222), .B0(n4154), .B1(n374), .Y(n5901) );
  AOI222XLTS U3230 ( .A0(n3257), .A1(n98), .B0(n3843), .B1(n247), .C0(n4312), 
        .C1(n3234), .Y(n5900) );
  AOI22X1TS U3231 ( .A0(n526), .A1(n3221), .B0(n4148), .B1(n370), .Y(n5905) );
  AOI222XLTS U3232 ( .A0(n3257), .A1(n99), .B0(n3837), .B1(n356), .C0(n4306), 
        .C1(n3234), .Y(n5904) );
  AOI22X1TS U3233 ( .A0(n458), .A1(n746), .B0(n4226), .B1(n728), .Y(n6045) );
  AOI222XLTS U3234 ( .A0(n299), .A1(n100), .B0(n3915), .B1(n761), .C0(n4384), 
        .C1(n3801), .Y(n6044) );
  AOI22X1TS U3235 ( .A0(n460), .A1(n748), .B0(n4223), .B1(n733), .Y(n6047) );
  AOI222XLTS U3236 ( .A0(n382), .A1(n101), .B0(n3912), .B1(n761), .C0(n4381), 
        .C1(n3801), .Y(n6046) );
  AOI22X1TS U3237 ( .A0(n468), .A1(n749), .B0(n4211), .B1(n732), .Y(n6055) );
  AOI222XLTS U3238 ( .A0(n299), .A1(n102), .B0(n3900), .B1(n760), .C0(n4369), 
        .C1(n3800), .Y(n6054) );
  AOI22X1TS U3239 ( .A0(n474), .A1(n738), .B0(n4202), .B1(n712), .Y(n6061) );
  AOI222XLTS U3240 ( .A0(n385), .A1(n103), .B0(n3891), .B1(n759), .C0(n4360), 
        .C1(n3799), .Y(n6060) );
  AOI22X1TS U3241 ( .A0(n496), .A1(n741), .B0(n4169), .B1(n712), .Y(n6083) );
  AOI222XLTS U3242 ( .A0(n3781), .A1(n104), .B0(n3858), .B1(n756), .C0(n4327), 
        .C1(n3804), .Y(n6082) );
  AOI22X1TS U3243 ( .A0(n511), .A1(n741), .B0(n4157), .B1(n706), .Y(n6091) );
  AOI222XLTS U3244 ( .A0(n382), .A1(n105), .B0(n3846), .B1(n755), .C0(n4315), 
        .C1(n3807), .Y(n6090) );
  AOI22X1TS U3245 ( .A0(n531), .A1(n742), .B0(n4148), .B1(n706), .Y(n6097) );
  AOI222XLTS U3246 ( .A0(n384), .A1(n106), .B0(n3837), .B1(n755), .C0(n4306), 
        .C1(n3805), .Y(n6096) );
  AOI22X1TS U3247 ( .A0(n537), .A1(n742), .B0(n4145), .B1(n705), .Y(n6099) );
  AOI222XLTS U3248 ( .A0(n344), .A1(n107), .B0(n3834), .B1(n754), .C0(n4303), 
        .C1(n3807), .Y(n6098) );
  AOI22X1TS U3249 ( .A0(n543), .A1(n743), .B0(n4142), .B1(n705), .Y(n6101) );
  AOI222XLTS U3250 ( .A0(n382), .A1(n108), .B0(n3831), .B1(n754), .C0(n4300), 
        .C1(n3807), .Y(n6100) );
  AOI22X1TS U3251 ( .A0(n507), .A1(n3222), .B0(n4163), .B1(n375), .Y(n5895) );
  AOI222XLTS U3252 ( .A0(n3256), .A1(n109), .B0(n3852), .B1(n357), .C0(n4321), 
        .C1(n3235), .Y(n5894) );
  AOI22X1TS U3253 ( .A0(n886), .A1(n175), .B0(n4106), .B1(n868), .Y(n5394) );
  AOI222XLTS U3254 ( .A0(n291), .A1(n110), .B0(n4263), .B1(n3196), .C0(n4420), 
        .C1(n3761), .Y(n5393) );
  AOI22X1TS U3255 ( .A0(n453), .A1(n919), .B0(n4076), .B1(n862), .Y(n5913) );
  AOI222XLTS U3256 ( .A0(n379), .A1(n111), .B0(n4233), .B1(n3193), .C0(n4390), 
        .C1(n3760), .Y(n5912) );
  AOI22X1TS U3257 ( .A0(n455), .A1(n919), .B0(n4073), .B1(n865), .Y(n5915) );
  AOI222XLTS U3258 ( .A0(n3752), .A1(n112), .B0(n4230), .B1(n3199), .C0(n4387), 
        .C1(n3759), .Y(n5914) );
  AOI22X1TS U3259 ( .A0(n457), .A1(n919), .B0(n4070), .B1(n868), .Y(n5917) );
  AOI222XLTS U3260 ( .A0(n298), .A1(n113), .B0(n4227), .B1(n3199), .C0(n4384), 
        .C1(n3759), .Y(n5916) );
  AOI22X1TS U3261 ( .A0(n461), .A1(n959), .B0(n4064), .B1(n865), .Y(n5921) );
  AOI222XLTS U3262 ( .A0(n291), .A1(n114), .B0(n4221), .B1(n3195), .C0(n4378), 
        .C1(n3759), .Y(n5920) );
  AOI22X1TS U3263 ( .A0(n463), .A1(n919), .B0(n4061), .B1(n861), .Y(n5923) );
  AOI222XLTS U3264 ( .A0(n380), .A1(n115), .B0(n4218), .B1(n3197), .C0(n4375), 
        .C1(n3758), .Y(n5922) );
  AOI22X1TS U3265 ( .A0(n467), .A1(n936), .B0(n4055), .B1(n861), .Y(n5927) );
  AOI222XLTS U3266 ( .A0(n292), .A1(n116), .B0(n4212), .B1(n3197), .C0(n4369), 
        .C1(n3758), .Y(n5926) );
  AOI22X1TS U3267 ( .A0(n471), .A1(n955), .B0(n4049), .B1(n860), .Y(n5931) );
  AOI222XLTS U3268 ( .A0(n378), .A1(n117), .B0(n4206), .B1(n1894), .C0(n4363), 
        .C1(n3757), .Y(n5930) );
  AOI22X1TS U3269 ( .A0(n473), .A1(n955), .B0(n4046), .B1(n860), .Y(n5933) );
  AOI222XLTS U3270 ( .A0(n381), .A1(n118), .B0(n4203), .B1(n1894), .C0(n4360), 
        .C1(n3757), .Y(n5932) );
  AOI22X1TS U3271 ( .A0(n475), .A1(n955), .B0(n4043), .B1(n860), .Y(n5935) );
  AOI222XLTS U3272 ( .A0(n291), .A1(n119), .B0(n4200), .B1(n1894), .C0(n4357), 
        .C1(n3757), .Y(n5934) );
  AOI22X1TS U3273 ( .A0(n477), .A1(n957), .B0(n4040), .B1(n859), .Y(n5937) );
  AOI222XLTS U3274 ( .A0(n259), .A1(n120), .B0(n4197), .B1(n1822), .C0(n4354), 
        .C1(n3757), .Y(n5936) );
  AOI22X1TS U3275 ( .A0(n479), .A1(n955), .B0(n4037), .B1(n859), .Y(n5939) );
  AOI222XLTS U3276 ( .A0(n379), .A1(n121), .B0(n4194), .B1(n1822), .C0(n4351), 
        .C1(n3756), .Y(n5938) );
  AOI22X1TS U3277 ( .A0(n483), .A1(n959), .B0(n4031), .B1(n859), .Y(n5943) );
  AOI222XLTS U3278 ( .A0(n292), .A1(n122), .B0(n4188), .B1(n1822), .C0(n4345), 
        .C1(n3756), .Y(n5942) );
  AOI22X1TS U3279 ( .A0(n485), .A1(n957), .B0(n4028), .B1(n858), .Y(n5945) );
  AOI222XLTS U3280 ( .A0(n380), .A1(n123), .B0(n4185), .B1(n1817), .C0(n4342), 
        .C1(n3756), .Y(n5944) );
  AOI22X1TS U3281 ( .A0(n487), .A1(n957), .B0(n4025), .B1(n858), .Y(n5947) );
  AOI222XLTS U3282 ( .A0(n291), .A1(n124), .B0(n4182), .B1(n1817), .C0(n4339), 
        .C1(n3755), .Y(n5946) );
  AOI22X1TS U3283 ( .A0(n489), .A1(n959), .B0(n4022), .B1(n858), .Y(n5949) );
  AOI222XLTS U3284 ( .A0(n296), .A1(n125), .B0(n4179), .B1(n1817), .C0(n4336), 
        .C1(n3755), .Y(n5948) );
  AOI22X1TS U3285 ( .A0(n491), .A1(n959), .B0(n4019), .B1(n858), .Y(n5951) );
  AOI222XLTS U3286 ( .A0(n380), .A1(n126), .B0(n4176), .B1(n1817), .C0(n4333), 
        .C1(n3755), .Y(n5950) );
  AOI22X1TS U3287 ( .A0(n495), .A1(n970), .B0(n4013), .B1(n860), .Y(n5955) );
  AOI222XLTS U3288 ( .A0(n296), .A1(n127), .B0(n4170), .B1(n1797), .C0(n4327), 
        .C1(n3754), .Y(n5954) );
  AOI22X1TS U3289 ( .A0(n501), .A1(n970), .B0(n4010), .B1(n857), .Y(n5957) );
  AOI222XLTS U3290 ( .A0(n298), .A1(n128), .B0(n4167), .B1(n1797), .C0(n4324), 
        .C1(n3754), .Y(n5956) );
  AOI22X1TS U3291 ( .A0(n505), .A1(n970), .B0(n4007), .B1(n857), .Y(n5959) );
  AOI222XLTS U3292 ( .A0(n340), .A1(n129), .B0(n4164), .B1(n1797), .C0(n4321), 
        .C1(n3754), .Y(n5958) );
  AOI22X1TS U3293 ( .A0(n510), .A1(n970), .B0(n4001), .B1(n856), .Y(n5963) );
  AOI22X1TS U3294 ( .A0(n512), .A1(n986), .B0(n3998), .B1(n856), .Y(n5965) );
  AOI222XLTS U3295 ( .A0(n381), .A1(n131), .B0(n4155), .B1(n1728), .C0(n4312), 
        .C1(n3762), .Y(n5964) );
  AOI22X1TS U3296 ( .A0(n515), .A1(n1402), .B0(n3995), .B1(n856), .Y(n5967) );
  AOI222XLTS U3297 ( .A0(n381), .A1(n132), .B0(n4152), .B1(n1728), .C0(n4309), 
        .C1(n3765), .Y(n5966) );
  AOI22X1TS U3298 ( .A0(n3941), .A1(n3465), .B0(n4410), .B1(n3691), .Y(n6211)
         );
  AOI222XLTS U3299 ( .A0(n4097), .A1(n3513), .B0(n159), .B1(n3503), .C0(n4254), 
        .C1(n3484), .Y(n6210) );
  AOI22X1TS U3300 ( .A0(n3938), .A1(n3464), .B0(n4407), .B1(n3691), .Y(n6213)
         );
  AOI222XLTS U3301 ( .A0(n4094), .A1(n3512), .B0(readRequesterAddress[4]), 
        .B1(n3503), .C0(n4251), .C1(n3484), .Y(n6212) );
  AOI22X1TS U3302 ( .A0(n3932), .A1(n3464), .B0(n4401), .B1(n3692), .Y(n6217)
         );
  AOI222XLTS U3303 ( .A0(n4088), .A1(n3512), .B0(readRequesterAddress[2]), 
        .B1(n3504), .C0(n4245), .C1(n3484), .Y(n6216) );
  AOI22X1TS U3304 ( .A0(n1598), .A1(n191), .B0(n4115), .B1(n866), .Y(n5388) );
  AOI222XLTS U3305 ( .A0(n378), .A1(n133), .B0(n4272), .B1(n1654), .C0(n4429), 
        .C1(n3761), .Y(n5387) );
  AOI22X1TS U3306 ( .A0(n886), .A1(n185), .B0(n4112), .B1(n867), .Y(n5390) );
  AOI222XLTS U3307 ( .A0(n296), .A1(n134), .B0(n4269), .B1(n3193), .C0(n4426), 
        .C1(n3761), .Y(n5389) );
  AOI22X1TS U3308 ( .A0(n886), .A1(n181), .B0(n4109), .B1(n870), .Y(n5392) );
  AOI222XLTS U3309 ( .A0(n298), .A1(n135), .B0(n4266), .B1(n3198), .C0(n4423), 
        .C1(n3761), .Y(n5391) );
  AOI22X1TS U3310 ( .A0(n871), .A1(n170), .B0(n4103), .B1(n862), .Y(n5396) );
  AOI222XLTS U3311 ( .A0(n296), .A1(n136), .B0(n4260), .B1(n3193), .C0(n4417), 
        .C1(n3760), .Y(n5395) );
  AOI22X1TS U3312 ( .A0(n886), .A1(n166), .B0(n4100), .B1(n862), .Y(n5398) );
  AOI222XLTS U3313 ( .A0(n292), .A1(n137), .B0(n4257), .B1(n3194), .C0(n4414), 
        .C1(n3760), .Y(n5397) );
  AOI22X1TS U3314 ( .A0(n459), .A1(n936), .B0(n4067), .B1(n866), .Y(n5919) );
  AOI222XLTS U3315 ( .A0(n259), .A1(n138), .B0(n4224), .B1(n6145), .C0(n4381), 
        .C1(n3759), .Y(n5918) );
  AOI22X1TS U3316 ( .A0(n493), .A1(n1402), .B0(n4016), .B1(n857), .Y(n5953) );
  AOI222XLTS U3317 ( .A0(n341), .A1(n139), .B0(n4173), .B1(n1797), .C0(n4330), 
        .C1(n3755), .Y(n5952) );
  AOI22X1TS U3318 ( .A0(n536), .A1(n986), .B0(n3989), .B1(n855), .Y(n5971) );
  AOI222XLTS U3319 ( .A0(n341), .A1(n140), .B0(n4146), .B1(n1654), .C0(n4303), 
        .C1(n3764), .Y(n5970) );
  AOI22X1TS U3320 ( .A0(n3935), .A1(n3464), .B0(n4404), .B1(n3692), .Y(n6215)
         );
  AOI222XLTS U3321 ( .A0(n4091), .A1(n3512), .B0(readRequesterAddress[3]), 
        .B1(n3504), .C0(n4248), .C1(n3483), .Y(n6214) );
  AOI22X1TS U3322 ( .A0(n3929), .A1(n3464), .B0(n4398), .B1(n3692), .Y(n6219)
         );
  AOI222XLTS U3323 ( .A0(n4085), .A1(n3512), .B0(readRequesterAddress[1]), 
        .B1(n3504), .C0(n4242), .C1(n3483), .Y(n6218) );
  AOI22X1TS U3324 ( .A0(n3926), .A1(n3470), .B0(n4395), .B1(n3692), .Y(n6225)
         );
  AOI222XLTS U3325 ( .A0(n4082), .A1(n3524), .B0(readRequesterAddress[0]), 
        .B1(n3504), .C0(n4239), .C1(n3492), .Y(n6224) );
  AOI22X1TS U3326 ( .A0(n451), .A1(n1402), .B0(n4079), .B1(n862), .Y(n5911) );
  AOI222XLTS U3327 ( .A0(n380), .A1(n141), .B0(n4236), .B1(n3194), .C0(n4393), 
        .C1(n3760), .Y(n5910) );
  AOI22X1TS U3328 ( .A0(n465), .A1(n936), .B0(n4058), .B1(n861), .Y(n5925) );
  AOI222XLTS U3329 ( .A0(n341), .A1(n142), .B0(n4215), .B1(n3192), .C0(n4372), 
        .C1(n3758), .Y(n5924) );
  AOI22X1TS U3330 ( .A0(n469), .A1(n936), .B0(n4052), .B1(n861), .Y(n5929) );
  AOI222XLTS U3331 ( .A0(n298), .A1(n143), .B0(n4209), .B1(n3192), .C0(n4366), 
        .C1(n3758), .Y(n5928) );
  AOI22X1TS U3332 ( .A0(n481), .A1(n957), .B0(n4034), .B1(n859), .Y(n5941) );
  AOI222XLTS U3333 ( .A0(n340), .A1(n144), .B0(n4191), .B1(n1822), .C0(n4348), 
        .C1(n3756), .Y(n5940) );
  AOI22X1TS U3334 ( .A0(n508), .A1(n986), .B0(n4004), .B1(n857), .Y(n5961) );
  AOI222XLTS U3335 ( .A0(n6306), .A1(n145), .B0(n4161), .B1(n1894), .C0(n4318), 
        .C1(n3754), .Y(n5960) );
  AOI22X1TS U3336 ( .A0(n526), .A1(n986), .B0(n3992), .B1(n856), .Y(n5969) );
  AOI222XLTS U3337 ( .A0(n340), .A1(n146), .B0(n4149), .B1(n1728), .C0(n4306), 
        .C1(n3765), .Y(n5968) );
  AOI22X1TS U3338 ( .A0(n541), .A1(n1402), .B0(n3986), .B1(n855), .Y(n5973) );
  AOI222XLTS U3339 ( .A0(n292), .A1(n147), .B0(n4143), .B1(n1654), .C0(n4300), 
        .C1(n3766), .Y(n5972) );
  AOI22XLTS U3340 ( .A0(n3820), .A1(n5569), .B0(n3815), .B1(n5568), .Y(n5570)
         );
  AOI222XLTS U3341 ( .A0(n3820), .A1(n5562), .B0(readIn_SOUTH), .B1(n5561), 
        .C0(n3828), .C1(n5560), .Y(n5563) );
  NAND2X1TS U3342 ( .A(n3814), .B(n6301), .Y(n5551) );
  AOI2BB2X1TS U3343 ( .B0(n5545), .B1(n5544), .A0N(n3260), .A1N(
        readOutbuffer[3]), .Y(n2566) );
  OAI22X1TS U3344 ( .A0(n441), .A1(n6235), .B0(n568), .B1(n6236), .Y(n2887) );
  CLKBUFX2TS U3345 ( .A(n5323), .Y(n568) );
  OAI22X1TS U3346 ( .A0(n6238), .A1(n441), .B0(n570), .B1(n6236), .Y(n2888) );
  OAI22X1TS U3347 ( .A0(n670), .A1(n4719), .B0(n5142), .B1(n3564), .Y(n5143)
         );
  NOR4XLTS U3348 ( .A(n5141), .B(n5140), .C(n5139), .D(n5138), .Y(n5142) );
  AO22X1TS U3349 ( .A0(n241), .A1(\requesterAddressbuffer[3][5] ), .B0(
        \requesterAddressbuffer[6][5] ), .B1(n5294), .Y(n5140) );
  OAI2BB2XLTS U3350 ( .B0(n6269), .B1(n3609), .A0N(
        \requesterAddressbuffer[0][5] ), .A1N(n288), .Y(n5141) );
  OAI22X1TS U3351 ( .A0(n670), .A1(n4720), .B0(n5150), .B1(n3564), .Y(n5151)
         );
  NOR4XLTS U3352 ( .A(n5149), .B(n5148), .C(n5147), .D(n5146), .Y(n5150) );
  AO22X1TS U3353 ( .A0(n293), .A1(\requesterAddressbuffer[3][4] ), .B0(
        \requesterAddressbuffer[6][4] ), .B1(n5294), .Y(n5148) );
  OAI2BB2XLTS U3354 ( .B0(n6270), .B1(n3609), .A0N(
        \requesterAddressbuffer[0][4] ), .A1N(n5295), .Y(n5149) );
  OAI22X1TS U3355 ( .A0(n669), .A1(n4721), .B0(n5166), .B1(n3563), .Y(n5167)
         );
  NOR4XLTS U3356 ( .A(n5165), .B(n5164), .C(n5163), .D(n5162), .Y(n5166) );
  AO22X1TS U3357 ( .A0(n241), .A1(\requesterAddressbuffer[3][2] ), .B0(
        \requesterAddressbuffer[6][2] ), .B1(n5294), .Y(n5164) );
  OAI2BB2XLTS U3358 ( .B0(n6260), .B1(n3608), .A0N(
        \requesterAddressbuffer[0][2] ), .A1N(n288), .Y(n5165) );
  OAI22X1TS U3359 ( .A0(n669), .A1(n4722), .B0(n5174), .B1(n3563), .Y(n5175)
         );
  NOR4XLTS U3360 ( .A(n5173), .B(n5172), .C(n5171), .D(n5170), .Y(n5174) );
  AO22X1TS U3361 ( .A0(n293), .A1(\requesterAddressbuffer[3][1] ), .B0(
        \requesterAddressbuffer[6][1] ), .B1(n450), .Y(n5172) );
  OAI2BB2XLTS U3362 ( .B0(n6261), .B1(n3608), .A0N(
        \requesterAddressbuffer[0][1] ), .A1N(n5295), .Y(n5173) );
  OAI22X1TS U3363 ( .A0(n669), .A1(n4846), .B0(n5158), .B1(n3563), .Y(n5159)
         );
  NOR4XLTS U3364 ( .A(n5157), .B(n5156), .C(n5155), .D(n5154), .Y(n5158) );
  AO22X1TS U3365 ( .A0(n241), .A1(\requesterAddressbuffer[3][3] ), .B0(
        \requesterAddressbuffer[6][3] ), .B1(n450), .Y(n5156) );
  OAI2BB2XLTS U3366 ( .B0(n6259), .B1(n3608), .A0N(
        \requesterAddressbuffer[0][3] ), .A1N(n288), .Y(n5157) );
  OAI22X1TS U3367 ( .A0(n669), .A1(n4845), .B0(n5182), .B1(n3563), .Y(n5183)
         );
  NOR4XLTS U3368 ( .A(n5181), .B(n5180), .C(n5179), .D(n5178), .Y(n5182) );
  AO22X1TS U3369 ( .A0(n293), .A1(\requesterAddressbuffer[3][0] ), .B0(
        \requesterAddressbuffer[6][0] ), .B1(n450), .Y(n5180) );
  OAI2BB2XLTS U3370 ( .B0(n6262), .B1(n3608), .A0N(
        \requesterAddressbuffer[0][0] ), .A1N(n5295), .Y(n5181) );
  OAI22X1TS U3371 ( .A0(n4431), .A1(n670), .B0(n4886), .B1(n3561), .Y(n4887)
         );
  NOR4XLTS U3372 ( .A(n4885), .B(n4884), .C(n4883), .D(n4882), .Y(n4886) );
  OAI22X1TS U3373 ( .A0(n4432), .A1(n3593), .B0(n4433), .B1(n3612), .Y(n4885)
         );
  OAI22X1TS U3374 ( .A0(n4434), .A1(n3640), .B0(n4435), .B1(n3655), .Y(n4884)
         );
  OAI22X1TS U3375 ( .A0(n4440), .A1(n679), .B0(n4894), .B1(n3575), .Y(n4895)
         );
  NOR4XLTS U3376 ( .A(n4893), .B(n4892), .C(n4891), .D(n4890), .Y(n4894) );
  OAI22X1TS U3377 ( .A0(n4445), .A1(n3593), .B0(n4441), .B1(n3622), .Y(n4893)
         );
  OAI22X1TS U3378 ( .A0(n4447), .A1(n3649), .B0(n4446), .B1(n3655), .Y(n4892)
         );
  OAI22X1TS U3379 ( .A0(n4449), .A1(n679), .B0(n4902), .B1(n3573), .Y(n4903)
         );
  NOR4XLTS U3380 ( .A(n4901), .B(n4900), .C(n4899), .D(n4898), .Y(n4902) );
  OAI22X1TS U3381 ( .A0(n4456), .A1(n3593), .B0(n4457), .B1(n6280), .Y(n4901)
         );
  OAI22X1TS U3382 ( .A0(n4452), .A1(n3649), .B0(n4454), .B1(n3655), .Y(n4900)
         );
  OAI22X1TS U3383 ( .A0(n4458), .A1(n679), .B0(n4910), .B1(n3570), .Y(n4911)
         );
  NOR4XLTS U3384 ( .A(n4909), .B(n4908), .C(n4907), .D(n4906), .Y(n4910) );
  OAI22X1TS U3385 ( .A0(n4465), .A1(n3593), .B0(n4459), .B1(n3619), .Y(n4909)
         );
  OAI22X1TS U3386 ( .A0(n4463), .A1(n3649), .B0(n4462), .B1(n3655), .Y(n4908)
         );
  OAI22X1TS U3387 ( .A0(n4467), .A1(n679), .B0(n4918), .B1(n3575), .Y(n4919)
         );
  NOR4XLTS U3388 ( .A(n4917), .B(n4916), .C(n4915), .D(n4914), .Y(n4918) );
  OAI22X1TS U3389 ( .A0(n4474), .A1(n3594), .B0(n4470), .B1(n3618), .Y(n4917)
         );
  OAI22X1TS U3390 ( .A0(n4472), .A1(n3648), .B0(n4471), .B1(n3656), .Y(n4916)
         );
  OAI22X1TS U3391 ( .A0(n4476), .A1(n678), .B0(n4926), .B1(n3572), .Y(n4927)
         );
  NOR4XLTS U3392 ( .A(n4925), .B(n4924), .C(n4923), .D(n4922), .Y(n4926) );
  OAI22X1TS U3393 ( .A0(n4481), .A1(n3594), .B0(n4477), .B1(n3621), .Y(n4925)
         );
  OAI22X1TS U3394 ( .A0(n4483), .A1(n3648), .B0(n4482), .B1(n3656), .Y(n4924)
         );
  OAI22X1TS U3395 ( .A0(n4485), .A1(n678), .B0(n4934), .B1(n3570), .Y(n4935)
         );
  NOR4XLTS U3396 ( .A(n4933), .B(n4932), .C(n4931), .D(n4930), .Y(n4934) );
  OAI22X1TS U3397 ( .A0(n4488), .A1(n3594), .B0(n4490), .B1(n3617), .Y(n4933)
         );
  OAI22X1TS U3398 ( .A0(n4487), .A1(n3648), .B0(n4492), .B1(n3656), .Y(n4932)
         );
  OAI22X1TS U3399 ( .A0(n4494), .A1(n678), .B0(n4942), .B1(n3571), .Y(n4943)
         );
  NOR4XLTS U3400 ( .A(n4941), .B(n4940), .C(n4939), .D(n4938), .Y(n4942) );
  OAI22X1TS U3401 ( .A0(n4497), .A1(n3594), .B0(n4495), .B1(n3622), .Y(n4941)
         );
  OAI22X1TS U3402 ( .A0(n4499), .A1(n3648), .B0(n4502), .B1(n3656), .Y(n4940)
         );
  OAI22X1TS U3403 ( .A0(n4503), .A1(n678), .B0(n4950), .B1(n3571), .Y(n4951)
         );
  NOR4XLTS U3404 ( .A(n4949), .B(n4948), .C(n4947), .D(n4946), .Y(n4950) );
  OAI22X1TS U3405 ( .A0(n4510), .A1(n3606), .B0(n4506), .B1(n3622), .Y(n4949)
         );
  OAI22X1TS U3406 ( .A0(n4511), .A1(n3647), .B0(n4504), .B1(n3668), .Y(n4948)
         );
  OAI22X1TS U3407 ( .A0(n4512), .A1(n677), .B0(n4958), .B1(n3572), .Y(n4959)
         );
  NOR4XLTS U3408 ( .A(n4957), .B(n4956), .C(n4955), .D(n4954), .Y(n4958) );
  OAI22X1TS U3409 ( .A0(n4513), .A1(n3603), .B0(n4516), .B1(n3616), .Y(n4957)
         );
  OAI22X1TS U3410 ( .A0(n4515), .A1(n3647), .B0(n4520), .B1(n3665), .Y(n4956)
         );
  OAI22X1TS U3411 ( .A0(n4521), .A1(n677), .B0(n4966), .B1(n3575), .Y(n4967)
         );
  NOR4XLTS U3412 ( .A(n4965), .B(n4964), .C(n4963), .D(n4962), .Y(n4966) );
  OAI22X1TS U3413 ( .A0(n4528), .A1(n3604), .B0(n4527), .B1(n3620), .Y(n4965)
         );
  OAI22X1TS U3414 ( .A0(n4526), .A1(n3647), .B0(n4524), .B1(n3667), .Y(n4964)
         );
  OAI22X1TS U3415 ( .A0(n4530), .A1(n677), .B0(n4974), .B1(n3569), .Y(n4975)
         );
  NOR4XLTS U3416 ( .A(n4973), .B(n4972), .C(n4971), .D(n4970), .Y(n4974) );
  OAI22X1TS U3417 ( .A0(n4537), .A1(n3601), .B0(n4536), .B1(n3620), .Y(n4973)
         );
  OAI22X1TS U3418 ( .A0(n4538), .A1(n3647), .B0(n4531), .B1(n3663), .Y(n4972)
         );
  OAI22X1TS U3419 ( .A0(n4539), .A1(n677), .B0(n4982), .B1(n3569), .Y(n4983)
         );
  NOR4XLTS U3420 ( .A(n4981), .B(n4980), .C(n4979), .D(n4978), .Y(n4982) );
  OAI22X1TS U3421 ( .A0(n4542), .A1(n3605), .B0(n4541), .B1(n3620), .Y(n4981)
         );
  OAI22X1TS U3422 ( .A0(n4546), .A1(n3646), .B0(n4543), .B1(n3666), .Y(n4980)
         );
  OAI22X1TS U3423 ( .A0(n4548), .A1(n676), .B0(n4990), .B1(n3569), .Y(n4991)
         );
  NOR4XLTS U3424 ( .A(n4989), .B(n4988), .C(n4987), .D(n4986), .Y(n4990) );
  OAI22X1TS U3425 ( .A0(n4551), .A1(n3603), .B0(n4549), .B1(n3623), .Y(n4989)
         );
  OAI22X1TS U3426 ( .A0(n4554), .A1(n3646), .B0(n4555), .B1(n6282), .Y(n4988)
         );
  OAI22X1TS U3427 ( .A0(n4557), .A1(n676), .B0(n4998), .B1(n3569), .Y(n4999)
         );
  NOR4XLTS U3428 ( .A(n4997), .B(n4996), .C(n4995), .D(n4994), .Y(n4998) );
  OAI22X1TS U3429 ( .A0(n4560), .A1(n3605), .B0(n4564), .B1(n3623), .Y(n4997)
         );
  OAI22X1TS U3430 ( .A0(n4558), .A1(n3646), .B0(n4565), .B1(n3665), .Y(n4996)
         );
  OAI22X1TS U3431 ( .A0(n4566), .A1(n676), .B0(n5006), .B1(n3568), .Y(n5007)
         );
  NOR4XLTS U3432 ( .A(n5005), .B(n5004), .C(n5003), .D(n5002), .Y(n5006) );
  OAI22X1TS U3433 ( .A0(n4569), .A1(n3604), .B0(n4568), .B1(n3623), .Y(n5005)
         );
  OAI22X1TS U3434 ( .A0(n4567), .A1(n3646), .B0(n4570), .B1(n3666), .Y(n5004)
         );
  OAI22X1TS U3435 ( .A0(n4575), .A1(n676), .B0(n5014), .B1(n3568), .Y(n5015)
         );
  NOR4XLTS U3436 ( .A(n5013), .B(n5012), .C(n5011), .D(n5010), .Y(n5014) );
  OAI22X1TS U3437 ( .A0(n4580), .A1(n3602), .B0(n4582), .B1(n3616), .Y(n5013)
         );
  OAI22X1TS U3438 ( .A0(n4579), .A1(n3645), .B0(n4583), .B1(n3664), .Y(n5012)
         );
  OAI22X1TS U3439 ( .A0(n4584), .A1(n675), .B0(n5022), .B1(n3568), .Y(n5023)
         );
  NOR4XLTS U3440 ( .A(n5021), .B(n5020), .C(n5019), .D(n5018), .Y(n5022) );
  OAI22X1TS U3441 ( .A0(n4587), .A1(n3602), .B0(n4591), .B1(n3613), .Y(n5021)
         );
  OAI22X1TS U3442 ( .A0(n4589), .A1(n3645), .B0(n4590), .B1(n3664), .Y(n5020)
         );
  OAI22X1TS U3443 ( .A0(n4593), .A1(n675), .B0(n5030), .B1(n3568), .Y(n5031)
         );
  NOR4XLTS U3444 ( .A(n5029), .B(n5028), .C(n5027), .D(n5026), .Y(n5030) );
  OAI22X1TS U3445 ( .A0(n4600), .A1(n3606), .B0(n4594), .B1(n3613), .Y(n5029)
         );
  OAI22X1TS U3446 ( .A0(n4597), .A1(n3645), .B0(n4598), .B1(n3667), .Y(n5028)
         );
  OAI22X1TS U3447 ( .A0(n4602), .A1(n675), .B0(n5038), .B1(n3567), .Y(n5039)
         );
  NOR4XLTS U3448 ( .A(n5037), .B(n5036), .C(n5035), .D(n5034), .Y(n5038) );
  OAI22X1TS U3449 ( .A0(n4607), .A1(n3607), .B0(n4606), .B1(n3613), .Y(n5037)
         );
  OAI22X1TS U3450 ( .A0(n4605), .A1(n3645), .B0(n4609), .B1(n3668), .Y(n5036)
         );
  OAI22X1TS U3451 ( .A0(n4611), .A1(n675), .B0(n5046), .B1(n3567), .Y(n5047)
         );
  NOR4XLTS U3452 ( .A(n5045), .B(n5044), .C(n5043), .D(n5042), .Y(n5046) );
  OAI22X1TS U3453 ( .A0(n4612), .A1(n3595), .B0(n4617), .B1(n3613), .Y(n5045)
         );
  OAI22X1TS U3454 ( .A0(n4616), .A1(n3644), .B0(n4619), .B1(n3657), .Y(n5044)
         );
  OAI22X1TS U3455 ( .A0(n4620), .A1(n674), .B0(n5054), .B1(n3567), .Y(n5055)
         );
  NOR4XLTS U3456 ( .A(n5053), .B(n5052), .C(n5051), .D(n5050), .Y(n5054) );
  OAI22X1TS U3457 ( .A0(n4625), .A1(n3595), .B0(n4624), .B1(n3612), .Y(n5053)
         );
  OAI22X1TS U3458 ( .A0(n4623), .A1(n3644), .B0(n4621), .B1(n3657), .Y(n5052)
         );
  OAI22X1TS U3459 ( .A0(n4629), .A1(n674), .B0(n5062), .B1(n3567), .Y(n5063)
         );
  NOR4XLTS U3460 ( .A(n5061), .B(n5060), .C(n5059), .D(n5058), .Y(n5062) );
  OAI22X1TS U3461 ( .A0(n4636), .A1(n3595), .B0(n4634), .B1(n3612), .Y(n5061)
         );
  OAI22X1TS U3462 ( .A0(n4632), .A1(n3644), .B0(n4635), .B1(n3657), .Y(n5060)
         );
  OAI22X1TS U3463 ( .A0(n4638), .A1(n674), .B0(n5070), .B1(n3566), .Y(n5071)
         );
  NOR4XLTS U3464 ( .A(n5069), .B(n5068), .C(n5067), .D(n5066), .Y(n5070) );
  OAI22X1TS U3465 ( .A0(n4645), .A1(n3595), .B0(n4640), .B1(n3612), .Y(n5069)
         );
  OAI22X1TS U3466 ( .A0(n4639), .A1(n3643), .B0(n4646), .B1(n3657), .Y(n5068)
         );
  OAI22X1TS U3467 ( .A0(n4647), .A1(n673), .B0(n5078), .B1(n3566), .Y(n5079)
         );
  NOR4XLTS U3468 ( .A(n5077), .B(n5076), .C(n5075), .D(n5074), .Y(n5078) );
  OAI22X1TS U3469 ( .A0(n4650), .A1(n3596), .B0(n4652), .B1(n3611), .Y(n5077)
         );
  OAI22X1TS U3470 ( .A0(n4654), .A1(n3643), .B0(n4651), .B1(n3658), .Y(n5076)
         );
  OAI22X1TS U3471 ( .A0(n4656), .A1(n673), .B0(n5086), .B1(n3566), .Y(n5087)
         );
  NOR4XLTS U3472 ( .A(n5085), .B(n5084), .C(n5083), .D(n5082), .Y(n5086) );
  OAI22X1TS U3473 ( .A0(n4659), .A1(n3596), .B0(n4662), .B1(n3611), .Y(n5085)
         );
  OAI22X1TS U3474 ( .A0(n4661), .A1(n3643), .B0(n4657), .B1(n3658), .Y(n5084)
         );
  OAI22X1TS U3475 ( .A0(n4665), .A1(n673), .B0(n5094), .B1(n3565), .Y(n5095)
         );
  NOR4XLTS U3476 ( .A(n5093), .B(n5092), .C(n5091), .D(n5090), .Y(n5094) );
  OAI22X1TS U3477 ( .A0(n4672), .A1(n3596), .B0(n4668), .B1(n3611), .Y(n5093)
         );
  OAI22X1TS U3478 ( .A0(n4671), .A1(n3643), .B0(n4669), .B1(n3658), .Y(n5092)
         );
  OAI22X1TS U3479 ( .A0(n4674), .A1(n673), .B0(n5102), .B1(n3565), .Y(n5103)
         );
  NOR4XLTS U3480 ( .A(n5101), .B(n5100), .C(n5099), .D(n5098), .Y(n5102) );
  OAI22X1TS U3481 ( .A0(n4675), .A1(n3596), .B0(n4679), .B1(n3611), .Y(n5101)
         );
  OAI22X1TS U3482 ( .A0(n4678), .A1(n3642), .B0(n4681), .B1(n3658), .Y(n5100)
         );
  OAI22X1TS U3483 ( .A0(n4683), .A1(n672), .B0(n5110), .B1(n3565), .Y(n5111)
         );
  NOR4XLTS U3484 ( .A(n5109), .B(n5108), .C(n5107), .D(n5106), .Y(n5110) );
  OAI22X1TS U3485 ( .A0(n4686), .A1(n3597), .B0(n4690), .B1(n3610), .Y(n5109)
         );
  OAI22X1TS U3486 ( .A0(n4688), .A1(n3642), .B0(n4685), .B1(n3659), .Y(n5108)
         );
  OAI22X1TS U3487 ( .A0(n4692), .A1(n672), .B0(n5118), .B1(n3565), .Y(n5119)
         );
  NOR4XLTS U3488 ( .A(n5117), .B(n5116), .C(n5115), .D(n5114), .Y(n5118) );
  OAI22X1TS U3489 ( .A0(n4699), .A1(n3597), .B0(n4695), .B1(n3610), .Y(n5117)
         );
  OAI22X1TS U3490 ( .A0(n4698), .A1(n3642), .B0(n4700), .B1(n3659), .Y(n5116)
         );
  OAI22X1TS U3491 ( .A0(n4701), .A1(n672), .B0(n5126), .B1(n3564), .Y(n5127)
         );
  NOR4XLTS U3492 ( .A(n5125), .B(n5124), .C(n5123), .D(n5122), .Y(n5126) );
  OAI22X1TS U3493 ( .A0(n4708), .A1(n3597), .B0(n4703), .B1(n3610), .Y(n5125)
         );
  OAI22X1TS U3494 ( .A0(n4702), .A1(n3642), .B0(n4704), .B1(n3659), .Y(n5124)
         );
  OAI22X1TS U3495 ( .A0(n4710), .A1(n672), .B0(n5134), .B1(n3564), .Y(n5135)
         );
  NOR4XLTS U3496 ( .A(n5133), .B(n5132), .C(n5131), .D(n5130), .Y(n5134) );
  OAI22X1TS U3497 ( .A0(n4715), .A1(n3597), .B0(n4714), .B1(n3610), .Y(n5133)
         );
  OAI22X1TS U3498 ( .A0(n4711), .A1(n3641), .B0(n4716), .B1(n3659), .Y(n5132)
         );
  OAI22X1TS U3499 ( .A0(n4723), .A1(n671), .B0(n5190), .B1(n3562), .Y(n5191)
         );
  NOR4XLTS U3500 ( .A(n5189), .B(n5188), .C(n5187), .D(n5186), .Y(n5190) );
  OAI22X1TS U3501 ( .A0(n4724), .A1(n3598), .B0(n4726), .B1(n3619), .Y(n5189)
         );
  OAI22X1TS U3502 ( .A0(n4730), .A1(n3641), .B0(n4728), .B1(n3660), .Y(n5188)
         );
  OAI22X1TS U3503 ( .A0(n4732), .A1(n671), .B0(n5198), .B1(n3562), .Y(n5199)
         );
  NOR4XLTS U3504 ( .A(n5197), .B(n5196), .C(n5195), .D(n5194), .Y(n5198) );
  OAI22X1TS U3505 ( .A0(n4736), .A1(n3598), .B0(n4737), .B1(n3619), .Y(n5197)
         );
  OAI22X1TS U3506 ( .A0(n4735), .A1(n3641), .B0(n4739), .B1(n3660), .Y(n5196)
         );
  OAI22X1TS U3507 ( .A0(n4741), .A1(n674), .B0(n5206), .B1(n3562), .Y(n5207)
         );
  NOR4XLTS U3508 ( .A(n5205), .B(n5204), .C(n5203), .D(n5202), .Y(n5206) );
  OAI22X1TS U3509 ( .A0(n4744), .A1(n3598), .B0(n4746), .B1(n3618), .Y(n5205)
         );
  OAI22X1TS U3510 ( .A0(n4748), .A1(n3641), .B0(n4742), .B1(n3660), .Y(n5204)
         );
  OAI22X1TS U3511 ( .A0(n4750), .A1(n671), .B0(n5214), .B1(n3562), .Y(n5215)
         );
  NOR4XLTS U3512 ( .A(n5213), .B(n5212), .C(n5211), .D(n5210), .Y(n5214) );
  OAI22X1TS U3513 ( .A0(n4755), .A1(n3598), .B0(n4751), .B1(n3609), .Y(n5213)
         );
  OAI22X1TS U3514 ( .A0(n4752), .A1(n3640), .B0(n4753), .B1(n3660), .Y(n5212)
         );
  OAI22X1TS U3515 ( .A0(n4759), .A1(n670), .B0(n5222), .B1(n3561), .Y(n5223)
         );
  NOR4XLTS U3516 ( .A(n5221), .B(n5220), .C(n5219), .D(n5218), .Y(n5222) );
  OAI22X1TS U3517 ( .A0(n4760), .A1(n3599), .B0(n4764), .B1(n3617), .Y(n5221)
         );
  OAI22X1TS U3518 ( .A0(n4766), .A1(n3640), .B0(n4762), .B1(n3661), .Y(n5220)
         );
  OAI22X1TS U3519 ( .A0(n4768), .A1(n671), .B0(n5231), .B1(n3561), .Y(n5232)
         );
  NOR4XLTS U3520 ( .A(n5230), .B(n5229), .C(n5228), .D(n5227), .Y(n5231) );
  OAI22X1TS U3521 ( .A0(n4774), .A1(n3599), .B0(n4769), .B1(n3609), .Y(n5230)
         );
  OAI22X1TS U3522 ( .A0(n4773), .A1(n3640), .B0(n4771), .B1(n3661), .Y(n5229)
         );
  OAI31X1TS U3523 ( .A0(n4843), .A1(n5322), .A2(n5321), .B0(n5320), .Y(n2450)
         );
  OAI221XLTS U3524 ( .A0(n5319), .A1(n5318), .B0(n5317), .B1(n5316), .C0(n4430), .Y(n5320) );
  OAI211X1TS U3525 ( .A0(n3592), .A1(n25), .B0(n4842), .C0(n5310), .Y(n5318)
         );
  OAI221XLTS U3526 ( .A0(n3601), .A1(n33), .B0(n3663), .B1(n19), .C0(n5308), 
        .Y(n5319) );
  OAI211X1TS U3527 ( .A0(n320), .A1(n605), .B0(n5241), .C0(n5240), .Y(n2441)
         );
  AOI22X1TS U3528 ( .A0(n544), .A1(n5239), .B0(n681), .B1(
        destinationAddressOut[13]), .Y(n5241) );
  AOI222XLTS U3529 ( .A0(n446), .A1(n4296), .B0(n637), .B1(n4140), .C0(n625), 
        .C1(destinationAddressIn_WEST[13]), .Y(n5240) );
  NAND4X1TS U3530 ( .A(n5238), .B(n5237), .C(n5236), .D(n5235), .Y(n5239) );
  OAI211X1TS U3531 ( .A0(n311), .A1(n605), .B0(n5248), .C0(n5247), .Y(n2442)
         );
  AOI22X1TS U3532 ( .A0(n545), .A1(n5246), .B0(n681), .B1(
        destinationAddressOut[12]), .Y(n5248) );
  AOI222XLTS U3533 ( .A0(n445), .A1(n4293), .B0(n637), .B1(n4137), .C0(n632), 
        .C1(destinationAddressIn_WEST[12]), .Y(n5247) );
  NAND4X1TS U3534 ( .A(n5245), .B(n5244), .C(n5243), .D(n5242), .Y(n5246) );
  OAI211X1TS U3535 ( .A0(n323), .A1(n605), .B0(n5255), .C0(n5254), .Y(n2443)
         );
  AOI22X1TS U3536 ( .A0(n545), .A1(n5253), .B0(n681), .B1(
        destinationAddressOut[11]), .Y(n5255) );
  AOI222XLTS U3537 ( .A0(n446), .A1(n4290), .B0(n637), .B1(n4134), .C0(n632), 
        .C1(destinationAddressIn_WEST[11]), .Y(n5254) );
  NAND4X1TS U3538 ( .A(n5252), .B(n5251), .C(n5250), .D(n5249), .Y(n5253) );
  OAI211X1TS U3539 ( .A0(n314), .A1(n606), .B0(n5262), .C0(n5261), .Y(n2444)
         );
  AOI22X1TS U3540 ( .A0(n544), .A1(n5260), .B0(n681), .B1(
        destinationAddressOut[10]), .Y(n5262) );
  AOI222XLTS U3541 ( .A0(n445), .A1(n4287), .B0(n637), .B1(n4131), .C0(n627), 
        .C1(destinationAddressIn_WEST[10]), .Y(n5261) );
  NAND4X1TS U3542 ( .A(n5259), .B(n5258), .C(n5257), .D(n5256), .Y(n5260) );
  OAI211X1TS U3543 ( .A0(n317), .A1(n606), .B0(n5269), .C0(n5268), .Y(n2445)
         );
  AOI22X1TS U3544 ( .A0(n545), .A1(n5267), .B0(n682), .B1(
        destinationAddressOut[9]), .Y(n5269) );
  AOI222XLTS U3545 ( .A0(n446), .A1(n4284), .B0(n636), .B1(n4128), .C0(n635), 
        .C1(destinationAddressIn_WEST[9]), .Y(n5268) );
  NAND4X1TS U3546 ( .A(n5266), .B(n5265), .C(n5264), .D(n5263), .Y(n5267) );
  OAI211X1TS U3547 ( .A0(n326), .A1(n606), .B0(n5276), .C0(n5275), .Y(n2446)
         );
  AOI22X1TS U3548 ( .A0(n544), .A1(n5274), .B0(n682), .B1(
        destinationAddressOut[8]), .Y(n5276) );
  AOI222XLTS U3549 ( .A0(n445), .A1(n4281), .B0(n636), .B1(n4125), .C0(n634), 
        .C1(destinationAddressIn_WEST[8]), .Y(n5275) );
  NAND4X1TS U3550 ( .A(n5273), .B(n5272), .C(n5271), .D(n5270), .Y(n5274) );
  OAI211X1TS U3551 ( .A0(n308), .A1(n607), .B0(n5283), .C0(n5282), .Y(n2447)
         );
  AOI22X1TS U3552 ( .A0(n544), .A1(n5281), .B0(n682), .B1(
        destinationAddressOut[7]), .Y(n5283) );
  AOI222XLTS U3553 ( .A0(n446), .A1(n4278), .B0(n636), .B1(n4122), .C0(n633), 
        .C1(destinationAddressIn_WEST[7]), .Y(n5282) );
  NAND4X1TS U3554 ( .A(n5280), .B(n5279), .C(n5278), .D(n5277), .Y(n5281) );
  OAI211X1TS U3555 ( .A0(n305), .A1(n607), .B0(n5293), .C0(n5292), .Y(n2448)
         );
  AOI22X1TS U3556 ( .A0(n545), .A1(n5288), .B0(n682), .B1(
        destinationAddressOut[6]), .Y(n5293) );
  AOI222XLTS U3557 ( .A0(n445), .A1(n4275), .B0(n636), .B1(n4119), .C0(n626), 
        .C1(destinationAddressIn_WEST[6]), .Y(n5292) );
  NAND4X1TS U3558 ( .A(n5287), .B(n5286), .C(n5285), .D(n5284), .Y(n5288) );
  OAI211X1TS U3559 ( .A0(n4237), .A1(n3547), .B0(n4889), .C0(n4888), .Y(n2397)
         );
  AOI22X1TS U3560 ( .A0(n5226), .A1(n452), .B0(n610), .B1(n3923), .Y(n4889) );
  AOI221X1TS U3561 ( .A0(n585), .A1(n4391), .B0(n649), .B1(n4080), .C0(n4887), 
        .Y(n4888) );
  OAI211X1TS U3562 ( .A0(n4234), .A1(n3547), .B0(n4897), .C0(n4896), .Y(n2398)
         );
  AOI22X1TS U3563 ( .A0(n5226), .A1(n454), .B0(n610), .B1(n3920), .Y(n4897) );
  AOI221X1TS U3564 ( .A0(n585), .A1(n4388), .B0(n648), .B1(n4077), .C0(n4895), 
        .Y(n4896) );
  OAI211X1TS U3565 ( .A0(n4231), .A1(n3547), .B0(n4905), .C0(n4904), .Y(n2399)
         );
  AOI22X1TS U3566 ( .A0(n582), .A1(n456), .B0(n610), .B1(n3917), .Y(n4905) );
  AOI221X1TS U3567 ( .A0(n585), .A1(n4385), .B0(n648), .B1(n4074), .C0(n4903), 
        .Y(n4904) );
  OAI211X1TS U3568 ( .A0(n4228), .A1(n3547), .B0(n4913), .C0(n4912), .Y(n2400)
         );
  AOI22X1TS U3569 ( .A0(n583), .A1(n458), .B0(n610), .B1(n3914), .Y(n4913) );
  AOI221X1TS U3570 ( .A0(n585), .A1(n4382), .B0(n651), .B1(n4071), .C0(n4911), 
        .Y(n4912) );
  OAI211X1TS U3571 ( .A0(n4225), .A1(n3557), .B0(n4921), .C0(n4920), .Y(n2401)
         );
  AOI22X1TS U3572 ( .A0(n571), .A1(n460), .B0(n611), .B1(n3911), .Y(n4921) );
  AOI221X1TS U3573 ( .A0(n586), .A1(n4379), .B0(n650), .B1(n4068), .C0(n4919), 
        .Y(n4920) );
  OAI211X1TS U3574 ( .A0(n4222), .A1(n3556), .B0(n4929), .C0(n4928), .Y(n2402)
         );
  AOI22X1TS U3575 ( .A0(n571), .A1(n462), .B0(n611), .B1(n3908), .Y(n4929) );
  AOI221X1TS U3576 ( .A0(n586), .A1(n4376), .B0(n5290), .B1(n4065), .C0(n4927), 
        .Y(n4928) );
  OAI211X1TS U3577 ( .A0(n4219), .A1(n3555), .B0(n4937), .C0(n4936), .Y(n2403)
         );
  AOI22X1TS U3578 ( .A0(n571), .A1(n464), .B0(n611), .B1(n3905), .Y(n4937) );
  AOI221X1TS U3579 ( .A0(n586), .A1(n4373), .B0(n5290), .B1(n4062), .C0(n4935), 
        .Y(n4936) );
  OAI211X1TS U3580 ( .A0(n4216), .A1(n3558), .B0(n4945), .C0(n4944), .Y(n2404)
         );
  AOI22X1TS U3581 ( .A0(n571), .A1(n466), .B0(n611), .B1(n3902), .Y(n4945) );
  AOI221X1TS U3582 ( .A0(n586), .A1(n4370), .B0(n5290), .B1(n4059), .C0(n4943), 
        .Y(n4944) );
  OAI211X1TS U3583 ( .A0(n4213), .A1(n3555), .B0(n4953), .C0(n4952), .Y(n2405)
         );
  AOI22X1TS U3584 ( .A0(n572), .A1(n468), .B0(n632), .B1(n3899), .Y(n4953) );
  AOI221X1TS U3585 ( .A0(n587), .A1(n4367), .B0(n646), .B1(n4056), .C0(n4951), 
        .Y(n4952) );
  OAI211X1TS U3586 ( .A0(n4210), .A1(n3559), .B0(n4961), .C0(n4960), .Y(n2406)
         );
  AOI22X1TS U3587 ( .A0(n572), .A1(n470), .B0(n634), .B1(n3896), .Y(n4961) );
  AOI221X1TS U3588 ( .A0(n587), .A1(n4364), .B0(n647), .B1(n4053), .C0(n4959), 
        .Y(n4960) );
  OAI211X1TS U3589 ( .A0(n4207), .A1(n3557), .B0(n4969), .C0(n4968), .Y(n2407)
         );
  AOI22X1TS U3590 ( .A0(n572), .A1(n472), .B0(n5289), .B1(n3893), .Y(n4969) );
  AOI221X1TS U3591 ( .A0(n587), .A1(n4361), .B0(n650), .B1(n4050), .C0(n4967), 
        .Y(n4968) );
  OAI211X1TS U3592 ( .A0(n4204), .A1(n3556), .B0(n4977), .C0(n4976), .Y(n2408)
         );
  AOI22X1TS U3593 ( .A0(n572), .A1(n474), .B0(n5289), .B1(n3890), .Y(n4977) );
  AOI221X1TS U3594 ( .A0(n587), .A1(n4358), .B0(n646), .B1(n4047), .C0(n4975), 
        .Y(n4976) );
  OAI211X1TS U3595 ( .A0(n4201), .A1(n3558), .B0(n4985), .C0(n4984), .Y(n2409)
         );
  AOI22X1TS U3596 ( .A0(n573), .A1(n476), .B0(n633), .B1(n3887), .Y(n4985) );
  AOI221X1TS U3597 ( .A0(n597), .A1(n4355), .B0(n645), .B1(n4044), .C0(n4983), 
        .Y(n4984) );
  OAI211X1TS U3598 ( .A0(n4198), .A1(n3558), .B0(n4993), .C0(n4992), .Y(n2410)
         );
  AOI22X1TS U3599 ( .A0(n573), .A1(n478), .B0(n625), .B1(n3884), .Y(n4993) );
  AOI221X1TS U3600 ( .A0(n597), .A1(n4352), .B0(n645), .B1(n4041), .C0(n4991), 
        .Y(n4992) );
  OAI211X1TS U3601 ( .A0(n4195), .A1(n3559), .B0(n5001), .C0(n5000), .Y(n2411)
         );
  AOI22X1TS U3602 ( .A0(n573), .A1(n480), .B0(n633), .B1(n3881), .Y(n5001) );
  AOI221X1TS U3603 ( .A0(n597), .A1(n4349), .B0(n645), .B1(n4038), .C0(n4999), 
        .Y(n5000) );
  OAI211X1TS U3604 ( .A0(n4192), .A1(n3560), .B0(n5009), .C0(n5008), .Y(n2412)
         );
  AOI22X1TS U3605 ( .A0(n573), .A1(n482), .B0(n627), .B1(n3878), .Y(n5009) );
  AOI221X1TS U3606 ( .A0(n597), .A1(n4346), .B0(n645), .B1(n4035), .C0(n5007), 
        .Y(n5008) );
  OAI211X1TS U3607 ( .A0(n4189), .A1(n3548), .B0(n5017), .C0(n5016), .Y(n2413)
         );
  AOI22X1TS U3608 ( .A0(n582), .A1(n484), .B0(n612), .B1(n3875), .Y(n5017) );
  AOI221X1TS U3609 ( .A0(n598), .A1(n4343), .B0(n644), .B1(n4032), .C0(n5015), 
        .Y(n5016) );
  OAI211X1TS U3610 ( .A0(n4186), .A1(n3548), .B0(n5025), .C0(n5024), .Y(n2414)
         );
  AOI22X1TS U3611 ( .A0(n581), .A1(n486), .B0(n612), .B1(n3872), .Y(n5025) );
  AOI221X1TS U3612 ( .A0(n598), .A1(n4340), .B0(n644), .B1(n4029), .C0(n5023), 
        .Y(n5024) );
  OAI211X1TS U3613 ( .A0(n4183), .A1(n3548), .B0(n5033), .C0(n5032), .Y(n2415)
         );
  AOI22X1TS U3614 ( .A0(n580), .A1(n488), .B0(n612), .B1(n3869), .Y(n5033) );
  AOI221X1TS U3615 ( .A0(n598), .A1(n4337), .B0(n644), .B1(n4026), .C0(n5031), 
        .Y(n5032) );
  OAI211X1TS U3616 ( .A0(n4180), .A1(n3548), .B0(n5041), .C0(n5040), .Y(n2416)
         );
  AOI22X1TS U3617 ( .A0(n581), .A1(n490), .B0(n612), .B1(n3866), .Y(n5041) );
  AOI221X1TS U3618 ( .A0(n598), .A1(n4334), .B0(n644), .B1(n4023), .C0(n5039), 
        .Y(n5040) );
  OAI211X1TS U3619 ( .A0(n4177), .A1(n3549), .B0(n5049), .C0(n5048), .Y(n2417)
         );
  AOI22X1TS U3620 ( .A0(n574), .A1(n492), .B0(n613), .B1(n3863), .Y(n5049) );
  AOI221X1TS U3621 ( .A0(n599), .A1(n4331), .B0(n643), .B1(n4020), .C0(n5047), 
        .Y(n5048) );
  OAI211X1TS U3622 ( .A0(n4174), .A1(n3549), .B0(n5057), .C0(n5056), .Y(n2418)
         );
  AOI22X1TS U3623 ( .A0(n574), .A1(n494), .B0(n613), .B1(n3860), .Y(n5057) );
  AOI221X1TS U3624 ( .A0(n599), .A1(n4328), .B0(n643), .B1(n4017), .C0(n5055), 
        .Y(n5056) );
  OAI211X1TS U3625 ( .A0(n4171), .A1(n3549), .B0(n5065), .C0(n5064), .Y(n2419)
         );
  AOI22X1TS U3626 ( .A0(n574), .A1(n496), .B0(n613), .B1(n3857), .Y(n5065) );
  AOI221X1TS U3627 ( .A0(n599), .A1(n4325), .B0(n643), .B1(n4014), .C0(n5063), 
        .Y(n5064) );
  OAI211X1TS U3628 ( .A0(n4168), .A1(n3549), .B0(n5073), .C0(n5072), .Y(n2420)
         );
  AOI22X1TS U3629 ( .A0(n574), .A1(n503), .B0(n613), .B1(n3854), .Y(n5073) );
  AOI221X1TS U3630 ( .A0(n599), .A1(n4322), .B0(n643), .B1(n4011), .C0(n5071), 
        .Y(n5072) );
  OAI211X1TS U3631 ( .A0(n4165), .A1(n3550), .B0(n5081), .C0(n5080), .Y(n2421)
         );
  AOI22X1TS U3632 ( .A0(n575), .A1(n507), .B0(n614), .B1(n3851), .Y(n5081) );
  AOI221X1TS U3633 ( .A0(n600), .A1(n4319), .B0(n642), .B1(n4008), .C0(n5079), 
        .Y(n5080) );
  OAI211X1TS U3634 ( .A0(n4162), .A1(n3550), .B0(n5089), .C0(n5088), .Y(n2422)
         );
  AOI22X1TS U3635 ( .A0(n575), .A1(n509), .B0(n614), .B1(n3848), .Y(n5089) );
  AOI221X1TS U3636 ( .A0(n600), .A1(n4316), .B0(n642), .B1(n4005), .C0(n5087), 
        .Y(n5088) );
  OAI211X1TS U3637 ( .A0(n4159), .A1(n3550), .B0(n5097), .C0(n5096), .Y(n2423)
         );
  AOI22X1TS U3638 ( .A0(n575), .A1(n511), .B0(n614), .B1(n3845), .Y(n5097) );
  AOI221X1TS U3639 ( .A0(n600), .A1(n4313), .B0(n642), .B1(n4002), .C0(n5095), 
        .Y(n5096) );
  OAI211X1TS U3640 ( .A0(n4156), .A1(n3550), .B0(n5105), .C0(n5104), .Y(n2424)
         );
  AOI22X1TS U3641 ( .A0(n575), .A1(n514), .B0(n614), .B1(n3842), .Y(n5105) );
  AOI221X1TS U3642 ( .A0(n600), .A1(n4310), .B0(n642), .B1(n3999), .C0(n5103), 
        .Y(n5104) );
  OAI211X1TS U3643 ( .A0(n4153), .A1(n3551), .B0(n5113), .C0(n5112), .Y(n2425)
         );
  AOI22X1TS U3644 ( .A0(n576), .A1(n516), .B0(n621), .B1(n3839), .Y(n5113) );
  AOI221X1TS U3645 ( .A0(n601), .A1(n4307), .B0(n641), .B1(n3996), .C0(n5111), 
        .Y(n5112) );
  OAI211X1TS U3646 ( .A0(n4150), .A1(n3551), .B0(n5121), .C0(n5120), .Y(n2426)
         );
  AOI22X1TS U3647 ( .A0(n576), .A1(n531), .B0(n621), .B1(n3836), .Y(n5121) );
  AOI221X1TS U3648 ( .A0(n601), .A1(n4304), .B0(n641), .B1(n3993), .C0(n5119), 
        .Y(n5120) );
  OAI211X1TS U3649 ( .A0(n4147), .A1(n3551), .B0(n5129), .C0(n5128), .Y(n2427)
         );
  AOI22X1TS U3650 ( .A0(n576), .A1(n537), .B0(n621), .B1(n3833), .Y(n5129) );
  AOI221X1TS U3651 ( .A0(n601), .A1(n4301), .B0(n641), .B1(n3990), .C0(n5127), 
        .Y(n5128) );
  OAI211X1TS U3652 ( .A0(n4144), .A1(n3551), .B0(n5137), .C0(n5136), .Y(n2428)
         );
  AOI22X1TS U3653 ( .A0(n576), .A1(n543), .B0(n621), .B1(n3830), .Y(n5137) );
  AOI221X1TS U3654 ( .A0(n601), .A1(n4298), .B0(n641), .B1(n3987), .C0(n5135), 
        .Y(n5136) );
  OAI211X1TS U3655 ( .A0(n4255), .A1(n3552), .B0(n5145), .C0(n5144), .Y(n2429)
         );
  AOI22X1TS U3656 ( .A0(n577), .A1(n159), .B0(n622), .B1(n3941), .Y(n5145) );
  AOI221X1TS U3657 ( .A0(n602), .A1(n4409), .B0(n640), .B1(n4098), .C0(n5143), 
        .Y(n5144) );
  OAI211X1TS U3658 ( .A0(n4252), .A1(n3552), .B0(n5153), .C0(n5152), .Y(n2430)
         );
  AOI22X1TS U3659 ( .A0(n577), .A1(n186), .B0(n622), .B1(n3938), .Y(n5153) );
  AOI221X1TS U3660 ( .A0(n602), .A1(n4406), .B0(n640), .B1(n4095), .C0(n5151), 
        .Y(n5152) );
  OAI211X1TS U3661 ( .A0(n4246), .A1(n3552), .B0(n5169), .C0(n5168), .Y(n2432)
         );
  AOI22X1TS U3662 ( .A0(n577), .A1(n176), .B0(n622), .B1(n3932), .Y(n5169) );
  AOI221X1TS U3663 ( .A0(n602), .A1(n4400), .B0(n640), .B1(n4089), .C0(n5167), 
        .Y(n5168) );
  OAI211X1TS U3664 ( .A0(n4243), .A1(n3553), .B0(n5177), .C0(n5176), .Y(n2433)
         );
  AOI22X1TS U3665 ( .A0(n578), .A1(n171), .B0(n623), .B1(n3929), .Y(n5177) );
  AOI221X1TS U3666 ( .A0(n603), .A1(n4397), .B0(n639), .B1(n4086), .C0(n5175), 
        .Y(n5176) );
  OAI211X1TS U3667 ( .A0(n4273), .A1(n3553), .B0(n5193), .C0(n5192), .Y(n2435)
         );
  AOI22X1TS U3668 ( .A0(n578), .A1(n192), .B0(n623), .B1(n3959), .Y(n5193) );
  AOI221X1TS U3669 ( .A0(n603), .A1(n4427), .B0(n639), .B1(n4116), .C0(n5191), 
        .Y(n5192) );
  OAI211X1TS U3670 ( .A0(n4270), .A1(n3553), .B0(n5201), .C0(n5200), .Y(n2436)
         );
  AOI22X1TS U3671 ( .A0(n578), .A1(n187), .B0(n623), .B1(n3956), .Y(n5201) );
  AOI221X1TS U3672 ( .A0(n603), .A1(n4424), .B0(n639), .B1(n4113), .C0(n5199), 
        .Y(n5200) );
  OAI211X1TS U3673 ( .A0(n4267), .A1(n3554), .B0(n5209), .C0(n5208), .Y(n2437)
         );
  AOI22X1TS U3674 ( .A0(n579), .A1(n181), .B0(n624), .B1(n3953), .Y(n5209) );
  AOI221X1TS U3675 ( .A0(n604), .A1(n4421), .B0(n638), .B1(n4110), .C0(n5207), 
        .Y(n5208) );
  OAI211X1TS U3676 ( .A0(n4264), .A1(n3554), .B0(n5217), .C0(n5216), .Y(n2438)
         );
  AOI22X1TS U3677 ( .A0(n579), .A1(n177), .B0(n624), .B1(n3950), .Y(n5217) );
  AOI221X1TS U3678 ( .A0(n604), .A1(n4418), .B0(n638), .B1(n4107), .C0(n5215), 
        .Y(n5216) );
  OAI211X1TS U3679 ( .A0(n4261), .A1(n3554), .B0(n5225), .C0(n5224), .Y(n2439)
         );
  AOI22X1TS U3680 ( .A0(n579), .A1(n172), .B0(n624), .B1(n3947), .Y(n5225) );
  AOI221X1TS U3681 ( .A0(n604), .A1(n4415), .B0(n638), .B1(n4104), .C0(n5223), 
        .Y(n5224) );
  OAI211X1TS U3682 ( .A0(n4258), .A1(n3554), .B0(n5234), .C0(n5233), .Y(n2440)
         );
  AOI22X1TS U3683 ( .A0(n579), .A1(n167), .B0(n624), .B1(n3944), .Y(n5234) );
  AOI221X1TS U3684 ( .A0(n604), .A1(n4412), .B0(n638), .B1(n4101), .C0(n5232), 
        .Y(n5233) );
  OAI211X1TS U3685 ( .A0(n4249), .A1(n3552), .B0(n5161), .C0(n5160), .Y(n2431)
         );
  AOI22X1TS U3686 ( .A0(n577), .A1(n182), .B0(n622), .B1(n3935), .Y(n5161) );
  AOI221X1TS U3687 ( .A0(n602), .A1(n4403), .B0(n640), .B1(n4092), .C0(n5159), 
        .Y(n5160) );
  OAI211X1TS U3688 ( .A0(n4240), .A1(n3553), .B0(n5185), .C0(n5184), .Y(n2434)
         );
  AOI22X1TS U3689 ( .A0(n578), .A1(n168), .B0(n623), .B1(n3926), .Y(n5185) );
  AOI221X1TS U3690 ( .A0(n603), .A1(n4394), .B0(n639), .B1(n4083), .C0(n5183), 
        .Y(n5184) );
  NOR2X1TS U3691 ( .A(reset), .B(n4842), .Y(n5303) );
  INVX2TS U3692 ( .A(readIn_SOUTH), .Y(n6242) );
  INVX2TS U3693 ( .A(writeIn_NORTH), .Y(n6244) );
  OAI31X1TS U3694 ( .A0(n4841), .A1(n5322), .A2(n5321), .B0(n5305), .Y(n2449)
         );
  OAI22X1TS U3695 ( .A0(n5304), .A1(n5303), .B0(n5302), .B1(n5301), .Y(n5305)
         );
  AOI31X1TS U3696 ( .A0(n5300), .A1(n5299), .A2(n5298), .B0(reset), .Y(n5304)
         );
  OAI22X1TS U3697 ( .A0(n3826), .A1(n5313), .B0(n3813), .B1(n5315), .Y(n5301)
         );
  OAI22X1TS U3698 ( .A0(n449), .A1(n6278), .B0(n9), .B1(n3566), .Y(n2889) );
  INVX2TS U3699 ( .A(destinationAddressIn_NORTH[7]), .Y(n6245) );
  INVX2TS U3700 ( .A(destinationAddressIn_NORTH[12]), .Y(n6250) );
  INVX2TS U3701 ( .A(destinationAddressIn_NORTH[10]), .Y(n6248) );
  INVX2TS U3702 ( .A(destinationAddressIn_NORTH[9]), .Y(n6247) );
  INVX2TS U3703 ( .A(destinationAddressIn_NORTH[13]), .Y(n6251) );
  INVX2TS U3704 ( .A(destinationAddressIn_NORTH[11]), .Y(n6249) );
  INVX2TS U3705 ( .A(destinationAddressIn_NORTH[8]), .Y(n6246) );
  NOR2X1TS U3706 ( .A(n6227), .B(n6228), .Y(n2883) );
  AOI21X1TS U3707 ( .A0(n348), .A1(n6226), .B0(n10), .Y(n6227) );
  XNOR2X1TS U3708 ( .A(n4852), .B(n6284), .Y(n6231) );
  XNOR2X1TS U3709 ( .A(n258), .B(n568), .Y(n4852) );
  OAI22X1TS U3710 ( .A0(n4438), .A1(n3682), .B0(n4439), .B1(n3581), .Y(n4882)
         );
  OAI22X1TS U3711 ( .A0(n4443), .A1(n3682), .B0(n4448), .B1(n3583), .Y(n4890)
         );
  OAI22X1TS U3712 ( .A0(n4450), .A1(n3682), .B0(n4453), .B1(n3583), .Y(n4898)
         );
  OAI22X1TS U3713 ( .A0(n4461), .A1(n3677), .B0(n4460), .B1(n3583), .Y(n4906)
         );
  OAI22X1TS U3714 ( .A0(n4475), .A1(n3682), .B0(n4468), .B1(n3583), .Y(n4914)
         );
  OAI22X1TS U3715 ( .A0(n4479), .A1(n3679), .B0(n4484), .B1(n3582), .Y(n4922)
         );
  OAI22X1TS U3716 ( .A0(n4486), .A1(n3677), .B0(n4491), .B1(n3582), .Y(n4930)
         );
  OAI22X1TS U3717 ( .A0(n4501), .A1(n3680), .B0(n4496), .B1(n3582), .Y(n4938)
         );
  OAI22X1TS U3718 ( .A0(n4508), .A1(n3681), .B0(n4505), .B1(n3582), .Y(n4946)
         );
  OAI22X1TS U3719 ( .A0(n4519), .A1(n3681), .B0(n4517), .B1(n3590), .Y(n4954)
         );
  OAI22X1TS U3720 ( .A0(n4522), .A1(n3681), .B0(n4523), .B1(n3590), .Y(n4962)
         );
  OAI22X1TS U3721 ( .A0(n4535), .A1(n3683), .B0(n4533), .B1(n3589), .Y(n4970)
         );
  OAI22X1TS U3722 ( .A0(n4540), .A1(n3678), .B0(n4544), .B1(n3588), .Y(n4978)
         );
  OAI22X1TS U3723 ( .A0(n4553), .A1(n3678), .B0(n4556), .B1(n3589), .Y(n4986)
         );
  OAI22X1TS U3724 ( .A0(n4562), .A1(n3681), .B0(n4559), .B1(n3591), .Y(n4994)
         );
  OAI22X1TS U3725 ( .A0(n4573), .A1(n3684), .B0(n4574), .B1(n3591), .Y(n5002)
         );
  OAI22X1TS U3726 ( .A0(n4578), .A1(n3670), .B0(n4581), .B1(n3592), .Y(n5010)
         );
  OAI22X1TS U3727 ( .A0(n4585), .A1(n3670), .B0(n4588), .B1(n3586), .Y(n5018)
         );
  OAI22X1TS U3728 ( .A0(n4596), .A1(n3670), .B0(n4601), .B1(n3586), .Y(n5026)
         );
  OAI22X1TS U3729 ( .A0(n4603), .A1(n3670), .B0(n4610), .B1(n3586), .Y(n5034)
         );
  OAI22X1TS U3730 ( .A0(n4618), .A1(n3671), .B0(n4613), .B1(n6279), .Y(n5042)
         );
  OAI22X1TS U3731 ( .A0(n4626), .A1(n3671), .B0(n4627), .B1(n3581), .Y(n5050)
         );
  OAI22X1TS U3732 ( .A0(n4630), .A1(n3671), .B0(n4631), .B1(n3581), .Y(n5058)
         );
  OAI22X1TS U3733 ( .A0(n4643), .A1(n3671), .B0(n4641), .B1(n3581), .Y(n5066)
         );
  OAI22X1TS U3734 ( .A0(n4648), .A1(n3672), .B0(n4655), .B1(n3580), .Y(n5074)
         );
  OAI22X1TS U3735 ( .A0(n4663), .A1(n3672), .B0(n4658), .B1(n3580), .Y(n5082)
         );
  OAI22X1TS U3736 ( .A0(n4670), .A1(n3672), .B0(n4666), .B1(n3580), .Y(n5090)
         );
  OAI22X1TS U3737 ( .A0(n4677), .A1(n3672), .B0(n4682), .B1(n3580), .Y(n5098)
         );
  OAI22X1TS U3738 ( .A0(n4684), .A1(n3673), .B0(n4687), .B1(n3579), .Y(n5106)
         );
  OAI22X1TS U3739 ( .A0(n4697), .A1(n3673), .B0(n4693), .B1(n3579), .Y(n5114)
         );
  OAI22X1TS U3740 ( .A0(n4709), .A1(n3673), .B0(n4705), .B1(n3579), .Y(n5122)
         );
  OAI22X1TS U3741 ( .A0(n4713), .A1(n3673), .B0(n4717), .B1(n3579), .Y(n5130)
         );
  OAI22X1TS U3742 ( .A0(n4727), .A1(n3674), .B0(n4725), .B1(n3578), .Y(n5186)
         );
  OAI22X1TS U3743 ( .A0(n4740), .A1(n3674), .B0(n4734), .B1(n3578), .Y(n5194)
         );
  OAI22X1TS U3744 ( .A0(n4749), .A1(n3674), .B0(n4745), .B1(n3578), .Y(n5202)
         );
  OAI22X1TS U3745 ( .A0(n4757), .A1(n3674), .B0(n4758), .B1(n3577), .Y(n5210)
         );
  OAI22X1TS U3746 ( .A0(n4763), .A1(n3675), .B0(n4767), .B1(n3578), .Y(n5218)
         );
  OAI22X1TS U3747 ( .A0(n4770), .A1(n3675), .B0(n4776), .B1(n3577), .Y(n5227)
         );
  OAI22X1TS U3748 ( .A0(n4436), .A1(n657), .B0(n4437), .B1(n3624), .Y(n4883)
         );
  OAI22X1TS U3749 ( .A0(n4444), .A1(n659), .B0(n4442), .B1(n3636), .Y(n4891)
         );
  OAI22X1TS U3750 ( .A0(n4455), .A1(n661), .B0(n4451), .B1(n3632), .Y(n4899)
         );
  OAI22X1TS U3751 ( .A0(n4466), .A1(n661), .B0(n4464), .B1(n3632), .Y(n4907)
         );
  OAI22X1TS U3752 ( .A0(n4469), .A1(n665), .B0(n4473), .B1(n3632), .Y(n4915)
         );
  OAI22X1TS U3753 ( .A0(n4478), .A1(n659), .B0(n4480), .B1(n3632), .Y(n4923)
         );
  OAI22X1TS U3754 ( .A0(n4493), .A1(n662), .B0(n4489), .B1(n3637), .Y(n4931)
         );
  OAI22X1TS U3755 ( .A0(n4500), .A1(n662), .B0(n4498), .B1(n3635), .Y(n4939)
         );
  OAI22X1TS U3756 ( .A0(n4507), .A1(n662), .B0(n4509), .B1(n3634), .Y(n4947)
         );
  OAI22X1TS U3757 ( .A0(n4518), .A1(n661), .B0(n4514), .B1(n3636), .Y(n4955)
         );
  OAI22X1TS U3758 ( .A0(n4525), .A1(n662), .B0(n4529), .B1(n3634), .Y(n4963)
         );
  OAI22X1TS U3759 ( .A0(n4532), .A1(n663), .B0(n4534), .B1(n3638), .Y(n4971)
         );
  OAI22X1TS U3760 ( .A0(n4545), .A1(n664), .B0(n4547), .B1(n3639), .Y(n4979)
         );
  OAI22X1TS U3761 ( .A0(n4552), .A1(n665), .B0(n4550), .B1(n3639), .Y(n4987)
         );
  OAI22X1TS U3762 ( .A0(n4563), .A1(n660), .B0(n4561), .B1(n3631), .Y(n4995)
         );
  OAI22X1TS U3763 ( .A0(n4571), .A1(n667), .B0(n4572), .B1(n3631), .Y(n5003)
         );
  OAI22X1TS U3764 ( .A0(n4576), .A1(n666), .B0(n4577), .B1(n3631), .Y(n5011)
         );
  OAI22X1TS U3765 ( .A0(n4586), .A1(n667), .B0(n4592), .B1(n3631), .Y(n5019)
         );
  OAI22X1TS U3766 ( .A0(n4599), .A1(n668), .B0(n4595), .B1(n3630), .Y(n5027)
         );
  OAI22X1TS U3767 ( .A0(n4608), .A1(n668), .B0(n4604), .B1(n3630), .Y(n5035)
         );
  OAI22X1TS U3768 ( .A0(n4614), .A1(n668), .B0(n4615), .B1(n3630), .Y(n5043)
         );
  OAI22X1TS U3769 ( .A0(n4622), .A1(n660), .B0(n4628), .B1(n3630), .Y(n5051)
         );
  OAI22X1TS U3770 ( .A0(n4633), .A1(n657), .B0(n4637), .B1(n3629), .Y(n5059)
         );
  OAI22X1TS U3771 ( .A0(n4644), .A1(n657), .B0(n4642), .B1(n3629), .Y(n5067)
         );
  OAI22X1TS U3772 ( .A0(n4653), .A1(n657), .B0(n4649), .B1(n3629), .Y(n5075)
         );
  OAI22X1TS U3773 ( .A0(n4660), .A1(n656), .B0(n4664), .B1(n3628), .Y(n5083)
         );
  OAI22X1TS U3774 ( .A0(n4673), .A1(n656), .B0(n4667), .B1(n3628), .Y(n5091)
         );
  OAI22X1TS U3775 ( .A0(n4680), .A1(n656), .B0(n4676), .B1(n3628), .Y(n5099)
         );
  OAI22X1TS U3776 ( .A0(n4691), .A1(n656), .B0(n4689), .B1(n3628), .Y(n5107)
         );
  OAI22X1TS U3777 ( .A0(n4696), .A1(n655), .B0(n4694), .B1(n3627), .Y(n5115)
         );
  OAI22X1TS U3778 ( .A0(n4706), .A1(n655), .B0(n4707), .B1(n3627), .Y(n5123)
         );
  OAI22X1TS U3779 ( .A0(n4718), .A1(n655), .B0(n4712), .B1(n3627), .Y(n5131)
         );
  OAI22X1TS U3780 ( .A0(n4729), .A1(n653), .B0(n4731), .B1(n3625), .Y(n5187)
         );
  OAI22X1TS U3781 ( .A0(n4738), .A1(n653), .B0(n4733), .B1(n3625), .Y(n5195)
         );
  OAI22X1TS U3782 ( .A0(n4747), .A1(n653), .B0(n4743), .B1(n3625), .Y(n5203)
         );
  OAI22X1TS U3783 ( .A0(n4756), .A1(n652), .B0(n4754), .B1(n3624), .Y(n5211)
         );
  OAI22X1TS U3784 ( .A0(n4765), .A1(n652), .B0(n4761), .B1(n3624), .Y(n5219)
         );
  OAI22X1TS U3785 ( .A0(n4772), .A1(n652), .B0(n4775), .B1(n3624), .Y(n5228)
         );
  NOR3X1TS U3786 ( .A(n9), .B(n258), .C(n193), .Y(n5307) );
  NOR3X1TS U3787 ( .A(n10), .B(n257), .C(n6278), .Y(n5297) );
  NAND3X1TS U3788 ( .A(n349), .B(n443), .C(n8), .Y(n5309) );
  AOI2BB2X1TS U3789 ( .B0(readOutbuffer[3]), .B1(n293), .A0N(n32), .A1N(n661), 
        .Y(n5310) );
  AOI222XLTS U3790 ( .A0(readOutbuffer[4]), .A1(n5307), .B0(readOutbuffer[7]), 
        .B1(n5306), .C0(readOutbuffer[2]), .C1(n239), .Y(n5308) );
  AOI221X1TS U3791 ( .A0(n5297), .A1(writeOutbuffer[1]), .B0(n239), .B1(
        writeOutbuffer[2]), .C0(n5296), .Y(n5298) );
  OAI22X1TS U3792 ( .A0(n6271), .A1(n652), .B0(n24), .B1(n3629), .Y(n5296) );
  OA22X1TS U3793 ( .A0(n3584), .A1(n4778), .B0(n3675), .B1(n4777), .Y(n5238)
         );
  OA22X1TS U3794 ( .A0(n3584), .A1(n4786), .B0(n3675), .B1(n4791), .Y(n5245)
         );
  OA22X1TS U3795 ( .A0(n3584), .A1(n4796), .B0(n3676), .B1(n4800), .Y(n5252)
         );
  OA22X1TS U3796 ( .A0(n3584), .A1(n4802), .B0(n3676), .B1(n4805), .Y(n5259)
         );
  OA22X1TS U3797 ( .A0(n3585), .A1(n4814), .B0(n3676), .B1(n4816), .Y(n5266)
         );
  OA22X1TS U3798 ( .A0(n3585), .A1(n4818), .B0(n3676), .B1(n4819), .Y(n5273)
         );
  OA22X1TS U3799 ( .A0(n3585), .A1(n4826), .B0(n3677), .B1(n4832), .Y(n5280)
         );
  OA22X1TS U3800 ( .A0(n3585), .A1(n4838), .B0(n3677), .B1(n4839), .Y(n5287)
         );
  OA22X1TS U3801 ( .A0(n3614), .A1(n4783), .B0(n3599), .B1(n4784), .Y(n5235)
         );
  OA22X1TS U3802 ( .A0(n3614), .A1(n4787), .B0(n3599), .B1(n4785), .Y(n5242)
         );
  OA22X1TS U3803 ( .A0(n3614), .A1(n4793), .B0(n3600), .B1(n4797), .Y(n5249)
         );
  OA22X1TS U3804 ( .A0(n3614), .A1(n4803), .B0(n3600), .B1(n4806), .Y(n5256)
         );
  OA22X1TS U3805 ( .A0(n3615), .A1(n4815), .B0(n3600), .B1(n4811), .Y(n5263)
         );
  OA22X1TS U3806 ( .A0(n3615), .A1(n4821), .B0(n3600), .B1(n4817), .Y(n5270)
         );
  OA22X1TS U3807 ( .A0(n3615), .A1(n4825), .B0(n3601), .B1(n4827), .Y(n5277)
         );
  OA22X1TS U3808 ( .A0(n3615), .A1(n4837), .B0(n3601), .B1(n4840), .Y(n5284)
         );
  OA22X1TS U3809 ( .A0(n3637), .A1(n4780), .B0(n663), .B1(n4782), .Y(n5237) );
  OA22X1TS U3810 ( .A0(n3635), .A1(n4790), .B0(n658), .B1(n4792), .Y(n5244) );
  OA22X1TS U3811 ( .A0(n3634), .A1(n4794), .B0(n664), .B1(n4798), .Y(n5251) );
  AOI2BB2X1TS U3812 ( .B0(n5306), .B1(n567), .A0N(n659), .A1N(n4808), .Y(n5258) );
  OA22X1TS U3813 ( .A0(n3633), .A1(n4813), .B0(n658), .B1(n4812), .Y(n5265) );
  OA22X1TS U3814 ( .A0(n3633), .A1(n4820), .B0(n658), .B1(n4822), .Y(n5272) );
  OA22X1TS U3815 ( .A0(n3633), .A1(n4830), .B0(n658), .B1(n4828), .Y(n5279) );
  OA22X1TS U3816 ( .A0(n3633), .A1(n4836), .B0(n659), .B1(n4834), .Y(n5286) );
  OA22X1TS U3817 ( .A0(n3661), .A1(n4779), .B0(n3649), .B1(n4781), .Y(n5236)
         );
  OA22X1TS U3818 ( .A0(n3661), .A1(n4789), .B0(n3650), .B1(n4788), .Y(n5243)
         );
  OA22X1TS U3819 ( .A0(n3662), .A1(n4799), .B0(n3654), .B1(n4795), .Y(n5250)
         );
  OA22X1TS U3820 ( .A0(n3662), .A1(n4801), .B0(n3651), .B1(n4807), .Y(n5257)
         );
  OA22X1TS U3821 ( .A0(n3662), .A1(n4809), .B0(n3652), .B1(n4810), .Y(n5264)
         );
  OA22X1TS U3822 ( .A0(n3662), .A1(n4823), .B0(n3650), .B1(n4824), .Y(n5271)
         );
  OA22X1TS U3823 ( .A0(n3663), .A1(n4829), .B0(n3650), .B1(n4831), .Y(n5278)
         );
  OA22X1TS U3824 ( .A0(n3663), .A1(n4833), .B0(n3653), .B1(n4835), .Y(n5285)
         );
  AOI22X1TS U3825 ( .A0(n450), .A1(writeOutbuffer[6]), .B0(writeOutbuffer[3]), 
        .B1(n241), .Y(n5300) );
  AOI22X1TS U3826 ( .A0(n5307), .A1(writeOutbuffer[4]), .B0(n288), .B1(
        writeOutbuffer[0]), .Y(n5299) );
  AOI21X1TS U3827 ( .A0(n3827), .A1(n5534), .B0(n5533), .Y(n5535) );
  AOI21XLTS U3828 ( .A0(n3815), .A1(n6298), .B0(n5538), .Y(n5545) );
  AOI32XLTS U3829 ( .A0(n5543), .A1(n5542), .A2(n3820), .B0(n5541), .B1(n5540), 
        .Y(n5544) );
  AOI21XLTS U3830 ( .A0(n3827), .A1(n220), .B0(n6310), .Y(n5525) );
  OAI221XLTS U3831 ( .A0(n334), .A1(n301), .B0(n5575), .B1(n156), .C0(n5574), 
        .Y(n2571) );
  OAI221XLTS U3832 ( .A0(n333), .A1(n305), .B0(n4840), .B1(n439), .C0(n5341), 
        .Y(n2458) );
  OAI221XLTS U3833 ( .A0(n334), .A1(n308), .B0(n4827), .B1(n438), .C0(n5340), 
        .Y(n2457) );
  OAI221XLTS U3834 ( .A0(n5576), .A1(n326), .B0(n4817), .B1(n439), .C0(n5339), 
        .Y(n2456) );
  OAI221XLTS U3835 ( .A0(n334), .A1(n317), .B0(n4811), .B1(n438), .C0(n5338), 
        .Y(n2455) );
  OAI221XLTS U3836 ( .A0(n5576), .A1(n314), .B0(n4806), .B1(n439), .C0(n5337), 
        .Y(n2454) );
  OAI221XLTS U3837 ( .A0(n334), .A1(n323), .B0(n4797), .B1(n438), .C0(n5336), 
        .Y(n2453) );
  OAI221XLTS U3838 ( .A0(n333), .A1(n311), .B0(n4785), .B1(n439), .C0(n5335), 
        .Y(n2452) );
  OAI221XLTS U3839 ( .A0(n333), .A1(n320), .B0(n4784), .B1(n438), .C0(n5334), 
        .Y(n2451) );
  AOI32XLTS U3840 ( .A0(n224), .A1(n5551), .A2(n5550), .B0(n3348), .B1(n148), 
        .Y(n2567) );
  AOI32XLTS U3841 ( .A0(n218), .A1(n5536), .A2(n5535), .B0(n259), .B1(n150), 
        .Y(n2565) );
  OAI221XLTS U3842 ( .A0(n338), .A1(n6244), .B0(n297), .B1(n154), .C0(n5579), 
        .Y(n2573) );
  OAI221XLTS U3843 ( .A0(n339), .A1(n303), .B0(n4839), .B1(n5580), .C0(n5386), 
        .Y(n2486) );
  OAI221XLTS U3844 ( .A0(n338), .A1(n6245), .B0(n4832), .B1(n290), .C0(n5385), 
        .Y(n2485) );
  OAI221XLTS U3845 ( .A0(n339), .A1(n6246), .B0(n4819), .B1(n5580), .C0(n5384), 
        .Y(n2484) );
  OAI221XLTS U3846 ( .A0(n338), .A1(n6247), .B0(n4816), .B1(n433), .C0(n5383), 
        .Y(n2483) );
  OAI221XLTS U3847 ( .A0(n339), .A1(n6248), .B0(n4805), .B1(n5580), .C0(n5382), 
        .Y(n2482) );
  OAI221XLTS U3848 ( .A0(n338), .A1(n6249), .B0(n4800), .B1(n290), .C0(n5381), 
        .Y(n2481) );
  OAI221XLTS U3849 ( .A0(n339), .A1(n6250), .B0(n4791), .B1(n433), .C0(n5380), 
        .Y(n2480) );
  OAI221XLTS U3850 ( .A0(n5581), .A1(n6251), .B0(n4777), .B1(n433), .C0(n5379), 
        .Y(n2479) );
  NOR3BX1TS U3851 ( .AN(n5537), .B(n5531), .C(n435), .Y(n6143) );
endmodule


module outputPortArbiter_2 ( clk, reset, selectBit_NORTH, 
        destinationAddressIn_NORTH, requesterAddressIn_NORTH, readIn_NORTH, 
        writeIn_NORTH, dataIn_NORTH, selectBit_SOUTH, 
        destinationAddressIn_SOUTH, requesterAddressIn_SOUTH, readIn_SOUTH, 
        writeIn_SOUTH, dataIn_SOUTH, selectBit_EAST, destinationAddressIn_EAST, 
        requesterAddressIn_EAST, readIn_EAST, writeIn_EAST, dataIn_EAST, 
        selectBit_WEST, destinationAddressIn_WEST, requesterAddressIn_WEST, 
        readIn_WEST, writeIn_WEST, dataIn_WEST, readReady, 
        readRequesterAddress, cacheDataOut, destinationAddressOut, 
        requesterAddressOut, readOut, writeOut, dataOut );
  input [13:0] destinationAddressIn_NORTH;
  input [5:0] requesterAddressIn_NORTH;
  input [31:0] dataIn_NORTH;
  input [13:0] destinationAddressIn_SOUTH;
  input [5:0] requesterAddressIn_SOUTH;
  input [31:0] dataIn_SOUTH;
  input [13:0] destinationAddressIn_EAST;
  input [5:0] requesterAddressIn_EAST;
  input [31:0] dataIn_EAST;
  input [13:0] destinationAddressIn_WEST;
  input [5:0] requesterAddressIn_WEST;
  input [31:0] dataIn_WEST;
  input [5:0] readRequesterAddress;
  input [31:0] cacheDataOut;
  output [13:0] destinationAddressOut;
  output [5:0] requesterAddressOut;
  output [31:0] dataOut;
  input clk, reset, selectBit_NORTH, readIn_NORTH, writeIn_NORTH,
         selectBit_SOUTH, readIn_SOUTH, writeIn_SOUTH, selectBit_EAST,
         readIn_EAST, writeIn_EAST, selectBit_WEST, readIn_WEST, writeIn_WEST,
         readReady;
  output readOut, writeOut;
  wire   N4718, n2888, n5327, n2886, n5326, n2889, n2883, n2887, n5323, n2569,
         n2567, n2566, n2578, n2638, n2624, n2617, n2577, n2544, n2541, n2540,
         n2537, n2535, n2703, n2692, n2691, n2689, n2511, n2507, n2731, n2574,
         n2499, n2496, n2493, n2770, n2768, n2764, n2754, n2748, n2746, n2739,
         n2486, n2484, n2482, n2480, n2802, n2834, n2833, n2832, n2829, n2825,
         n2814, n2811, n2807, n2806, n2457, n2455, n2453, n2570, n2565, n2573,
         n2568, n2564, n2563, n2575, n2882, n2881, n2879, n2610, n2609, n2608,
         n2607, n2606, n2605, n2604, n2603, n2602, n2601, n2600, n2599, n2598,
         n2597, n2596, n2595, n2594, n2593, n2592, n2591, n2590, n2589, n2588,
         n2587, n2586, n2585, n2584, n2583, n2582, n2581, n2580, n2579, n2561,
         n2560, n2559, n2557, n2556, n2555, n2554, n2552, n2551, n2550, n2549,
         n2642, n2640, n2639, n2637, n2635, n2634, n2633, n2631, n2628, n2627,
         n2626, n2625, n2623, n2620, n2618, n2616, n2615, n2614, n2612, n2611,
         n2870, n2869, n2868, n2867, n2866, n2865, n2674, n2672, n2671, n2670,
         n2669, n2668, n2667, n2666, n2665, n2664, n2662, n2661, n2660, n2657,
         n2656, n2655, n2654, n2653, n2652, n2651, n2650, n2649, n2648, n2647,
         n2646, n2645, n2644, n2576, n2534, n2533, n2532, n2531, n2530, n2529,
         n2528, n2527, n2526, n2525, n2524, n2523, n2522, n2521, n2860, n2859,
         n2706, n2705, n2700, n2698, n2696, n2695, n2694, n2690, n2687, n2686,
         n2685, n2684, n2677, n2675, n2736, n2734, n2733, n2725, n2723, n2720,
         n2718, n2715, n2713, n2504, n2498, n2497, n2494, n2850,
         \requesterAddressbuffer[2][2] , n2849, \requesterAddressbuffer[2][3] ,
         n2847, \requesterAddressbuffer[2][5] , n2769, n2760, n2743, n2492,
         n2491, n2489, n2488, n2487, n2485, n2483, n2481, n2846, n2845, n2844,
         n2843, n2842, n2841, n2801, n2799, n2798, n2796, n2795, n2793, n2791,
         n2790, n2789, n2788, n2787, n2786, n2785, n2784, n2781, n2779, n2778,
         n2777, n2776, n2774, n2773, n2772, n2771, n2572, n2478, n2477, n2476,
         n2475, n2474, n2473, n2472, n2471, n2470, n2469, n2468, n2467, n2466,
         n2465, n2840, \requesterAddressbuffer[0][0] , n2839,
         \requesterAddressbuffer[0][1] , n2838, \requesterAddressbuffer[0][2] ,
         n2836, \requesterAddressbuffer[0][4] , n2571, n2464, n2460, n2458,
         n2454, n2451, n2880, n2878, n2877, n2562, n2558, n2553, n2876,
         \requesterAddressbuffer[6][0] , n2875, \requesterAddressbuffer[6][1] ,
         n2874, \requesterAddressbuffer[6][2] , n2873,
         \requesterAddressbuffer[6][3] , n2872, \requesterAddressbuffer[6][4] ,
         n2871, \requesterAddressbuffer[6][5] , n2641, n2636, n2632, n2630,
         n2629, n2622, n2621, n2619, n2613, n2548, n2547, n2546, n2545, n2543,
         n2542, n2539, n2538, n2536, n2673, n2663, n2659, n2658, n2643, n2864,
         n2863, n2862, n2861, n2704, n2702, n2701, n2699, n2697, n2693, n2688,
         n2683, n2682, n2681, n2680, n2679, n2678, n2676, n2520, n2519, n2518,
         n2517, n2516, n2515, n2514, n2513, n2512, n2510, n2509, n2508, n2858,
         \requesterAddressbuffer[3][0] , n2857, \requesterAddressbuffer[3][1] ,
         n2856, \requesterAddressbuffer[3][2] , n2855,
         \requesterAddressbuffer[3][3] , n2854, \requesterAddressbuffer[3][4] ,
         n2853, \requesterAddressbuffer[3][5] , n2738, n2737, n2735, n2732,
         n2730, n2729, n2728, n2727, n2726, n2724, n2722, n2721, n2719, n2717,
         n2716, n2714, n2712, n2711, n2710, n2709, n2708, n2707, n2506, n2505,
         n2503, n2502, n2501, n2500, n2495, n2852,
         \requesterAddressbuffer[2][0] , n2851, \requesterAddressbuffer[2][1] ,
         n2848, \requesterAddressbuffer[2][4] , n2767, n2766, n2765, n2763,
         n2762, n2761, n2759, n2758, n2757, n2756, n2755, n2753, n2752, n2751,
         n2750, n2749, n2747, n2745, n2744, n2742, n2741, n2740, n2490, n2479,
         n2800, n2797, n2794, n2792, n2783, n2782, n2780, n2775, n2837,
         \requesterAddressbuffer[0][3] , n2835, \requesterAddressbuffer[0][5] ,
         n2831, n2830, n2828, n2827, n2826, n2824, n2823, n2822, n2821, n2820,
         n2819, n2818, n2817, n2816, n2815, n2813, n2812, n2810, n2809, n2808,
         n2805, n2804, n2803, n2463, n2462, n2461, n2459, n2456, n2452, n2885,
         n2449, n2434, n2431, n2450, n2448, n2447, n2446, n2445, n2444, n2443,
         n2442, n2441, n2440, n2439, n2438, n2437, n2436, n2435, n2433, n2432,
         n2430, n2429, n2428, n2427, n2426, n2425, n2424, n2423, n2422, n2421,
         n2420, n2419, n2418, n2417, n2416, n2415, n2414, n2413, n2412, n2411,
         n2410, n2409, n2408, n2407, n2406, n2405, n2404, n2403, n2402, n2401,
         n2400, n2399, n2398, n2397, n2884, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n500, n501, n502, n503, n504, n505, n507, n508, n509,
         n511, n514, n516, n517, n534, n536, n537, n541, n543, n544, n545,
         n546, n548, n551, n554, n555, n556, n557, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n584, n594, n607, n608,
         n609, n610, n611, n612, n613, n614, n622, n623, n624, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n711, n712, n714, n715, n716, n717, n729,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n886, n919, n936, n955, n957, n970,
         n986, n1005, n1402, n1537, n1586, n1653, n1654, n1728, n1764, n1817,
         n1822, n1894, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5324, n5325, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349;
  wire   [0:7] readOutbuffer;
  wire   [0:7] writeOutbuffer;

  DFFNSRX2TS \destinationAddressbuffer_reg[2][6]  ( .D(n2486), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4827) );
  DFFNSRX2TS \destinationAddressbuffer_reg[2][8]  ( .D(n2484), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4807) );
  DFFNSRX2TS \destinationAddressbuffer_reg[2][10]  ( .D(n2482), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4793) );
  DFFNSRX2TS \destinationAddressbuffer_reg[2][12]  ( .D(n2480), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4779) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][7]  ( .D(n2457), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4815) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][9]  ( .D(n2455), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4799) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][11]  ( .D(n2453), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4785) );
  DFFNSRX2TS \destinationAddressbuffer_reg[2][7]  ( .D(n2485), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4820) );
  DFFNSRX2TS \destinationAddressbuffer_reg[2][9]  ( .D(n2483), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4804) );
  DFFNSRX2TS \destinationAddressbuffer_reg[2][11]  ( .D(n2481), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4788) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][6]  ( .D(n2458), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4828) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][10]  ( .D(n2454), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4794) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][13]  ( .D(n2451), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4772) );
  DFFNSRX2TS \destinationAddressbuffer_reg[2][13]  ( .D(n2479), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4765) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][8]  ( .D(n2456), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4805) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][12]  ( .D(n2452), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4773) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][7]  ( .D(n2499), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4819) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][10]  ( .D(n2496), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4795) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][13]  ( .D(n2493), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4769) );
  DFFNSRX2TS \destinationAddressbuffer_reg[5][6]  ( .D(n2528), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4822) );
  DFFNSRX2TS \destinationAddressbuffer_reg[5][7]  ( .D(n2527), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4816) );
  DFFNSRX2TS \destinationAddressbuffer_reg[5][8]  ( .D(n2526), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4810) );
  DFFNSRX2TS \destinationAddressbuffer_reg[5][9]  ( .D(n2525), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4800) );
  DFFNSRX2TS \destinationAddressbuffer_reg[5][10]  ( .D(n2524), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4796) );
  DFFNSRX2TS \destinationAddressbuffer_reg[5][11]  ( .D(n2523), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4786) );
  DFFNSRX2TS \destinationAddressbuffer_reg[5][12]  ( .D(n2522), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4780) );
  DFFNSRX2TS \destinationAddressbuffer_reg[5][13]  ( .D(n2521), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4770) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][8]  ( .D(n2498), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4812) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][9]  ( .D(n2497), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4798) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][12]  ( .D(n2494), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4776) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][6]  ( .D(n2500), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4823) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][11]  ( .D(n2495), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4783) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][9]  ( .D(n2511), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4803) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][13]  ( .D(n2507), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4771) );
  DFFNSRX2TS \destinationAddressbuffer_reg[6][10]  ( .D(n2538), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4789) );
  DFFNSRX2TS \destinationAddressbuffer_reg[6][12]  ( .D(n2536), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4777) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][6]  ( .D(n2514), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4825) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][7]  ( .D(n2513), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4813) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][8]  ( .D(n2512), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4809) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][10]  ( .D(n2510), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4791) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][11]  ( .D(n2509), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4781) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][12]  ( .D(n2508), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4775) );
  DFFNSRX2TS \dataoutbuffer_reg[4][3]  ( .D(n2703), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4678) );
  DFFNSRX2TS \dataoutbuffer_reg[4][14]  ( .D(n2692), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4579) );
  DFFNSRX2TS \dataoutbuffer_reg[4][15]  ( .D(n2691), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4570) );
  DFFNSRX2TS \dataoutbuffer_reg[4][17]  ( .D(n2689), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4552) );
  DFFNSRX2TS \dataoutbuffer_reg[4][0]  ( .D(n2706), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4702) );
  DFFNSRX2TS \dataoutbuffer_reg[4][1]  ( .D(n2705), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4691) );
  DFFNSRX2TS \dataoutbuffer_reg[4][6]  ( .D(n2700), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4650) );
  DFFNSRX2TS \dataoutbuffer_reg[4][8]  ( .D(n2698), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4628) );
  DFFNSRX2TS \dataoutbuffer_reg[4][10]  ( .D(n2696), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4612) );
  DFFNSRX2TS \dataoutbuffer_reg[4][11]  ( .D(n2695), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4605) );
  DFFNSRX2TS \dataoutbuffer_reg[4][12]  ( .D(n2694), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4594) );
  DFFNSRX2TS \dataoutbuffer_reg[4][16]  ( .D(n2690), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4556) );
  DFFNSRX2TS \dataoutbuffer_reg[4][19]  ( .D(n2687), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4529) );
  DFFNSRX2TS \dataoutbuffer_reg[4][20]  ( .D(n2686), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4524) );
  DFFNSRX2TS \dataoutbuffer_reg[4][21]  ( .D(n2685), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4515) );
  DFFNSRX2TS \dataoutbuffer_reg[4][22]  ( .D(n2684), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4504) );
  DFFNSRX2TS \dataoutbuffer_reg[4][29]  ( .D(n2677), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4445) );
  DFFNSRX2TS \dataoutbuffer_reg[4][31]  ( .D(n2675), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4421) );
  DFFNSRX2TS \dataoutbuffer_reg[4][2]  ( .D(n2704), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4683) );
  DFFNSRX2TS \dataoutbuffer_reg[4][4]  ( .D(n2702), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4667) );
  DFFNSRX2TS \dataoutbuffer_reg[4][5]  ( .D(n2701), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4656) );
  DFFNSRX2TS \dataoutbuffer_reg[4][7]  ( .D(n2699), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4640) );
  DFFNSRX2TS \dataoutbuffer_reg[4][9]  ( .D(n2697), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4622) );
  DFFNSRX2TS \dataoutbuffer_reg[4][13]  ( .D(n2693), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4582) );
  DFFNSRX2TS \dataoutbuffer_reg[4][18]  ( .D(n2688), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4537) );
  DFFNSRX2TS \dataoutbuffer_reg[4][23]  ( .D(n2683), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4494) );
  DFFNSRX2TS \dataoutbuffer_reg[4][24]  ( .D(n2682), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4483) );
  DFFNSRX2TS \dataoutbuffer_reg[4][25]  ( .D(n2681), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4478) );
  DFFNSRX2TS \dataoutbuffer_reg[4][26]  ( .D(n2680), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4465) );
  DFFNSRX2TS \dataoutbuffer_reg[4][27]  ( .D(n2679), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4458) );
  DFFNSRX2TS \dataoutbuffer_reg[4][28]  ( .D(n2678), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4447) );
  DFFNSRX2TS \dataoutbuffer_reg[4][30]  ( .D(n2676), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4429) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][0]  ( .D(n2520), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4757) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][1]  ( .D(n2519), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4752) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][2]  ( .D(n2518), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4739) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][3]  ( .D(n2517), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4734) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][5]  ( .D(n2515), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4714) );
  DFFNSRX2TS \requesterAddressbuffer_reg[2][2]  ( .D(n2850), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][2] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[2][3]  ( .D(n2849), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][3] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[2][5]  ( .D(n2847), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][5] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[0][0]  ( .D(n2840), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][0] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[0][1]  ( .D(n2839), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][1] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[0][2]  ( .D(n2838), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][2] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[0][4]  ( .D(n2836), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][4] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[2][0]  ( .D(n2852), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][0] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[2][1]  ( .D(n2851), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][1] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[2][4]  ( .D(n2848), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][4] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[0][3]  ( .D(n2837), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][3] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[0][5]  ( .D(n2835), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][5] ) );
  DFFNSRX2TS \readOutbuffer_reg[3]  ( .D(n2566), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[3]) );
  DFFNSRX2TS \readOutbuffer_reg[6]  ( .D(n2569), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n18) );
  DFFNSRX2TS \readOutbuffer_reg[5]  ( .D(n2568), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n19) );
  DFFNSRX2TS \readOutbuffer_reg[1]  ( .D(n2564), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n16) );
  DFFNSRX2TS \writeOutbuffer_reg[5]  ( .D(n2576), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n17) );
  DFFNSRX2TS \writeOutbuffer_reg[2]  ( .D(n2573), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[2]), .QN(n101) );
  DFFNSRX2TS \dataoutbuffer_reg[2][0]  ( .D(n2770), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n95), .QN(n4701) );
  DFFNSRX2TS \dataoutbuffer_reg[2][2]  ( .D(n2768), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n94), .QN(n4685) );
  DFFNSRX2TS \dataoutbuffer_reg[2][6]  ( .D(n2764), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n93), .QN(n4651) );
  DFFNSRX2TS \dataoutbuffer_reg[2][16]  ( .D(n2754), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n92), .QN(n4561) );
  DFFNSRX2TS \dataoutbuffer_reg[2][22]  ( .D(n2748), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n91), .QN(n4507) );
  DFFNSRX2TS \dataoutbuffer_reg[2][24]  ( .D(n2746), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n90), .QN(n4489) );
  DFFNSRX2TS \dataoutbuffer_reg[2][31]  ( .D(n2739), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n89), .QN(n4426) );
  DFFNSRX2TS \dataoutbuffer_reg[0][0]  ( .D(n2834), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n57), .QN(n4703) );
  DFFNSRX2TS \dataoutbuffer_reg[0][1]  ( .D(n2833), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n56), .QN(n4696) );
  DFFNSRX2TS \dataoutbuffer_reg[0][2]  ( .D(n2832), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n55), .QN(n4687) );
  DFFNSRX2TS \dataoutbuffer_reg[0][5]  ( .D(n2829), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n54), .QN(n4660) );
  DFFNSRX2TS \dataoutbuffer_reg[0][9]  ( .D(n2825), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n53), .QN(n4624) );
  DFFNSRX2TS \dataoutbuffer_reg[0][20]  ( .D(n2814), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n52), .QN(n4525) );
  DFFNSRX2TS \dataoutbuffer_reg[0][23]  ( .D(n2811), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n51), .QN(n4498) );
  DFFNSRX2TS \dataoutbuffer_reg[0][27]  ( .D(n2807), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n50), .QN(n4462) );
  DFFNSRX2TS \dataoutbuffer_reg[0][28]  ( .D(n2806), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n49), .QN(n4453) );
  DFFNSRX2TS \dataoutbuffer_reg[2][1]  ( .D(n2769), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n88), .QN(n4697) );
  DFFNSRX2TS \dataoutbuffer_reg[2][10]  ( .D(n2760), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n87), .QN(n4614) );
  DFFNSRX2TS \dataoutbuffer_reg[2][27]  ( .D(n2743), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n86), .QN(n4463) );
  DFFNSRX2TS \destinationAddressbuffer_reg[2][0]  ( .D(n2492), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n85), .QN(n4758) );
  DFFNSRX2TS \destinationAddressbuffer_reg[2][1]  ( .D(n2491), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n84), .QN(n4751) );
  DFFNSRX2TS \destinationAddressbuffer_reg[2][3]  ( .D(n2489), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n83), .QN(n4737) );
  DFFNSRX2TS \destinationAddressbuffer_reg[2][4]  ( .D(n2488), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n82), .QN(n4728) );
  DFFNSRX2TS \destinationAddressbuffer_reg[2][5]  ( .D(n2487), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n81), .QN(n4715) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][0]  ( .D(n2464), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n48), .QN(n4762) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][4]  ( .D(n2460), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n47), .QN(n4724) );
  DFFNSRX2TS \dataoutbuffer_reg[2][3]  ( .D(n2767), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n80), .QN(n4672) );
  DFFNSRX2TS \dataoutbuffer_reg[2][4]  ( .D(n2766), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n79), .QN(n4665) );
  DFFNSRX2TS \dataoutbuffer_reg[2][5]  ( .D(n2765), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n78), .QN(n4658) );
  DFFNSRX2TS \dataoutbuffer_reg[2][7]  ( .D(n2763), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n77), .QN(n4636) );
  DFFNSRX2TS \dataoutbuffer_reg[2][8]  ( .D(n2762), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n76), .QN(n4631) );
  DFFNSRX2TS \dataoutbuffer_reg[2][9]  ( .D(n2761), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n75), .QN(n4618) );
  DFFNSRX2TS \dataoutbuffer_reg[2][11]  ( .D(n2759), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n74), .QN(n4606) );
  DFFNSRX2TS \dataoutbuffer_reg[2][12]  ( .D(n2758), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n73), .QN(n4591) );
  DFFNSRX2TS \dataoutbuffer_reg[2][13]  ( .D(n2757), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n72), .QN(n4584) );
  DFFNSRX2TS \dataoutbuffer_reg[2][14]  ( .D(n2756), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n71), .QN(n4573) );
  DFFNSRX2TS \dataoutbuffer_reg[2][15]  ( .D(n2755), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n70), .QN(n4566) );
  DFFNSRX2TS \dataoutbuffer_reg[2][17]  ( .D(n2753), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n69), .QN(n4550) );
  DFFNSRX2TS \dataoutbuffer_reg[2][18]  ( .D(n2752), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n68), .QN(n4541) );
  DFFNSRX2TS \dataoutbuffer_reg[2][19]  ( .D(n2751), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n67), .QN(n4528) );
  DFFNSRX2TS \dataoutbuffer_reg[2][20]  ( .D(n2750), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n66), .QN(n4523) );
  DFFNSRX2TS \dataoutbuffer_reg[2][21]  ( .D(n2749), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n65), .QN(n4510) );
  DFFNSRX2TS \dataoutbuffer_reg[2][23]  ( .D(n2747), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n64), .QN(n4496) );
  DFFNSRX2TS \dataoutbuffer_reg[2][25]  ( .D(n2745), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n63), .QN(n4474) );
  DFFNSRX2TS \dataoutbuffer_reg[2][26]  ( .D(n2744), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n62), .QN(n4467) );
  DFFNSRX2TS \dataoutbuffer_reg[2][28]  ( .D(n2742), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n61), .QN(n4449) );
  DFFNSRX2TS \dataoutbuffer_reg[2][29]  ( .D(n2741), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n60), .QN(n4438) );
  DFFNSRX2TS \dataoutbuffer_reg[2][30]  ( .D(n2740), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n59), .QN(n4431) );
  DFFNSRX2TS \destinationAddressbuffer_reg[2][2]  ( .D(n2490), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n58), .QN(n4745) );
  DFFNSRX2TS \dataoutbuffer_reg[0][3]  ( .D(n2831), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n46), .QN(n4674) );
  DFFNSRX2TS \dataoutbuffer_reg[0][4]  ( .D(n2830), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n45), .QN(n4663) );
  DFFNSRX2TS \dataoutbuffer_reg[0][6]  ( .D(n2828), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n44), .QN(n4647) );
  DFFNSRX2TS \dataoutbuffer_reg[0][7]  ( .D(n2827), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n43), .QN(n4638) );
  DFFNSRX2TS \dataoutbuffer_reg[0][8]  ( .D(n2826), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n42), .QN(n4633) );
  DFFNSRX2TS \dataoutbuffer_reg[0][10]  ( .D(n2824), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n41), .QN(n4613) );
  DFFNSRX2TS \dataoutbuffer_reg[0][11]  ( .D(n2823), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n40), .QN(n4600) );
  DFFNSRX2TS \dataoutbuffer_reg[0][12]  ( .D(n2822), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n39), .QN(n4595) );
  DFFNSRX2TS \dataoutbuffer_reg[0][13]  ( .D(n2821), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n38), .QN(n4588) );
  DFFNSRX2TS \dataoutbuffer_reg[0][14]  ( .D(n2820), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n37), .QN(n4575) );
  DFFNSRX2TS \dataoutbuffer_reg[0][15]  ( .D(n2819), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n36), .QN(n4568) );
  DFFNSRX2TS \dataoutbuffer_reg[0][16]  ( .D(n2818), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n35), .QN(n4557) );
  DFFNSRX2TS \dataoutbuffer_reg[0][17]  ( .D(n2817), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n34), .QN(n4548) );
  DFFNSRX2TS \dataoutbuffer_reg[0][18]  ( .D(n2816), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n33), .QN(n4539) );
  DFFNSRX2TS \dataoutbuffer_reg[0][19]  ( .D(n2815), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n32), .QN(n4530) );
  DFFNSRX2TS \dataoutbuffer_reg[0][21]  ( .D(n2813), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n31), .QN(n4516) );
  DFFNSRX2TS \dataoutbuffer_reg[0][22]  ( .D(n2812), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n30), .QN(n4501) );
  DFFNSRX2TS \dataoutbuffer_reg[0][24]  ( .D(n2810), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n29), .QN(n4485) );
  DFFNSRX2TS \dataoutbuffer_reg[0][25]  ( .D(n2809), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n28), .QN(n4476) );
  DFFNSRX2TS \dataoutbuffer_reg[0][26]  ( .D(n2808), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n27), .QN(n4469) );
  DFFNSRX2TS \dataoutbuffer_reg[0][29]  ( .D(n2805), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n26), .QN(n4444) );
  DFFNSRX2TS \dataoutbuffer_reg[0][30]  ( .D(n2804), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n25), .QN(n4433) );
  DFFNSRX2TS \dataoutbuffer_reg[0][31]  ( .D(n2803), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n24), .QN(n4420) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][1]  ( .D(n2463), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n23), .QN(n4748) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][2]  ( .D(n2462), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n22), .QN(n4743) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][3]  ( .D(n2461), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n21), .QN(n4732) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][5]  ( .D(n2459), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n20), .QN(n4712) );
  DFFNSRX2TS \writeOutbuffer_reg[0]  ( .D(n2571), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[0]), .QN(n103) );
  DFFNSRX2TS \writeOutbuffer_reg[3]  ( .D(n2574), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[3]), .QN(n102) );
  DFFNSRX2TS \writeOutbuffer_reg[4]  ( .D(n2575), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[4]), .QN(n100) );
  DFFNSRX2TS \readOutbuffer_reg[7]  ( .D(n2570), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[7]), .QN(n98) );
  DFFNSRX2TS \readOutbuffer_reg[2]  ( .D(n2565), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[2]), .QN(n99) );
  DFFNSRX2TS \readOutbuffer_reg[4]  ( .D(n2567), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[4]), .QN(n97) );
  DFFNSRX2TS \read_reg_reg[0]  ( .D(n2889), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n4), .QN(n7) );
  DFFNSRX2TS full_reg_reg ( .D(N4718), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        n4832), .QN(n96) );
  DFFNSRX2TS \write_reg_reg[1]  ( .D(n2887), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n393), .QN(n5323) );
  DFFNSRX2TS writeOut_reg ( .D(n2449), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        writeOut), .QN(n4829) );
  DFFNSRX2TS \requesterAddressOut_reg[0]  ( .D(n2434), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[0]), .QN(n4833) );
  DFFNSRX2TS \requesterAddressOut_reg[3]  ( .D(n2431), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[3]), .QN(n4834) );
  DFFNSRX2TS readOut_reg ( .D(n2450), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        readOut), .QN(n4831) );
  DFFNSRX2TS \destinationAddressOut_reg[0]  ( .D(n2440), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[0]), .QN(n4756) );
  DFFNSRX2TS \destinationAddressOut_reg[1]  ( .D(n2439), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[1]), .QN(n4747) );
  DFFNSRX2TS \destinationAddressOut_reg[2]  ( .D(n2438), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[2]), .QN(n4738) );
  DFFNSRX2TS \destinationAddressOut_reg[3]  ( .D(n2437), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[3]), .QN(n4729) );
  DFFNSRX2TS \destinationAddressOut_reg[4]  ( .D(n2436), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[4]), .QN(n4720) );
  DFFNSRX2TS \destinationAddressOut_reg[5]  ( .D(n2435), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[5]), .QN(n4711) );
  DFFNSRX2TS \requesterAddressOut_reg[1]  ( .D(n2433), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[1]), .QN(n4710) );
  DFFNSRX2TS \requesterAddressOut_reg[2]  ( .D(n2432), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[2]), .QN(n4709) );
  DFFNSRX2TS \requesterAddressOut_reg[4]  ( .D(n2430), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[4]), .QN(n4708) );
  DFFNSRX2TS \requesterAddressOut_reg[5]  ( .D(n2429), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[5]), .QN(n4707) );
  DFFNSRX2TS \dataOut_reg[0]  ( .D(n2428), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[0]), .QN(n4698) );
  DFFNSRX2TS \dataOut_reg[1]  ( .D(n2427), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[1]), .QN(n4689) );
  DFFNSRX2TS \dataOut_reg[2]  ( .D(n2426), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[2]), .QN(n4680) );
  DFFNSRX2TS \dataOut_reg[3]  ( .D(n2425), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[3]), .QN(n4671) );
  DFFNSRX2TS \dataOut_reg[4]  ( .D(n2424), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[4]), .QN(n4662) );
  DFFNSRX2TS \dataOut_reg[5]  ( .D(n2423), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[5]), .QN(n4653) );
  DFFNSRX2TS \dataOut_reg[6]  ( .D(n2422), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[6]), .QN(n4644) );
  DFFNSRX2TS \dataOut_reg[7]  ( .D(n2421), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[7]), .QN(n4635) );
  DFFNSRX2TS \dataOut_reg[8]  ( .D(n2420), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[8]), .QN(n4626) );
  DFFNSRX2TS \dataOut_reg[9]  ( .D(n2419), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[9]), .QN(n4617) );
  DFFNSRX2TS \dataOut_reg[10]  ( .D(n2418), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[10]), .QN(n4608) );
  DFFNSRX2TS \dataOut_reg[11]  ( .D(n2417), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[11]), .QN(n4599) );
  DFFNSRX2TS \dataOut_reg[12]  ( .D(n2416), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[12]), .QN(n4590) );
  DFFNSRX2TS \dataOut_reg[13]  ( .D(n2415), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[13]), .QN(n4581) );
  DFFNSRX2TS \dataOut_reg[14]  ( .D(n2414), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[14]), .QN(n4572) );
  DFFNSRX2TS \dataOut_reg[15]  ( .D(n2413), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[15]), .QN(n4563) );
  DFFNSRX2TS \dataOut_reg[16]  ( .D(n2412), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[16]), .QN(n4554) );
  DFFNSRX2TS \dataOut_reg[17]  ( .D(n2411), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[17]), .QN(n4545) );
  DFFNSRX2TS \dataOut_reg[18]  ( .D(n2410), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[18]), .QN(n4536) );
  DFFNSRX2TS \dataOut_reg[19]  ( .D(n2409), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[19]), .QN(n4527) );
  DFFNSRX2TS \dataOut_reg[20]  ( .D(n2408), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[20]), .QN(n4518) );
  DFFNSRX2TS \dataOut_reg[21]  ( .D(n2407), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[21]), .QN(n4509) );
  DFFNSRX2TS \dataOut_reg[22]  ( .D(n2406), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[22]), .QN(n4500) );
  DFFNSRX2TS \dataOut_reg[23]  ( .D(n2405), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[23]), .QN(n4491) );
  DFFNSRX2TS \dataOut_reg[24]  ( .D(n2404), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[24]), .QN(n4482) );
  DFFNSRX2TS \dataOut_reg[25]  ( .D(n2403), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[25]), .QN(n4473) );
  DFFNSRX2TS \dataOut_reg[26]  ( .D(n2402), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[26]), .QN(n4464) );
  DFFNSRX2TS \dataOut_reg[27]  ( .D(n2401), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[27]), .QN(n4455) );
  DFFNSRX2TS \dataOut_reg[28]  ( .D(n2400), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[28]), .QN(n4446) );
  DFFNSRX2TS \dataOut_reg[29]  ( .D(n2399), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[29]), .QN(n4437) );
  DFFNSRX2TS \dataOut_reg[30]  ( .D(n2398), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[30]), .QN(n4428) );
  DFFNSRX2TS \dataOut_reg[31]  ( .D(n2397), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[31]), .QN(n4419) );
  DFFNSRX2TS \destinationAddressOut_reg[6]  ( .D(n2448), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[6]) );
  DFFNSRX2TS \destinationAddressOut_reg[7]  ( .D(n2447), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[7]) );
  DFFNSRX2TS \destinationAddressOut_reg[8]  ( .D(n2446), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[8]) );
  DFFNSRX2TS \destinationAddressOut_reg[9]  ( .D(n2445), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[9]) );
  DFFNSRX2TS \destinationAddressOut_reg[10]  ( .D(n2444), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[10]) );
  DFFNSRX2TS \destinationAddressOut_reg[11]  ( .D(n2443), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[11]) );
  DFFNSRX2TS \destinationAddressOut_reg[12]  ( .D(n2442), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[12]) );
  DFFNSRX2TS \destinationAddressOut_reg[13]  ( .D(n2441), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[13]) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][13]  ( .D(n2549), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4768) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][6]  ( .D(n2472), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4826) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][7]  ( .D(n2471), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4814) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][8]  ( .D(n2470), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4806) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][9]  ( .D(n2469), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4802) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][10]  ( .D(n2468), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4790) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][11]  ( .D(n2467), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4784) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][12]  ( .D(n2466), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4774) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][13]  ( .D(n2465), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4766) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][4]  ( .D(n2530), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4726) );
  DFFNSRXLTS \dataoutbuffer_reg[5][0]  ( .D(n2674), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4706) );
  DFFNSRXLTS \dataoutbuffer_reg[5][2]  ( .D(n2672), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4684) );
  DFFNSRXLTS \dataoutbuffer_reg[5][3]  ( .D(n2671), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4679) );
  DFFNSRXLTS \dataoutbuffer_reg[5][4]  ( .D(n2670), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4668) );
  DFFNSRXLTS \dataoutbuffer_reg[5][5]  ( .D(n2669), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4661) );
  DFFNSRXLTS \dataoutbuffer_reg[5][6]  ( .D(n2668), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4648) );
  DFFNSRXLTS \dataoutbuffer_reg[5][7]  ( .D(n2667), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4641) );
  DFFNSRXLTS \dataoutbuffer_reg[5][8]  ( .D(n2666), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4632) );
  DFFNSRXLTS \dataoutbuffer_reg[5][9]  ( .D(n2665), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4621) );
  DFFNSRXLTS \dataoutbuffer_reg[5][10]  ( .D(n2664), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4610) );
  DFFNSRXLTS \dataoutbuffer_reg[5][12]  ( .D(n2662), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4596) );
  DFFNSRXLTS \dataoutbuffer_reg[5][13]  ( .D(n2661), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4587) );
  DFFNSRXLTS \dataoutbuffer_reg[5][14]  ( .D(n2660), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4574) );
  DFFNSRXLTS \dataoutbuffer_reg[5][17]  ( .D(n2657), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4551) );
  DFFNSRXLTS \dataoutbuffer_reg[5][18]  ( .D(n2656), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4540) );
  DFFNSRXLTS \dataoutbuffer_reg[5][19]  ( .D(n2655), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4533) );
  DFFNSRXLTS \dataoutbuffer_reg[5][20]  ( .D(n2654), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4520) );
  DFFNSRXLTS \dataoutbuffer_reg[5][21]  ( .D(n2653), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4513) );
  DFFNSRXLTS \dataoutbuffer_reg[5][22]  ( .D(n2652), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4506) );
  DFFNSRXLTS \dataoutbuffer_reg[5][23]  ( .D(n2651), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4495) );
  DFFNSRXLTS \dataoutbuffer_reg[5][24]  ( .D(n2650), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4488) );
  DFFNSRXLTS \dataoutbuffer_reg[5][25]  ( .D(n2649), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4481) );
  DFFNSRXLTS \dataoutbuffer_reg[5][26]  ( .D(n2648), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4466) );
  DFFNSRXLTS \dataoutbuffer_reg[5][27]  ( .D(n2647), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4457) );
  DFFNSRXLTS \dataoutbuffer_reg[5][28]  ( .D(n2646), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4454) );
  DFFNSRXLTS \dataoutbuffer_reg[5][29]  ( .D(n2645), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4443) );
  DFFNSRXLTS \dataoutbuffer_reg[5][30]  ( .D(n2644), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4432) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][0]  ( .D(n2534), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4760) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][1]  ( .D(n2533), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4753) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][2]  ( .D(n2532), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4744) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][3]  ( .D(n2531), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4735) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][5]  ( .D(n2529), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4717) );
  DFFNSRXLTS \dataoutbuffer_reg[5][1]  ( .D(n2673), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4694) );
  DFFNSRXLTS \dataoutbuffer_reg[5][11]  ( .D(n2663), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4602) );
  DFFNSRXLTS \dataoutbuffer_reg[5][15]  ( .D(n2659), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4564) );
  DFFNSRXLTS \dataoutbuffer_reg[5][16]  ( .D(n2658), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4559) );
  DFFNSRXLTS \dataoutbuffer_reg[5][31]  ( .D(n2643), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4424) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][4]  ( .D(n2558), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4721) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][4]  ( .D(n2516), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4725) );
  DFFNSRXLTS \dataoutbuffer_reg[6][4]  ( .D(n2638), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4669) );
  DFFNSRXLTS \dataoutbuffer_reg[6][18]  ( .D(n2624), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4543) );
  DFFNSRXLTS \dataoutbuffer_reg[1][0]  ( .D(n2802), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4705) );
  DFFNSRXLTS \dataoutbuffer_reg[7][1]  ( .D(n2609), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4695) );
  DFFNSRXLTS \dataoutbuffer_reg[7][2]  ( .D(n2608), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4682) );
  DFFNSRXLTS \dataoutbuffer_reg[7][3]  ( .D(n2607), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4677) );
  DFFNSRXLTS \dataoutbuffer_reg[7][4]  ( .D(n2606), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4664) );
  DFFNSRXLTS \dataoutbuffer_reg[7][5]  ( .D(n2605), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4655) );
  DFFNSRXLTS \dataoutbuffer_reg[7][6]  ( .D(n2604), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4652) );
  DFFNSRXLTS \dataoutbuffer_reg[7][7]  ( .D(n2603), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4637) );
  DFFNSRXLTS \dataoutbuffer_reg[7][8]  ( .D(n2602), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4630) );
  DFFNSRXLTS \dataoutbuffer_reg[7][9]  ( .D(n2601), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4625) );
  DFFNSRXLTS \dataoutbuffer_reg[7][10]  ( .D(n2600), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4616) );
  DFFNSRXLTS \dataoutbuffer_reg[7][11]  ( .D(n2599), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4603) );
  DFFNSRXLTS \dataoutbuffer_reg[7][12]  ( .D(n2598), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4592) );
  DFFNSRXLTS \dataoutbuffer_reg[7][16]  ( .D(n2594), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4560) );
  DFFNSRXLTS \dataoutbuffer_reg[7][17]  ( .D(n2593), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4549) );
  DFFNSRXLTS \dataoutbuffer_reg[7][18]  ( .D(n2592), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4538) );
  DFFNSRXLTS \dataoutbuffer_reg[7][19]  ( .D(n2591), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4535) );
  DFFNSRXLTS \dataoutbuffer_reg[7][20]  ( .D(n2590), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4522) );
  DFFNSRXLTS \dataoutbuffer_reg[7][21]  ( .D(n2589), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4517) );
  DFFNSRXLTS \dataoutbuffer_reg[7][22]  ( .D(n2588), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4502) );
  DFFNSRXLTS \dataoutbuffer_reg[7][23]  ( .D(n2587), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4497) );
  DFFNSRXLTS \dataoutbuffer_reg[7][24]  ( .D(n2586), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4486) );
  DFFNSRXLTS \dataoutbuffer_reg[7][25]  ( .D(n2585), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4477) );
  DFFNSRXLTS \dataoutbuffer_reg[7][26]  ( .D(n2584), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4468) );
  DFFNSRXLTS \dataoutbuffer_reg[7][27]  ( .D(n2583), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4461) );
  DFFNSRXLTS \dataoutbuffer_reg[7][28]  ( .D(n2582), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4452) );
  DFFNSRXLTS \dataoutbuffer_reg[7][29]  ( .D(n2581), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4439) );
  DFFNSRXLTS \dataoutbuffer_reg[7][30]  ( .D(n2580), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4430) );
  DFFNSRXLTS \dataoutbuffer_reg[7][31]  ( .D(n2579), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4425) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][1]  ( .D(n2561), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4749) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][2]  ( .D(n2560), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4742) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][3]  ( .D(n2559), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4731) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][5]  ( .D(n2557), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4719) );
  DFFNSRXLTS \dataoutbuffer_reg[6][0]  ( .D(n2642), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4704) );
  DFFNSRXLTS \dataoutbuffer_reg[6][2]  ( .D(n2640), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4688) );
  DFFNSRXLTS \dataoutbuffer_reg[6][3]  ( .D(n2639), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4673) );
  DFFNSRXLTS \dataoutbuffer_reg[6][5]  ( .D(n2637), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4657) );
  DFFNSRXLTS \dataoutbuffer_reg[6][9]  ( .D(n2633), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4623) );
  DFFNSRXLTS \dataoutbuffer_reg[6][14]  ( .D(n2628), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4578) );
  DFFNSRXLTS \dataoutbuffer_reg[6][28]  ( .D(n2614), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4450) );
  DFFNSRXLTS \dataoutbuffer_reg[6][30]  ( .D(n2612), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4434) );
  DFFNSRXLTS \dataoutbuffer_reg[1][1]  ( .D(n2801), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4693) );
  DFFNSRXLTS \dataoutbuffer_reg[1][3]  ( .D(n2799), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4675) );
  DFFNSRXLTS \dataoutbuffer_reg[1][4]  ( .D(n2798), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4670) );
  DFFNSRXLTS \dataoutbuffer_reg[1][6]  ( .D(n2796), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4646) );
  DFFNSRXLTS \dataoutbuffer_reg[1][7]  ( .D(n2795), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4643) );
  DFFNSRXLTS \dataoutbuffer_reg[1][9]  ( .D(n2793), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4619) );
  DFFNSRXLTS \dataoutbuffer_reg[1][11]  ( .D(n2791), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4601) );
  DFFNSRXLTS \dataoutbuffer_reg[1][12]  ( .D(n2790), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4598) );
  DFFNSRXLTS \dataoutbuffer_reg[1][13]  ( .D(n2789), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4589) );
  DFFNSRXLTS \dataoutbuffer_reg[1][14]  ( .D(n2788), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4576) );
  DFFNSRXLTS \dataoutbuffer_reg[1][15]  ( .D(n2787), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4569) );
  DFFNSRXLTS \dataoutbuffer_reg[1][16]  ( .D(n2786), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4562) );
  DFFNSRXLTS \dataoutbuffer_reg[1][17]  ( .D(n2785), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4547) );
  DFFNSRXLTS \dataoutbuffer_reg[1][18]  ( .D(n2784), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4544) );
  DFFNSRXLTS \dataoutbuffer_reg[1][21]  ( .D(n2781), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4511) );
  DFFNSRXLTS \dataoutbuffer_reg[1][23]  ( .D(n2779), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4493) );
  DFFNSRXLTS \dataoutbuffer_reg[1][24]  ( .D(n2778), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4484) );
  DFFNSRXLTS \dataoutbuffer_reg[1][25]  ( .D(n2777), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4479) );
  DFFNSRXLTS \dataoutbuffer_reg[1][26]  ( .D(n2776), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4472) );
  DFFNSRXLTS \dataoutbuffer_reg[1][28]  ( .D(n2774), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4448) );
  DFFNSRXLTS \dataoutbuffer_reg[1][29]  ( .D(n2773), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4441) );
  DFFNSRXLTS \dataoutbuffer_reg[1][30]  ( .D(n2772), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4436) );
  DFFNSRXLTS \dataoutbuffer_reg[1][31]  ( .D(n2771), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4427) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][0]  ( .D(n2478), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4764) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][1]  ( .D(n2477), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4755) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][2]  ( .D(n2476), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4746) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][3]  ( .D(n2475), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4733) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][5]  ( .D(n2473), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4713) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][0]  ( .D(n2562), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4763) );
  DFFNSRXLTS \dataoutbuffer_reg[6][1]  ( .D(n2641), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4692) );
  DFFNSRXLTS \dataoutbuffer_reg[6][6]  ( .D(n2636), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4645) );
  DFFNSRXLTS \dataoutbuffer_reg[6][10]  ( .D(n2632), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4609) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][0]  ( .D(n2548), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4759) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][1]  ( .D(n2547), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4750) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][2]  ( .D(n2546), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4741) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][3]  ( .D(n2545), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4730) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][5]  ( .D(n2543), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4716) );
  DFFNSRXLTS \dataoutbuffer_reg[1][2]  ( .D(n2800), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4681) );
  DFFNSRXLTS \dataoutbuffer_reg[1][5]  ( .D(n2797), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4654) );
  DFFNSRXLTS \dataoutbuffer_reg[1][8]  ( .D(n2794), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4629) );
  DFFNSRXLTS \dataoutbuffer_reg[1][10]  ( .D(n2792), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4615) );
  DFFNSRXLTS \dataoutbuffer_reg[1][19]  ( .D(n2783), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4532) );
  DFFNSRXLTS \dataoutbuffer_reg[1][20]  ( .D(n2782), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4521) );
  DFFNSRXLTS \dataoutbuffer_reg[1][22]  ( .D(n2780), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4505) );
  DFFNSRXLTS \dataoutbuffer_reg[1][27]  ( .D(n2775), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4456) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][4]  ( .D(n2544), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4727) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][10]  ( .D(n2552), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n480), .QN(n4792) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][4]  ( .D(n2474), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4722) );
  DFFNSRXLTS \dataoutbuffer_reg[3][7]  ( .D(n2731), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n6313), .QN(n4642) );
  DFFNSRXLTS \dataoutbuffer_reg[3][2]  ( .D(n2736), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n6300), .QN(n4686) );
  DFFNSRXLTS \dataoutbuffer_reg[3][4]  ( .D(n2734), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n6299), .QN(n4666) );
  DFFNSRXLTS \dataoutbuffer_reg[3][5]  ( .D(n2733), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n6298), .QN(n4659) );
  DFFNSRXLTS \dataoutbuffer_reg[3][13]  ( .D(n2725), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6297), .QN(n4585) );
  DFFNSRXLTS \dataoutbuffer_reg[3][15]  ( .D(n2723), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6296), .QN(n4567) );
  DFFNSRXLTS \dataoutbuffer_reg[3][18]  ( .D(n2720), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6295), .QN(n4542) );
  DFFNSRXLTS \dataoutbuffer_reg[3][20]  ( .D(n2718), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6294), .QN(n4526) );
  DFFNSRXLTS \dataoutbuffer_reg[3][23]  ( .D(n2715), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6293), .QN(n4499) );
  DFFNSRXLTS \dataoutbuffer_reg[3][25]  ( .D(n2713), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6292), .QN(n4475) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][2]  ( .D(n2504), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n6291), .QN(n4740) );
  DFFNSRXLTS \dataoutbuffer_reg[3][0]  ( .D(n2738), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n6276), .QN(n4699) );
  DFFNSRXLTS \dataoutbuffer_reg[3][1]  ( .D(n2737), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n6275), .QN(n4690) );
  DFFNSRXLTS \dataoutbuffer_reg[3][3]  ( .D(n2735), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n6274), .QN(n4676) );
  DFFNSRXLTS \dataoutbuffer_reg[3][6]  ( .D(n2732), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n6273), .QN(n4649) );
  DFFNSRXLTS \dataoutbuffer_reg[3][8]  ( .D(n2730), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n6272), .QN(n4627) );
  DFFNSRXLTS \dataoutbuffer_reg[3][9]  ( .D(n2729), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n6271), .QN(n4620) );
  DFFNSRXLTS \dataoutbuffer_reg[3][10]  ( .D(n2728), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6270), .QN(n4611) );
  DFFNSRXLTS \dataoutbuffer_reg[3][11]  ( .D(n2727), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6269), .QN(n4604) );
  DFFNSRXLTS \dataoutbuffer_reg[3][12]  ( .D(n2726), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6268), .QN(n4593) );
  DFFNSRXLTS \dataoutbuffer_reg[3][14]  ( .D(n2724), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6267), .QN(n4577) );
  DFFNSRXLTS \dataoutbuffer_reg[3][16]  ( .D(n2722), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6266), .QN(n4555) );
  DFFNSRXLTS \dataoutbuffer_reg[3][17]  ( .D(n2721), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6265), .QN(n4546) );
  DFFNSRXLTS \dataoutbuffer_reg[3][19]  ( .D(n2719), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6264), .QN(n4534) );
  DFFNSRXLTS \dataoutbuffer_reg[3][21]  ( .D(n2717), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6263), .QN(n4514) );
  DFFNSRXLTS \dataoutbuffer_reg[3][22]  ( .D(n2716), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6262), .QN(n4503) );
  DFFNSRXLTS \dataoutbuffer_reg[3][24]  ( .D(n2714), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6261), .QN(n4487) );
  DFFNSRXLTS \dataoutbuffer_reg[3][26]  ( .D(n2712), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6260), .QN(n4471) );
  DFFNSRXLTS \dataoutbuffer_reg[3][27]  ( .D(n2711), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6259), .QN(n4460) );
  DFFNSRXLTS \dataoutbuffer_reg[3][28]  ( .D(n2710), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6258), .QN(n4451) );
  DFFNSRXLTS \dataoutbuffer_reg[3][29]  ( .D(n2709), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6257), .QN(n4440) );
  DFFNSRXLTS \dataoutbuffer_reg[3][30]  ( .D(n2708), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6256), .QN(n4435) );
  DFFNSRXLTS \dataoutbuffer_reg[3][31]  ( .D(n2707), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6255), .QN(n4422) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][0]  ( .D(n2506), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n6254), .QN(n4761) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][1]  ( .D(n2505), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n6253), .QN(n4754) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][3]  ( .D(n2503), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n6252), .QN(n4736) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][4]  ( .D(n2502), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n6251), .QN(n4723) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][5]  ( .D(n2501), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n6250), .QN(n4718) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][0]  ( .D(n2858), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][0] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][1]  ( .D(n2857), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][1] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][2]  ( .D(n2856), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][2] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][3]  ( .D(n2855), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][3] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][5]  ( .D(n2853), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][5] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][4]  ( .D(n2854), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][4] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[6][1]  ( .D(n2875), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][1] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[6][2]  ( .D(n2874), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][2] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[6][3]  ( .D(n2873), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][3] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[6][4]  ( .D(n2872), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][4] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[6][5]  ( .D(n2871), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][5] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[6][0]  ( .D(n2876), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][0] ) );
  DFFNSRXLTS \writeOutbuffer_reg[7]  ( .D(n2578), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n6315) );
  DFFNSRXLTS \requesterAddressbuffer_reg[7][0]  ( .D(n2882), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6311) );
  DFFNSRXLTS \requesterAddressbuffer_reg[7][1]  ( .D(n2881), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6310) );
  DFFNSRXLTS \requesterAddressbuffer_reg[7][3]  ( .D(n2879), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6309) );
  DFFNSRXLTS \requesterAddressbuffer_reg[5][0]  ( .D(n2870), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6308) );
  DFFNSRXLTS \requesterAddressbuffer_reg[5][1]  ( .D(n2869), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6307) );
  DFFNSRXLTS \requesterAddressbuffer_reg[5][2]  ( .D(n2868), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6306) );
  DFFNSRXLTS \requesterAddressbuffer_reg[5][3]  ( .D(n2867), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6305) );
  DFFNSRXLTS \requesterAddressbuffer_reg[5][4]  ( .D(n2866), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6304) );
  DFFNSRXLTS \requesterAddressbuffer_reg[5][5]  ( .D(n2865), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6303) );
  DFFNSRXLTS \requesterAddressbuffer_reg[7][2]  ( .D(n2880), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6283) );
  DFFNSRXLTS \requesterAddressbuffer_reg[7][4]  ( .D(n2878), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6282) );
  DFFNSRXLTS \requesterAddressbuffer_reg[7][5]  ( .D(n2877), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6281) );
  DFFNSRXLTS \readOutbuffer_reg[0]  ( .D(n2563), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n6312) );
  DFFNSRXLTS \requesterAddressbuffer_reg[4][4]  ( .D(n2860), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6302) );
  DFFNSRXLTS \requesterAddressbuffer_reg[4][5]  ( .D(n2859), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6301) );
  DFFNSRXLTS \requesterAddressbuffer_reg[4][0]  ( .D(n2864), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6280) );
  DFFNSRXLTS \requesterAddressbuffer_reg[4][1]  ( .D(n2863), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6279) );
  DFFNSRXLTS \requesterAddressbuffer_reg[4][2]  ( .D(n2862), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6278) );
  DFFNSRXLTS \requesterAddressbuffer_reg[4][3]  ( .D(n2861), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6277) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][0]  ( .D(n2846), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6290) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][1]  ( .D(n2845), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6289) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][2]  ( .D(n2844), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6288) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][3]  ( .D(n2843), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6287) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][4]  ( .D(n2842), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6286) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][5]  ( .D(n2841), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6285) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][7]  ( .D(n2541), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4817) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][8]  ( .D(n2540), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4811) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][11]  ( .D(n2537), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4787) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][13]  ( .D(n2535), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4767) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][6]  ( .D(n2556), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4824) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][7]  ( .D(n2555), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4818) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][8]  ( .D(n2554), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4808) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][11]  ( .D(n2551), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4782) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][12]  ( .D(n2550), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4778) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][9]  ( .D(n2553), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4801) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][6]  ( .D(n2542), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4821) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][9]  ( .D(n2539), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4797) );
  DFFNSRXLTS \writeOutbuffer_reg[6]  ( .D(n2577), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[6]), .QN(n6314) );
  DFFNSRXLTS \writeOutbuffer_reg[1]  ( .D(n2572), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[1]), .QN(n6284) );
  DFFNSRX2TS \read_reg_reg[1]  ( .D(n2883), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n5), .QN(n388) );
  DFFNSRX2TS \read_reg_reg[2]  ( .D(n2884), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n3), .QN(n385) );
  DFFNSRXLTS \dataoutbuffer_reg[7][15]  ( .D(n2595), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4565) );
  DFFNSRXLTS \dataoutbuffer_reg[7][14]  ( .D(n2596), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4580) );
  DFFNSRXLTS \dataoutbuffer_reg[7][13]  ( .D(n2597), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4583) );
  DFFNSRXLTS \dataoutbuffer_reg[7][0]  ( .D(n2610), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4700) );
  DFFNSRXLTS \dataoutbuffer_reg[6][31]  ( .D(n2611), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4423) );
  DFFNSRXLTS \dataoutbuffer_reg[6][29]  ( .D(n2613), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4442) );
  DFFNSRXLTS \dataoutbuffer_reg[6][27]  ( .D(n2615), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4459) );
  DFFNSRXLTS \dataoutbuffer_reg[6][26]  ( .D(n2616), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4470) );
  DFFNSRXLTS \dataoutbuffer_reg[6][25]  ( .D(n2617), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4480) );
  DFFNSRXLTS \dataoutbuffer_reg[6][24]  ( .D(n2618), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4490) );
  DFFNSRXLTS \dataoutbuffer_reg[6][23]  ( .D(n2619), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4492) );
  DFFNSRXLTS \dataoutbuffer_reg[6][22]  ( .D(n2620), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4508) );
  DFFNSRXLTS \dataoutbuffer_reg[6][21]  ( .D(n2621), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4512) );
  DFFNSRXLTS \dataoutbuffer_reg[6][20]  ( .D(n2622), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4519) );
  DFFNSRXLTS \dataoutbuffer_reg[6][19]  ( .D(n2623), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4531) );
  DFFNSRXLTS \dataoutbuffer_reg[6][17]  ( .D(n2625), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4553) );
  DFFNSRXLTS \dataoutbuffer_reg[6][16]  ( .D(n2626), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4558) );
  DFFNSRXLTS \dataoutbuffer_reg[6][15]  ( .D(n2627), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4571) );
  DFFNSRXLTS \dataoutbuffer_reg[6][13]  ( .D(n2629), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4586) );
  DFFNSRXLTS \dataoutbuffer_reg[6][12]  ( .D(n2630), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4597) );
  DFFNSRXLTS \dataoutbuffer_reg[6][11]  ( .D(n2631), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4607) );
  DFFNSRXLTS \dataoutbuffer_reg[6][8]  ( .D(n2634), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4634) );
  DFFNSRXLTS \dataoutbuffer_reg[6][7]  ( .D(n2635), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4639) );
  DFFNSRXLTS empty_reg_reg ( .D(n2885), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        n6248), .QN(n4830) );
  DFFNSRXLTS \write_reg_reg[0]  ( .D(n2888), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n9), .QN(n5327) );
  DFFNSRXLTS \write_reg_reg[2]  ( .D(n2886), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n6), .QN(n5326) );
  INVX2TS U2 ( .A(selectBit_NORTH), .Y(n6246) );
  XOR2X4TS U3 ( .A(n5314), .B(n189), .Y(n5388) );
  CLKINVX2TS U4 ( .A(n5312), .Y(n6328) );
  NOR2XLTS U5 ( .A(n5323), .B(n5312), .Y(n5313) );
  AOI222X1TS U6 ( .A0(n4103), .A1(n3339), .B0(n3318), .B1(n160), .C0(n3948), 
        .C1(n3298), .Y(n5423) );
  NOR2BXLTS U7 ( .AN(n5520), .B(n238), .Y(n6118) );
  CLKBUFX2TS U8 ( .A(n3469), .Y(n3465) );
  CLKBUFX2TS U9 ( .A(n3470), .Y(n3467) );
  INVX2TS U10 ( .A(n5388), .Y(n6335) );
  NOR2X2TS U11 ( .A(n6244), .B(n481), .Y(n5316) );
  AOI21X1TS U12 ( .A0(n392), .A1(n170), .B0(n474), .Y(n5548) );
  NAND2X1TS U13 ( .A(n6328), .B(n173), .Y(n5515) );
  AOI21X1TS U14 ( .A0(n225), .A1(n201), .B0(n475), .Y(n5555) );
  XNOR2X1TS U15 ( .A(n173), .B(n5316), .Y(n5314) );
  CLKBUFX2TS U16 ( .A(n774), .Y(n763) );
  CLKBUFX2TS U17 ( .A(n3469), .Y(n3468) );
  CLKBUFX2TS U18 ( .A(n775), .Y(n761) );
  CLKBUFX2TS U19 ( .A(n753), .Y(n750) );
  CLKBUFX2TS U20 ( .A(n775), .Y(n762) );
  NAND2BX1TS U21 ( .AN(n5366), .B(n5387), .Y(n5535) );
  AOI2BB1X1TS U22 ( .A0N(n467), .A1N(n5413), .B0(n5536), .Y(n5538) );
  OA21XLTS U23 ( .A0(n5437), .A1(n5436), .B0(n5544), .Y(n5543) );
  CLKBUFX2TS U24 ( .A(n5548), .Y(n104) );
  AOI21X1TS U25 ( .A0(n5532), .A1(n5389), .B0(n6337), .Y(n5530) );
  CLKBUFX2TS U26 ( .A(n837), .Y(n836) );
  AOI222XLTS U27 ( .A0(n4284), .A1(n3465), .B0(n4129), .B1(n3442), .C0(n3973), 
        .C1(n6343), .Y(n5461) );
  AOI222XLTS U28 ( .A0(n4278), .A1(n3467), .B0(n4123), .B1(n3440), .C0(n3967), 
        .C1(n3724), .Y(n5463) );
  AOI222XLTS U29 ( .A0(n3899), .A1(n804), .B0(n405), .B1(n779), .C0(n4212), 
        .C1(n768), .Y(n5973) );
  AOI222XLTS U30 ( .A0(n3884), .A1(n800), .B0(n415), .B1(n782), .C0(n4197), 
        .C1(n772), .Y(n5983) );
  AOI222XLTS U31 ( .A0(n3878), .A1(n799), .B0(n419), .B1(n782), .C0(n4191), 
        .C1(n777), .Y(n5987) );
  AOI222XLTS U32 ( .A0(n3875), .A1(n799), .B0(n421), .B1(n783), .C0(n4188), 
        .C1(n772), .Y(n5989) );
  AOI222XLTS U33 ( .A0(n3848), .A1(n796), .B0(n439), .B1(n785), .C0(n4161), 
        .C1(n766), .Y(n6007) );
  AOI222XLTS U34 ( .A0(n3842), .A1(n796), .B0(n443), .B1(n785), .C0(n4155), 
        .C1(n765), .Y(n6011) );
  AOI222XLTS U35 ( .A0(n3833), .A1(n795), .B0(n449), .B1(n786), .C0(n4146), 
        .C1(n765), .Y(n6017) );
  AOI222XLTS U36 ( .A0(n3824), .A1(n795), .B0(n455), .B1(n786), .C0(n4137), 
        .C1(n764), .Y(n6023) );
  OAI211X1TS U37 ( .A0(n4713), .A1(n813), .B0(n5355), .C0(n5354), .Y(n2473) );
  AOI222XLTS U38 ( .A0(n3948), .A1(n801), .B0(n790), .B1(n162), .C0(n4260), 
        .C1(n774), .Y(n5354) );
  AOI222XLTS U39 ( .A0(n3911), .A1(n806), .B0(n397), .B1(n780), .C0(n4224), 
        .C1(n769), .Y(n5965) );
  AOI222XLTS U40 ( .A0(n3908), .A1(n806), .B0(n400), .B1(n779), .C0(n4221), 
        .C1(n769), .Y(n5967) );
  AOI222XLTS U41 ( .A0(n3905), .A1(n804), .B0(n402), .B1(n780), .C0(n4218), 
        .C1(n769), .Y(n5969) );
  AOI222XLTS U42 ( .A0(n3902), .A1(n805), .B0(n403), .B1(n779), .C0(n4215), 
        .C1(n769), .Y(n5971) );
  AOI222XLTS U43 ( .A0(n3896), .A1(n805), .B0(n407), .B1(n781), .C0(n4209), 
        .C1(n768), .Y(n5975) );
  AOI222XLTS U44 ( .A0(n3893), .A1(n800), .B0(n409), .B1(n781), .C0(n4206), 
        .C1(n768), .Y(n5977) );
  AOI222XLTS U45 ( .A0(n3890), .A1(n800), .B0(n411), .B1(n780), .C0(n4203), 
        .C1(n768), .Y(n5979) );
  AOI222XLTS U46 ( .A0(n3887), .A1(n800), .B0(n414), .B1(n782), .C0(n4200), 
        .C1(n772), .Y(n5981) );
  AOI222XLTS U47 ( .A0(n3881), .A1(n799), .B0(n418), .B1(n780), .C0(n4194), 
        .C1(n771), .Y(n5985) );
  AOI222XLTS U48 ( .A0(n3872), .A1(n798), .B0(n423), .B1(n781), .C0(n4185), 
        .C1(n773), .Y(n5991) );
  AOI222XLTS U49 ( .A0(n3869), .A1(n798), .B0(n425), .B1(n783), .C0(n4182), 
        .C1(n771), .Y(n5993) );
  AOI222XLTS U50 ( .A0(n3866), .A1(n798), .B0(n428), .B1(n779), .C0(n4179), 
        .C1(n772), .Y(n5995) );
  AOI222XLTS U51 ( .A0(n3863), .A1(n798), .B0(n430), .B1(n782), .C0(n4176), 
        .C1(n767), .Y(n5997) );
  AOI222XLTS U52 ( .A0(n3860), .A1(n797), .B0(n431), .B1(n781), .C0(n4173), 
        .C1(n767), .Y(n5999) );
  AOI222XLTS U53 ( .A0(n3857), .A1(n797), .B0(n434), .B1(n784), .C0(n4170), 
        .C1(n767), .Y(n6001) );
  AOI222XLTS U54 ( .A0(n3854), .A1(n797), .B0(n436), .B1(n783), .C0(n4167), 
        .C1(n766), .Y(n6003) );
  AOI222XLTS U55 ( .A0(n3851), .A1(n797), .B0(n438), .B1(n785), .C0(n4164), 
        .C1(n766), .Y(n6005) );
  AOI222XLTS U56 ( .A0(n3845), .A1(n799), .B0(n441), .B1(n784), .C0(n4158), 
        .C1(n766), .Y(n6009) );
  AOI222XLTS U57 ( .A0(n3839), .A1(n796), .B0(n445), .B1(n784), .C0(n4152), 
        .C1(n765), .Y(n6013) );
  AOI222XLTS U58 ( .A0(n3836), .A1(n796), .B0(n448), .B1(n784), .C0(n4149), 
        .C1(n767), .Y(n6015) );
  AOI222XLTS U59 ( .A0(n3830), .A1(n795), .B0(n451), .B1(n786), .C0(n4143), 
        .C1(n765), .Y(n6019) );
  AOI222XLTS U60 ( .A0(n3827), .A1(n795), .B0(n453), .B1(n785), .C0(n4140), 
        .C1(n764), .Y(n6021) );
  AOI222XLTS U61 ( .A0(n3821), .A1(n794), .B0(n457), .B1(n786), .C0(n4134), 
        .C1(n764), .Y(n6025) );
  AOI222XLTS U62 ( .A0(n4068), .A1(n3528), .B0(n398), .B1(n3509), .C0(n4224), 
        .C1(n3501), .Y(n5581) );
  AOI222XLTS U63 ( .A0(n4065), .A1(n3528), .B0(n400), .B1(n3509), .C0(n4221), 
        .C1(n3506), .Y(n5583) );
  AOI222XLTS U64 ( .A0(n4062), .A1(n3527), .B0(n402), .B1(n3520), .C0(n4218), 
        .C1(n3503), .Y(n5585) );
  AOI222XLTS U65 ( .A0(n4059), .A1(n3527), .B0(n404), .B1(n3520), .C0(n4215), 
        .C1(n3505), .Y(n5587) );
  AOI222XLTS U66 ( .A0(n4056), .A1(n3527), .B0(n406), .B1(n3520), .C0(n4212), 
        .C1(n3501), .Y(n5589) );
  AOI222XLTS U67 ( .A0(n4053), .A1(n3527), .B0(n408), .B1(n3518), .C0(n4209), 
        .C1(n3505), .Y(n5591) );
  AOI222XLTS U68 ( .A0(n4050), .A1(n3526), .B0(n409), .B1(n3519), .C0(n4206), 
        .C1(n3507), .Y(n5593) );
  AOI222XLTS U69 ( .A0(n4047), .A1(n3526), .B0(n412), .B1(n3518), .C0(n4203), 
        .C1(n3503), .Y(n5595) );
  AOI222XLTS U70 ( .A0(n4044), .A1(n3526), .B0(n414), .B1(n3516), .C0(n4200), 
        .C1(n3502), .Y(n5597) );
  AOI222XLTS U71 ( .A0(n4041), .A1(n3526), .B0(n416), .B1(n3522), .C0(n4197), 
        .C1(n3502), .Y(n5599) );
  AOI222XLTS U72 ( .A0(n4038), .A1(n3525), .B0(n418), .B1(n3519), .C0(n4194), 
        .C1(n3501), .Y(n5601) );
  AOI222XLTS U73 ( .A0(n4035), .A1(n3525), .B0(n420), .B1(n3521), .C0(n4191), 
        .C1(n3506), .Y(n5603) );
  AOI222XLTS U74 ( .A0(n4032), .A1(n3525), .B0(n422), .B1(n3516), .C0(n4188), 
        .C1(n3504), .Y(n5605) );
  AOI222XLTS U75 ( .A0(n4029), .A1(n3539), .B0(n423), .B1(n3521), .C0(n4185), 
        .C1(n3502), .Y(n5607) );
  AOI222XLTS U76 ( .A0(n4026), .A1(n6214), .B0(n426), .B1(n3510), .C0(n4182), 
        .C1(n3504), .Y(n5609) );
  AOI222XLTS U77 ( .A0(n4023), .A1(n6214), .B0(n428), .B1(n3510), .C0(n4179), 
        .C1(n3502), .Y(n5611) );
  AOI222XLTS U78 ( .A0(n4011), .A1(n3535), .B0(n436), .B1(n3511), .C0(n4167), 
        .C1(n3498), .Y(n5619) );
  AOI222XLTS U79 ( .A0(n4008), .A1(n3537), .B0(n438), .B1(n3511), .C0(n4164), 
        .C1(n3498), .Y(n5621) );
  AOI222XLTS U80 ( .A0(n4005), .A1(n3536), .B0(n440), .B1(n3511), .C0(n4161), 
        .C1(n3498), .Y(n5623) );
  AOI222XLTS U81 ( .A0(n4002), .A1(n3534), .B0(n442), .B1(n3512), .C0(n4158), 
        .C1(n3498), .Y(n5625) );
  AOI222XLTS U82 ( .A0(n3999), .A1(n3537), .B0(n444), .B1(n3512), .C0(n4155), 
        .C1(n3497), .Y(n5627) );
  AOI222XLTS U83 ( .A0(n3996), .A1(n3534), .B0(n446), .B1(n3512), .C0(n4152), 
        .C1(n3497), .Y(n5629) );
  AOI222XLTS U84 ( .A0(n3993), .A1(n3536), .B0(n448), .B1(n3512), .C0(n4149), 
        .C1(n3497), .Y(n5631) );
  AOI222XLTS U85 ( .A0(n3990), .A1(n3536), .B0(n450), .B1(n3513), .C0(n4146), 
        .C1(n3497), .Y(n5633) );
  AOI222XLTS U86 ( .A0(n3987), .A1(n3536), .B0(n451), .B1(n3513), .C0(n4143), 
        .C1(n3496), .Y(n5635) );
  AOI222XLTS U87 ( .A0(n3984), .A1(n3533), .B0(n454), .B1(n3513), .C0(n4140), 
        .C1(n3496), .Y(n5637) );
  AOI222XLTS U88 ( .A0(n3981), .A1(n3524), .B0(n456), .B1(n3513), .C0(n4137), 
        .C1(n3496), .Y(n5639) );
  AOI222XLTS U89 ( .A0(n3978), .A1(n3524), .B0(n458), .B1(n3514), .C0(n4134), 
        .C1(n3496), .Y(n5641) );
  AOI222XLTS U90 ( .A0(n3818), .A1(n794), .B0(n460), .B1(n783), .C0(n4131), 
        .C1(n764), .Y(n6027) );
  AOI222XLTS U91 ( .A0(n4281), .A1(n3467), .B0(n4126), .B1(n3441), .C0(n3970), 
        .C1(n3724), .Y(n5462) );
  AOI222XLTS U92 ( .A0(n4275), .A1(n3467), .B0(n4120), .B1(n3440), .C0(n3964), 
        .C1(n3720), .Y(n5464) );
  INVX2TS U93 ( .A(n5535), .Y(n6333) );
  CLKBUFX2TS U94 ( .A(n475), .Y(n695) );
  OA22X1TS U95 ( .A0(n5538), .A1(n128), .B0(n226), .B1(n169), .Y(n478) );
  OR2X2TS U96 ( .A(n6221), .B(n216), .Y(n1) );
  NOR2BX1TS U97 ( .AN(n5548), .B(n5515), .Y(n6180) );
  AND3XLTS U98 ( .A(n5545), .B(n5517), .C(n5520), .Y(n6117) );
  INVX2TS U99 ( .A(n5435), .Y(n386) );
  INVX1TS U100 ( .A(n237), .Y(n238) );
  INVXLTS U101 ( .A(n5544), .Y(n6336) );
  AND3X2TS U102 ( .A(n200), .B(n5544), .C(n5548), .Y(n6182) );
  AND2XLTS U103 ( .A(n5548), .B(n6336), .Y(n6179) );
  AOI221X2TS U104 ( .A0(n6332), .A1(n5389), .B0(n249), .B1(n5459), .C0(n5522), 
        .Y(n5524) );
  AOI21X2TS U105 ( .A0(n6333), .A1(n5389), .B0(n6341), .Y(n5512) );
  NOR2X1TS U106 ( .A(n236), .B(n6327), .Y(n5389) );
  CLKINVX1TS U107 ( .A(n188), .Y(n189) );
  INVX1TS U108 ( .A(n5317), .Y(n188) );
  INVX2TS U109 ( .A(n235), .Y(n236) );
  OA21X1TS U110 ( .A0(n5528), .A1(n5413), .B0(n5512), .Y(n5508) );
  INVX2TS U111 ( .A(n115), .Y(n117) );
  INVX2TS U112 ( .A(n110), .Y(n111) );
  XOR2XLTS U113 ( .A(n4861), .B(n189), .Y(n4853) );
  OAI21X2TS U114 ( .A0(n5483), .A1(n204), .B0(n5414), .Y(n5536) );
  NAND3X1TS U115 ( .A(n5460), .B(n5435), .C(n6335), .Y(n5414) );
  NAND3X1TS U116 ( .A(n5482), .B(n5388), .C(n6334), .Y(n5531) );
  AND3XLTS U117 ( .A(n5460), .B(n5388), .C(n6334), .Y(n5522) );
  CLKBUFX2TS U118 ( .A(n3505), .Y(n3495) );
  CLKBUFX2TS U119 ( .A(n3503), .Y(n3499) );
  CLKBUFX2TS U120 ( .A(n6117), .Y(n759) );
  CLKBUFX2TS U121 ( .A(n6349), .Y(n3783) );
  CLKBUFX2TS U122 ( .A(n6163), .Y(n3293) );
  CLKBUFX2TS U123 ( .A(n6343), .Y(n3724) );
  OA22X1TS U124 ( .A0(n5550), .A1(n127), .B0(n224), .B1(n227), .Y(n475) );
  CLKBUFX2TS U125 ( .A(n6103), .Y(n715) );
  CLKBUFX2TS U126 ( .A(n6133), .Y(n844) );
  OA22X1TS U127 ( .A0(n5556), .A1(n127), .B0(n224), .B1(n5484), .Y(n477) );
  OA22X1TS U128 ( .A0(n5543), .A1(n128), .B0(n5484), .B1(n169), .Y(n474) );
  CLKBUFX2TS U129 ( .A(n6120), .Y(n808) );
  XOR2X2TS U130 ( .A(n5318), .B(n6), .Y(n5435) );
  OAI21X1TS U131 ( .A0(n5313), .A1(n466), .B0(n6326), .Y(n5437) );
  NAND2X1TS U132 ( .A(n470), .B(n5392), .Y(n5527) );
  NOR2BX1TS U133 ( .AN(n5343), .B(n6231), .Y(n5482) );
  CLKBUFX2TS U134 ( .A(n3342), .Y(n3336) );
  CLKBUFX2TS U135 ( .A(n3293), .Y(n3286) );
  AOI21X1TS U136 ( .A0(n202), .A1(n223), .B0(n6347), .Y(n5319) );
  CLKBUFX2TS U137 ( .A(n3532), .Y(n3530) );
  CLKBUFX2TS U138 ( .A(n3505), .Y(n3494) );
  CLKBUFX2TS U139 ( .A(n3308), .Y(n3297) );
  OA21XLTS U140 ( .A0(n6327), .A1(n5436), .B0(n5517), .Y(n5516) );
  NAND3X1TS U141 ( .A(n389), .B(n5482), .C(n6334), .Y(n5517) );
  INVX2TS U142 ( .A(n107), .Y(n108) );
  NOR3X1TS U143 ( .A(n5551), .B(n5552), .C(n5549), .Y(n5550) );
  CLKBUFX2TS U144 ( .A(n3308), .Y(n3298) );
  CLKBUFX2TS U145 ( .A(n3341), .Y(n3335) );
  CLKBUFX2TS U146 ( .A(n3408), .Y(n3403) );
  NAND2X1TS U147 ( .A(n5524), .B(n192), .Y(n5571) );
  INVX2TS U148 ( .A(n12), .Y(n192) );
  AOI222XLTS U149 ( .A0(n3840), .A1(n3711), .B0(n445), .B1(n3447), .C0(n3996), 
        .C1(n3429), .Y(n5693) );
  AOI222XLTS U150 ( .A0(n3843), .A1(n3711), .B0(n443), .B1(n3447), .C0(n3999), 
        .C1(n3429), .Y(n5691) );
  AOI222XLTS U151 ( .A0(n3852), .A1(n3712), .B0(n437), .B1(n3448), .C0(n4008), 
        .C1(n3430), .Y(n5685) );
  AOI222XLTS U152 ( .A0(n3855), .A1(n3712), .B0(n435), .B1(n3448), .C0(n4011), 
        .C1(n3430), .Y(n5683) );
  AOI222XLTS U153 ( .A0(n3858), .A1(n3713), .B0(n433), .B1(n3448), .C0(n4014), 
        .C1(n3431), .Y(n5681) );
  AOI222XLTS U154 ( .A0(n3864), .A1(n3713), .B0(n429), .B1(n3456), .C0(n4020), 
        .C1(n3431), .Y(n5677) );
  AOI222XLTS U155 ( .A0(n3867), .A1(n3713), .B0(n427), .B1(n3453), .C0(n4023), 
        .C1(n3432), .Y(n5675) );
  AOI222XLTS U156 ( .A0(n3870), .A1(n3714), .B0(n425), .B1(n3454), .C0(n4026), 
        .C1(n3432), .Y(n5673) );
  AOI222XLTS U157 ( .A0(n3876), .A1(n3714), .B0(n421), .B1(n3457), .C0(n4032), 
        .C1(n3432), .Y(n5669) );
  AOI222XLTS U158 ( .A0(n3879), .A1(n3714), .B0(n420), .B1(n3457), .C0(n4035), 
        .C1(n3433), .Y(n5667) );
  AOI222XLTS U159 ( .A0(n3882), .A1(n3715), .B0(n417), .B1(n3454), .C0(n4038), 
        .C1(n3433), .Y(n5665) );
  AOI222XLTS U160 ( .A0(n3885), .A1(n3715), .B0(n415), .B1(n3449), .C0(n4041), 
        .C1(n3433), .Y(n5663) );
  AOI222XLTS U161 ( .A0(n3888), .A1(n3715), .B0(n413), .B1(n3449), .C0(n4044), 
        .C1(n3433), .Y(n5661) );
  AOI222XLTS U162 ( .A0(n3891), .A1(n3716), .B0(n411), .B1(n3449), .C0(n4047), 
        .C1(n3434), .Y(n5659) );
  AOI222XLTS U163 ( .A0(n3894), .A1(n3716), .B0(n410), .B1(n3449), .C0(n4050), 
        .C1(n3434), .Y(n5657) );
  AOI222XLTS U164 ( .A0(n3897), .A1(n3716), .B0(n407), .B1(n3450), .C0(n4053), 
        .C1(n3434), .Y(n5655) );
  AOI222XLTS U165 ( .A0(n3900), .A1(n3716), .B0(n405), .B1(n3450), .C0(n4056), 
        .C1(n3434), .Y(n5653) );
  AOI222XLTS U166 ( .A0(n3906), .A1(n3717), .B0(n401), .B1(n3450), .C0(n4062), 
        .C1(n3435), .Y(n5649) );
  AOI222XLTS U167 ( .A0(n3912), .A1(n3717), .B0(n397), .B1(n3451), .C0(n4068), 
        .C1(n3435), .Y(n5645) );
  AOI222XLTS U168 ( .A0(n3975), .A1(n3524), .B0(n459), .B1(n3514), .C0(n4131), 
        .C1(n3495), .Y(n5643) );
  AOI222XLTS U169 ( .A0(n4014), .A1(n3533), .B0(n434), .B1(n3511), .C0(n4170), 
        .C1(n3499), .Y(n5617) );
  AOI222XLTS U170 ( .A0(n4017), .A1(n3535), .B0(n432), .B1(n3510), .C0(n4173), 
        .C1(n3499), .Y(n5615) );
  AOI222XLTS U171 ( .A0(n4020), .A1(n3535), .B0(n430), .B1(n3510), .C0(n4176), 
        .C1(n3499), .Y(n5613) );
  AOI222XLTS U172 ( .A0(n794), .A1(n3929), .B0(n787), .B1(n162), .C0(n770), 
        .C1(n4242), .Y(n6107) );
  AOI222XLTS U173 ( .A0(n3849), .A1(n3712), .B0(n440), .B1(n3448), .C0(n4005), 
        .C1(n3430), .Y(n5687) );
  AOI222XLTS U174 ( .A0(n3837), .A1(n3711), .B0(n447), .B1(n3447), .C0(n3993), 
        .C1(n3431), .Y(n5695) );
  AOI222XLTS U175 ( .A0(n3822), .A1(n3710), .B0(n457), .B1(n3445), .C0(n3978), 
        .C1(n3428), .Y(n5705) );
  AOI222XLTS U176 ( .A0(n3909), .A1(n3717), .B0(n399), .B1(n3451), .C0(n4065), 
        .C1(n3435), .Y(n5647) );
  AOI222XLTS U177 ( .A0(n3903), .A1(n3717), .B0(n403), .B1(n3450), .C0(n4059), 
        .C1(n3435), .Y(n5651) );
  AOI222XLTS U178 ( .A0(n3861), .A1(n3713), .B0(n431), .B1(n3456), .C0(n4017), 
        .C1(n3431), .Y(n5679) );
  AOI222XLTS U179 ( .A0(n3846), .A1(n3712), .B0(n441), .B1(n3447), .C0(n4002), 
        .C1(n3430), .Y(n5689) );
  AOI222XLTS U180 ( .A0(n3834), .A1(n3711), .B0(n449), .B1(n3446), .C0(n3990), 
        .C1(n3429), .Y(n5697) );
  AOI222XLTS U181 ( .A0(n3828), .A1(n3710), .B0(n453), .B1(n3446), .C0(n3984), 
        .C1(n3428), .Y(n5701) );
  AOI222XLTS U182 ( .A0(n3825), .A1(n3710), .B0(n455), .B1(n3446), .C0(n3981), 
        .C1(n3428), .Y(n5703) );
  AOI222XLTS U183 ( .A0(n3819), .A1(n3715), .B0(n459), .B1(n3445), .C0(n3975), 
        .C1(n3428), .Y(n5707) );
  AOI222XLTS U184 ( .A0(n3873), .A1(n3714), .B0(n424), .B1(n3457), .C0(n4029), 
        .C1(n3432), .Y(n5671) );
  AOI222XLTS U185 ( .A0(n3831), .A1(n3710), .B0(n452), .B1(n3446), .C0(n3987), 
        .C1(n3429), .Y(n5699) );
  AOI222XLTS U186 ( .A0(n4067), .A1(n3401), .B0(n398), .B1(n3378), .C0(n4224), 
        .C1(n247), .Y(n5709) );
  AOI222XLTS U187 ( .A0(n4022), .A1(n3397), .B0(n427), .B1(n3390), .C0(n4179), 
        .C1(n323), .Y(n5739) );
  AOI222XLTS U188 ( .A0(n4019), .A1(n3397), .B0(n429), .B1(n3380), .C0(n4176), 
        .C1(n248), .Y(n5741) );
  AOI222XLTS U189 ( .A0(n4007), .A1(n3396), .B0(n437), .B1(n3382), .C0(n4164), 
        .C1(n244), .Y(n5749) );
  AOI222XLTS U190 ( .A0(n3977), .A1(n3393), .B0(n458), .B1(n3383), .C0(n4134), 
        .C1(n333), .Y(n5769) );
  AOI222XLTS U191 ( .A0(n4064), .A1(n3401), .B0(n399), .B1(n3390), .C0(n4221), 
        .C1(n244), .Y(n5711) );
  AOI222XLTS U192 ( .A0(n4061), .A1(n3400), .B0(n401), .B1(n3378), .C0(n4218), 
        .C1(n321), .Y(n5713) );
  AOI222XLTS U193 ( .A0(n4058), .A1(n3400), .B0(n404), .B1(n3389), .C0(n4215), 
        .C1(n323), .Y(n5715) );
  AOI222XLTS U194 ( .A0(n4055), .A1(n3400), .B0(n406), .B1(n3390), .C0(n4212), 
        .C1(n247), .Y(n5717) );
  AOI222XLTS U195 ( .A0(n4052), .A1(n3400), .B0(n408), .B1(n3379), .C0(n4209), 
        .C1(n243), .Y(n5719) );
  AOI222XLTS U196 ( .A0(n4049), .A1(n3399), .B0(n410), .B1(n3379), .C0(n4206), 
        .C1(n322), .Y(n5721) );
  AOI222XLTS U197 ( .A0(n4046), .A1(n3399), .B0(n412), .B1(n3378), .C0(n4203), 
        .C1(n322), .Y(n5723) );
  AOI222XLTS U198 ( .A0(n4043), .A1(n3399), .B0(n413), .B1(n3380), .C0(n4200), 
        .C1(n248), .Y(n5725) );
  AOI222XLTS U199 ( .A0(n4040), .A1(n3399), .B0(n416), .B1(n3380), .C0(n4197), 
        .C1(n244), .Y(n5727) );
  AOI222XLTS U200 ( .A0(n4037), .A1(n3398), .B0(n417), .B1(n3378), .C0(n4194), 
        .C1(n323), .Y(n5729) );
  AOI222XLTS U201 ( .A0(n4034), .A1(n3398), .B0(n419), .B1(n3380), .C0(n4191), 
        .C1(n321), .Y(n5731) );
  AOI222XLTS U202 ( .A0(n4031), .A1(n3398), .B0(n422), .B1(n3381), .C0(n4188), 
        .C1(n248), .Y(n5733) );
  AOI222XLTS U203 ( .A0(n4028), .A1(n3397), .B0(n424), .B1(n3379), .C0(n4185), 
        .C1(n243), .Y(n5735) );
  AOI222XLTS U204 ( .A0(n4025), .A1(n3397), .B0(n426), .B1(n3381), .C0(n4182), 
        .C1(n321), .Y(n5737) );
  AOI222XLTS U205 ( .A0(n4016), .A1(n3396), .B0(n432), .B1(n3379), .C0(n4173), 
        .C1(n243), .Y(n5743) );
  AOI222XLTS U206 ( .A0(n4013), .A1(n3396), .B0(n433), .B1(n3389), .C0(n4170), 
        .C1(n323), .Y(n5745) );
  AOI222XLTS U207 ( .A0(n4010), .A1(n3396), .B0(n435), .B1(n3381), .C0(n4167), 
        .C1(n248), .Y(n5747) );
  AOI222XLTS U208 ( .A0(n4004), .A1(n3395), .B0(n439), .B1(n3382), .C0(n4161), 
        .C1(n322), .Y(n5751) );
  AOI222XLTS U209 ( .A0(n4001), .A1(n3398), .B0(n442), .B1(n3387), .C0(n4158), 
        .C1(n322), .Y(n5753) );
  AOI222XLTS U210 ( .A0(n3998), .A1(n3395), .B0(n444), .B1(n3382), .C0(n4155), 
        .C1(n305), .Y(n5755) );
  AOI222XLTS U211 ( .A0(n3995), .A1(n3395), .B0(n446), .B1(n3387), .C0(n4152), 
        .C1(n304), .Y(n5757) );
  AOI222XLTS U212 ( .A0(n3992), .A1(n3395), .B0(n447), .B1(n3391), .C0(n4149), 
        .C1(n321), .Y(n5759) );
  AOI222XLTS U213 ( .A0(n3989), .A1(n3394), .B0(n450), .B1(n3383), .C0(n4146), 
        .C1(n332), .Y(n5761) );
  AOI222XLTS U214 ( .A0(n3986), .A1(n3394), .B0(n452), .B1(n3383), .C0(n4143), 
        .C1(n332), .Y(n5763) );
  AOI222XLTS U215 ( .A0(n3983), .A1(n3394), .B0(n454), .B1(n3382), .C0(n4140), 
        .C1(n247), .Y(n5765) );
  AOI222XLTS U216 ( .A0(n3980), .A1(n3394), .B0(n456), .B1(n3383), .C0(n4137), 
        .C1(n243), .Y(n5767) );
  AOI222XLTS U217 ( .A0(n3974), .A1(n3393), .B0(n460), .B1(n3381), .C0(n4131), 
        .C1(n334), .Y(n5771) );
  AOI222XLTS U218 ( .A0(n3799), .A1(n3369), .B0(n3813), .B1(n334), .C0(n3805), 
        .C1(n6182), .Y(n5575) );
  AOI222XLTS U219 ( .A0(n3972), .A1(n3376), .B0(n4285), .B1(n333), .C0(n4128), 
        .C1(n3405), .Y(n5438) );
  INVX2TS U220 ( .A(n5568), .Y(n181) );
  INVX2TS U221 ( .A(n5568), .Y(n186) );
  INVX2TS U222 ( .A(n3768), .Y(n378) );
  AND2X2TS U223 ( .A(n5538), .B(n5541), .Y(n2) );
  CLKINVX2TS U224 ( .A(n3769), .Y(n335) );
  INVX2TS U225 ( .A(n171), .Y(n127) );
  CLKINVX2TS U226 ( .A(n172), .Y(n126) );
  CLKINVX2TS U227 ( .A(n6180), .Y(n376) );
  CLKINVX1TS U228 ( .A(n6180), .Y(n242) );
  OAI22X1TS U229 ( .A0(n5508), .A1(n127), .B0(n227), .B1(n6321), .Y(n5565) );
  INVX2TS U230 ( .A(n373), .Y(n220) );
  AOI221X1TS U231 ( .A0(n225), .A1(n5344), .B0(n6325), .B1(n249), .C0(n223), 
        .Y(n5528) );
  CLKBUFX2TS U232 ( .A(n3294), .Y(n3285) );
  OR3X1TS U233 ( .A(n302), .B(n216), .C(n388), .Y(n8) );
  XOR2X1TS U234 ( .A(n5344), .B(n219), .Y(n10) );
  AND2X2TS U235 ( .A(n300), .B(n171), .Y(n11) );
  AO21X2TS U236 ( .A0(n201), .A1(n5390), .B0(n220), .Y(n12) );
  OR2X1TS U237 ( .A(n5509), .B(n6348), .Y(n13) );
  OR2X2TS U238 ( .A(n4832), .B(n5310), .Y(n14) );
  INVX2TS U239 ( .A(n5522), .Y(n195) );
  INVX2TS U240 ( .A(n5528), .Y(n187) );
  INVX2TS U241 ( .A(n5545), .Y(n199) );
  NOR2BX1TS U242 ( .AN(n165), .B(n5387), .Y(n5545) );
  CLKINVX2TS U243 ( .A(n293), .Y(n294) );
  OR2X2TS U244 ( .A(n6230), .B(n9), .Y(n15) );
  CLKINVX2TS U245 ( .A(n5555), .Y(n107) );
  INVXLTS U246 ( .A(n5562), .Y(n105) );
  INVXLTS U247 ( .A(n105), .Y(n106) );
  AOI21X1TS U248 ( .A0(n392), .A1(n225), .B0(n477), .Y(n5562) );
  CLKBUFX2TS U249 ( .A(n5541), .Y(n109) );
  AOI21X1TS U250 ( .A0(n202), .A1(n5446), .B0(n478), .Y(n5541) );
  CLKBUFX2TS U251 ( .A(n13), .Y(n110) );
  CLKBUFX2TS U252 ( .A(n13), .Y(n384) );
  INVXLTS U253 ( .A(n110), .Y(n112) );
  INVX2TS U254 ( .A(n384), .Y(n125) );
  INVXLTS U255 ( .A(n110), .Y(n113) );
  INVXLTS U256 ( .A(n384), .Y(n114) );
  INVX2TS U257 ( .A(n125), .Y(n115) );
  INVXLTS U258 ( .A(n115), .Y(n116) );
  INVXLTS U259 ( .A(n115), .Y(n118) );
  INVXLTS U260 ( .A(n115), .Y(n119) );
  INVXLTS U261 ( .A(n13), .Y(n120) );
  INVXLTS U262 ( .A(n384), .Y(n121) );
  INVXLTS U263 ( .A(n13), .Y(n122) );
  INVXLTS U264 ( .A(n110), .Y(n123) );
  INVXLTS U265 ( .A(n384), .Y(n124) );
  CLKINVX1TS U266 ( .A(n171), .Y(n128) );
  INVXLTS U267 ( .A(n6325), .Y(n129) );
  INVXLTS U268 ( .A(n159), .Y(n130) );
  CLKBUFX2TS U269 ( .A(readReady), .Y(n131) );
  CLKBUFX2TS U270 ( .A(selectBit_WEST), .Y(n132) );
  CLKBUFX2TS U271 ( .A(selectBit_NORTH), .Y(n133) );
  INVXLTS U272 ( .A(readRequesterAddress[0]), .Y(n134) );
  INVXLTS U273 ( .A(n134), .Y(n135) );
  INVXLTS U274 ( .A(n134), .Y(n136) );
  INVXLTS U275 ( .A(n134), .Y(n137) );
  INVXLTS U276 ( .A(n134), .Y(n138) );
  INVXLTS U277 ( .A(readRequesterAddress[1]), .Y(n139) );
  INVXLTS U278 ( .A(n139), .Y(n140) );
  INVXLTS U279 ( .A(n139), .Y(n141) );
  INVXLTS U280 ( .A(n139), .Y(n142) );
  INVXLTS U281 ( .A(n139), .Y(n143) );
  INVXLTS U282 ( .A(readRequesterAddress[2]), .Y(n144) );
  INVXLTS U283 ( .A(n144), .Y(n145) );
  INVXLTS U284 ( .A(n144), .Y(n146) );
  INVXLTS U285 ( .A(n144), .Y(n147) );
  INVXLTS U286 ( .A(n144), .Y(n148) );
  INVXLTS U287 ( .A(readRequesterAddress[3]), .Y(n149) );
  INVXLTS U288 ( .A(n149), .Y(n150) );
  INVXLTS U289 ( .A(n149), .Y(n151) );
  INVXLTS U290 ( .A(n149), .Y(n152) );
  INVXLTS U291 ( .A(n149), .Y(n153) );
  INVXLTS U292 ( .A(readRequesterAddress[4]), .Y(n154) );
  INVXLTS U293 ( .A(n154), .Y(n155) );
  INVXLTS U294 ( .A(n154), .Y(n156) );
  INVXLTS U295 ( .A(n154), .Y(n157) );
  INVXLTS U296 ( .A(n154), .Y(n158) );
  INVXLTS U297 ( .A(readRequesterAddress[5]), .Y(n159) );
  INVXLTS U298 ( .A(n159), .Y(n160) );
  INVXLTS U299 ( .A(n159), .Y(n161) );
  INVXLTS U300 ( .A(n159), .Y(n162) );
  INVXLTS U301 ( .A(n3), .Y(n163) );
  INVXLTS U302 ( .A(n5), .Y(n164) );
  INVXLTS U303 ( .A(n10), .Y(n165) );
  INVXLTS U304 ( .A(n10), .Y(n166) );
  INVXLTS U305 ( .A(n5390), .Y(n167) );
  INVXLTS U306 ( .A(n167), .Y(n168) );
  INVXLTS U307 ( .A(n5446), .Y(n169) );
  INVXLTS U308 ( .A(n169), .Y(n170) );
  INVXLTS U309 ( .A(n14), .Y(n171) );
  INVX1TS U310 ( .A(n14), .Y(n172) );
  INVXLTS U311 ( .A(n219), .Y(n173) );
  INVX1TS U312 ( .A(n380), .Y(n174) );
  CLKINVX1TS U313 ( .A(n174), .Y(n175) );
  CLKINVX1TS U314 ( .A(n174), .Y(n176) );
  CLKINVX1TS U315 ( .A(n174), .Y(n177) );
  CLKINVX1TS U316 ( .A(n174), .Y(n178) );
  INVXLTS U317 ( .A(n379), .Y(n179) );
  CLKINVX1TS U318 ( .A(n182), .Y(n180) );
  INVX2TS U319 ( .A(n186), .Y(n182) );
  CLKINVX1TS U320 ( .A(n182), .Y(n183) );
  CLKINVX1TS U321 ( .A(n182), .Y(n184) );
  CLKINVX1TS U322 ( .A(n182), .Y(n185) );
  INVX2TS U323 ( .A(n5568), .Y(n380) );
  INVX2TS U324 ( .A(n5565), .Y(n190) );
  INVXLTS U325 ( .A(n190), .Y(n191) );
  INVXLTS U326 ( .A(n12), .Y(n193) );
  CLKBUFX2TS U327 ( .A(n5520), .Y(n194) );
  INVXLTS U328 ( .A(n195), .Y(n196) );
  CLKBUFX2TS U329 ( .A(n5508), .Y(n197) );
  INVXLTS U330 ( .A(n6329), .Y(n198) );
  INVXLTS U331 ( .A(n199), .Y(n200) );
  INVXLTS U332 ( .A(n15), .Y(n201) );
  INVXLTS U333 ( .A(n15), .Y(n202) );
  CLKBUFX2TS U334 ( .A(n5527), .Y(n203) );
  NOR3X1TS U335 ( .A(n6338), .B(n5528), .C(n5527), .Y(n6148) );
  CLKINVX1TS U336 ( .A(n6333), .Y(n204) );
  INVXLTS U337 ( .A(n8), .Y(n205) );
  INVXLTS U338 ( .A(n8), .Y(n206) );
  INVXLTS U339 ( .A(n1), .Y(n207) );
  INVXLTS U340 ( .A(n5565), .Y(n208) );
  INVXLTS U341 ( .A(n335), .Y(n209) );
  INVXLTS U342 ( .A(n336), .Y(n210) );
  INVX1TS U343 ( .A(n6234), .Y(n211) );
  CLKINVX1TS U344 ( .A(n211), .Y(n212) );
  NOR3X1TS U345 ( .A(n187), .B(n218), .C(n5312), .Y(n5557) );
  INVXLTS U346 ( .A(n4839), .Y(n213) );
  INVXLTS U347 ( .A(n6233), .Y(n214) );
  INVXLTS U348 ( .A(n214), .Y(n215) );
  INVXLTS U349 ( .A(n385), .Y(n216) );
  INVXLTS U350 ( .A(n388), .Y(n217) );
  INVXLTS U351 ( .A(n393), .Y(n218) );
  INVXLTS U352 ( .A(n218), .Y(n219) );
  INVXLTS U353 ( .A(n220), .Y(n221) );
  INVXLTS U354 ( .A(n220), .Y(n222) );
  INVXLTS U355 ( .A(n6321), .Y(n223) );
  INVXLTS U356 ( .A(n5494), .Y(n224) );
  INVXLTS U357 ( .A(n224), .Y(n225) );
  INVXLTS U358 ( .A(n11), .Y(n226) );
  INVXLTS U359 ( .A(n11), .Y(n227) );
  INVXLTS U360 ( .A(n335), .Y(n228) );
  INVXLTS U361 ( .A(n5565), .Y(n229) );
  INVXLTS U362 ( .A(n335), .Y(n230) );
  INVXLTS U363 ( .A(n335), .Y(n231) );
  INVXLTS U364 ( .A(n337), .Y(n232) );
  INVXLTS U365 ( .A(n232), .Y(n233) );
  CLKBUFX2TS U366 ( .A(n4868), .Y(n234) );
  INVX2TS U367 ( .A(n6232), .Y(n235) );
  INVXLTS U368 ( .A(n5515), .Y(n237) );
  INVX2TS U369 ( .A(n292), .Y(n329) );
  INVX2TS U370 ( .A(n329), .Y(n239) );
  INVX1TS U371 ( .A(n239), .Y(n240) );
  CLKINVX2TS U372 ( .A(n239), .Y(n241) );
  INVXLTS U373 ( .A(n242), .Y(n243) );
  INVXLTS U374 ( .A(n242), .Y(n244) );
  INVXLTS U375 ( .A(n5283), .Y(n245) );
  INVXLTS U376 ( .A(n245), .Y(n246) );
  INVXLTS U377 ( .A(n376), .Y(n247) );
  INVXLTS U378 ( .A(n376), .Y(n248) );
  INVXLTS U379 ( .A(n6), .Y(n249) );
  INVXLTS U380 ( .A(n5570), .Y(n250) );
  INVXLTS U381 ( .A(n258), .Y(n251) );
  INVXLTS U382 ( .A(n291), .Y(n252) );
  INVXLTS U383 ( .A(n3665), .Y(n253) );
  INVXLTS U384 ( .A(n5566), .Y(n254) );
  INVXLTS U385 ( .A(n254), .Y(n255) );
  INVXLTS U386 ( .A(n254), .Y(n256) );
  INVXLTS U387 ( .A(n221), .Y(n257) );
  INVXLTS U388 ( .A(n339), .Y(n258) );
  INVXLTS U389 ( .A(n258), .Y(n259) );
  INVXLTS U390 ( .A(n258), .Y(n260) );
  INVXLTS U391 ( .A(n258), .Y(n261) );
  INVXLTS U392 ( .A(n6235), .Y(n262) );
  INVXLTS U393 ( .A(n262), .Y(n263) );
  INVXLTS U394 ( .A(n262), .Y(n264) );
  INVXLTS U395 ( .A(n6236), .Y(n265) );
  INVXLTS U396 ( .A(n265), .Y(n266) );
  INVXLTS U397 ( .A(n265), .Y(n267) );
  INVXLTS U398 ( .A(n6237), .Y(n268) );
  INVXLTS U399 ( .A(n268), .Y(n269) );
  INVXLTS U400 ( .A(n268), .Y(n270) );
  INVXLTS U401 ( .A(n6242), .Y(n271) );
  INVXLTS U402 ( .A(n271), .Y(n272) );
  INVXLTS U403 ( .A(n271), .Y(n273) );
  INVXLTS U404 ( .A(n6240), .Y(n274) );
  INVXLTS U405 ( .A(n274), .Y(n275) );
  INVXLTS U406 ( .A(n274), .Y(n276) );
  INVXLTS U407 ( .A(n6239), .Y(n277) );
  INVXLTS U408 ( .A(n277), .Y(n278) );
  INVXLTS U409 ( .A(n277), .Y(n279) );
  INVXLTS U410 ( .A(n6243), .Y(n280) );
  INVXLTS U411 ( .A(n280), .Y(n281) );
  INVXLTS U412 ( .A(n280), .Y(n282) );
  INVXLTS U413 ( .A(n6241), .Y(n283) );
  INVXLTS U414 ( .A(n283), .Y(n284) );
  INVXLTS U415 ( .A(n283), .Y(n285) );
  INVXLTS U416 ( .A(n6238), .Y(n286) );
  INVXLTS U417 ( .A(n286), .Y(n287) );
  INVXLTS U418 ( .A(n286), .Y(n288) );
  INVXLTS U419 ( .A(n5578), .Y(n289) );
  INVXLTS U420 ( .A(n289), .Y(n290) );
  INVXLTS U421 ( .A(n289), .Y(n291) );
  INVXLTS U422 ( .A(n289), .Y(n292) );
  INVX2TS U423 ( .A(n5571), .Y(n293) );
  INVXLTS U424 ( .A(n293), .Y(n295) );
  INVXLTS U425 ( .A(n340), .Y(n296) );
  INVXLTS U426 ( .A(n296), .Y(n297) );
  INVXLTS U427 ( .A(n296), .Y(n298) );
  INVXLTS U428 ( .A(n296), .Y(n299) );
  INVXLTS U429 ( .A(n9), .Y(n300) );
  INVXLTS U430 ( .A(n7), .Y(n301) );
  INVXLTS U431 ( .A(n7), .Y(n302) );
  INVXLTS U432 ( .A(n242), .Y(n303) );
  INVXLTS U433 ( .A(n320), .Y(n304) );
  INVXLTS U434 ( .A(n242), .Y(n305) );
  INVXLTS U435 ( .A(n342), .Y(n306) );
  INVXLTS U436 ( .A(n309), .Y(n307) );
  INVXLTS U437 ( .A(n342), .Y(n308) );
  INVXLTS U438 ( .A(n344), .Y(n309) );
  INVXLTS U439 ( .A(n309), .Y(n310) );
  INVXLTS U440 ( .A(n309), .Y(n311) );
  INVXLTS U441 ( .A(n309), .Y(n312) );
  INVXLTS U442 ( .A(n2), .Y(n313) );
  INVXLTS U443 ( .A(n313), .Y(n314) );
  INVXLTS U444 ( .A(n313), .Y(n315) );
  INVXLTS U445 ( .A(n313), .Y(n316) );
  INVXLTS U446 ( .A(n5578), .Y(n317) );
  INVXLTS U447 ( .A(n239), .Y(n318) );
  INVXLTS U448 ( .A(n5578), .Y(n319) );
  INVXLTS U449 ( .A(n6180), .Y(n320) );
  INVXLTS U450 ( .A(n320), .Y(n321) );
  INVXLTS U451 ( .A(n320), .Y(n322) );
  INVXLTS U452 ( .A(n320), .Y(n323) );
  INVX2TS U453 ( .A(n289), .Y(n324) );
  INVX2TS U454 ( .A(n324), .Y(n325) );
  INVXLTS U455 ( .A(n324), .Y(n326) );
  INVXLTS U456 ( .A(n324), .Y(n327) );
  INVXLTS U457 ( .A(n324), .Y(n328) );
  INVX2TS U458 ( .A(n6180), .Y(n330) );
  INVXLTS U459 ( .A(n330), .Y(n331) );
  INVXLTS U460 ( .A(n330), .Y(n332) );
  INVXLTS U461 ( .A(n330), .Y(n333) );
  INVXLTS U462 ( .A(n330), .Y(n334) );
  INVXLTS U463 ( .A(n190), .Y(n336) );
  INVXLTS U464 ( .A(n336), .Y(n337) );
  INVXLTS U465 ( .A(n336), .Y(n338) );
  INVXLTS U466 ( .A(n373), .Y(n339) );
  INVXLTS U467 ( .A(n373), .Y(n340) );
  INVXLTS U468 ( .A(n222), .Y(n341) );
  INVXLTS U469 ( .A(n2), .Y(n342) );
  CLKINVX1TS U470 ( .A(n342), .Y(n343) );
  CLKINVX1TS U471 ( .A(n342), .Y(n344) );
  OAI21X1TS U498 ( .A0(n5391), .A1(n128), .B0(n471), .Y(n470) );
  AOI21X1TS U499 ( .A0(n5485), .A1(n5353), .B0(n476), .Y(n5520) );
  CLKBUFX2TS U500 ( .A(n5580), .Y(n371) );
  CLKBUFX2TS U501 ( .A(n5580), .Y(n372) );
  NAND3X1TS U502 ( .A(n5482), .B(n5435), .C(n389), .Y(n5544) );
  NAND2XLTS U503 ( .A(n5550), .B(n5555), .Y(n5578) );
  OAI22X1TS U504 ( .A0(n5524), .A1(n127), .B0(n226), .B1(n167), .Y(n373) );
  OAI22X1TS U505 ( .A0(n5524), .A1(n14), .B0(n226), .B1(n167), .Y(n5570) );
  AOI32X1TS U506 ( .A0(n6232), .A1(n6234), .A2(n133), .B0(n4835), .B1(
        selectBit_SOUTH), .Y(n4836) );
  XNOR2X1TS U507 ( .A(selectBit_NORTH), .B(selectBit_EAST), .Y(n4835) );
  NAND2XLTS U508 ( .A(n5549), .B(n5555), .Y(n6200) );
  INVX1TS U509 ( .A(selectBit_SOUTH), .Y(n6234) );
  NAND2X1TS U510 ( .A(n6327), .B(selectBit_EAST), .Y(n5483) );
  OAI2BB1X1TS U511 ( .A0N(n4868), .A1N(selectBit_EAST), .B0(n4836), .Y(n4839)
         );
  CLKBUFX2TS U512 ( .A(n5576), .Y(n374) );
  CLKBUFX2TS U513 ( .A(n5576), .Y(n375) );
  OAI22X1TS U514 ( .A0(n6246), .A1(n212), .B0(n4868), .B1(n6232), .Y(n5317) );
  NOR2X1TS U515 ( .A(n212), .B(n5311), .Y(n5511) );
  CLKINVX2TS U516 ( .A(n3768), .Y(n377) );
  INVX1TS U517 ( .A(n186), .Y(n379) );
  NOR3BX1TS U518 ( .AN(n109), .B(n5536), .C(n6329), .Y(n6163) );
  CLKINVX2TS U519 ( .A(n3739), .Y(n381) );
  CLKINVX2TS U520 ( .A(n3739), .Y(n382) );
  OAI22X1TS U521 ( .A0(n197), .A1(n128), .B0(n227), .B1(n6321), .Y(n383) );
  NOR3BX1TS U522 ( .AN(n193), .B(n5521), .C(n196), .Y(n6133) );
  NOR3BX1TS U523 ( .AN(n5482), .B(n386), .C(n389), .Y(n5558) );
  NOR3BX1TS U524 ( .AN(n5460), .B(n386), .C(n389), .Y(n5549) );
  NAND3X1TS U525 ( .A(n6335), .B(n5460), .C(n6334), .Y(n5509) );
  INVX3TS U526 ( .A(n5435), .Y(n6334) );
  CLKBUFX2TS U527 ( .A(n6228), .Y(n387) );
  INVX1TS U528 ( .A(n5388), .Y(n389) );
  OR2X2TS U529 ( .A(n5301), .B(n6247), .Y(n5279) );
  INVX2TS U530 ( .A(n5279), .Y(n390) );
  INVX2TS U531 ( .A(n5279), .Y(n391) );
  CLKBUFX2TS U532 ( .A(n5485), .Y(n392) );
  OAI31XLTS U533 ( .A0(n5485), .A1(n6328), .A2(n129), .B0(n172), .Y(n5484) );
  INVX2TS U534 ( .A(n3719), .Y(n394) );
  INVX1TS U535 ( .A(n6200), .Y(n6343) );
  INVX2TS U536 ( .A(n5291), .Y(n395) );
  INVX2TS U537 ( .A(n3680), .Y(n396) );
  CLKBUFX2TS U538 ( .A(cacheDataOut[31]), .Y(n397) );
  CLKBUFX2TS U539 ( .A(cacheDataOut[31]), .Y(n398) );
  CLKBUFX2TS U540 ( .A(cacheDataOut[30]), .Y(n399) );
  CLKBUFX2TS U541 ( .A(cacheDataOut[30]), .Y(n400) );
  CLKBUFX2TS U542 ( .A(cacheDataOut[29]), .Y(n401) );
  CLKBUFX2TS U543 ( .A(cacheDataOut[29]), .Y(n402) );
  CLKBUFX2TS U544 ( .A(cacheDataOut[28]), .Y(n403) );
  CLKBUFX2TS U545 ( .A(cacheDataOut[28]), .Y(n404) );
  CLKBUFX2TS U546 ( .A(cacheDataOut[27]), .Y(n405) );
  CLKBUFX2TS U547 ( .A(cacheDataOut[27]), .Y(n406) );
  CLKBUFX2TS U548 ( .A(cacheDataOut[26]), .Y(n407) );
  CLKBUFX2TS U549 ( .A(cacheDataOut[26]), .Y(n408) );
  CLKBUFX2TS U550 ( .A(cacheDataOut[25]), .Y(n409) );
  CLKBUFX2TS U551 ( .A(cacheDataOut[25]), .Y(n410) );
  CLKBUFX2TS U552 ( .A(cacheDataOut[24]), .Y(n411) );
  CLKBUFX2TS U553 ( .A(cacheDataOut[24]), .Y(n412) );
  CLKBUFX2TS U554 ( .A(cacheDataOut[23]), .Y(n413) );
  CLKBUFX2TS U555 ( .A(cacheDataOut[23]), .Y(n414) );
  CLKBUFX2TS U556 ( .A(cacheDataOut[22]), .Y(n415) );
  CLKBUFX2TS U557 ( .A(cacheDataOut[22]), .Y(n416) );
  CLKBUFX2TS U558 ( .A(cacheDataOut[21]), .Y(n417) );
  CLKBUFX2TS U559 ( .A(cacheDataOut[21]), .Y(n418) );
  CLKBUFX2TS U560 ( .A(cacheDataOut[20]), .Y(n419) );
  CLKBUFX2TS U561 ( .A(cacheDataOut[20]), .Y(n420) );
  CLKBUFX2TS U562 ( .A(cacheDataOut[19]), .Y(n421) );
  CLKBUFX2TS U563 ( .A(cacheDataOut[19]), .Y(n422) );
  CLKBUFX2TS U564 ( .A(cacheDataOut[18]), .Y(n423) );
  CLKBUFX2TS U565 ( .A(cacheDataOut[18]), .Y(n424) );
  CLKBUFX2TS U566 ( .A(cacheDataOut[17]), .Y(n425) );
  CLKBUFX2TS U567 ( .A(cacheDataOut[17]), .Y(n426) );
  CLKBUFX2TS U568 ( .A(cacheDataOut[16]), .Y(n427) );
  CLKBUFX2TS U569 ( .A(cacheDataOut[16]), .Y(n428) );
  CLKBUFX2TS U570 ( .A(cacheDataOut[15]), .Y(n429) );
  CLKBUFX2TS U571 ( .A(cacheDataOut[15]), .Y(n430) );
  CLKBUFX2TS U572 ( .A(cacheDataOut[14]), .Y(n431) );
  CLKBUFX2TS U573 ( .A(cacheDataOut[14]), .Y(n432) );
  CLKBUFX2TS U574 ( .A(cacheDataOut[13]), .Y(n433) );
  CLKBUFX2TS U575 ( .A(cacheDataOut[13]), .Y(n434) );
  CLKBUFX2TS U576 ( .A(cacheDataOut[12]), .Y(n435) );
  CLKBUFX2TS U577 ( .A(cacheDataOut[12]), .Y(n436) );
  CLKBUFX2TS U578 ( .A(cacheDataOut[11]), .Y(n437) );
  CLKBUFX2TS U579 ( .A(cacheDataOut[11]), .Y(n438) );
  CLKBUFX2TS U580 ( .A(cacheDataOut[10]), .Y(n439) );
  CLKBUFX2TS U581 ( .A(cacheDataOut[10]), .Y(n440) );
  CLKBUFX2TS U582 ( .A(cacheDataOut[9]), .Y(n441) );
  CLKBUFX2TS U583 ( .A(cacheDataOut[9]), .Y(n442) );
  CLKBUFX2TS U584 ( .A(cacheDataOut[8]), .Y(n443) );
  CLKBUFX2TS U585 ( .A(cacheDataOut[8]), .Y(n444) );
  CLKBUFX2TS U586 ( .A(cacheDataOut[7]), .Y(n445) );
  CLKBUFX2TS U587 ( .A(cacheDataOut[7]), .Y(n446) );
  CLKBUFX2TS U588 ( .A(cacheDataOut[6]), .Y(n447) );
  CLKBUFX2TS U589 ( .A(cacheDataOut[6]), .Y(n448) );
  CLKBUFX2TS U590 ( .A(cacheDataOut[5]), .Y(n449) );
  CLKBUFX2TS U591 ( .A(cacheDataOut[5]), .Y(n450) );
  CLKBUFX2TS U592 ( .A(cacheDataOut[4]), .Y(n451) );
  CLKBUFX2TS U593 ( .A(cacheDataOut[4]), .Y(n452) );
  CLKBUFX2TS U594 ( .A(cacheDataOut[3]), .Y(n453) );
  CLKBUFX2TS U595 ( .A(cacheDataOut[3]), .Y(n454) );
  CLKBUFX2TS U596 ( .A(cacheDataOut[2]), .Y(n455) );
  CLKBUFX2TS U597 ( .A(cacheDataOut[2]), .Y(n456) );
  CLKBUFX2TS U598 ( .A(cacheDataOut[1]), .Y(n457) );
  CLKBUFX2TS U599 ( .A(cacheDataOut[1]), .Y(n458) );
  CLKBUFX2TS U600 ( .A(cacheDataOut[0]), .Y(n459) );
  CLKBUFX2TS U601 ( .A(cacheDataOut[0]), .Y(n460) );
  CLKBUFX2TS U602 ( .A(n6217), .Y(n461) );
  CLKBUFX2TS U603 ( .A(n6217), .Y(n462) );
  CLKBUFX2TS U604 ( .A(n5572), .Y(n463) );
  CLKBUFX2TS U605 ( .A(n5572), .Y(n464) );
  NOR3X1TS U606 ( .A(n6331), .B(n6337), .C(n203), .Y(n5572) );
  INVX2TS U607 ( .A(n5437), .Y(n6327) );
  AND2XLTS U608 ( .A(n5508), .B(n5319), .Y(n465) );
  OR2XLTS U609 ( .A(n5527), .B(n467), .Y(n472) );
  CLKINVX2TS U610 ( .A(n5565), .Y(n6347) );
  NOR3XLTS U611 ( .A(n5535), .B(n6341), .C(n6348), .Y(n5563) );
  AND3XLTS U612 ( .A(n5541), .B(n6333), .C(n5414), .Y(n6166) );
  AND2XLTS U613 ( .A(n5541), .B(n6340), .Y(n6164) );
  INVXLTS U614 ( .A(n5319), .Y(n6348) );
  INVX1TS U615 ( .A(n5572), .Y(n6346) );
  CLKBUFX2TS U616 ( .A(n6211), .Y(n3490) );
  CLKINVX2TS U617 ( .A(n5532), .Y(n6331) );
  NOR2X1TS U618 ( .A(n5531), .B(n5527), .Y(n6150) );
  INVX2TS U619 ( .A(n3221), .Y(n471) );
  AND2XLTS U620 ( .A(n5559), .B(n5562), .Y(n6214) );
  AND2XLTS U621 ( .A(n5562), .B(n5557), .Y(n6212) );
  NOR2XLTS U622 ( .A(n5343), .B(n6231), .Y(n5460) );
  AND2XLTS U623 ( .A(n392), .B(n172), .Y(n5495) );
  NAND2XLTS U624 ( .A(n172), .B(n4418), .Y(n6228) );
  INVXLTS U625 ( .A(selectBit_WEST), .Y(n6231) );
  OAI31XLTS U626 ( .A0(n4831), .A1(n5310), .A2(n5309), .B0(n5308), .Y(n2450)
         );
  OAI31XLTS U627 ( .A0(n4829), .A1(n5310), .A2(n5309), .B0(n5293), .Y(n2449)
         );
  INVXLTS U628 ( .A(n187), .Y(n466) );
  INVX2TS U629 ( .A(n466), .Y(n467) );
  INVXLTS U630 ( .A(n6349), .Y(n468) );
  INVXLTS U631 ( .A(n6349), .Y(n469) );
  INVXLTS U632 ( .A(n3192), .Y(n1728) );
  INVXLTS U633 ( .A(n1894), .Y(n1764) );
  INVXLTS U634 ( .A(n1822), .Y(n1817) );
  INVXLTS U635 ( .A(n3359), .Y(n3355) );
  INVXLTS U636 ( .A(n3359), .Y(n3354) );
  CLKBUFX2TS U637 ( .A(n828), .Y(n824) );
  CLKBUFX2TS U638 ( .A(n694), .Y(n691) );
  CLKBUFX2TS U639 ( .A(n694), .Y(n690) );
  CLKBUFX2TS U640 ( .A(n3360), .Y(n3357) );
  CLKBUFX2TS U641 ( .A(n828), .Y(n826) );
  CLKBUFX2TS U642 ( .A(n3426), .Y(n3423) );
  CLKBUFX2TS U643 ( .A(n3557), .Y(n3554) );
  CLKBUFX2TS U644 ( .A(n3360), .Y(n3358) );
  CLKBUFX2TS U645 ( .A(n3426), .Y(n3424) );
  CLKBUFX2TS U646 ( .A(n3557), .Y(n3555) );
  NAND3XLTS U647 ( .A(n106), .B(n6326), .C(n5556), .Y(n5580) );
  NOR2XLTS U648 ( .A(n6329), .B(n165), .Y(n5459) );
  CLKAND2X2TS U649 ( .A(n193), .B(n5459), .Y(n6135) );
  AND2XLTS U650 ( .A(n196), .B(n193), .Y(n473) );
  CLKBUFX2TS U651 ( .A(n677), .Y(n672) );
  NAND3XLTS U652 ( .A(n194), .B(n238), .C(n5516), .Y(n5568) );
  NAND3XLTS U653 ( .A(n104), .B(n5515), .C(n5543), .Y(n5576) );
  NOR2XLTS U654 ( .A(n166), .B(n5387), .Y(n5532) );
  NAND2XLTS U655 ( .A(n5387), .B(n5366), .Y(n5521) );
  NAND2XLTS U656 ( .A(n5511), .B(n165), .Y(n5413) );
  AND2XLTS U657 ( .A(n5551), .B(n108), .Y(n6197) );
  AND2XLTS U658 ( .A(n5552), .B(n5555), .Y(n6195) );
  NOR2X1TS U659 ( .A(n393), .B(n6), .Y(n5353) );
  XOR2XLTS U660 ( .A(n300), .B(n6244), .Y(n5343) );
  NOR2X1TS U661 ( .A(n6246), .B(n300), .Y(n5344) );
  AOI21XLTS U662 ( .A0(n212), .A1(n5311), .B0(n5511), .Y(n5387) );
  AOI32XLTS U663 ( .A0(n104), .A1(n5547), .A2(n5546), .B0(n3425), .B1(n19), 
        .Y(n2568) );
  AOI32XLTS U664 ( .A0(n5545), .A1(n5544), .A2(n3808), .B0(n5543), .B1(n5542), 
        .Y(n5546) );
  AOI32XLTS U665 ( .A0(n194), .A1(n5519), .A2(n5518), .B0(n824), .B1(n16), .Y(
        n2564) );
  AOI32XLTS U666 ( .A0(n5545), .A1(n5517), .A2(n3809), .B0(n5516), .B1(n5542), 
        .Y(n5518) );
  AND2XLTS U667 ( .A(n4868), .B(n4866), .Y(n5310) );
  INVXLTS U668 ( .A(n5344), .Y(n6325) );
  AND2XLTS U669 ( .A(n4867), .B(n236), .Y(n4866) );
  INVXLTS U670 ( .A(n5521), .Y(n6332) );
  OAI32XLTS U671 ( .A0(n3811), .A1(n196), .A2(n5521), .B0(n6330), .B1(n215), 
        .Y(n5523) );
  NOR2X1TS U672 ( .A(n6230), .B(n5327), .Y(n5485) );
  NOR2X1TS U673 ( .A(n249), .B(n5323), .Y(n5494) );
  NOR2X1TS U674 ( .A(n6), .B(n173), .Y(n5390) );
  NOR2X1TS U675 ( .A(n393), .B(n249), .Y(n5446) );
  NOR2X1TS U676 ( .A(n301), .B(n481), .Y(n4841) );
  NOR3X1TS U677 ( .A(n385), .B(n4), .C(n164), .Y(n5282) );
  OAI211XLTS U678 ( .A0(n4087), .A1(n3777), .B0(n6094), .C0(n6093), .Y(n2835)
         );
  OAI211XLTS U679 ( .A0(n4084), .A1(n3777), .B0(n6096), .C0(n6095), .Y(n2836)
         );
  OAI211XLTS U680 ( .A0(n4081), .A1(n3776), .B0(n6098), .C0(n6097), .Y(n2837)
         );
  OAI211XLTS U681 ( .A0(n4078), .A1(n3776), .B0(n6100), .C0(n6099), .Y(n2838)
         );
  OAI211XLTS U682 ( .A0(n4075), .A1(n3776), .B0(n6102), .C0(n6101), .Y(n2839)
         );
  OAI211XLTS U683 ( .A0(n4072), .A1(n3776), .B0(n6106), .C0(n6105), .Y(n2840)
         );
  OAI211XLTS U684 ( .A0(n3781), .A1(n3979), .B0(n6090), .C0(n6089), .Y(n2833)
         );
  OAI211XLTS U685 ( .A0(n3783), .A1(n3976), .B0(n6092), .C0(n6091), .Y(n2834)
         );
  OAI211XLTS U686 ( .A0(n3770), .A1(n4105), .B0(n5332), .C0(n5331), .Y(n2459)
         );
  OAI211XLTS U687 ( .A0(n3770), .A1(n4099), .B0(n5336), .C0(n5335), .Y(n2461)
         );
  OAI211XLTS U688 ( .A0(n3770), .A1(n4096), .B0(n5338), .C0(n5337), .Y(n2462)
         );
  OAI211XLTS U689 ( .A0(n3771), .A1(n4093), .B0(n5340), .C0(n5339), .Y(n2463)
         );
  OAI211XLTS U690 ( .A0(n3771), .A1(n4069), .B0(n6030), .C0(n6029), .Y(n2803)
         );
  OAI211XLTS U691 ( .A0(n3771), .A1(n4066), .B0(n6032), .C0(n6031), .Y(n2804)
         );
  OAI211XLTS U692 ( .A0(n3772), .A1(n4063), .B0(n6034), .C0(n6033), .Y(n2805)
         );
  OAI211XLTS U693 ( .A0(n3772), .A1(n4054), .B0(n6040), .C0(n6039), .Y(n2808)
         );
  OAI211XLTS U694 ( .A0(n3773), .A1(n4051), .B0(n6042), .C0(n6041), .Y(n2809)
         );
  OAI211XLTS U695 ( .A0(n3773), .A1(n4048), .B0(n6044), .C0(n6043), .Y(n2810)
         );
  OAI211XLTS U696 ( .A0(n3773), .A1(n4042), .B0(n6048), .C0(n6047), .Y(n2812)
         );
  OAI211XLTS U697 ( .A0(n3774), .A1(n4039), .B0(n6050), .C0(n6049), .Y(n2813)
         );
  OAI211XLTS U698 ( .A0(n3774), .A1(n4033), .B0(n6054), .C0(n6053), .Y(n2815)
         );
  OAI211XLTS U699 ( .A0(n3774), .A1(n4030), .B0(n6056), .C0(n6055), .Y(n2816)
         );
  OAI211XLTS U700 ( .A0(n3775), .A1(n4027), .B0(n6058), .C0(n6057), .Y(n2817)
         );
  OAI211XLTS U701 ( .A0(n3775), .A1(n4024), .B0(n6060), .C0(n6059), .Y(n2818)
         );
  OAI211XLTS U702 ( .A0(n3775), .A1(n4021), .B0(n6062), .C0(n6061), .Y(n2819)
         );
  OAI211XLTS U703 ( .A0(n3775), .A1(n4018), .B0(n6064), .C0(n6063), .Y(n2820)
         );
  OAI211XLTS U704 ( .A0(n3780), .A1(n4015), .B0(n6066), .C0(n6065), .Y(n2821)
         );
  OAI211XLTS U705 ( .A0(n3779), .A1(n4012), .B0(n6068), .C0(n6067), .Y(n2822)
         );
  OAI211XLTS U706 ( .A0(n3782), .A1(n4009), .B0(n6070), .C0(n6069), .Y(n2823)
         );
  OAI211XLTS U707 ( .A0(n3778), .A1(n4006), .B0(n6072), .C0(n6071), .Y(n2824)
         );
  OAI211XLTS U708 ( .A0(n3777), .A1(n4000), .B0(n6076), .C0(n6075), .Y(n2826)
         );
  OAI211XLTS U709 ( .A0(n3780), .A1(n3997), .B0(n6078), .C0(n6077), .Y(n2827)
         );
  OAI211XLTS U710 ( .A0(n3779), .A1(n3994), .B0(n6080), .C0(n6079), .Y(n2828)
         );
  OAI211XLTS U711 ( .A0(n3778), .A1(n3988), .B0(n6084), .C0(n6083), .Y(n2830)
         );
  OAI211XLTS U712 ( .A0(n3781), .A1(n3985), .B0(n6086), .C0(n6085), .Y(n2831)
         );
  OAI211XLTS U713 ( .A0(n3770), .A1(n4102), .B0(n5334), .C0(n5333), .Y(n2460)
         );
  OAI211XLTS U714 ( .A0(n3771), .A1(n4090), .B0(n5342), .C0(n5341), .Y(n2464)
         );
  OAI211XLTS U715 ( .A0(n3772), .A1(n4060), .B0(n6036), .C0(n6035), .Y(n2806)
         );
  OAI211XLTS U716 ( .A0(n3772), .A1(n4057), .B0(n6038), .C0(n6037), .Y(n2807)
         );
  OAI211XLTS U717 ( .A0(n3773), .A1(n4045), .B0(n6046), .C0(n6045), .Y(n2811)
         );
  OAI211XLTS U718 ( .A0(n3774), .A1(n4036), .B0(n6052), .C0(n6051), .Y(n2814)
         );
  OAI211XLTS U719 ( .A0(n3778), .A1(n4003), .B0(n6074), .C0(n6073), .Y(n2825)
         );
  OAI211XLTS U720 ( .A0(n3783), .A1(n3991), .B0(n6082), .C0(n6081), .Y(n2829)
         );
  OAI211XLTS U721 ( .A0(n3781), .A1(n3982), .B0(n6088), .C0(n6087), .Y(n2832)
         );
  OAI32XLTS U722 ( .A0(n3810), .A1(n6341), .A2(n204), .B0(n5509), .B1(n3804), 
        .Y(n5510) );
  AOI22XLTS U723 ( .A0(n5514), .A1(n5513), .B0(n190), .B1(n6312), .Y(n2563) );
  AOI31XLTS U724 ( .A0(n5512), .A1(n198), .A2(readIn_SOUTH), .B0(n5510), .Y(
        n5513) );
  OAI22XLTS U725 ( .A0(n466), .A1(n215), .B0(n467), .B1(n3817), .Y(n5529) );
  AOI21XLTS U726 ( .A0(n3815), .A1(n5524), .B0(n5523), .Y(n5525) );
  NAND2XLTS U727 ( .A(n3803), .B(n196), .Y(n5526) );
  AOI21XLTS U728 ( .A0(n3815), .A1(n5538), .B0(n5537), .Y(n5539) );
  AOI2BB2XLTS U729 ( .B0(readReady), .B1(selectBit_WEST), .A0N(n4867), .A1N(
        n6244), .Y(n4861) );
  NAND2XLTS U730 ( .A(n5311), .B(selectBit_SOUTH), .Y(n5312) );
  OAI211XLTS U731 ( .A0(n3931), .A1(n6200), .B0(n6186), .C0(n6185), .Y(n2871)
         );
  AOI22XLTS U732 ( .A0(n3445), .A1(n130), .B0(n3439), .B1(n4085), .Y(n6186) );
  OAI211XLTS U733 ( .A0(n3928), .A1(n6200), .B0(n6188), .C0(n6187), .Y(n2872)
         );
  OAI211XLTS U734 ( .A0(n3925), .A1(n394), .B0(n6190), .C0(n6189), .Y(n2873)
         );
  OAI211XLTS U735 ( .A0(n3922), .A1(n394), .B0(n6192), .C0(n6191), .Y(n2874)
         );
  OAI211XLTS U736 ( .A0(n3919), .A1(n394), .B0(n6194), .C0(n6193), .Y(n2875)
         );
  OAI211XLTS U737 ( .A0(n3916), .A1(n394), .B0(n6199), .C0(n6198), .Y(n2876)
         );
  AOI22XLTS U738 ( .A0(n3444), .A1(n136), .B0(n3438), .B1(n4070), .Y(n6199) );
  OAI211XLTS U739 ( .A0(n3344), .A1(n6277), .B0(n6158), .C0(n6157), .Y(n2861)
         );
  OAI211XLTS U740 ( .A0(n3343), .A1(n6278), .B0(n6160), .C0(n6159), .Y(n2862)
         );
  OAI211XLTS U741 ( .A0(n3343), .A1(n6279), .B0(n6162), .C0(n6161), .Y(n2863)
         );
  OAI211XLTS U742 ( .A0(n3344), .A1(n6280), .B0(n6168), .C0(n6167), .Y(n2864)
         );
  OAI211XLTS U743 ( .A0(n3344), .A1(n6301), .B0(n6154), .C0(n6153), .Y(n2859)
         );
  OAI211XLTS U744 ( .A0(n3343), .A1(n6302), .B0(n6156), .C0(n6155), .Y(n2860)
         );
  OAI211XLTS U745 ( .A0(n811), .A1(n6287), .B0(n6112), .C0(n6111), .Y(n2843)
         );
  OAI211XLTS U746 ( .A0(n810), .A1(n6288), .B0(n6114), .C0(n6113), .Y(n2844)
         );
  OAI211XLTS U747 ( .A0(n810), .A1(n6289), .B0(n6116), .C0(n6115), .Y(n2845)
         );
  OAI211XLTS U748 ( .A0(n811), .A1(n6285), .B0(n6108), .C0(n6107), .Y(n2841)
         );
  OAI211XLTS U749 ( .A0(n810), .A1(n6286), .B0(n6110), .C0(n6109), .Y(n2842)
         );
  OAI211XLTS U750 ( .A0(n811), .A1(n6290), .B0(n6122), .C0(n6121), .Y(n2846)
         );
  OAI211XLTS U751 ( .A0(n3541), .A1(n6309), .B0(n6206), .C0(n6205), .Y(n2879)
         );
  OAI211XLTS U752 ( .A0(n3540), .A1(n6310), .B0(n6210), .C0(n6209), .Y(n2881)
         );
  OAI211XLTS U753 ( .A0(n3541), .A1(n6281), .B0(n6202), .C0(n6201), .Y(n2877)
         );
  OAI211XLTS U754 ( .A0(n3540), .A1(n6282), .B0(n6204), .C0(n6203), .Y(n2878)
         );
  OAI211XLTS U755 ( .A0(n3540), .A1(n6283), .B0(n6208), .C0(n6207), .Y(n2880)
         );
  OAI211XLTS U756 ( .A0(n3541), .A1(n6311), .B0(n6216), .C0(n6215), .Y(n2882)
         );
  OAI211XLTS U757 ( .A0(n3410), .A1(n6305), .B0(n6174), .C0(n6173), .Y(n2867)
         );
  OAI211XLTS U758 ( .A0(n3409), .A1(n6306), .B0(n6176), .C0(n6175), .Y(n2868)
         );
  OAI211XLTS U759 ( .A0(n3409), .A1(n6307), .B0(n6178), .C0(n6177), .Y(n2869)
         );
  OAI211XLTS U760 ( .A0(n3410), .A1(n6303), .B0(n6170), .C0(n6169), .Y(n2865)
         );
  OAI211XLTS U761 ( .A0(n3409), .A1(n6304), .B0(n6172), .C0(n6171), .Y(n2866)
         );
  OAI211XLTS U762 ( .A0(n3410), .A1(n6308), .B0(n6184), .C0(n6183), .Y(n2870)
         );
  OAI211XLTS U763 ( .A0(n1764), .A1(n3823), .B0(n5962), .C0(n5961), .Y(n2769)
         );
  OAI211XLTS U764 ( .A0(n1764), .A1(n3820), .B0(n5964), .C0(n5963), .Y(n2770)
         );
  OAI211XLTS U765 ( .A0(n970), .A1(n3940), .B0(n5382), .C0(n5381), .Y(n2490)
         );
  OAI211XLTS U766 ( .A0(n970), .A1(n3946), .B0(n5378), .C0(n5377), .Y(n2488)
         );
  OAI211XLTS U767 ( .A0(n970), .A1(n3943), .B0(n5380), .C0(n5379), .Y(n2489)
         );
  OAI211XLTS U768 ( .A0(n970), .A1(n3949), .B0(n5376), .C0(n5375), .Y(n2487)
         );
  OAI211XLTS U769 ( .A0(n986), .A1(n3910), .B0(n5904), .C0(n5903), .Y(n2740)
         );
  OAI211XLTS U770 ( .A0(n1005), .A1(n3907), .B0(n5906), .C0(n5905), .Y(n2741)
         );
  OAI211XLTS U771 ( .A0(n1005), .A1(n3904), .B0(n5908), .C0(n5907), .Y(n2742)
         );
  OAI211XLTS U772 ( .A0(n1005), .A1(n3898), .B0(n5912), .C0(n5911), .Y(n2744)
         );
  OAI211XLTS U773 ( .A0(n1402), .A1(n3895), .B0(n5914), .C0(n5913), .Y(n2745)
         );
  OAI211XLTS U774 ( .A0(n1402), .A1(n3889), .B0(n5918), .C0(n5917), .Y(n2747)
         );
  OAI211XLTS U775 ( .A0(n1537), .A1(n3883), .B0(n5922), .C0(n5921), .Y(n2749)
         );
  OAI211XLTS U776 ( .A0(n1537), .A1(n3880), .B0(n5924), .C0(n5923), .Y(n2750)
         );
  OAI211XLTS U777 ( .A0(n1537), .A1(n3877), .B0(n5926), .C0(n5925), .Y(n2751)
         );
  OAI211XLTS U778 ( .A0(n1537), .A1(n3874), .B0(n5928), .C0(n5927), .Y(n2752)
         );
  OAI211XLTS U779 ( .A0(n1586), .A1(n3871), .B0(n5930), .C0(n5929), .Y(n2753)
         );
  OAI211XLTS U780 ( .A0(n1586), .A1(n3865), .B0(n5934), .C0(n5933), .Y(n2755)
         );
  OAI211XLTS U781 ( .A0(n1586), .A1(n3862), .B0(n5936), .C0(n5935), .Y(n2756)
         );
  OAI211XLTS U782 ( .A0(n1653), .A1(n3859), .B0(n5938), .C0(n5937), .Y(n2757)
         );
  OAI211XLTS U783 ( .A0(n1653), .A1(n3856), .B0(n5940), .C0(n5939), .Y(n2758)
         );
  OAI211XLTS U784 ( .A0(n1653), .A1(n3853), .B0(n5942), .C0(n5941), .Y(n2759)
         );
  OAI211XLTS U785 ( .A0(n1654), .A1(n3847), .B0(n5946), .C0(n5945), .Y(n2761)
         );
  OAI211XLTS U786 ( .A0(n1654), .A1(n3844), .B0(n5948), .C0(n5947), .Y(n2762)
         );
  OAI211XLTS U787 ( .A0(n1654), .A1(n3841), .B0(n5950), .C0(n5949), .Y(n2763)
         );
  OAI211XLTS U788 ( .A0(n1728), .A1(n3835), .B0(n5954), .C0(n5953), .Y(n2765)
         );
  OAI211XLTS U789 ( .A0(n1728), .A1(n3832), .B0(n5956), .C0(n5955), .Y(n2766)
         );
  OAI211XLTS U790 ( .A0(n1728), .A1(n3829), .B0(n5958), .C0(n5957), .Y(n2767)
         );
  OAI211XLTS U791 ( .A0(n986), .A1(n3937), .B0(n5384), .C0(n5383), .Y(n2491)
         );
  OAI211XLTS U792 ( .A0(n986), .A1(n3934), .B0(n5386), .C0(n5385), .Y(n2492)
         );
  OAI211XLTS U793 ( .A0(n1005), .A1(n3901), .B0(n5910), .C0(n5909), .Y(n2743)
         );
  OAI211XLTS U794 ( .A0(n1653), .A1(n3850), .B0(n5944), .C0(n5943), .Y(n2760)
         );
  OAI211XLTS U795 ( .A0(n986), .A1(n3913), .B0(n5902), .C0(n5901), .Y(n2739)
         );
  OAI211XLTS U796 ( .A0(n1402), .A1(n3892), .B0(n5916), .C0(n5915), .Y(n2746)
         );
  OAI211XLTS U797 ( .A0(n1402), .A1(n3886), .B0(n5920), .C0(n5919), .Y(n2748)
         );
  OAI211XLTS U798 ( .A0(n1586), .A1(n3868), .B0(n5932), .C0(n5931), .Y(n2754)
         );
  OAI211XLTS U799 ( .A0(n1654), .A1(n3838), .B0(n5952), .C0(n5951), .Y(n2764)
         );
  OAI211XLTS U800 ( .A0(n1728), .A1(n3826), .B0(n5960), .C0(n5959), .Y(n2768)
         );
  OAI211XLTS U801 ( .A0(n3928), .A1(n1764), .B0(n6126), .C0(n6125), .Y(n2848)
         );
  OAI211XLTS U802 ( .A0(n3931), .A1(n1764), .B0(n6124), .C0(n6123), .Y(n2847)
         );
  OAI211XLTS U803 ( .A0(n3919), .A1(n1817), .B0(n6132), .C0(n6131), .Y(n2851)
         );
  OAI211XLTS U804 ( .A0(n3916), .A1(n1817), .B0(n6137), .C0(n6136), .Y(n2852)
         );
  OAI211XLTS U805 ( .A0(n3925), .A1(n1817), .B0(n6128), .C0(n6127), .Y(n2849)
         );
  OAI211XLTS U806 ( .A0(n3922), .A1(n1817), .B0(n6130), .C0(n6129), .Y(n2850)
         );
  OAI211XLTS U807 ( .A0(n4087), .A1(n3745), .B0(n6139), .C0(n6138), .Y(n2853)
         );
  OAI211XLTS U808 ( .A0(n4081), .A1(n3746), .B0(n6143), .C0(n6142), .Y(n2855)
         );
  OAI211XLTS U809 ( .A0(n4078), .A1(n3746), .B0(n6145), .C0(n6144), .Y(n2856)
         );
  OAI211XLTS U810 ( .A0(n4075), .A1(n3746), .B0(n6147), .C0(n6146), .Y(n2857)
         );
  OAI211XLTS U811 ( .A0(n4072), .A1(n3746), .B0(n6152), .C0(n6151), .Y(n2858)
         );
  OAI211XLTS U812 ( .A0(n4084), .A1(n3745), .B0(n6141), .C0(n6140), .Y(n2854)
         );
  OAI211XLTS U813 ( .A0(n4725), .A1(n3356), .B0(n5426), .C0(n5425), .Y(n2516)
         );
  INVXLTS U814 ( .A(n3358), .Y(n3356) );
  OAI211XLTS U815 ( .A0(n4714), .A1(n3346), .B0(n5424), .C0(n5423), .Y(n2515)
         );
  OAI211XLTS U816 ( .A0(n4429), .A1(n3354), .B0(n5776), .C0(n5775), .Y(n2676)
         );
  OAI211XLTS U817 ( .A0(n4447), .A1(n3354), .B0(n5780), .C0(n5779), .Y(n2678)
         );
  OAI211XLTS U818 ( .A0(n4458), .A1(n3353), .B0(n5782), .C0(n5781), .Y(n2679)
         );
  OAI211XLTS U819 ( .A0(n4465), .A1(n3353), .B0(n5784), .C0(n5783), .Y(n2680)
         );
  OAI211XLTS U820 ( .A0(n4478), .A1(n3353), .B0(n5786), .C0(n5785), .Y(n2681)
         );
  OAI211XLTS U821 ( .A0(n4483), .A1(n3353), .B0(n5788), .C0(n5787), .Y(n2682)
         );
  OAI211XLTS U822 ( .A0(n4494), .A1(n3352), .B0(n5790), .C0(n5789), .Y(n2683)
         );
  OAI211XLTS U823 ( .A0(n4537), .A1(n3351), .B0(n5800), .C0(n5799), .Y(n2688)
         );
  OAI211XLTS U824 ( .A0(n4582), .A1(n3350), .B0(n5810), .C0(n5809), .Y(n2693)
         );
  OAI211XLTS U825 ( .A0(n4622), .A1(n3349), .B0(n5818), .C0(n5817), .Y(n2697)
         );
  OAI211XLTS U826 ( .A0(n4640), .A1(n3348), .B0(n5822), .C0(n5821), .Y(n2699)
         );
  OAI211XLTS U827 ( .A0(n4656), .A1(n3348), .B0(n5826), .C0(n5825), .Y(n2701)
         );
  OAI211XLTS U828 ( .A0(n4667), .A1(n3348), .B0(n5828), .C0(n5827), .Y(n2702)
         );
  OAI211XLTS U829 ( .A0(n4683), .A1(n3347), .B0(n5832), .C0(n5831), .Y(n2704)
         );
  OAI211XLTS U830 ( .A0(n4421), .A1(n3354), .B0(n5774), .C0(n5773), .Y(n2675)
         );
  OAI211XLTS U831 ( .A0(n4445), .A1(n3354), .B0(n5778), .C0(n5777), .Y(n2677)
         );
  OAI211XLTS U832 ( .A0(n4504), .A1(n3352), .B0(n5792), .C0(n5791), .Y(n2684)
         );
  OAI211XLTS U833 ( .A0(n4515), .A1(n3352), .B0(n5794), .C0(n5793), .Y(n2685)
         );
  OAI211XLTS U834 ( .A0(n4524), .A1(n3352), .B0(n5796), .C0(n5795), .Y(n2686)
         );
  OAI211XLTS U835 ( .A0(n4529), .A1(n3351), .B0(n5798), .C0(n5797), .Y(n2687)
         );
  OAI211XLTS U836 ( .A0(n4556), .A1(n3351), .B0(n5804), .C0(n5803), .Y(n2690)
         );
  OAI211XLTS U837 ( .A0(n4594), .A1(n3349), .B0(n5812), .C0(n5811), .Y(n2694)
         );
  OAI211XLTS U838 ( .A0(n4605), .A1(n3349), .B0(n5814), .C0(n5813), .Y(n2695)
         );
  OAI211XLTS U839 ( .A0(n4612), .A1(n3349), .B0(n5816), .C0(n5815), .Y(n2696)
         );
  OAI211XLTS U840 ( .A0(n4628), .A1(n3348), .B0(n5820), .C0(n5819), .Y(n2698)
         );
  OAI211XLTS U841 ( .A0(n4650), .A1(n3350), .B0(n5824), .C0(n5823), .Y(n2700)
         );
  OAI211XLTS U842 ( .A0(n4691), .A1(n3347), .B0(n5834), .C0(n5833), .Y(n2705)
         );
  OAI211XLTS U843 ( .A0(n4702), .A1(n3347), .B0(n5836), .C0(n5835), .Y(n2706)
         );
  OAI211XLTS U844 ( .A0(n4552), .A1(n3351), .B0(n5802), .C0(n5801), .Y(n2689)
         );
  OAI211XLTS U845 ( .A0(n4570), .A1(n3350), .B0(n5806), .C0(n5805), .Y(n2691)
         );
  OAI211XLTS U846 ( .A0(n4579), .A1(n3350), .B0(n5808), .C0(n5807), .Y(n2692)
         );
  OAI211XLTS U847 ( .A0(n4678), .A1(n3347), .B0(n5830), .C0(n5829), .Y(n2703)
         );
  OAI211XLTS U848 ( .A0(n4734), .A1(n3355), .B0(n5428), .C0(n5427), .Y(n2517)
         );
  OAI211XLTS U849 ( .A0(n4739), .A1(n3355), .B0(n5430), .C0(n5429), .Y(n2518)
         );
  OAI211XLTS U850 ( .A0(n4752), .A1(n3355), .B0(n5432), .C0(n5431), .Y(n2519)
         );
  OAI211XLTS U851 ( .A0(n4757), .A1(n3355), .B0(n5434), .C0(n5433), .Y(n2520)
         );
  OAI211XLTS U852 ( .A0(n4456), .A1(n820), .B0(n5974), .C0(n5973), .Y(n2775)
         );
  OAI211XLTS U853 ( .A0(n4505), .A1(n819), .B0(n5984), .C0(n5983), .Y(n2780)
         );
  OAI211XLTS U854 ( .A0(n4521), .A1(n819), .B0(n5988), .C0(n5987), .Y(n2782)
         );
  OAI211XLTS U855 ( .A0(n4532), .A1(n818), .B0(n5990), .C0(n5989), .Y(n2783)
         );
  OAI211XLTS U856 ( .A0(n4615), .A1(n816), .B0(n6008), .C0(n6007), .Y(n2792)
         );
  OAI211XLTS U857 ( .A0(n4629), .A1(n815), .B0(n6012), .C0(n6011), .Y(n2794)
         );
  OAI211XLTS U858 ( .A0(n4654), .A1(n815), .B0(n6018), .C0(n6017), .Y(n2797)
         );
  OAI211XLTS U859 ( .A0(n4681), .A1(n814), .B0(n6024), .C0(n6023), .Y(n2800)
         );
  OAI211XLTS U860 ( .A0(n4427), .A1(n821), .B0(n5966), .C0(n5965), .Y(n2771)
         );
  OAI211XLTS U861 ( .A0(n4436), .A1(n821), .B0(n5968), .C0(n5967), .Y(n2772)
         );
  OAI211XLTS U862 ( .A0(n4441), .A1(n821), .B0(n5970), .C0(n5969), .Y(n2773)
         );
  OAI211XLTS U863 ( .A0(n4448), .A1(n821), .B0(n5972), .C0(n5971), .Y(n2774)
         );
  OAI211XLTS U864 ( .A0(n4472), .A1(n820), .B0(n5976), .C0(n5975), .Y(n2776)
         );
  OAI211XLTS U865 ( .A0(n4479), .A1(n820), .B0(n5978), .C0(n5977), .Y(n2777)
         );
  OAI211XLTS U866 ( .A0(n4484), .A1(n820), .B0(n5980), .C0(n5979), .Y(n2778)
         );
  OAI211XLTS U867 ( .A0(n4493), .A1(n819), .B0(n5982), .C0(n5981), .Y(n2779)
         );
  OAI211XLTS U868 ( .A0(n4511), .A1(n819), .B0(n5986), .C0(n5985), .Y(n2781)
         );
  OAI211XLTS U869 ( .A0(n4544), .A1(n818), .B0(n5992), .C0(n5991), .Y(n2784)
         );
  OAI211XLTS U870 ( .A0(n4547), .A1(n818), .B0(n5994), .C0(n5993), .Y(n2785)
         );
  OAI211XLTS U871 ( .A0(n4562), .A1(n818), .B0(n5996), .C0(n5995), .Y(n2786)
         );
  OAI211XLTS U872 ( .A0(n4569), .A1(n817), .B0(n5998), .C0(n5997), .Y(n2787)
         );
  OAI211XLTS U873 ( .A0(n4576), .A1(n817), .B0(n6000), .C0(n5999), .Y(n2788)
         );
  OAI211XLTS U874 ( .A0(n4589), .A1(n817), .B0(n6002), .C0(n6001), .Y(n2789)
         );
  OAI211XLTS U875 ( .A0(n4598), .A1(n816), .B0(n6004), .C0(n6003), .Y(n2790)
         );
  OAI211XLTS U876 ( .A0(n4601), .A1(n816), .B0(n6006), .C0(n6005), .Y(n2791)
         );
  OAI211XLTS U877 ( .A0(n4619), .A1(n816), .B0(n6010), .C0(n6009), .Y(n2793)
         );
  OAI211XLTS U878 ( .A0(n4643), .A1(n815), .B0(n6014), .C0(n6013), .Y(n2795)
         );
  OAI211XLTS U879 ( .A0(n4646), .A1(n817), .B0(n6016), .C0(n6015), .Y(n2796)
         );
  OAI211XLTS U880 ( .A0(n4670), .A1(n815), .B0(n6020), .C0(n6019), .Y(n2798)
         );
  OAI211XLTS U881 ( .A0(n4675), .A1(n814), .B0(n6022), .C0(n6021), .Y(n2799)
         );
  OAI211XLTS U882 ( .A0(n4693), .A1(n814), .B0(n6026), .C0(n6025), .Y(n2801)
         );
  OAI211XLTS U883 ( .A0(n4705), .A1(n814), .B0(n6028), .C0(n6027), .Y(n2802)
         );
  OAI211XLTS U884 ( .A0(n4733), .A1(n822), .B0(n5359), .C0(n5358), .Y(n2475)
         );
  OAI211XLTS U885 ( .A0(n4746), .A1(n822), .B0(n5361), .C0(n5360), .Y(n2476)
         );
  OAI211XLTS U886 ( .A0(n4755), .A1(n822), .B0(n5363), .C0(n5362), .Y(n2477)
         );
  OAI211XLTS U887 ( .A0(n4764), .A1(n822), .B0(n5365), .C0(n5364), .Y(n2478)
         );
  OAI211XLTS U888 ( .A0(n4730), .A1(n689), .B0(n5475), .C0(n5474), .Y(n2545)
         );
  OAI211XLTS U889 ( .A0(n4741), .A1(n689), .B0(n5477), .C0(n5476), .Y(n2546)
         );
  OAI211XLTS U890 ( .A0(n4750), .A1(n688), .B0(n5479), .C0(n5478), .Y(n2547)
         );
  OAI211XLTS U891 ( .A0(n4759), .A1(n688), .B0(n5481), .C0(n5480), .Y(n2548)
         );
  OAI211XLTS U892 ( .A0(n4442), .A1(n687), .B0(n5650), .C0(n5649), .Y(n2613)
         );
  OAI211XLTS U893 ( .A0(n4492), .A1(n686), .B0(n5662), .C0(n5661), .Y(n2619)
         );
  OAI211XLTS U894 ( .A0(n4512), .A1(n685), .B0(n5666), .C0(n5665), .Y(n2621)
         );
  OAI211XLTS U895 ( .A0(n4519), .A1(n685), .B0(n5668), .C0(n5667), .Y(n2622)
         );
  OAI211XLTS U896 ( .A0(n4586), .A1(n683), .B0(n5682), .C0(n5681), .Y(n2629)
         );
  OAI211XLTS U897 ( .A0(n4597), .A1(n683), .B0(n5684), .C0(n5683), .Y(n2630)
         );
  OAI211XLTS U898 ( .A0(n4609), .A1(n682), .B0(n5687), .C0(n5688), .Y(n2632)
         );
  OAI211XLTS U899 ( .A0(n4645), .A1(n681), .B0(n5695), .C0(n5696), .Y(n2636)
         );
  OAI211XLTS U900 ( .A0(n4692), .A1(n680), .B0(n5706), .C0(n5705), .Y(n2641)
         );
  AOI22XLTS U901 ( .A0(n4133), .A1(n3458), .B0(n4290), .B1(n329), .Y(n5706) );
  OAI211XLTS U902 ( .A0(n4423), .A1(n688), .B0(n5645), .C0(n5646), .Y(n2611)
         );
  OAI211XLTS U903 ( .A0(n4434), .A1(n688), .B0(n5647), .C0(n5648), .Y(n2612)
         );
  OAI211XLTS U904 ( .A0(n4450), .A1(n687), .B0(n5651), .C0(n5652), .Y(n2614)
         );
  OAI211XLTS U905 ( .A0(n4459), .A1(n687), .B0(n5654), .C0(n5653), .Y(n2615)
         );
  OAI211XLTS U906 ( .A0(n4470), .A1(n687), .B0(n5656), .C0(n5655), .Y(n2616)
         );
  OAI211XLTS U907 ( .A0(n4490), .A1(n686), .B0(n5660), .C0(n5659), .Y(n2618)
         );
  OAI211XLTS U908 ( .A0(n4508), .A1(n686), .B0(n5664), .C0(n5663), .Y(n2620)
         );
  OAI211XLTS U909 ( .A0(n4531), .A1(n685), .B0(n5670), .C0(n5669), .Y(n2623)
         );
  OAI211XLTS U910 ( .A0(n4553), .A1(n684), .B0(n5674), .C0(n5673), .Y(n2625)
         );
  OAI211XLTS U911 ( .A0(n4558), .A1(n684), .B0(n5676), .C0(n5675), .Y(n2626)
         );
  OAI211XLTS U912 ( .A0(n4571), .A1(n684), .B0(n5678), .C0(n5677), .Y(n2627)
         );
  OAI211XLTS U913 ( .A0(n4578), .A1(n683), .B0(n5679), .C0(n5680), .Y(n2628)
         );
  OAI211XLTS U914 ( .A0(n4607), .A1(n683), .B0(n5686), .C0(n5685), .Y(n2631)
         );
  OAI211XLTS U915 ( .A0(n4623), .A1(n682), .B0(n5689), .C0(n5690), .Y(n2633)
         );
  OAI211XLTS U916 ( .A0(n4634), .A1(n682), .B0(n5692), .C0(n5691), .Y(n2634)
         );
  OAI211XLTS U917 ( .A0(n4639), .A1(n682), .B0(n5694), .C0(n5693), .Y(n2635)
         );
  OAI211XLTS U918 ( .A0(n4657), .A1(n681), .B0(n5698), .C0(n5697), .Y(n2637)
         );
  OAI211XLTS U919 ( .A0(n4673), .A1(n681), .B0(n5702), .C0(n5701), .Y(n2639)
         );
  OAI211XLTS U920 ( .A0(n4688), .A1(n680), .B0(n5704), .C0(n5703), .Y(n2640)
         );
  OAI211XLTS U921 ( .A0(n4704), .A1(n685), .B0(n5708), .C0(n5707), .Y(n2642)
         );
  AOI22XLTS U922 ( .A0(n4130), .A1(n3458), .B0(n4287), .B1(n329), .Y(n5708) );
  OAI211XLTS U923 ( .A0(n4480), .A1(n686), .B0(n5658), .C0(n5657), .Y(n2617)
         );
  OAI211XLTS U924 ( .A0(n4543), .A1(n684), .B0(n5671), .C0(n5672), .Y(n2624)
         );
  OAI211XLTS U925 ( .A0(n4669), .A1(n681), .B0(n5700), .C0(n5699), .Y(n2638)
         );
  OAI211XLTS U926 ( .A0(n4716), .A1(n680), .B0(n5471), .C0(n5470), .Y(n2543)
         );
  OAI211XLTS U927 ( .A0(n4727), .A1(n689), .B0(n5473), .C0(n5472), .Y(n2544)
         );
  OAI211XLTS U928 ( .A0(n4719), .A1(n3543), .B0(n5497), .C0(n5496), .Y(n2557)
         );
  OAI211XLTS U929 ( .A0(n4425), .A1(n3551), .B0(n5582), .C0(n5581), .Y(n2579)
         );
  OAI211XLTS U930 ( .A0(n4430), .A1(n3551), .B0(n5584), .C0(n5583), .Y(n2580)
         );
  OAI211XLTS U931 ( .A0(n4439), .A1(n3551), .B0(n5586), .C0(n5585), .Y(n2581)
         );
  OAI211XLTS U932 ( .A0(n4452), .A1(n3551), .B0(n5588), .C0(n5587), .Y(n2582)
         );
  OAI211XLTS U933 ( .A0(n4461), .A1(n3550), .B0(n5590), .C0(n5589), .Y(n2583)
         );
  OAI211XLTS U934 ( .A0(n4468), .A1(n3550), .B0(n5592), .C0(n5591), .Y(n2584)
         );
  OAI211XLTS U935 ( .A0(n4477), .A1(n3550), .B0(n5594), .C0(n5593), .Y(n2585)
         );
  OAI211XLTS U936 ( .A0(n4486), .A1(n3550), .B0(n5596), .C0(n5595), .Y(n2586)
         );
  OAI211XLTS U937 ( .A0(n4497), .A1(n3549), .B0(n5598), .C0(n5597), .Y(n2587)
         );
  OAI211XLTS U938 ( .A0(n4502), .A1(n3549), .B0(n5600), .C0(n5599), .Y(n2588)
         );
  OAI211XLTS U939 ( .A0(n4517), .A1(n3549), .B0(n5602), .C0(n5601), .Y(n2589)
         );
  OAI211XLTS U940 ( .A0(n4522), .A1(n3549), .B0(n5604), .C0(n5603), .Y(n2590)
         );
  OAI211XLTS U941 ( .A0(n4535), .A1(n3548), .B0(n5606), .C0(n5605), .Y(n2591)
         );
  OAI211XLTS U942 ( .A0(n4538), .A1(n3548), .B0(n5608), .C0(n5607), .Y(n2592)
         );
  OAI211XLTS U943 ( .A0(n4549), .A1(n3548), .B0(n5610), .C0(n5609), .Y(n2593)
         );
  OAI211XLTS U944 ( .A0(n4560), .A1(n3548), .B0(n5612), .C0(n5611), .Y(n2594)
         );
  OAI211XLTS U945 ( .A0(n4565), .A1(n3547), .B0(n5614), .C0(n5613), .Y(n2595)
         );
  OAI211XLTS U946 ( .A0(n4580), .A1(n3547), .B0(n5616), .C0(n5615), .Y(n2596)
         );
  OAI211XLTS U947 ( .A0(n4583), .A1(n3547), .B0(n5618), .C0(n5617), .Y(n2597)
         );
  OAI211XLTS U948 ( .A0(n4592), .A1(n3546), .B0(n5620), .C0(n5619), .Y(n2598)
         );
  OAI211XLTS U949 ( .A0(n4603), .A1(n3546), .B0(n5622), .C0(n5621), .Y(n2599)
         );
  OAI211XLTS U950 ( .A0(n4616), .A1(n3546), .B0(n5624), .C0(n5623), .Y(n2600)
         );
  OAI211XLTS U951 ( .A0(n4625), .A1(n3546), .B0(n5626), .C0(n5625), .Y(n2601)
         );
  OAI211XLTS U952 ( .A0(n4630), .A1(n3545), .B0(n5628), .C0(n5627), .Y(n2602)
         );
  OAI211XLTS U953 ( .A0(n4637), .A1(n3545), .B0(n5630), .C0(n5629), .Y(n2603)
         );
  OAI211XLTS U954 ( .A0(n4652), .A1(n3547), .B0(n5632), .C0(n5631), .Y(n2604)
         );
  OAI211XLTS U955 ( .A0(n4655), .A1(n3545), .B0(n5634), .C0(n5633), .Y(n2605)
         );
  OAI211XLTS U956 ( .A0(n4664), .A1(n3545), .B0(n5636), .C0(n5635), .Y(n2606)
         );
  OAI211XLTS U957 ( .A0(n4677), .A1(n3544), .B0(n5638), .C0(n5637), .Y(n2607)
         );
  OAI211XLTS U958 ( .A0(n4682), .A1(n3544), .B0(n5640), .C0(n5639), .Y(n2608)
         );
  OAI211XLTS U959 ( .A0(n4695), .A1(n3544), .B0(n5642), .C0(n5641), .Y(n2609)
         );
  OAI211XLTS U960 ( .A0(n4700), .A1(n3544), .B0(n5644), .C0(n5643), .Y(n2610)
         );
  OAI211XLTS U961 ( .A0(n4763), .A1(n3552), .B0(n5507), .C0(n5506), .Y(n2562)
         );
  OAI211XLTS U962 ( .A0(n4731), .A1(n3552), .B0(n5501), .C0(n5500), .Y(n2559)
         );
  OAI211XLTS U963 ( .A0(n4742), .A1(n3552), .B0(n5503), .C0(n5502), .Y(n2560)
         );
  OAI211XLTS U964 ( .A0(n4749), .A1(n3552), .B0(n5505), .C0(n5504), .Y(n2561)
         );
  OAI211XLTS U965 ( .A0(n4717), .A1(n3412), .B0(n5448), .C0(n5447), .Y(n2529)
         );
  OAI211XLTS U966 ( .A0(n4424), .A1(n3420), .B0(n5710), .C0(n5709), .Y(n2643)
         );
  OAI211XLTS U967 ( .A0(n4559), .A1(n3417), .B0(n5740), .C0(n5739), .Y(n2658)
         );
  OAI211XLTS U968 ( .A0(n4564), .A1(n3416), .B0(n5742), .C0(n5741), .Y(n2659)
         );
  OAI211XLTS U969 ( .A0(n4602), .A1(n3415), .B0(n5750), .C0(n5749), .Y(n2663)
         );
  OAI211XLTS U970 ( .A0(n4694), .A1(n3413), .B0(n5770), .C0(n5769), .Y(n2673)
         );
  OAI211XLTS U971 ( .A0(n4432), .A1(n3420), .B0(n5712), .C0(n5711), .Y(n2644)
         );
  OAI211XLTS U972 ( .A0(n4443), .A1(n3420), .B0(n5714), .C0(n5713), .Y(n2645)
         );
  OAI211XLTS U973 ( .A0(n4454), .A1(n3420), .B0(n5716), .C0(n5715), .Y(n2646)
         );
  OAI211XLTS U974 ( .A0(n4457), .A1(n3419), .B0(n5718), .C0(n5717), .Y(n2647)
         );
  OAI211XLTS U975 ( .A0(n4466), .A1(n3419), .B0(n5720), .C0(n5719), .Y(n2648)
         );
  OAI211XLTS U976 ( .A0(n4481), .A1(n3419), .B0(n5722), .C0(n5721), .Y(n2649)
         );
  OAI211XLTS U977 ( .A0(n4488), .A1(n3419), .B0(n5724), .C0(n5723), .Y(n2650)
         );
  OAI211XLTS U978 ( .A0(n4495), .A1(n3418), .B0(n5726), .C0(n5725), .Y(n2651)
         );
  OAI211XLTS U979 ( .A0(n4506), .A1(n3418), .B0(n5728), .C0(n5727), .Y(n2652)
         );
  OAI211XLTS U980 ( .A0(n4513), .A1(n3418), .B0(n5730), .C0(n5729), .Y(n2653)
         );
  OAI211XLTS U981 ( .A0(n4520), .A1(n3418), .B0(n5732), .C0(n5731), .Y(n2654)
         );
  OAI211XLTS U982 ( .A0(n4533), .A1(n3417), .B0(n5734), .C0(n5733), .Y(n2655)
         );
  OAI211XLTS U983 ( .A0(n4540), .A1(n3417), .B0(n5736), .C0(n5735), .Y(n2656)
         );
  OAI211XLTS U984 ( .A0(n4551), .A1(n3417), .B0(n5738), .C0(n5737), .Y(n2657)
         );
  OAI211XLTS U985 ( .A0(n4574), .A1(n3416), .B0(n5744), .C0(n5743), .Y(n2660)
         );
  OAI211XLTS U986 ( .A0(n4587), .A1(n3416), .B0(n5746), .C0(n5745), .Y(n2661)
         );
  OAI211XLTS U987 ( .A0(n4596), .A1(n3415), .B0(n5748), .C0(n5747), .Y(n2662)
         );
  OAI211XLTS U988 ( .A0(n4610), .A1(n3415), .B0(n5752), .C0(n5751), .Y(n2664)
         );
  OAI211XLTS U989 ( .A0(n4621), .A1(n3415), .B0(n5754), .C0(n5753), .Y(n2665)
         );
  OAI211XLTS U990 ( .A0(n4632), .A1(n3414), .B0(n5756), .C0(n5755), .Y(n2666)
         );
  OAI211XLTS U991 ( .A0(n4641), .A1(n3414), .B0(n5758), .C0(n5757), .Y(n2667)
         );
  OAI211XLTS U992 ( .A0(n4648), .A1(n3416), .B0(n5760), .C0(n5759), .Y(n2668)
         );
  OAI211XLTS U993 ( .A0(n4661), .A1(n3414), .B0(n5762), .C0(n5761), .Y(n2669)
         );
  OAI211XLTS U994 ( .A0(n4668), .A1(n3414), .B0(n5764), .C0(n5763), .Y(n2670)
         );
  OAI211XLTS U995 ( .A0(n4679), .A1(n3413), .B0(n5766), .C0(n5765), .Y(n2671)
         );
  OAI211XLTS U996 ( .A0(n4684), .A1(n3413), .B0(n5768), .C0(n5767), .Y(n2672)
         );
  OAI211XLTS U997 ( .A0(n4706), .A1(n3413), .B0(n5772), .C0(n5771), .Y(n2674)
         );
  OAI211XLTS U998 ( .A0(n4721), .A1(n3553), .B0(n5499), .C0(n5498), .Y(n2558)
         );
  INVXLTS U999 ( .A(n3554), .Y(n3553) );
  OAI211XLTS U1000 ( .A0(n4735), .A1(n3421), .B0(n5452), .C0(n5451), .Y(n2531)
         );
  OAI211XLTS U1001 ( .A0(n4744), .A1(n3421), .B0(n5454), .C0(n5453), .Y(n2532)
         );
  OAI211XLTS U1002 ( .A0(n4753), .A1(n3421), .B0(n5456), .C0(n5455), .Y(n2533)
         );
  OAI211XLTS U1003 ( .A0(n4760), .A1(n3421), .B0(n5458), .C0(n5457), .Y(n2534)
         );
  OAI211XLTS U1004 ( .A0(n4726), .A1(n3422), .B0(n5450), .C0(n5449), .Y(n2530)
         );
  INVXLTS U1005 ( .A(n3423), .Y(n3422) );
  OAI211XLTS U1006 ( .A0(n3740), .A1(n4102), .B0(n5404), .C0(n5403), .Y(n2502)
         );
  OAI211XLTS U1007 ( .A0(n3740), .A1(n4099), .B0(n5406), .C0(n5405), .Y(n2503)
         );
  OAI211XLTS U1008 ( .A0(n3740), .A1(n4096), .B0(n5408), .C0(n5407), .Y(n2504)
         );
  OAI211XLTS U1009 ( .A0(n3740), .A1(n4105), .B0(n5402), .C0(n5401), .Y(n2501)
         );
  OAI211XLTS U1010 ( .A0(n3745), .A1(n3979), .B0(n5898), .C0(n5897), .Y(n2737)
         );
  OAI211XLTS U1011 ( .A0(n3745), .A1(n3976), .B0(n5900), .C0(n5899), .Y(n2738)
         );
  OAI211XLTS U1012 ( .A0(n3750), .A1(n4093), .B0(n5410), .C0(n5409), .Y(n2505)
         );
  OAI211XLTS U1013 ( .A0(n3748), .A1(n4090), .B0(n5412), .C0(n5411), .Y(n2506)
         );
  OAI211XLTS U1014 ( .A0(n3752), .A1(n4069), .B0(n5838), .C0(n5837), .Y(n2707)
         );
  OAI211XLTS U1015 ( .A0(n3747), .A1(n4066), .B0(n5840), .C0(n5839), .Y(n2708)
         );
  OAI211XLTS U1016 ( .A0(n3747), .A1(n4063), .B0(n5842), .C0(n5841), .Y(n2709)
         );
  OAI211XLTS U1017 ( .A0(n3753), .A1(n4060), .B0(n5844), .C0(n5843), .Y(n2710)
         );
  OAI211XLTS U1018 ( .A0(n3750), .A1(n4057), .B0(n5846), .C0(n5845), .Y(n2711)
         );
  OAI211XLTS U1019 ( .A0(n3749), .A1(n4054), .B0(n5848), .C0(n5847), .Y(n2712)
         );
  OAI211XLTS U1020 ( .A0(n3748), .A1(n4048), .B0(n5852), .C0(n5851), .Y(n2714)
         );
  OAI211XLTS U1021 ( .A0(n3750), .A1(n4042), .B0(n5856), .C0(n5855), .Y(n2716)
         );
  OAI211XLTS U1022 ( .A0(n3751), .A1(n4039), .B0(n5858), .C0(n5857), .Y(n2717)
         );
  OAI211XLTS U1023 ( .A0(n3751), .A1(n4033), .B0(n5862), .C0(n5861), .Y(n2719)
         );
  OAI211XLTS U1024 ( .A0(n3741), .A1(n4027), .B0(n5866), .C0(n5865), .Y(n2721)
         );
  OAI211XLTS U1025 ( .A0(n3741), .A1(n4024), .B0(n5868), .C0(n5867), .Y(n2722)
         );
  OAI211XLTS U1026 ( .A0(n3741), .A1(n4018), .B0(n5872), .C0(n5871), .Y(n2724)
         );
  OAI211XLTS U1027 ( .A0(n3742), .A1(n4012), .B0(n5876), .C0(n5875), .Y(n2726)
         );
  OAI211XLTS U1028 ( .A0(n3742), .A1(n4009), .B0(n5878), .C0(n5877), .Y(n2727)
         );
  OAI211XLTS U1029 ( .A0(n3742), .A1(n4006), .B0(n5880), .C0(n5879), .Y(n2728)
         );
  OAI211XLTS U1030 ( .A0(n3743), .A1(n4003), .B0(n5882), .C0(n5881), .Y(n2729)
         );
  OAI211XLTS U1031 ( .A0(n3743), .A1(n4000), .B0(n5884), .C0(n5883), .Y(n2730)
         );
  OAI211XLTS U1032 ( .A0(n3743), .A1(n3994), .B0(n5888), .C0(n5887), .Y(n2732)
         );
  OAI211XLTS U1033 ( .A0(n3744), .A1(n3985), .B0(n5894), .C0(n5893), .Y(n2735)
         );
  OAI211XLTS U1034 ( .A0(n3750), .A1(n4051), .B0(n5850), .C0(n5849), .Y(n2713)
         );
  OAI211XLTS U1035 ( .A0(n3749), .A1(n4045), .B0(n5854), .C0(n5853), .Y(n2715)
         );
  OAI211XLTS U1036 ( .A0(n3752), .A1(n4036), .B0(n5860), .C0(n5859), .Y(n2718)
         );
  OAI211XLTS U1037 ( .A0(n3751), .A1(n4030), .B0(n5864), .C0(n5863), .Y(n2720)
         );
  OAI211XLTS U1038 ( .A0(n3741), .A1(n4021), .B0(n5870), .C0(n5869), .Y(n2723)
         );
  OAI211XLTS U1039 ( .A0(n3742), .A1(n4015), .B0(n5874), .C0(n5873), .Y(n2725)
         );
  OAI211XLTS U1040 ( .A0(n3744), .A1(n3991), .B0(n5890), .C0(n5889), .Y(n2733)
         );
  OAI211XLTS U1041 ( .A0(n3744), .A1(n3988), .B0(n5892), .C0(n5891), .Y(n2734)
         );
  OAI211XLTS U1042 ( .A0(n3744), .A1(n3982), .B0(n5896), .C0(n5895), .Y(n2736)
         );
  OAI211XLTS U1043 ( .A0(n3743), .A1(n3997), .B0(n5886), .C0(n5885), .Y(n2731)
         );
  OAI2BB1XLTS U1044 ( .A0N(n4839), .A1N(n4867), .B0(n4838), .Y(n4850) );
  AOI32XLTS U1045 ( .A0(n131), .A1(n6231), .A2(n213), .B0(n132), .B1(n4837), 
        .Y(n4838) );
  XNOR2XLTS U1046 ( .A(n6230), .B(n213), .Y(n4837) );
  AOI32XLTS U1047 ( .A0(n106), .A1(n5561), .A2(n5560), .B0(n3556), .B1(n98), 
        .Y(n2570) );
  AOI22XLTS U1048 ( .A0(n3808), .A1(n5559), .B0(n3803), .B1(n5558), .Y(n5560)
         );
  AOI32XLTS U1049 ( .A0(n108), .A1(n5554), .A2(n5553), .B0(n692), .B1(n18), 
        .Y(n2569) );
  NAND2XLTS U1050 ( .A(n3802), .B(n5549), .Y(n5554) );
  NAND2XLTS U1051 ( .A(n200), .B(n235), .Y(n5436) );
  NAND3XLTS U1052 ( .A(n4866), .B(n6246), .C(n211), .Y(n5301) );
  NAND3XLTS U1053 ( .A(n234), .B(n4867), .C(n235), .Y(n5302) );
  NAND3XLTS U1054 ( .A(n4866), .B(n212), .C(n133), .Y(n5300) );
  NAND4XLTS U1055 ( .A(n132), .B(n234), .C(n6230), .D(n236), .Y(n5303) );
  NAND4XLTS U1056 ( .A(n131), .B(n234), .C(n236), .D(n6231), .Y(n5299) );
  CLKBUFX2TS U1057 ( .A(n5327), .Y(n481) );
  NOR3X1TS U1058 ( .A(n217), .B(n3), .C(n302), .Y(n5283) );
  OAI2BB2XLTS U1059 ( .B0(n6285), .B1(n3588), .A0N(
        \requesterAddressbuffer[2][5] ), .A1N(n206), .Y(n5126) );
  OAI2BB2XLTS U1060 ( .B0(n6286), .B1(n3588), .A0N(
        \requesterAddressbuffer[2][4] ), .A1N(n206), .Y(n5134) );
  OAI2BB2XLTS U1061 ( .B0(n6288), .B1(n3587), .A0N(
        \requesterAddressbuffer[2][2] ), .A1N(n205), .Y(n5150) );
  OAI2BB2XLTS U1062 ( .B0(n6289), .B1(n3587), .A0N(
        \requesterAddressbuffer[2][1] ), .A1N(n205), .Y(n5158) );
  OAI2BB2XLTS U1063 ( .B0(n6287), .B1(n3587), .A0N(
        \requesterAddressbuffer[2][3] ), .A1N(n206), .Y(n5142) );
  OAI2BB2XLTS U1064 ( .B0(n6290), .B1(n3587), .A0N(
        \requesterAddressbuffer[2][0] ), .A1N(n206), .Y(n5166) );
  NAND2X1TS U1065 ( .A(n5), .B(n301), .Y(n6221) );
  CLKBUFX2TS U1066 ( .A(n3749), .Y(n3741) );
  CLKBUFX2TS U1067 ( .A(n3749), .Y(n3742) );
  CLKBUFX2TS U1068 ( .A(n3748), .Y(n3744) );
  CLKBUFX2TS U1069 ( .A(n3748), .Y(n3743) );
  CLKBUFX2TS U1070 ( .A(n3747), .Y(n3745) );
  CLKBUFX2TS U1071 ( .A(n3747), .Y(n3746) );
  CLKBUFX2TS U1072 ( .A(n3752), .Y(n3750) );
  CLKBUFX2TS U1073 ( .A(n3753), .Y(n3747) );
  CLKBUFX2TS U1074 ( .A(n3753), .Y(n3749) );
  CLKBUFX2TS U1075 ( .A(n3753), .Y(n3748) );
  CLKBUFX2TS U1076 ( .A(n3708), .Y(n3697) );
  CLKBUFX2TS U1077 ( .A(n3707), .Y(n3698) );
  CLKBUFX2TS U1078 ( .A(n3705), .Y(n3699) );
  CLKBUFX2TS U1079 ( .A(n3705), .Y(n3700) );
  CLKBUFX2TS U1080 ( .A(n3706), .Y(n3701) );
  CLKBUFX2TS U1081 ( .A(n3706), .Y(n3702) );
  CLKBUFX2TS U1082 ( .A(n3705), .Y(n3703) );
  CLKBUFX2TS U1083 ( .A(n3705), .Y(n3704) );
  CLKBUFX2TS U1084 ( .A(n3719), .Y(n3717) );
  CLKBUFX2TS U1085 ( .A(n3721), .Y(n3713) );
  CLKBUFX2TS U1086 ( .A(n3721), .Y(n3712) );
  CLKBUFX2TS U1087 ( .A(n3722), .Y(n3711) );
  CLKBUFX2TS U1088 ( .A(n3720), .Y(n3715) );
  CLKBUFX2TS U1089 ( .A(n3719), .Y(n3716) );
  CLKBUFX2TS U1090 ( .A(n3720), .Y(n3714) );
  CLKBUFX2TS U1091 ( .A(n3722), .Y(n3710) );
  CLKBUFX2TS U1092 ( .A(n3794), .Y(n3786) );
  CLKBUFX2TS U1093 ( .A(n3795), .Y(n3785) );
  CLKBUFX2TS U1094 ( .A(n3792), .Y(n3791) );
  CLKBUFX2TS U1095 ( .A(n3792), .Y(n3790) );
  CLKBUFX2TS U1096 ( .A(n3793), .Y(n3789) );
  CLKBUFX2TS U1097 ( .A(n3793), .Y(n3788) );
  CLKBUFX2TS U1098 ( .A(n3794), .Y(n3787) );
  CLKBUFX2TS U1099 ( .A(n3795), .Y(n3784) );
  CLKBUFX2TS U1100 ( .A(n3778), .Y(n3775) );
  CLKBUFX2TS U1101 ( .A(n3780), .Y(n3771) );
  CLKBUFX2TS U1102 ( .A(n3780), .Y(n3772) );
  CLKBUFX2TS U1103 ( .A(n3779), .Y(n3773) );
  CLKBUFX2TS U1104 ( .A(n3779), .Y(n3774) );
  CLKBUFX2TS U1105 ( .A(n3751), .Y(n3740) );
  CLKBUFX2TS U1106 ( .A(n3752), .Y(n3751) );
  CLKBUFX2TS U1107 ( .A(n3777), .Y(n3776) );
  CLKBUFX2TS U1108 ( .A(n3798), .Y(n3792) );
  CLKBUFX2TS U1109 ( .A(n3798), .Y(n3793) );
  CLKBUFX2TS U1110 ( .A(n3798), .Y(n3794) );
  CLKBUFX2TS U1111 ( .A(n3797), .Y(n3795) );
  CLKBUFX2TS U1112 ( .A(n3797), .Y(n3796) );
  CLKBUFX2TS U1113 ( .A(n3723), .Y(n3721) );
  CLKBUFX2TS U1114 ( .A(n6342), .Y(n3707) );
  CLKBUFX2TS U1115 ( .A(n3709), .Y(n3706) );
  CLKBUFX2TS U1116 ( .A(n3709), .Y(n3705) );
  CLKBUFX2TS U1117 ( .A(n3724), .Y(n3718) );
  CLKBUFX2TS U1118 ( .A(n3724), .Y(n3719) );
  CLKBUFX2TS U1119 ( .A(n3723), .Y(n3720) );
  CLKBUFX2TS U1120 ( .A(n3723), .Y(n3722) );
  CLKBUFX2TS U1121 ( .A(n3783), .Y(n3778) );
  CLKBUFX2TS U1122 ( .A(n3782), .Y(n3780) );
  CLKBUFX2TS U1123 ( .A(n3782), .Y(n3779) );
  CLKBUFX2TS U1124 ( .A(n3783), .Y(n3777) );
  CLKBUFX2TS U1125 ( .A(n837), .Y(n835) );
  CLKBUFX2TS U1126 ( .A(n6346), .Y(n3752) );
  CLKBUFX2TS U1127 ( .A(n6346), .Y(n3753) );
  CLKBUFX2TS U1128 ( .A(n3375), .Y(n3361) );
  CLKBUFX2TS U1129 ( .A(n3375), .Y(n3362) );
  CLKBUFX2TS U1130 ( .A(n753), .Y(n749) );
  CLKBUFX2TS U1131 ( .A(n754), .Y(n748) );
  CLKBUFX2TS U1132 ( .A(n754), .Y(n747) );
  CLKBUFX2TS U1133 ( .A(n755), .Y(n746) );
  CLKBUFX2TS U1134 ( .A(n755), .Y(n745) );
  CLKBUFX2TS U1135 ( .A(n758), .Y(n743) );
  CLKBUFX2TS U1136 ( .A(n3370), .Y(n3368) );
  CLKBUFX2TS U1137 ( .A(n3373), .Y(n3366) );
  CLKBUFX2TS U1138 ( .A(n3373), .Y(n3365) );
  CLKBUFX2TS U1139 ( .A(n3372), .Y(n3367) );
  CLKBUFX2TS U1140 ( .A(n3374), .Y(n3364) );
  CLKBUFX2TS U1141 ( .A(n3374), .Y(n3363) );
  CLKBUFX2TS U1142 ( .A(n3485), .Y(n3481) );
  CLKBUFX2TS U1143 ( .A(n3486), .Y(n3480) );
  CLKBUFX2TS U1144 ( .A(n3486), .Y(n3479) );
  CLKBUFX2TS U1145 ( .A(n3487), .Y(n3478) );
  CLKBUFX2TS U1146 ( .A(n3487), .Y(n3477) );
  CLKBUFX2TS U1147 ( .A(n3488), .Y(n3476) );
  CLKBUFX2TS U1148 ( .A(n3488), .Y(n3475) );
  CLKBUFX2TS U1149 ( .A(n842), .Y(n829) );
  CLKBUFX2TS U1150 ( .A(n3736), .Y(n3726) );
  CLKBUFX2TS U1151 ( .A(n842), .Y(n830) );
  CLKBUFX2TS U1152 ( .A(n840), .Y(n833) );
  CLKBUFX2TS U1153 ( .A(n3736), .Y(n3733) );
  CLKBUFX2TS U1154 ( .A(n3734), .Y(n3732) );
  CLKBUFX2TS U1155 ( .A(n3734), .Y(n3731) );
  CLKBUFX2TS U1156 ( .A(n3734), .Y(n3730) );
  CLKBUFX2TS U1157 ( .A(n3735), .Y(n3729) );
  CLKBUFX2TS U1158 ( .A(n3735), .Y(n3728) );
  CLKBUFX2TS U1159 ( .A(n3736), .Y(n3727) );
  CLKBUFX2TS U1160 ( .A(n840), .Y(n834) );
  CLKBUFX2TS U1161 ( .A(n841), .Y(n832) );
  CLKBUFX2TS U1162 ( .A(n841), .Y(n831) );
  CLKBUFX2TS U1163 ( .A(n3708), .Y(n3696) );
  CLKBUFX2TS U1164 ( .A(n6342), .Y(n3708) );
  CLKBUFX2TS U1165 ( .A(n806), .Y(n793) );
  CLKBUFX2TS U1166 ( .A(n3340), .Y(n3326) );
  CLKBUFX2TS U1167 ( .A(n3407), .Y(n3392) );
  CLKBUFX2TS U1168 ( .A(n3340), .Y(n3327) );
  CLKBUFX2TS U1169 ( .A(n3407), .Y(n3393) );
  CLKBUFX2TS U1170 ( .A(n806), .Y(n794) );
  CLKBUFX2TS U1171 ( .A(n803), .Y(n801) );
  CLKBUFX2TS U1172 ( .A(n803), .Y(n800) );
  CLKBUFX2TS U1173 ( .A(n804), .Y(n798) );
  CLKBUFX2TS U1174 ( .A(n804), .Y(n797) );
  CLKBUFX2TS U1175 ( .A(n802), .Y(n799) );
  CLKBUFX2TS U1176 ( .A(n805), .Y(n796) );
  CLKBUFX2TS U1177 ( .A(n805), .Y(n795) );
  CLKBUFX2TS U1178 ( .A(n3342), .Y(n3334) );
  CLKBUFX2TS U1179 ( .A(n3337), .Y(n3333) );
  CLKBUFX2TS U1180 ( .A(n3337), .Y(n3332) );
  CLKBUFX2TS U1181 ( .A(n3339), .Y(n3329) );
  CLKBUFX2TS U1182 ( .A(n3407), .Y(n3402) );
  CLKBUFX2TS U1183 ( .A(n3370), .Y(n3369) );
  CLKBUFX2TS U1184 ( .A(n3404), .Y(n3401) );
  CLKBUFX2TS U1185 ( .A(n3404), .Y(n3400) );
  CLKBUFX2TS U1186 ( .A(n3405), .Y(n3399) );
  CLKBUFX2TS U1187 ( .A(n3406), .Y(n3397) );
  CLKBUFX2TS U1188 ( .A(n3406), .Y(n3396) );
  CLKBUFX2TS U1189 ( .A(n3405), .Y(n3398) );
  CLKBUFX2TS U1190 ( .A(n3406), .Y(n3395) );
  CLKBUFX2TS U1191 ( .A(n3406), .Y(n3394) );
  CLKBUFX2TS U1192 ( .A(n936), .Y(n860) );
  CLKBUFX2TS U1193 ( .A(n936), .Y(n861) );
  CLKBUFX2TS U1194 ( .A(n3258), .Y(n3244) );
  CLKBUFX2TS U1195 ( .A(n3258), .Y(n3245) );
  CLKBUFX2TS U1196 ( .A(n3338), .Y(n3331) );
  CLKBUFX2TS U1197 ( .A(n3338), .Y(n3330) );
  CLKBUFX2TS U1198 ( .A(n3339), .Y(n3328) );
  CLKBUFX2TS U1199 ( .A(n3485), .Y(n3482) );
  CLKBUFX2TS U1200 ( .A(n919), .Y(n862) );
  CLKBUFX2TS U1201 ( .A(n3257), .Y(n3246) );
  CLKBUFX2TS U1202 ( .A(n886), .Y(n865) );
  CLKBUFX2TS U1203 ( .A(n870), .Y(n869) );
  CLKBUFX2TS U1204 ( .A(n886), .Y(n864) );
  CLKBUFX2TS U1205 ( .A(n870), .Y(n868) );
  CLKBUFX2TS U1206 ( .A(n871), .Y(n866) );
  CLKBUFX2TS U1207 ( .A(n871), .Y(n867) );
  CLKBUFX2TS U1208 ( .A(n919), .Y(n863) );
  CLKBUFX2TS U1209 ( .A(n3309), .Y(n3295) );
  CLKBUFX2TS U1210 ( .A(n3309), .Y(n3296) );
  CLKBUFX2TS U1211 ( .A(n3253), .Y(n3252) );
  CLKBUFX2TS U1212 ( .A(n3254), .Y(n3251) );
  CLKBUFX2TS U1213 ( .A(n3254), .Y(n3250) );
  CLKBUFX2TS U1214 ( .A(n3256), .Y(n3249) );
  CLKBUFX2TS U1215 ( .A(n3257), .Y(n3247) );
  CLKBUFX2TS U1216 ( .A(n3256), .Y(n3248) );
  CLKBUFX2TS U1217 ( .A(n3764), .Y(n3755) );
  CLKBUFX2TS U1218 ( .A(n3761), .Y(n3760) );
  CLKBUFX2TS U1219 ( .A(n3305), .Y(n3304) );
  CLKBUFX2TS U1220 ( .A(n3306), .Y(n3301) );
  CLKBUFX2TS U1221 ( .A(n3307), .Y(n3300) );
  CLKBUFX2TS U1222 ( .A(n3761), .Y(n3759) );
  CLKBUFX2TS U1223 ( .A(n3767), .Y(n3758) );
  CLKBUFX2TS U1224 ( .A(n3763), .Y(n3757) );
  CLKBUFX2TS U1225 ( .A(n3764), .Y(n3756) );
  CLKBUFX2TS U1226 ( .A(n3305), .Y(n3303) );
  CLKBUFX2TS U1227 ( .A(n3306), .Y(n3302) );
  CLKBUFX2TS U1228 ( .A(n3307), .Y(n3299) );
  CLKBUFX2TS U1229 ( .A(n3781), .Y(n3770) );
  CLKBUFX2TS U1230 ( .A(n3782), .Y(n3781) );
  INVX2TS U1231 ( .A(n3239), .Y(n3236) );
  INVX2TS U1232 ( .A(n3240), .Y(n3235) );
  INVX2TS U1233 ( .A(n3238), .Y(n3237) );
  CLKBUFX2TS U1234 ( .A(n740), .Y(n716) );
  CLKBUFX2TS U1235 ( .A(n738), .Y(n729) );
  CLKBUFX2TS U1236 ( .A(n737), .Y(n732) );
  CLKBUFX2TS U1237 ( .A(n738), .Y(n717) );
  CLKBUFX2TS U1238 ( .A(n737), .Y(n733) );
  CLKBUFX2TS U1239 ( .A(n736), .Y(n734) );
  CLKBUFX2TS U1240 ( .A(n736), .Y(n735) );
  CLKBUFX2TS U1241 ( .A(n3243), .Y(n3238) );
  CLKBUFX2TS U1242 ( .A(n3243), .Y(n3239) );
  CLKBUFX2TS U1243 ( .A(n3243), .Y(n3240) );
  CLKBUFX2TS U1244 ( .A(n3195), .Y(n1822) );
  CLKBUFX2TS U1245 ( .A(n3195), .Y(n3192) );
  CLKBUFX2TS U1246 ( .A(n3195), .Y(n1894) );
  CLKBUFX2TS U1247 ( .A(n955), .Y(n886) );
  CLKBUFX2TS U1248 ( .A(n3310), .Y(n3308) );
  CLKBUFX2TS U1249 ( .A(n3767), .Y(n3761) );
  CLKBUFX2TS U1250 ( .A(n3767), .Y(n3762) );
  CLKBUFX2TS U1251 ( .A(n6135), .Y(n870) );
  CLKBUFX2TS U1252 ( .A(n3766), .Y(n3763) );
  CLKBUFX2TS U1253 ( .A(n955), .Y(n871) );
  CLKBUFX2TS U1254 ( .A(n3766), .Y(n3764) );
  CLKBUFX2TS U1255 ( .A(n955), .Y(n919) );
  CLKBUFX2TS U1256 ( .A(n3310), .Y(n3309) );
  CLKBUFX2TS U1257 ( .A(n3310), .Y(n3305) );
  CLKBUFX2TS U1258 ( .A(n6164), .Y(n3306) );
  CLKBUFX2TS U1259 ( .A(n3310), .Y(n3307) );
  CLKBUFX2TS U1260 ( .A(n808), .Y(n803) );
  CLKBUFX2TS U1261 ( .A(n759), .Y(n753) );
  CLKBUFX2TS U1262 ( .A(n759), .Y(n754) );
  CLKBUFX2TS U1263 ( .A(n807), .Y(n804) );
  CLKBUFX2TS U1264 ( .A(n758), .Y(n756) );
  CLKBUFX2TS U1265 ( .A(n759), .Y(n755) );
  CLKBUFX2TS U1266 ( .A(n807), .Y(n805) );
  CLKBUFX2TS U1267 ( .A(n3260), .Y(n3253) );
  CLKBUFX2TS U1268 ( .A(n3260), .Y(n3254) );
  CLKBUFX2TS U1269 ( .A(n3260), .Y(n3255) );
  CLKBUFX2TS U1270 ( .A(n3377), .Y(n3370) );
  CLKBUFX2TS U1271 ( .A(n6182), .Y(n3404) );
  CLKBUFX2TS U1272 ( .A(n3377), .Y(n3371) );
  CLKBUFX2TS U1273 ( .A(n6345), .Y(n3734) );
  CLKBUFX2TS U1274 ( .A(n3376), .Y(n3373) );
  CLKBUFX2TS U1275 ( .A(n6182), .Y(n3405) );
  CLKBUFX2TS U1276 ( .A(n3377), .Y(n3372) );
  CLKBUFX2TS U1277 ( .A(n3738), .Y(n3735) );
  CLKBUFX2TS U1278 ( .A(n3408), .Y(n3406) );
  CLKBUFX2TS U1279 ( .A(n3376), .Y(n3374) );
  CLKBUFX2TS U1280 ( .A(n3738), .Y(n3736) );
  CLKBUFX2TS U1281 ( .A(n3408), .Y(n3407) );
  CLKBUFX2TS U1282 ( .A(n3376), .Y(n3375) );
  CLKBUFX2TS U1283 ( .A(n3489), .Y(n3486) );
  CLKBUFX2TS U1284 ( .A(n3489), .Y(n3487) );
  CLKBUFX2TS U1285 ( .A(n3489), .Y(n3488) );
  CLKBUFX2TS U1286 ( .A(n807), .Y(n806) );
  CLKBUFX2TS U1287 ( .A(n758), .Y(n757) );
  CLKBUFX2TS U1288 ( .A(n955), .Y(n936) );
  CLKBUFX2TS U1289 ( .A(n3259), .Y(n3258) );
  CLKBUFX2TS U1290 ( .A(n3259), .Y(n3257) );
  CLKBUFX2TS U1291 ( .A(n3259), .Y(n3256) );
  CLKBUFX2TS U1292 ( .A(n3490), .Y(n3485) );
  CLKBUFX2TS U1293 ( .A(n3342), .Y(n3337) );
  CLKBUFX2TS U1294 ( .A(n3341), .Y(n3340) );
  CLKBUFX2TS U1295 ( .A(n844), .Y(n838) );
  CLKBUFX2TS U1296 ( .A(n844), .Y(n839) );
  CLKBUFX2TS U1297 ( .A(n3341), .Y(n3339) );
  CLKBUFX2TS U1298 ( .A(n843), .Y(n840) );
  CLKBUFX2TS U1299 ( .A(n843), .Y(n841) );
  CLKBUFX2TS U1300 ( .A(n843), .Y(n842) );
  CLKBUFX2TS U1301 ( .A(n3341), .Y(n3338) );
  CLKBUFX2TS U1302 ( .A(n343), .Y(n3739) );
  CLKBUFX2TS U1303 ( .A(n6349), .Y(n3782) );
  CLKBUFX2TS U1304 ( .A(n465), .Y(n3798) );
  CLKBUFX2TS U1305 ( .A(n465), .Y(n3797) );
  CLKBUFX2TS U1306 ( .A(n6343), .Y(n3723) );
  CLKBUFX2TS U1307 ( .A(n6342), .Y(n3709) );
  CLKBUFX2TS U1308 ( .A(n3291), .Y(n3278) );
  CLKBUFX2TS U1309 ( .A(n844), .Y(n837) );
  CLKBUFX2TS U1310 ( .A(n3291), .Y(n3279) );
  CLKBUFX2TS U1311 ( .A(n3288), .Y(n3284) );
  CLKBUFX2TS U1312 ( .A(n3290), .Y(n3281) );
  CLKBUFX2TS U1313 ( .A(n3469), .Y(n3464) );
  CLKBUFX2TS U1314 ( .A(n3471), .Y(n3463) );
  CLKBUFX2TS U1315 ( .A(n3472), .Y(n3461) );
  CLKBUFX2TS U1316 ( .A(n3472), .Y(n3460) );
  CLKBUFX2TS U1317 ( .A(n3473), .Y(n3458) );
  CLKBUFX2TS U1318 ( .A(n3289), .Y(n3283) );
  CLKBUFX2TS U1319 ( .A(n3289), .Y(n3282) );
  CLKBUFX2TS U1320 ( .A(n3290), .Y(n3280) );
  CLKBUFX2TS U1321 ( .A(n3471), .Y(n3462) );
  CLKBUFX2TS U1322 ( .A(n3473), .Y(n3459) );
  CLKBUFX2TS U1323 ( .A(n3210), .Y(n3196) );
  CLKBUFX2TS U1324 ( .A(n712), .Y(n696) );
  CLKBUFX2TS U1325 ( .A(n3737), .Y(n3725) );
  CLKBUFX2TS U1326 ( .A(n3738), .Y(n3737) );
  CLKBUFX2TS U1327 ( .A(n3210), .Y(n3197) );
  CLKBUFX2TS U1328 ( .A(n712), .Y(n697) );
  CLKBUFX2TS U1329 ( .A(n708), .Y(n701) );
  CLKBUFX2TS U1330 ( .A(n708), .Y(n700) );
  CLKBUFX2TS U1331 ( .A(n711), .Y(n699) );
  CLKBUFX2TS U1332 ( .A(n3208), .Y(n3204) );
  CLKBUFX2TS U1333 ( .A(n3207), .Y(n3203) );
  CLKBUFX2TS U1334 ( .A(n3207), .Y(n3202) );
  CLKBUFX2TS U1335 ( .A(n3208), .Y(n3201) );
  CLKBUFX2TS U1336 ( .A(n3208), .Y(n3200) );
  CLKBUFX2TS U1337 ( .A(n3209), .Y(n3198) );
  CLKBUFX2TS U1338 ( .A(n706), .Y(n704) );
  CLKBUFX2TS U1339 ( .A(n707), .Y(n703) );
  CLKBUFX2TS U1340 ( .A(n707), .Y(n702) );
  CLKBUFX2TS U1341 ( .A(n711), .Y(n698) );
  CLKBUFX2TS U1342 ( .A(n3209), .Y(n3199) );
  CLKBUFX2TS U1343 ( .A(n752), .Y(n751) );
  CLKBUFX2TS U1344 ( .A(n3484), .Y(n3483) );
  CLKBUFX2TS U1345 ( .A(n3532), .Y(n3529) );
  CLKBUFX2TS U1346 ( .A(n3533), .Y(n3528) );
  CLKBUFX2TS U1347 ( .A(n3533), .Y(n3527) );
  CLKBUFX2TS U1348 ( .A(n3534), .Y(n3526) );
  CLKBUFX2TS U1349 ( .A(n3537), .Y(n3524) );
  CLKBUFX2TS U1350 ( .A(n3537), .Y(n3523) );
  CLKBUFX2TS U1351 ( .A(n3534), .Y(n3525) );
  CLKBUFX2TS U1352 ( .A(n3469), .Y(n3466) );
  CLKBUFX2TS U1353 ( .A(n3506), .Y(n3492) );
  CLKBUFX2TS U1354 ( .A(n3506), .Y(n3493) );
  CLKBUFX2TS U1355 ( .A(n3442), .Y(n3427) );
  CLKBUFX2TS U1356 ( .A(n771), .Y(n769) );
  CLKBUFX2TS U1357 ( .A(n771), .Y(n768) );
  CLKBUFX2TS U1358 ( .A(n6118), .Y(n766) );
  CLKBUFX2TS U1359 ( .A(n773), .Y(n767) );
  CLKBUFX2TS U1360 ( .A(n773), .Y(n765) );
  CLKBUFX2TS U1361 ( .A(n3437), .Y(n3435) );
  CLKBUFX2TS U1362 ( .A(n3438), .Y(n3433) );
  CLKBUFX2TS U1363 ( .A(n3439), .Y(n3431) );
  CLKBUFX2TS U1364 ( .A(n3439), .Y(n3430) );
  CLKBUFX2TS U1365 ( .A(n3440), .Y(n3428) );
  CLKBUFX2TS U1366 ( .A(n3503), .Y(n3498) );
  CLKBUFX2TS U1367 ( .A(n3504), .Y(n3497) );
  CLKBUFX2TS U1368 ( .A(n3504), .Y(n3496) );
  CLKBUFX2TS U1369 ( .A(n773), .Y(n764) );
  CLKBUFX2TS U1370 ( .A(n3437), .Y(n3434) );
  CLKBUFX2TS U1371 ( .A(n3438), .Y(n3432) );
  CLKBUFX2TS U1372 ( .A(n3440), .Y(n3429) );
  CLKBUFX2TS U1373 ( .A(n3765), .Y(n3754) );
  CLKBUFX2TS U1374 ( .A(n3766), .Y(n3765) );
  INVX2TS U1375 ( .A(n3241), .Y(n3227) );
  INVX2TS U1376 ( .A(n3242), .Y(n3228) );
  INVX2TS U1377 ( .A(n3241), .Y(n3234) );
  CLKBUFX2TS U1378 ( .A(n3243), .Y(n3241) );
  INVX2TS U1379 ( .A(n3242), .Y(n3233) );
  CLKBUFX2TS U1380 ( .A(n472), .Y(n3242) );
  INVX2TS U1381 ( .A(n3242), .Y(n3232) );
  INVX2TS U1382 ( .A(n3242), .Y(n3231) );
  INVX2TS U1383 ( .A(n3241), .Y(n3229) );
  INVX2TS U1384 ( .A(n3241), .Y(n3230) );
  INVX2TS U1385 ( .A(n3194), .Y(n1537) );
  INVX2TS U1386 ( .A(n3193), .Y(n970) );
  CLKBUFX2TS U1387 ( .A(n3194), .Y(n3193) );
  INVX2TS U1388 ( .A(n3195), .Y(n1005) );
  INVX2TS U1389 ( .A(n3194), .Y(n1653) );
  INVX2TS U1390 ( .A(n3193), .Y(n986) );
  INVX2TS U1391 ( .A(n3193), .Y(n1402) );
  INVX2TS U1392 ( .A(n3193), .Y(n1586) );
  INVX2TS U1393 ( .A(n3194), .Y(n1654) );
  INVX2TS U1394 ( .A(n3272), .Y(n3262) );
  INVX2TS U1395 ( .A(n3272), .Y(n3261) );
  INVX2TS U1396 ( .A(n3273), .Y(n3263) );
  INVX2TS U1397 ( .A(n3273), .Y(n3264) );
  INVX2TS U1398 ( .A(n3274), .Y(n3265) );
  INVX2TS U1399 ( .A(n3275), .Y(n3266) );
  INVX2TS U1400 ( .A(n3275), .Y(n3267) );
  INVX2TS U1401 ( .A(n3276), .Y(n3269) );
  INVX2TS U1402 ( .A(n3276), .Y(n3268) );
  INVX2TS U1403 ( .A(n3274), .Y(n3271) );
  INVX2TS U1404 ( .A(n693), .Y(n688) );
  INVX2TS U1405 ( .A(n693), .Y(n687) );
  INVX2TS U1406 ( .A(n690), .Y(n683) );
  INVX2TS U1407 ( .A(n690), .Y(n682) );
  INVX2TS U1408 ( .A(n691), .Y(n685) );
  INVX2TS U1409 ( .A(n694), .Y(n686) );
  INVX2TS U1410 ( .A(n691), .Y(n684) );
  INVX2TS U1411 ( .A(n690), .Y(n681) );
  INVX2TS U1412 ( .A(n824), .Y(n820) );
  INVX2TS U1413 ( .A(n824), .Y(n819) );
  INVX2TS U1414 ( .A(n824), .Y(n818) );
  INVX2TS U1415 ( .A(n3425), .Y(n3419) );
  INVX2TS U1416 ( .A(n3426), .Y(n3418) );
  INVX2TS U1417 ( .A(n3424), .Y(n3417) );
  INVX2TS U1418 ( .A(n3555), .Y(n3550) );
  INVX2TS U1419 ( .A(n3556), .Y(n3549) );
  INVX2TS U1420 ( .A(n3557), .Y(n3548) );
  INVX2TS U1421 ( .A(n3357), .Y(n3353) );
  INVX2TS U1422 ( .A(n3357), .Y(n3352) );
  INVX2TS U1423 ( .A(n3357), .Y(n3351) );
  INVX2TS U1424 ( .A(n476), .Y(n812) );
  INVX2TS U1425 ( .A(n3424), .Y(n3411) );
  INVX2TS U1426 ( .A(n3555), .Y(n3542) );
  INVX2TS U1427 ( .A(n3360), .Y(n3345) );
  INVX2TS U1428 ( .A(n828), .Y(n813) );
  INVX2TS U1429 ( .A(n3424), .Y(n3412) );
  INVX2TS U1430 ( .A(n3555), .Y(n3543) );
  INVX2TS U1431 ( .A(n478), .Y(n3346) );
  INVX2TS U1432 ( .A(n826), .Y(n816) );
  INVX2TS U1433 ( .A(n826), .Y(n817) );
  INVX2TS U1434 ( .A(n826), .Y(n815) );
  INVX2TS U1435 ( .A(n3358), .Y(n3349) );
  INVX2TS U1436 ( .A(n3358), .Y(n3348) );
  INVX2TS U1437 ( .A(n3423), .Y(n3415) );
  INVX2TS U1438 ( .A(n3423), .Y(n3416) );
  INVX2TS U1439 ( .A(n3423), .Y(n3414) );
  INVX2TS U1440 ( .A(n3424), .Y(n3413) );
  INVX2TS U1441 ( .A(n3554), .Y(n3546) );
  INVX2TS U1442 ( .A(n3554), .Y(n3547) );
  INVX2TS U1443 ( .A(n3554), .Y(n3545) );
  INVX2TS U1444 ( .A(n3555), .Y(n3544) );
  INVX2TS U1445 ( .A(n476), .Y(n814) );
  INVX2TS U1446 ( .A(n3358), .Y(n3350) );
  INVX2TS U1447 ( .A(n478), .Y(n3347) );
  INVX2TS U1448 ( .A(n470), .Y(n3270) );
  INVX2TS U1449 ( .A(n691), .Y(n689) );
  INVX2TS U1450 ( .A(n827), .Y(n810) );
  INVX2TS U1451 ( .A(n3425), .Y(n3409) );
  INVX2TS U1452 ( .A(n3359), .Y(n3343) );
  INVX2TS U1453 ( .A(n3556), .Y(n3540) );
  INVX2TS U1454 ( .A(n827), .Y(n811) );
  INVX2TS U1455 ( .A(n3359), .Y(n3344) );
  INVX2TS U1456 ( .A(n3425), .Y(n3410) );
  INVX2TS U1457 ( .A(n3556), .Y(n3541) );
  CLKBUFX2TS U1458 ( .A(n741), .Y(n740) );
  CLKBUFX2TS U1459 ( .A(n741), .Y(n739) );
  CLKBUFX2TS U1460 ( .A(n742), .Y(n738) );
  CLKBUFX2TS U1461 ( .A(n742), .Y(n737) );
  CLKBUFX2TS U1462 ( .A(n742), .Y(n736) );
  CLKBUFX2TS U1463 ( .A(n3225), .Y(n3213) );
  CLKBUFX2TS U1464 ( .A(n3224), .Y(n3215) );
  CLKBUFX2TS U1465 ( .A(n857), .Y(n846) );
  CLKBUFX2TS U1466 ( .A(n3225), .Y(n3214) );
  CLKBUFX2TS U1467 ( .A(n855), .Y(n847) );
  CLKBUFX2TS U1468 ( .A(n854), .Y(n849) );
  CLKBUFX2TS U1469 ( .A(n854), .Y(n850) );
  CLKBUFX2TS U1470 ( .A(n3221), .Y(n3220) );
  CLKBUFX2TS U1471 ( .A(n3223), .Y(n3218) );
  CLKBUFX2TS U1472 ( .A(n3222), .Y(n3219) );
  CLKBUFX2TS U1473 ( .A(n3224), .Y(n3216) );
  CLKBUFX2TS U1474 ( .A(n855), .Y(n848) );
  CLKBUFX2TS U1475 ( .A(n853), .Y(n851) );
  CLKBUFX2TS U1476 ( .A(n853), .Y(n852) );
  CLKBUFX2TS U1477 ( .A(n3223), .Y(n3217) );
  CLKBUFX2TS U1478 ( .A(n3456), .Y(n3445) );
  CLKBUFX2TS U1479 ( .A(n790), .Y(n780) );
  CLKBUFX2TS U1480 ( .A(n789), .Y(n782) );
  CLKBUFX2TS U1481 ( .A(n790), .Y(n781) );
  CLKBUFX2TS U1482 ( .A(n788), .Y(n784) );
  CLKBUFX2TS U1483 ( .A(n788), .Y(n785) );
  CLKBUFX2TS U1484 ( .A(n787), .Y(n786) );
  CLKBUFX2TS U1485 ( .A(n3323), .Y(n3312) );
  CLKBUFX2TS U1486 ( .A(n3322), .Y(n3316) );
  CLKBUFX2TS U1487 ( .A(n3390), .Y(n3378) );
  CLKBUFX2TS U1488 ( .A(n3389), .Y(n3380) );
  CLKBUFX2TS U1489 ( .A(n6181), .Y(n3379) );
  CLKBUFX2TS U1490 ( .A(n3388), .Y(n3382) );
  CLKBUFX2TS U1491 ( .A(n3388), .Y(n3383) );
  CLKBUFX2TS U1492 ( .A(n3389), .Y(n3381) );
  CLKBUFX2TS U1493 ( .A(n3454), .Y(n3450) );
  CLKBUFX2TS U1494 ( .A(n3455), .Y(n3448) );
  CLKBUFX2TS U1495 ( .A(n3455), .Y(n3447) );
  CLKBUFX2TS U1496 ( .A(n3520), .Y(n3509) );
  CLKBUFX2TS U1497 ( .A(n3518), .Y(n3510) );
  CLKBUFX2TS U1498 ( .A(n3518), .Y(n3511) );
  CLKBUFX2TS U1499 ( .A(n3517), .Y(n3512) );
  CLKBUFX2TS U1500 ( .A(n3517), .Y(n3513) );
  CLKBUFX2TS U1501 ( .A(n3516), .Y(n3514) );
  CLKBUFX2TS U1502 ( .A(n3516), .Y(n3515) );
  CLKBUFX2TS U1503 ( .A(n789), .Y(n783) );
  CLKBUFX2TS U1504 ( .A(n3324), .Y(n3315) );
  CLKBUFX2TS U1505 ( .A(n6165), .Y(n3314) );
  CLKBUFX2TS U1506 ( .A(n3323), .Y(n3313) );
  CLKBUFX2TS U1507 ( .A(n3322), .Y(n3317) );
  CLKBUFX2TS U1508 ( .A(n3454), .Y(n3449) );
  CLKBUFX2TS U1509 ( .A(n3456), .Y(n3446) );
  CLKBUFX2TS U1510 ( .A(n3453), .Y(n3451) );
  CLKBUFX2TS U1511 ( .A(n3321), .Y(n3320) );
  CLKBUFX2TS U1512 ( .A(n3321), .Y(n3318) );
  CLKBUFX2TS U1513 ( .A(n3321), .Y(n3319) );
  CLKBUFX2TS U1514 ( .A(n3387), .Y(n3386) );
  CLKBUFX2TS U1515 ( .A(n3388), .Y(n3384) );
  CLKBUFX2TS U1516 ( .A(n3387), .Y(n3385) );
  CLKBUFX2TS U1517 ( .A(n3453), .Y(n3452) );
  CLKBUFX2TS U1518 ( .A(n3584), .Y(n3572) );
  CLKBUFX2TS U1519 ( .A(n3584), .Y(n3580) );
  CLKBUFX2TS U1520 ( .A(n3581), .Y(n3579) );
  CLKBUFX2TS U1521 ( .A(n3581), .Y(n3578) );
  CLKBUFX2TS U1522 ( .A(n3582), .Y(n3577) );
  CLKBUFX2TS U1523 ( .A(n3582), .Y(n3576) );
  CLKBUFX2TS U1524 ( .A(n3583), .Y(n3575) );
  CLKBUFX2TS U1525 ( .A(n3584), .Y(n3573) );
  CLKBUFX2TS U1526 ( .A(n3583), .Y(n3574) );
  CLKBUFX2TS U1527 ( .A(n3569), .Y(n3558) );
  CLKBUFX2TS U1528 ( .A(n3567), .Y(n3559) );
  CLKBUFX2TS U1529 ( .A(n3567), .Y(n3560) );
  CLKBUFX2TS U1530 ( .A(n3566), .Y(n3561) );
  CLKBUFX2TS U1531 ( .A(n3565), .Y(n3564) );
  CLKBUFX2TS U1532 ( .A(n3566), .Y(n3562) );
  CLKBUFX2TS U1533 ( .A(n3565), .Y(n3563) );
  CLKBUFX2TS U1534 ( .A(n3678), .Y(n3666) );
  CLKBUFX2TS U1535 ( .A(n3678), .Y(n3667) );
  CLKBUFX2TS U1536 ( .A(n3650), .Y(n3643) );
  CLKBUFX2TS U1537 ( .A(n3645), .Y(n3642) );
  CLKBUFX2TS U1538 ( .A(n3645), .Y(n3641) );
  CLKBUFX2TS U1539 ( .A(n3679), .Y(n3668) );
  CLKBUFX2TS U1540 ( .A(n3677), .Y(n3669) );
  CLKBUFX2TS U1541 ( .A(n3646), .Y(n3639) );
  CLKBUFX2TS U1542 ( .A(n3677), .Y(n3670) );
  CLKBUFX2TS U1543 ( .A(n3647), .Y(n3638) );
  CLKBUFX2TS U1544 ( .A(n3676), .Y(n3671) );
  CLKBUFX2TS U1545 ( .A(n3648), .Y(n3635) );
  CLKBUFX2TS U1546 ( .A(n3647), .Y(n3637) );
  CLKBUFX2TS U1547 ( .A(n3648), .Y(n3636) );
  CLKBUFX2TS U1548 ( .A(n3646), .Y(n3640) );
  CLKBUFX2TS U1549 ( .A(n3676), .Y(n3672) );
  CLKBUFX2TS U1550 ( .A(n3675), .Y(n3673) );
  CLKBUFX2TS U1551 ( .A(n3675), .Y(n3674) );
  CLKBUFX2TS U1552 ( .A(n3211), .Y(n3210) );
  CLKBUFX2TS U1553 ( .A(n3211), .Y(n3208) );
  CLKBUFX2TS U1554 ( .A(n3211), .Y(n3209) );
  CLKBUFX2TS U1555 ( .A(n3442), .Y(n3441) );
  CLKBUFX2TS U1556 ( .A(n6149), .Y(n3221) );
  CLKBUFX2TS U1557 ( .A(n776), .Y(n775) );
  CLKBUFX2TS U1558 ( .A(n776), .Y(n771) );
  CLKBUFX2TS U1559 ( .A(n6118), .Y(n772) );
  CLKBUFX2TS U1560 ( .A(n776), .Y(n774) );
  CLKBUFX2TS U1561 ( .A(n3293), .Y(n3287) );
  CLKBUFX2TS U1562 ( .A(n3293), .Y(n3288) );
  CLKBUFX2TS U1563 ( .A(n3292), .Y(n3291) );
  CLKBUFX2TS U1564 ( .A(n3443), .Y(n3439) );
  CLKBUFX2TS U1565 ( .A(n3474), .Y(n3472) );
  CLKBUFX2TS U1566 ( .A(n3507), .Y(n3506) );
  CLKBUFX2TS U1567 ( .A(n3539), .Y(n3533) );
  CLKBUFX2TS U1568 ( .A(n3508), .Y(n3501) );
  CLKBUFX2TS U1569 ( .A(n3508), .Y(n3502) );
  CLKBUFX2TS U1570 ( .A(n3538), .Y(n3535) );
  CLKBUFX2TS U1571 ( .A(n3538), .Y(n3536) );
  CLKBUFX2TS U1572 ( .A(n3507), .Y(n3504) );
  CLKBUFX2TS U1573 ( .A(n3538), .Y(n3537) );
  CLKBUFX2TS U1574 ( .A(n3508), .Y(n3503) );
  CLKBUFX2TS U1575 ( .A(n3539), .Y(n3534) );
  CLKBUFX2TS U1576 ( .A(n776), .Y(n773) );
  CLKBUFX2TS U1577 ( .A(n3292), .Y(n3289) );
  CLKBUFX2TS U1578 ( .A(n3292), .Y(n3290) );
  CLKBUFX2TS U1579 ( .A(n6197), .Y(n3469) );
  CLKBUFX2TS U1580 ( .A(n3443), .Y(n3437) );
  CLKBUFX2TS U1581 ( .A(n6197), .Y(n3470) );
  CLKBUFX2TS U1582 ( .A(n3443), .Y(n3438) );
  CLKBUFX2TS U1583 ( .A(n3474), .Y(n3471) );
  CLKBUFX2TS U1584 ( .A(n3442), .Y(n3440) );
  CLKBUFX2TS U1585 ( .A(n3474), .Y(n3473) );
  CLKBUFX2TS U1586 ( .A(n3539), .Y(n3532) );
  CLKBUFX2TS U1587 ( .A(n3507), .Y(n3505) );
  CLKBUFX2TS U1588 ( .A(n6164), .Y(n3311) );
  CLKBUFX2TS U1589 ( .A(n6135), .Y(n957) );
  CLKBUFX2TS U1590 ( .A(n715), .Y(n705) );
  CLKBUFX2TS U1591 ( .A(n714), .Y(n708) );
  CLKBUFX2TS U1592 ( .A(n3208), .Y(n3206) );
  CLKBUFX2TS U1593 ( .A(n809), .Y(n802) );
  CLKBUFX2TS U1594 ( .A(n6120), .Y(n809) );
  CLKBUFX2TS U1595 ( .A(n760), .Y(n752) );
  CLKBUFX2TS U1596 ( .A(n6117), .Y(n760) );
  CLKBUFX2TS U1597 ( .A(n3212), .Y(n3207) );
  CLKBUFX2TS U1598 ( .A(n3491), .Y(n3484) );
  CLKBUFX2TS U1599 ( .A(n6211), .Y(n3491) );
  CLKBUFX2TS U1600 ( .A(n715), .Y(n706) );
  CLKBUFX2TS U1601 ( .A(n715), .Y(n707) );
  CLKBUFX2TS U1602 ( .A(n714), .Y(n711) );
  CLKBUFX2TS U1603 ( .A(n714), .Y(n712) );
  CLKBUFX2TS U1604 ( .A(n6133), .Y(n845) );
  CLKBUFX2TS U1605 ( .A(n6133), .Y(n843) );
  CLKBUFX2TS U1606 ( .A(n6150), .Y(n3260) );
  CLKBUFX2TS U1607 ( .A(n6150), .Y(n3259) );
  CLKBUFX2TS U1608 ( .A(n6135), .Y(n955) );
  CLKBUFX2TS U1609 ( .A(n6164), .Y(n3310) );
  CLKBUFX2TS U1610 ( .A(n6347), .Y(n3769) );
  CLKBUFX2TS U1611 ( .A(n6179), .Y(n3377) );
  CLKBUFX2TS U1612 ( .A(n6182), .Y(n3408) );
  CLKBUFX2TS U1613 ( .A(n6179), .Y(n3376) );
  CLKBUFX2TS U1614 ( .A(n6211), .Y(n3489) );
  CLKBUFX2TS U1615 ( .A(n6120), .Y(n807) );
  CLKBUFX2TS U1616 ( .A(n6117), .Y(n758) );
  CLKBUFX2TS U1617 ( .A(n293), .Y(n3767) );
  CLKBUFX2TS U1618 ( .A(n293), .Y(n3766) );
  CLKBUFX2TS U1619 ( .A(n380), .Y(n3768) );
  CLKBUFX2TS U1620 ( .A(n6345), .Y(n3738) );
  INVX2TS U1621 ( .A(n5563), .Y(n6349) );
  CLKBUFX2TS U1622 ( .A(n6166), .Y(n3342) );
  CLKBUFX2TS U1623 ( .A(n6166), .Y(n3341) );
  INVX2TS U1624 ( .A(n5580), .Y(n6342) );
  INVX2TS U1625 ( .A(n290), .Y(n6344) );
  CLKBUFX2TS U1626 ( .A(n473), .Y(n3194) );
  CLKBUFX2TS U1627 ( .A(n472), .Y(n3243) );
  CLKBUFX2TS U1628 ( .A(n473), .Y(n3195) );
  CLKBUFX2TS U1629 ( .A(n693), .Y(n692) );
  CLKBUFX2TS U1630 ( .A(n3212), .Y(n3205) );
  CLKBUFX2TS U1631 ( .A(n3443), .Y(n3436) );
  CLKBUFX2TS U1632 ( .A(n3538), .Y(n3531) );
  CLKBUFX2TS U1633 ( .A(n3508), .Y(n3500) );
  CLKBUFX2TS U1634 ( .A(n3277), .Y(n3272) );
  CLKBUFX2TS U1635 ( .A(n3277), .Y(n3276) );
  CLKBUFX2TS U1636 ( .A(n3277), .Y(n3273) );
  CLKBUFX2TS U1637 ( .A(n3277), .Y(n3274) );
  CLKBUFX2TS U1638 ( .A(n470), .Y(n3275) );
  CLKBUFX2TS U1639 ( .A(n828), .Y(n827) );
  CLKBUFX2TS U1640 ( .A(n3426), .Y(n3425) );
  CLKBUFX2TS U1641 ( .A(n3360), .Y(n3359) );
  CLKBUFX2TS U1642 ( .A(n3557), .Y(n3556) );
  INVX2TS U1643 ( .A(n5459), .Y(n6330) );
  INVX2TS U1644 ( .A(n695), .Y(n678) );
  INVX2TS U1645 ( .A(n695), .Y(n679) );
  INVX2TS U1646 ( .A(n695), .Y(n680) );
  INVX2TS U1647 ( .A(n826), .Y(n822) );
  INVX2TS U1648 ( .A(n827), .Y(n821) );
  INVX2TS U1649 ( .A(n474), .Y(n3421) );
  INVX2TS U1650 ( .A(n474), .Y(n3420) );
  INVX2TS U1651 ( .A(n477), .Y(n3552) );
  INVX2TS U1652 ( .A(n477), .Y(n3551) );
  CLKBUFX2TS U1653 ( .A(n859), .Y(n854) );
  CLKBUFX2TS U1654 ( .A(n792), .Y(n790) );
  CLKBUFX2TS U1655 ( .A(n792), .Y(n788) );
  CLKBUFX2TS U1656 ( .A(n6119), .Y(n787) );
  CLKBUFX2TS U1657 ( .A(n858), .Y(n857) );
  CLKBUFX2TS U1658 ( .A(n3226), .Y(n3225) );
  CLKBUFX2TS U1659 ( .A(n3226), .Y(n3222) );
  CLKBUFX2TS U1660 ( .A(n3226), .Y(n3224) );
  CLKBUFX2TS U1661 ( .A(n3325), .Y(n3321) );
  CLKBUFX2TS U1662 ( .A(n6181), .Y(n3389) );
  CLKBUFX2TS U1663 ( .A(n3391), .Y(n3388) );
  CLKBUFX2TS U1664 ( .A(n3391), .Y(n3387) );
  CLKBUFX2TS U1665 ( .A(n6196), .Y(n3455) );
  CLKBUFX2TS U1666 ( .A(n3521), .Y(n3520) );
  CLKBUFX2TS U1667 ( .A(n3521), .Y(n3519) );
  CLKBUFX2TS U1668 ( .A(n3522), .Y(n3518) );
  CLKBUFX2TS U1669 ( .A(n3522), .Y(n3517) );
  CLKBUFX2TS U1670 ( .A(n3522), .Y(n3516) );
  CLKBUFX2TS U1671 ( .A(n792), .Y(n789) );
  CLKBUFX2TS U1672 ( .A(n858), .Y(n856) );
  CLKBUFX2TS U1673 ( .A(n859), .Y(n855) );
  CLKBUFX2TS U1674 ( .A(n859), .Y(n853) );
  CLKBUFX2TS U1675 ( .A(n3226), .Y(n3223) );
  CLKBUFX2TS U1676 ( .A(n6165), .Y(n3323) );
  CLKBUFX2TS U1677 ( .A(n3325), .Y(n3322) );
  CLKBUFX2TS U1678 ( .A(n6196), .Y(n3453) );
  CLKBUFX2TS U1679 ( .A(n6196), .Y(n3454) );
  CLKBUFX2TS U1680 ( .A(n6196), .Y(n3456) );
  CLKBUFX2TS U1681 ( .A(n6104), .Y(n741) );
  CLKBUFX2TS U1682 ( .A(n6104), .Y(n742) );
  CLKBUFX2TS U1683 ( .A(n3457), .Y(n3444) );
  CLKBUFX2TS U1684 ( .A(n3453), .Y(n3457) );
  INVX2TS U1685 ( .A(n676), .Y(n661) );
  INVX2TS U1686 ( .A(n677), .Y(n662) );
  INVX2TS U1687 ( .A(n675), .Y(n671) );
  INVX2TS U1688 ( .A(n675), .Y(n670) );
  INVX2TS U1689 ( .A(n672), .Y(n669) );
  INVX2TS U1690 ( .A(n672), .Y(n668) );
  INVX2TS U1691 ( .A(n672), .Y(n667) );
  INVX2TS U1692 ( .A(n676), .Y(n665) );
  INVX2TS U1693 ( .A(n676), .Y(n664) );
  INVX2TS U1694 ( .A(n676), .Y(n666) );
  INVX2TS U1695 ( .A(n672), .Y(n663) );
  CLKBUFX2TS U1696 ( .A(n791), .Y(n779) );
  CLKBUFX2TS U1697 ( .A(n792), .Y(n791) );
  CLKBUFX2TS U1698 ( .A(n6165), .Y(n3324) );
  CLKBUFX2TS U1699 ( .A(n6181), .Y(n3390) );
  CLKBUFX2TS U1700 ( .A(n578), .Y(n566) );
  CLKBUFX2TS U1701 ( .A(n576), .Y(n574) );
  CLKBUFX2TS U1702 ( .A(n575), .Y(n573) );
  CLKBUFX2TS U1703 ( .A(n575), .Y(n572) );
  CLKBUFX2TS U1704 ( .A(n576), .Y(n571) );
  CLKBUFX2TS U1705 ( .A(n576), .Y(n570) );
  CLKBUFX2TS U1706 ( .A(n578), .Y(n567) );
  CLKBUFX2TS U1707 ( .A(n577), .Y(n569) );
  CLKBUFX2TS U1708 ( .A(n577), .Y(n568) );
  INVX2TS U1709 ( .A(n514), .Y(n511) );
  INVX2TS U1710 ( .A(n516), .Y(n509) );
  INVX2TS U1711 ( .A(n517), .Y(n508) );
  CLKBUFX2TS U1712 ( .A(n3586), .Y(n3581) );
  CLKBUFX2TS U1713 ( .A(n3585), .Y(n3582) );
  CLKBUFX2TS U1714 ( .A(n3585), .Y(n3584) );
  CLKBUFX2TS U1715 ( .A(n3585), .Y(n3583) );
  CLKBUFX2TS U1716 ( .A(n3570), .Y(n3569) );
  CLKBUFX2TS U1717 ( .A(n3570), .Y(n3568) );
  CLKBUFX2TS U1718 ( .A(n3571), .Y(n3567) );
  CLKBUFX2TS U1719 ( .A(n3571), .Y(n3566) );
  CLKBUFX2TS U1720 ( .A(n3571), .Y(n3565) );
  CLKBUFX2TS U1721 ( .A(n494), .Y(n482) );
  CLKBUFX2TS U1722 ( .A(n5214), .Y(n483) );
  CLKBUFX2TS U1723 ( .A(n493), .Y(n484) );
  CLKBUFX2TS U1724 ( .A(n493), .Y(n485) );
  CLKBUFX2TS U1725 ( .A(n491), .Y(n486) );
  CLKBUFX2TS U1726 ( .A(n492), .Y(n487) );
  CLKBUFX2TS U1727 ( .A(n491), .Y(n490) );
  CLKBUFX2TS U1728 ( .A(n492), .Y(n488) );
  CLKBUFX2TS U1729 ( .A(n491), .Y(n489) );
  CLKBUFX2TS U1730 ( .A(n561), .Y(n537) );
  CLKBUFX2TS U1731 ( .A(n561), .Y(n541) );
  CLKBUFX2TS U1732 ( .A(n556), .Y(n543) );
  CLKBUFX2TS U1733 ( .A(n556), .Y(n544) );
  CLKBUFX2TS U1734 ( .A(n555), .Y(n545) );
  CLKBUFX2TS U1735 ( .A(n554), .Y(n551) );
  CLKBUFX2TS U1736 ( .A(n555), .Y(n546) );
  CLKBUFX2TS U1737 ( .A(n554), .Y(n548) );
  INVX2TS U1738 ( .A(reset), .Y(n4418) );
  CLKBUFX2TS U1739 ( .A(n3661), .Y(n3656) );
  CLKBUFX2TS U1740 ( .A(n3662), .Y(n3655) );
  CLKBUFX2TS U1741 ( .A(n3694), .Y(n3681) );
  CLKBUFX2TS U1742 ( .A(n3662), .Y(n3654) );
  CLKBUFX2TS U1743 ( .A(n3693), .Y(n3682) );
  CLKBUFX2TS U1744 ( .A(n3615), .Y(n3604) );
  CLKBUFX2TS U1745 ( .A(n3661), .Y(n3653) );
  CLKBUFX2TS U1746 ( .A(n3693), .Y(n3683) );
  CLKBUFX2TS U1747 ( .A(n3615), .Y(n3605) );
  CLKBUFX2TS U1748 ( .A(n3663), .Y(n3652) );
  CLKBUFX2TS U1749 ( .A(n3692), .Y(n3684) );
  CLKBUFX2TS U1750 ( .A(n3614), .Y(n3606) );
  CLKBUFX2TS U1751 ( .A(n3663), .Y(n3651) );
  CLKBUFX2TS U1752 ( .A(n3692), .Y(n3685) );
  CLKBUFX2TS U1753 ( .A(n3614), .Y(n3607) );
  CLKBUFX2TS U1754 ( .A(n3691), .Y(n3686) );
  CLKBUFX2TS U1755 ( .A(n3613), .Y(n3608) );
  CLKBUFX2TS U1756 ( .A(n3601), .Y(n3587) );
  CLKBUFX2TS U1757 ( .A(n3601), .Y(n3588) );
  CLKBUFX2TS U1758 ( .A(n3629), .Y(n3625) );
  CLKBUFX2TS U1759 ( .A(n3603), .Y(n3595) );
  CLKBUFX2TS U1760 ( .A(n3629), .Y(n3624) );
  CLKBUFX2TS U1761 ( .A(n3630), .Y(n3623) );
  CLKBUFX2TS U1762 ( .A(n3598), .Y(n3594) );
  CLKBUFX2TS U1763 ( .A(n3630), .Y(n3622) );
  CLKBUFX2TS U1764 ( .A(n3598), .Y(n3593) );
  CLKBUFX2TS U1765 ( .A(n3631), .Y(n3621) );
  CLKBUFX2TS U1766 ( .A(n3599), .Y(n3592) );
  CLKBUFX2TS U1767 ( .A(n3631), .Y(n3620) );
  CLKBUFX2TS U1768 ( .A(n3599), .Y(n3591) );
  CLKBUFX2TS U1769 ( .A(n3600), .Y(n3590) );
  CLKBUFX2TS U1770 ( .A(n3600), .Y(n3589) );
  CLKBUFX2TS U1771 ( .A(n3661), .Y(n3657) );
  CLKBUFX2TS U1772 ( .A(n3613), .Y(n3609) );
  CLKBUFX2TS U1773 ( .A(n3691), .Y(n3687) );
  CLKBUFX2TS U1774 ( .A(n3612), .Y(n3611) );
  CLKBUFX2TS U1775 ( .A(n3679), .Y(n3678) );
  CLKBUFX2TS U1776 ( .A(n3650), .Y(n3645) );
  CLKBUFX2TS U1777 ( .A(n3680), .Y(n3677) );
  CLKBUFX2TS U1778 ( .A(n3680), .Y(n3676) );
  CLKBUFX2TS U1779 ( .A(n3649), .Y(n3647) );
  CLKBUFX2TS U1780 ( .A(n3649), .Y(n3648) );
  CLKBUFX2TS U1781 ( .A(n3649), .Y(n3646) );
  CLKBUFX2TS U1782 ( .A(n3680), .Y(n3675) );
  CLKBUFX2TS U1783 ( .A(n6319), .Y(n3644) );
  CLKBUFX2TS U1784 ( .A(n3612), .Y(n3610) );
  CLKBUFX2TS U1785 ( .A(n3660), .Y(n3658) );
  CLKBUFX2TS U1786 ( .A(n3690), .Y(n3688) );
  CLKBUFX2TS U1787 ( .A(n3660), .Y(n3659) );
  CLKBUFX2TS U1788 ( .A(n3690), .Y(n3689) );
  NAND2X1TS U1789 ( .A(n5508), .B(n5319), .Y(n5566) );
  AND2X2TS U1790 ( .A(n5558), .B(n5562), .Y(n6211) );
  AND2X2TS U1791 ( .A(n5520), .B(n6339), .Y(n6120) );
  CLKBUFX2TS U1792 ( .A(n6148), .Y(n3211) );
  CLKBUFX2TS U1793 ( .A(n475), .Y(n693) );
  CLKBUFX2TS U1794 ( .A(n475), .Y(n694) );
  CLKBUFX2TS U1795 ( .A(n6148), .Y(n3212) );
  CLKBUFX2TS U1796 ( .A(n6163), .Y(n3294) );
  CLKBUFX2TS U1797 ( .A(n777), .Y(n770) );
  CLKBUFX2TS U1798 ( .A(n6118), .Y(n777) );
  CLKBUFX2TS U1799 ( .A(n6163), .Y(n3292) );
  CLKBUFX2TS U1800 ( .A(n6118), .Y(n776) );
  CLKBUFX2TS U1801 ( .A(n6195), .Y(n3442) );
  CLKBUFX2TS U1802 ( .A(n6214), .Y(n3538) );
  CLKBUFX2TS U1803 ( .A(n6212), .Y(n3508) );
  CLKBUFX2TS U1804 ( .A(n6195), .Y(n3443) );
  CLKBUFX2TS U1805 ( .A(n6197), .Y(n3474) );
  CLKBUFX2TS U1806 ( .A(n6214), .Y(n3539) );
  CLKBUFX2TS U1807 ( .A(n6212), .Y(n3507) );
  INVX2TS U1808 ( .A(n5509), .Y(n6341) );
  CLKBUFX2TS U1809 ( .A(n6103), .Y(n714) );
  INVX2TS U1810 ( .A(n5576), .Y(n6345) );
  INVX2TS U1811 ( .A(n5530), .Y(n6338) );
  INVX2TS U1812 ( .A(n5531), .Y(n6337) );
  CLKBUFX2TS U1813 ( .A(n474), .Y(n3426) );
  CLKBUFX2TS U1814 ( .A(n476), .Y(n828) );
  CLKBUFX2TS U1815 ( .A(n477), .Y(n3557) );
  CLKBUFX2TS U1816 ( .A(n478), .Y(n3360) );
  INVX2TS U1817 ( .A(n5414), .Y(n6340) );
  CLKBUFX2TS U1818 ( .A(n470), .Y(n3277) );
  INVX2TS U1819 ( .A(n5517), .Y(n6339) );
  CLKBUFX2TS U1820 ( .A(n536), .Y(n514) );
  CLKBUFX2TS U1821 ( .A(n536), .Y(n516) );
  CLKBUFX2TS U1822 ( .A(n536), .Y(n517) );
  AND2X2TS U1823 ( .A(n5469), .B(n5353), .Y(n6104) );
  CLKBUFX2TS U1824 ( .A(n578), .Y(n575) );
  CLKBUFX2TS U1825 ( .A(n5278), .Y(n576) );
  CLKBUFX2TS U1826 ( .A(n580), .Y(n578) );
  CLKBUFX2TS U1827 ( .A(n580), .Y(n577) );
  CLKBUFX2TS U1828 ( .A(n6181), .Y(n3391) );
  CLKBUFX2TS U1829 ( .A(n6213), .Y(n3521) );
  CLKBUFX2TS U1830 ( .A(n6213), .Y(n3522) );
  CLKBUFX2TS U1831 ( .A(n6119), .Y(n792) );
  CLKBUFX2TS U1832 ( .A(n6134), .Y(n858) );
  CLKBUFX2TS U1833 ( .A(n6134), .Y(n859) );
  CLKBUFX2TS U1834 ( .A(n6149), .Y(n3226) );
  CLKBUFX2TS U1835 ( .A(n6165), .Y(n3325) );
  CLKBUFX2TS U1836 ( .A(n675), .Y(n673) );
  CLKBUFX2TS U1837 ( .A(n675), .Y(n674) );
  CLKBUFX2TS U1838 ( .A(n579), .Y(n565) );
  CLKBUFX2TS U1839 ( .A(n580), .Y(n579) );
  INVX2TS U1840 ( .A(n534), .Y(n496) );
  CLKBUFX2TS U1841 ( .A(n536), .Y(n534) );
  INVX2TS U1842 ( .A(n479), .Y(n500) );
  INVX2TS U1843 ( .A(n534), .Y(n501) );
  INVX2TS U1844 ( .A(n479), .Y(n502) );
  INVX2TS U1845 ( .A(n479), .Y(n503) );
  INVX2TS U1846 ( .A(n534), .Y(n504) );
  INVX2TS U1847 ( .A(n534), .Y(n505) );
  INVX2TS U1848 ( .A(n517), .Y(n507) );
  CLKBUFX2TS U1849 ( .A(n563), .Y(n561) );
  CLKBUFX2TS U1850 ( .A(n563), .Y(n557) );
  CLKBUFX2TS U1851 ( .A(n5214), .Y(n493) );
  CLKBUFX2TS U1852 ( .A(n564), .Y(n556) );
  CLKBUFX2TS U1853 ( .A(n564), .Y(n555) );
  CLKBUFX2TS U1854 ( .A(n495), .Y(n492) );
  CLKBUFX2TS U1855 ( .A(n564), .Y(n554) );
  CLKBUFX2TS U1856 ( .A(n495), .Y(n491) );
  CLKBUFX2TS U1857 ( .A(n6249), .Y(n3586) );
  CLKBUFX2TS U1858 ( .A(n6249), .Y(n3585) );
  CLKBUFX2TS U1859 ( .A(n5279), .Y(n3570) );
  CLKBUFX2TS U1860 ( .A(n5279), .Y(n3571) );
  CLKBUFX2TS U1861 ( .A(n5214), .Y(n494) );
  CLKBUFX2TS U1862 ( .A(n563), .Y(n562) );
  CLKBUFX2TS U1863 ( .A(n4262), .Y(n4263) );
  CLKBUFX2TS U1864 ( .A(n4265), .Y(n4266) );
  CLKBUFX2TS U1865 ( .A(n4262), .Y(n4264) );
  CLKBUFX2TS U1866 ( .A(n4265), .Y(n4267) );
  INVX2TS U1867 ( .A(n3810), .Y(n3808) );
  CLKBUFX2TS U1868 ( .A(n3665), .Y(n3661) );
  CLKBUFX2TS U1869 ( .A(n3617), .Y(n3616) );
  CLKBUFX2TS U1870 ( .A(n3633), .Y(n3629) );
  CLKBUFX2TS U1871 ( .A(n3665), .Y(n3662) );
  CLKBUFX2TS U1872 ( .A(n3633), .Y(n3630) );
  CLKBUFX2TS U1873 ( .A(n6317), .Y(n3598) );
  CLKBUFX2TS U1874 ( .A(n3694), .Y(n3693) );
  CLKBUFX2TS U1875 ( .A(n3617), .Y(n3615) );
  CLKBUFX2TS U1876 ( .A(n3633), .Y(n3631) );
  CLKBUFX2TS U1877 ( .A(n3602), .Y(n3599) );
  CLKBUFX2TS U1878 ( .A(n1), .Y(n3663) );
  CLKBUFX2TS U1879 ( .A(n3695), .Y(n3692) );
  CLKBUFX2TS U1880 ( .A(n3618), .Y(n3614) );
  CLKBUFX2TS U1881 ( .A(n3695), .Y(n3691) );
  CLKBUFX2TS U1882 ( .A(n3618), .Y(n3613) );
  CLKBUFX2TS U1883 ( .A(n3602), .Y(n3600) );
  CLKBUFX2TS U1884 ( .A(n1), .Y(n3664) );
  CLKBUFX2TS U1885 ( .A(n3602), .Y(n3601) );
  CLKBUFX2TS U1886 ( .A(n3618), .Y(n3612) );
  CLKBUFX2TS U1887 ( .A(n614), .Y(n608) );
  CLKBUFX2TS U1888 ( .A(n614), .Y(n607) );
  CLKBUFX2TS U1889 ( .A(n622), .Y(n594) );
  CLKBUFX2TS U1890 ( .A(n622), .Y(n584) );
  CLKBUFX2TS U1891 ( .A(n623), .Y(n582) );
  CLKBUFX2TS U1892 ( .A(n623), .Y(n581) );
  CLKBUFX2TS U1893 ( .A(n3632), .Y(n3619) );
  CLKBUFX2TS U1894 ( .A(n6318), .Y(n3632) );
  INVX2TS U1895 ( .A(n5353), .Y(n6321) );
  CLKBUFX2TS U1896 ( .A(n3665), .Y(n3660) );
  CLKBUFX2TS U1897 ( .A(n3695), .Y(n3690) );
  CLKBUFX2TS U1898 ( .A(n6320), .Y(n3679) );
  CLKBUFX2TS U1899 ( .A(n6320), .Y(n3680) );
  CLKBUFX2TS U1900 ( .A(n6319), .Y(n3650) );
  CLKBUFX2TS U1901 ( .A(n6319), .Y(n3649) );
  CLKBUFX2TS U1902 ( .A(n3628), .Y(n3626) );
  CLKBUFX2TS U1903 ( .A(n3628), .Y(n3627) );
  CLKBUFX2TS U1904 ( .A(n3597), .Y(n3596) );
  OAI21X1TS U1905 ( .A0(n6328), .A1(n166), .B0(n238), .Y(n5366) );
  NOR2X1TS U1906 ( .A(n5558), .B(n5559), .Y(n5556) );
  NOR2X1TS U1907 ( .A(n4853), .B(n6324), .Y(n4858) );
  OAI2BB1X1TS U1908 ( .A0N(n5317), .A1N(n5316), .B0(n5315), .Y(n5318) );
  OAI21X1TS U1909 ( .A0(n5316), .A1(n5317), .B0(n393), .Y(n5315) );
  NOR2X1TS U1910 ( .A(n5392), .B(n126), .Y(n6149) );
  INVX2TS U1911 ( .A(n4852), .Y(n6324) );
  OA22X1TS U1912 ( .A0(n5516), .A1(n126), .B0(n5484), .B1(n6321), .Y(n476) );
  OR2X2TS U1913 ( .A(n4858), .B(n4857), .Y(n4859) );
  INVX2TS U1914 ( .A(n5557), .Y(n6326) );
  INVX2TS U1915 ( .A(n5511), .Y(n6329) );
  AOI21X1TS U1916 ( .A0(n168), .A1(n6327), .B0(n6338), .Y(n5391) );
  XNOR2X1TS U1917 ( .A(n6316), .B(n6229), .Y(n4856) );
  NAND2X1TS U1918 ( .A(n168), .B(n5485), .Y(n5392) );
  NOR2BX1TS U1919 ( .AN(n201), .B(n14), .Y(n5469) );
  AND2X2TS U1920 ( .A(n5469), .B(n168), .Y(n6134) );
  AND2X2TS U1921 ( .A(n5495), .B(n225), .Y(n6213) );
  AND2X2TS U1922 ( .A(n5495), .B(n223), .Y(n6119) );
  AND2X2TS U1923 ( .A(n5469), .B(n5494), .Y(n6196) );
  AND2X2TS U1924 ( .A(n5495), .B(n170), .Y(n6181) );
  AND2X2TS U1925 ( .A(n5469), .B(n5446), .Y(n6165) );
  CLKBUFX2TS U1926 ( .A(n677), .Y(n676) );
  CLKBUFX2TS U1927 ( .A(n677), .Y(n675) );
  CLKBUFX2TS U1928 ( .A(n5278), .Y(n580) );
  CLKBUFX2TS U1929 ( .A(n479), .Y(n536) );
  NAND2X1TS U1930 ( .A(n126), .B(n4418), .Y(n6227) );
  CLKBUFX2TS U1931 ( .A(n3811), .Y(n3810) );
  CLKBUFX2TS U1932 ( .A(destinationAddressIn_SOUTH[6]), .Y(n4262) );
  CLKBUFX2TS U1933 ( .A(destinationAddressIn_SOUTH[7]), .Y(n4265) );
  CLKBUFX2TS U1934 ( .A(n5277), .Y(n563) );
  CLKBUFX2TS U1935 ( .A(n5277), .Y(n564) );
  CLKBUFX2TS U1936 ( .A(n5214), .Y(n495) );
  CLKBUFX2TS U1937 ( .A(n4289), .Y(n4290) );
  CLKBUFX2TS U1938 ( .A(n4400), .Y(n4401) );
  CLKBUFX2TS U1939 ( .A(n4373), .Y(n4374) );
  CLKBUFX2TS U1940 ( .A(n4355), .Y(n4356) );
  CLKBUFX2TS U1941 ( .A(n4349), .Y(n4350) );
  CLKBUFX2TS U1942 ( .A(n4346), .Y(n4347) );
  CLKBUFX2TS U1943 ( .A(n4325), .Y(n4326) );
  CLKBUFX2TS U1944 ( .A(n4322), .Y(n4323) );
  CLKBUFX2TS U1945 ( .A(n4316), .Y(n4317) );
  CLKBUFX2TS U1946 ( .A(n4304), .Y(n4305) );
  CLKBUFX2TS U1947 ( .A(n4379), .Y(n4380) );
  CLKBUFX2TS U1948 ( .A(n4376), .Y(n4377) );
  CLKBUFX2TS U1949 ( .A(n4370), .Y(n4371) );
  CLKBUFX2TS U1950 ( .A(n4367), .Y(n4368) );
  CLKBUFX2TS U1951 ( .A(n4364), .Y(n4365) );
  CLKBUFX2TS U1952 ( .A(n4358), .Y(n4359) );
  CLKBUFX2TS U1953 ( .A(n4352), .Y(n4353) );
  CLKBUFX2TS U1954 ( .A(n4343), .Y(n4344) );
  CLKBUFX2TS U1955 ( .A(n4334), .Y(n4335) );
  CLKBUFX2TS U1956 ( .A(n4319), .Y(n4320) );
  CLKBUFX2TS U1957 ( .A(n4313), .Y(n4314) );
  CLKBUFX2TS U1958 ( .A(n4310), .Y(n4311) );
  CLKBUFX2TS U1959 ( .A(n4307), .Y(n4308) );
  CLKBUFX2TS U1960 ( .A(n4301), .Y(n4302) );
  CLKBUFX2TS U1961 ( .A(n4292), .Y(n4293) );
  CLKBUFX2TS U1962 ( .A(n4415), .Y(n4416) );
  CLKBUFX2TS U1963 ( .A(n4409), .Y(n4410) );
  CLKBUFX2TS U1964 ( .A(n4406), .Y(n4407) );
  CLKBUFX2TS U1965 ( .A(n4403), .Y(n4404) );
  CLKBUFX2TS U1966 ( .A(n4286), .Y(n4287) );
  CLKBUFX2TS U1967 ( .A(n4337), .Y(n4338) );
  CLKBUFX2TS U1968 ( .A(n4331), .Y(n4332) );
  CLKBUFX2TS U1969 ( .A(n4328), .Y(n4329) );
  CLKBUFX2TS U1970 ( .A(n4295), .Y(n4296) );
  CLKBUFX2TS U1971 ( .A(n4412), .Y(n4413) );
  CLKBUFX2TS U1972 ( .A(n4361), .Y(n4362) );
  CLKBUFX2TS U1973 ( .A(n4340), .Y(n4341) );
  CLKBUFX2TS U1974 ( .A(n4298), .Y(n4299) );
  CLKBUFX2TS U1975 ( .A(n4397), .Y(n4398) );
  CLKBUFX2TS U1976 ( .A(n4394), .Y(n4395) );
  CLKBUFX2TS U1977 ( .A(n4388), .Y(n4389) );
  CLKBUFX2TS U1978 ( .A(n4391), .Y(n4392) );
  CLKBUFX2TS U1979 ( .A(n4385), .Y(n4386) );
  CLKBUFX2TS U1980 ( .A(n4382), .Y(n4383) );
  INVX2TS U1981 ( .A(n3913), .Y(n3911) );
  INVX2TS U1982 ( .A(n3910), .Y(n3908) );
  INVX2TS U1983 ( .A(n3907), .Y(n3905) );
  INVX2TS U1984 ( .A(n3904), .Y(n3902) );
  INVX2TS U1985 ( .A(n3901), .Y(n3899) );
  INVX2TS U1986 ( .A(n3898), .Y(n3896) );
  INVX2TS U1987 ( .A(n3895), .Y(n3893) );
  INVX2TS U1988 ( .A(n3892), .Y(n3890) );
  INVX2TS U1989 ( .A(n3889), .Y(n3887) );
  INVX2TS U1990 ( .A(n3886), .Y(n3884) );
  INVX2TS U1991 ( .A(n3883), .Y(n3881) );
  INVX2TS U1992 ( .A(n3880), .Y(n3878) );
  INVX2TS U1993 ( .A(n3877), .Y(n3875) );
  INVX2TS U1994 ( .A(n3874), .Y(n3872) );
  INVX2TS U1995 ( .A(n3871), .Y(n3869) );
  INVX2TS U1996 ( .A(n3868), .Y(n3866) );
  INVX2TS U1997 ( .A(n3865), .Y(n3863) );
  INVX2TS U1998 ( .A(n3862), .Y(n3860) );
  INVX2TS U1999 ( .A(n3859), .Y(n3857) );
  INVX2TS U2000 ( .A(n3856), .Y(n3854) );
  INVX2TS U2001 ( .A(n3853), .Y(n3851) );
  INVX2TS U2002 ( .A(n3850), .Y(n3848) );
  INVX2TS U2003 ( .A(n3847), .Y(n3845) );
  INVX2TS U2004 ( .A(n3844), .Y(n3842) );
  INVX2TS U2005 ( .A(n3841), .Y(n3839) );
  INVX2TS U2006 ( .A(n3838), .Y(n3836) );
  INVX2TS U2007 ( .A(n3835), .Y(n3833) );
  INVX2TS U2008 ( .A(n3832), .Y(n3830) );
  INVX2TS U2009 ( .A(n3829), .Y(n3827) );
  INVX2TS U2010 ( .A(n3826), .Y(n3824) );
  INVX2TS U2011 ( .A(n3823), .Y(n3821) );
  INVX2TS U2012 ( .A(n3820), .Y(n3818) );
  INVX2TS U2013 ( .A(n3934), .Y(n3932) );
  INVX2TS U2014 ( .A(n3949), .Y(n3947) );
  INVX2TS U2015 ( .A(n3943), .Y(n3941) );
  INVX2TS U2016 ( .A(n3940), .Y(n3938) );
  INVX2TS U2017 ( .A(n3937), .Y(n3935) );
  INVX2TS U2018 ( .A(n3946), .Y(n3944) );
  INVX2TS U2019 ( .A(n3931), .Y(n3929) );
  INVX2TS U2020 ( .A(n3928), .Y(n3926) );
  INVX2TS U2021 ( .A(n3922), .Y(n3920) );
  INVX2TS U2022 ( .A(n3925), .Y(n3923) );
  INVX2TS U2023 ( .A(n3919), .Y(n3917) );
  INVX2TS U2024 ( .A(n3916), .Y(n3914) );
  INVX2TS U2025 ( .A(n6217), .Y(n6249) );
  INVX2TS U2026 ( .A(n4084), .Y(n4082) );
  INVX2TS U2027 ( .A(n4087), .Y(n4085) );
  INVX2TS U2028 ( .A(n4078), .Y(n4076) );
  INVX2TS U2029 ( .A(n4081), .Y(n4079) );
  INVX2TS U2030 ( .A(n4075), .Y(n4073) );
  INVX2TS U2031 ( .A(n4072), .Y(n4070) );
  INVX2TS U2032 ( .A(n4237), .Y(n4235) );
  INVX2TS U2033 ( .A(n4234), .Y(n4232) );
  INVX2TS U2034 ( .A(n4231), .Y(n4229) );
  INVX2TS U2035 ( .A(n4228), .Y(n4226) );
  INVX2TS U2036 ( .A(n4243), .Y(n4241) );
  INVX2TS U2037 ( .A(n4240), .Y(n4238) );
  INVX2TS U2038 ( .A(n3804), .Y(n3803) );
  CLKBUFX2TS U2039 ( .A(n4415), .Y(n4417) );
  CLKBUFX2TS U2040 ( .A(n4412), .Y(n4414) );
  CLKBUFX2TS U2041 ( .A(n4409), .Y(n4411) );
  CLKBUFX2TS U2042 ( .A(n4403), .Y(n4405) );
  CLKBUFX2TS U2043 ( .A(n4400), .Y(n4402) );
  CLKBUFX2TS U2044 ( .A(n4406), .Y(n4408) );
  CLKBUFX2TS U2045 ( .A(n4376), .Y(n4378) );
  CLKBUFX2TS U2046 ( .A(n4373), .Y(n4375) );
  CLKBUFX2TS U2047 ( .A(n4364), .Y(n4366) );
  CLKBUFX2TS U2048 ( .A(n4361), .Y(n4363) );
  CLKBUFX2TS U2049 ( .A(n4349), .Y(n4351) );
  CLKBUFX2TS U2050 ( .A(n4343), .Y(n4345) );
  CLKBUFX2TS U2051 ( .A(n4340), .Y(n4342) );
  CLKBUFX2TS U2052 ( .A(n4337), .Y(n4339) );
  CLKBUFX2TS U2053 ( .A(n4331), .Y(n4333) );
  CLKBUFX2TS U2054 ( .A(n4328), .Y(n4330) );
  CLKBUFX2TS U2055 ( .A(n4325), .Y(n4327) );
  CLKBUFX2TS U2056 ( .A(n4322), .Y(n4324) );
  CLKBUFX2TS U2057 ( .A(n4319), .Y(n4321) );
  CLKBUFX2TS U2058 ( .A(n4316), .Y(n4318) );
  CLKBUFX2TS U2059 ( .A(n4310), .Y(n4312) );
  CLKBUFX2TS U2060 ( .A(n4298), .Y(n4300) );
  CLKBUFX2TS U2061 ( .A(n4295), .Y(n4297) );
  CLKBUFX2TS U2062 ( .A(n4370), .Y(n4372) );
  CLKBUFX2TS U2063 ( .A(n4367), .Y(n4369) );
  CLKBUFX2TS U2064 ( .A(n4355), .Y(n4357) );
  CLKBUFX2TS U2065 ( .A(n4346), .Y(n4348) );
  CLKBUFX2TS U2066 ( .A(n4313), .Y(n4315) );
  CLKBUFX2TS U2067 ( .A(n4301), .Y(n4303) );
  CLKBUFX2TS U2068 ( .A(n4289), .Y(n4291) );
  CLKBUFX2TS U2069 ( .A(n4379), .Y(n4381) );
  CLKBUFX2TS U2070 ( .A(n4358), .Y(n4360) );
  CLKBUFX2TS U2071 ( .A(n4352), .Y(n4354) );
  CLKBUFX2TS U2072 ( .A(n4334), .Y(n4336) );
  CLKBUFX2TS U2073 ( .A(n4304), .Y(n4306) );
  CLKBUFX2TS U2074 ( .A(n4292), .Y(n4294) );
  CLKBUFX2TS U2075 ( .A(n4286), .Y(n4288) );
  CLKBUFX2TS U2076 ( .A(n4307), .Y(n4309) );
  INVX2TS U2077 ( .A(n4009), .Y(n4007) );
  INVX2TS U2078 ( .A(n3979), .Y(n3977) );
  INVX2TS U2079 ( .A(n4066), .Y(n4064) );
  INVX2TS U2080 ( .A(n4063), .Y(n4061) );
  INVX2TS U2081 ( .A(n4060), .Y(n4058) );
  INVX2TS U2082 ( .A(n4057), .Y(n4055) );
  INVX2TS U2083 ( .A(n4054), .Y(n4052) );
  INVX2TS U2084 ( .A(n4051), .Y(n4049) );
  INVX2TS U2085 ( .A(n4045), .Y(n4043) );
  INVX2TS U2086 ( .A(n4039), .Y(n4037) );
  INVX2TS U2087 ( .A(n4036), .Y(n4034) );
  INVX2TS U2088 ( .A(n4033), .Y(n4031) );
  INVX2TS U2089 ( .A(n4030), .Y(n4028) );
  INVX2TS U2090 ( .A(n4015), .Y(n4013) );
  INVX2TS U2091 ( .A(n4012), .Y(n4010) );
  INVX2TS U2092 ( .A(n4006), .Y(n4004) );
  INVX2TS U2093 ( .A(n4003), .Y(n4001) );
  INVX2TS U2094 ( .A(n4000), .Y(n3998) );
  INVX2TS U2095 ( .A(n3997), .Y(n3995) );
  INVX2TS U2096 ( .A(n3991), .Y(n3989) );
  INVX2TS U2097 ( .A(n3988), .Y(n3986) );
  INVX2TS U2098 ( .A(n4069), .Y(n4067) );
  INVX2TS U2099 ( .A(n4048), .Y(n4046) );
  INVX2TS U2100 ( .A(n4042), .Y(n4040) );
  INVX2TS U2101 ( .A(n4024), .Y(n4022) );
  INVX2TS U2102 ( .A(n3994), .Y(n3992) );
  INVX2TS U2103 ( .A(n3982), .Y(n3980) );
  INVX2TS U2104 ( .A(n3976), .Y(n3974) );
  INVX2TS U2105 ( .A(n4027), .Y(n4025) );
  INVX2TS U2106 ( .A(n4021), .Y(n4019) );
  INVX2TS U2107 ( .A(n4018), .Y(n4016) );
  INVX2TS U2108 ( .A(n3985), .Y(n3983) );
  INVX2TS U2109 ( .A(n4105), .Y(n4103) );
  INVX2TS U2110 ( .A(n4102), .Y(n4100) );
  INVX2TS U2111 ( .A(n4099), .Y(n4097) );
  INVX2TS U2112 ( .A(n4096), .Y(n4094) );
  INVX2TS U2113 ( .A(n4093), .Y(n4091) );
  INVX2TS U2114 ( .A(n4090), .Y(n4088) );
  INVX2TS U2115 ( .A(n3817), .Y(n3815) );
  CLKBUFX2TS U2116 ( .A(n3968), .Y(n3969) );
  CLKBUFX2TS U2117 ( .A(n3956), .Y(n3957) );
  CLKBUFX2TS U2118 ( .A(n3950), .Y(n3951) );
  CLKBUFX2TS U2119 ( .A(n3965), .Y(n3966) );
  CLKBUFX2TS U2120 ( .A(n3959), .Y(n3960) );
  CLKBUFX2TS U2121 ( .A(n3971), .Y(n3972) );
  CLKBUFX2TS U2122 ( .A(n3962), .Y(n3963) );
  CLKBUFX2TS U2123 ( .A(n3953), .Y(n3954) );
  CLKBUFX2TS U2124 ( .A(n4280), .Y(n4281) );
  CLKBUFX2TS U2125 ( .A(n4274), .Y(n4275) );
  CLKBUFX2TS U2126 ( .A(n4271), .Y(n4272) );
  CLKBUFX2TS U2127 ( .A(n4283), .Y(n4284) );
  CLKBUFX2TS U2128 ( .A(n4277), .Y(n4278) );
  CLKBUFX2TS U2129 ( .A(n4268), .Y(n4269) );
  CLKBUFX2TS U2130 ( .A(n4127), .Y(n4128) );
  CLKBUFX2TS U2131 ( .A(n4124), .Y(n4125) );
  CLKBUFX2TS U2132 ( .A(n4118), .Y(n4119) );
  CLKBUFX2TS U2133 ( .A(n4112), .Y(n4113) );
  CLKBUFX2TS U2134 ( .A(n4106), .Y(n4107) );
  CLKBUFX2TS U2135 ( .A(n4121), .Y(n4122) );
  CLKBUFX2TS U2136 ( .A(n4115), .Y(n4116) );
  CLKBUFX2TS U2137 ( .A(n4109), .Y(n4110) );
  CLKBUFX2TS U2138 ( .A(n4124), .Y(n4126) );
  CLKBUFX2TS U2139 ( .A(n4106), .Y(n4108) );
  CLKBUFX2TS U2140 ( .A(n3968), .Y(n3970) );
  CLKBUFX2TS U2141 ( .A(n3962), .Y(n3964) );
  CLKBUFX2TS U2142 ( .A(n3950), .Y(n3952) );
  CLKBUFX2TS U2143 ( .A(n4118), .Y(n4120) );
  CLKBUFX2TS U2144 ( .A(n4115), .Y(n4117) );
  CLKBUFX2TS U2145 ( .A(n3959), .Y(n3961) );
  CLKBUFX2TS U2146 ( .A(n3971), .Y(n3973) );
  CLKBUFX2TS U2147 ( .A(n4127), .Y(n4129) );
  CLKBUFX2TS U2148 ( .A(n3965), .Y(n3967) );
  CLKBUFX2TS U2149 ( .A(n4121), .Y(n4123) );
  CLKBUFX2TS U2150 ( .A(n3956), .Y(n3958) );
  CLKBUFX2TS U2151 ( .A(n4112), .Y(n4114) );
  CLKBUFX2TS U2152 ( .A(n3953), .Y(n3955) );
  CLKBUFX2TS U2153 ( .A(n4109), .Y(n4111) );
  CLKBUFX2TS U2154 ( .A(n4280), .Y(n4282) );
  CLKBUFX2TS U2155 ( .A(n4268), .Y(n4270) );
  CLKBUFX2TS U2156 ( .A(n4277), .Y(n4279) );
  CLKBUFX2TS U2157 ( .A(n4271), .Y(n4273) );
  CLKBUFX2TS U2158 ( .A(n4283), .Y(n4285) );
  CLKBUFX2TS U2159 ( .A(n4274), .Y(n4276) );
  CLKBUFX2TS U2160 ( .A(n4394), .Y(n4396) );
  CLKBUFX2TS U2161 ( .A(n4385), .Y(n4387) );
  CLKBUFX2TS U2162 ( .A(n4382), .Y(n4384) );
  CLKBUFX2TS U2163 ( .A(n4397), .Y(n4399) );
  CLKBUFX2TS U2164 ( .A(n4391), .Y(n4393) );
  CLKBUFX2TS U2165 ( .A(n4388), .Y(n4390) );
  INVX2TS U2166 ( .A(n3801), .Y(n3799) );
  INVX2TS U2167 ( .A(n3814), .Y(n3812) );
  INVX2TS U2168 ( .A(n3807), .Y(n3805) );
  INVX2TS U2169 ( .A(n3859), .Y(n3858) );
  INVX2TS U2170 ( .A(n3907), .Y(n3906) );
  INVX2TS U2171 ( .A(n3883), .Y(n3882) );
  INVX2TS U2172 ( .A(n3856), .Y(n3855) );
  INVX2TS U2173 ( .A(n3850), .Y(n3849) );
  INVX2TS U2174 ( .A(n3838), .Y(n3837) );
  INVX2TS U2175 ( .A(n3913), .Y(n3912) );
  INVX2TS U2176 ( .A(n3910), .Y(n3909) );
  INVX2TS U2177 ( .A(n3898), .Y(n3897) );
  INVX2TS U2178 ( .A(n3892), .Y(n3891) );
  INVX2TS U2179 ( .A(n3886), .Y(n3885) );
  INVX2TS U2180 ( .A(n3877), .Y(n3876) );
  INVX2TS U2181 ( .A(n3868), .Y(n3867) );
  INVX2TS U2182 ( .A(n3853), .Y(n3852) );
  INVX2TS U2183 ( .A(n3844), .Y(n3843) );
  INVX2TS U2184 ( .A(n3904), .Y(n3903) );
  INVX2TS U2185 ( .A(n3901), .Y(n3900) );
  INVX2TS U2186 ( .A(n3889), .Y(n3888) );
  INVX2TS U2187 ( .A(n3880), .Y(n3879) );
  INVX2TS U2188 ( .A(n3847), .Y(n3846) );
  INVX2TS U2189 ( .A(n3835), .Y(n3834) );
  INVX2TS U2190 ( .A(n3826), .Y(n3825) );
  INVX2TS U2191 ( .A(n3823), .Y(n3822) );
  INVX2TS U2192 ( .A(n3820), .Y(n3819) );
  INVX2TS U2193 ( .A(n3841), .Y(n3840) );
  INVX2TS U2194 ( .A(n3871), .Y(n3870) );
  INVX2TS U2195 ( .A(n3865), .Y(n3864) );
  INVX2TS U2196 ( .A(n3862), .Y(n3861) );
  INVX2TS U2197 ( .A(n3829), .Y(n3828) );
  INVX2TS U2198 ( .A(n3895), .Y(n3894) );
  INVX2TS U2199 ( .A(n3874), .Y(n3873) );
  INVX2TS U2200 ( .A(n3832), .Y(n3831) );
  INVX2TS U2201 ( .A(n3949), .Y(n3948) );
  INVX2TS U2202 ( .A(n3946), .Y(n3945) );
  INVX2TS U2203 ( .A(n3943), .Y(n3942) );
  INVX2TS U2204 ( .A(n3937), .Y(n3936) );
  INVX2TS U2205 ( .A(n3934), .Y(n3933) );
  INVX2TS U2206 ( .A(n3940), .Y(n3939) );
  INVX2TS U2207 ( .A(n3801), .Y(n3800) );
  INVX2TS U2208 ( .A(n4258), .Y(n4257) );
  INVX2TS U2209 ( .A(n4246), .Y(n4245) );
  INVX2TS U2210 ( .A(n4261), .Y(n4260) );
  INVX2TS U2211 ( .A(n4255), .Y(n4254) );
  INVX2TS U2212 ( .A(n4252), .Y(n4251) );
  INVX2TS U2213 ( .A(n4249), .Y(n4248) );
  INVX2TS U2214 ( .A(n4222), .Y(n4221) );
  INVX2TS U2215 ( .A(n4219), .Y(n4218) );
  INVX2TS U2216 ( .A(n4216), .Y(n4215) );
  INVX2TS U2217 ( .A(n4213), .Y(n4212) );
  INVX2TS U2218 ( .A(n4210), .Y(n4209) );
  INVX2TS U2219 ( .A(n4207), .Y(n4206) );
  INVX2TS U2220 ( .A(n4201), .Y(n4200) );
  INVX2TS U2221 ( .A(n4195), .Y(n4194) );
  INVX2TS U2222 ( .A(n4192), .Y(n4191) );
  INVX2TS U2223 ( .A(n4189), .Y(n4188) );
  INVX2TS U2224 ( .A(n4186), .Y(n4185) );
  INVX2TS U2225 ( .A(n4183), .Y(n4182) );
  INVX2TS U2226 ( .A(n4177), .Y(n4176) );
  INVX2TS U2227 ( .A(n4174), .Y(n4173) );
  INVX2TS U2228 ( .A(n4171), .Y(n4170) );
  INVX2TS U2229 ( .A(n4168), .Y(n4167) );
  INVX2TS U2230 ( .A(n4165), .Y(n4164) );
  INVX2TS U2231 ( .A(n4162), .Y(n4161) );
  INVX2TS U2232 ( .A(n4159), .Y(n4158) );
  INVX2TS U2233 ( .A(n4156), .Y(n4155) );
  INVX2TS U2234 ( .A(n4153), .Y(n4152) );
  INVX2TS U2235 ( .A(n4147), .Y(n4146) );
  INVX2TS U2236 ( .A(n4144), .Y(n4143) );
  INVX2TS U2237 ( .A(n4141), .Y(n4140) );
  INVX2TS U2238 ( .A(n4135), .Y(n4134) );
  INVX2TS U2239 ( .A(n4225), .Y(n4224) );
  INVX2TS U2240 ( .A(n4204), .Y(n4203) );
  INVX2TS U2241 ( .A(n4198), .Y(n4197) );
  INVX2TS U2242 ( .A(n4180), .Y(n4179) );
  INVX2TS U2243 ( .A(n4150), .Y(n4149) );
  INVX2TS U2244 ( .A(n4138), .Y(n4137) );
  INVX2TS U2245 ( .A(n4132), .Y(n4131) );
  INVX2TS U2246 ( .A(n3814), .Y(n3813) );
  INVX2TS U2247 ( .A(n4243), .Y(n4242) );
  INVX2TS U2248 ( .A(n4240), .Y(n4239) );
  INVX2TS U2249 ( .A(n4234), .Y(n4233) );
  INVX2TS U2250 ( .A(n4237), .Y(n4236) );
  INVX2TS U2251 ( .A(n4231), .Y(n4230) );
  INVX2TS U2252 ( .A(n4228), .Y(n4227) );
  INVX2TS U2253 ( .A(n3807), .Y(n3806) );
  INVX2TS U2254 ( .A(n4069), .Y(n4068) );
  INVX2TS U2255 ( .A(n4066), .Y(n4065) );
  INVX2TS U2256 ( .A(n4063), .Y(n4062) );
  INVX2TS U2257 ( .A(n4060), .Y(n4059) );
  INVX2TS U2258 ( .A(n4057), .Y(n4056) );
  INVX2TS U2259 ( .A(n4054), .Y(n4053) );
  INVX2TS U2260 ( .A(n4048), .Y(n4047) );
  INVX2TS U2261 ( .A(n4045), .Y(n4044) );
  INVX2TS U2262 ( .A(n4042), .Y(n4041) );
  INVX2TS U2263 ( .A(n4039), .Y(n4038) );
  INVX2TS U2264 ( .A(n4036), .Y(n4035) );
  INVX2TS U2265 ( .A(n4033), .Y(n4032) );
  INVX2TS U2266 ( .A(n4027), .Y(n4026) );
  INVX2TS U2267 ( .A(n4024), .Y(n4023) );
  INVX2TS U2268 ( .A(n4021), .Y(n4020) );
  INVX2TS U2269 ( .A(n4018), .Y(n4017) );
  INVX2TS U2270 ( .A(n4015), .Y(n4014) );
  INVX2TS U2271 ( .A(n4012), .Y(n4011) );
  INVX2TS U2272 ( .A(n4009), .Y(n4008) );
  INVX2TS U2273 ( .A(n4006), .Y(n4005) );
  INVX2TS U2274 ( .A(n4003), .Y(n4002) );
  INVX2TS U2275 ( .A(n4000), .Y(n3999) );
  INVX2TS U2276 ( .A(n3997), .Y(n3996) );
  INVX2TS U2277 ( .A(n3994), .Y(n3993) );
  INVX2TS U2278 ( .A(n3991), .Y(n3990) );
  INVX2TS U2279 ( .A(n3985), .Y(n3984) );
  INVX2TS U2280 ( .A(n3982), .Y(n3981) );
  INVX2TS U2281 ( .A(n3979), .Y(n3978) );
  INVX2TS U2282 ( .A(n3976), .Y(n3975) );
  INVX2TS U2283 ( .A(n4051), .Y(n4050) );
  INVX2TS U2284 ( .A(n4030), .Y(n4029) );
  INVX2TS U2285 ( .A(n3988), .Y(n3987) );
  INVX2TS U2286 ( .A(n4090), .Y(n4089) );
  INVX2TS U2287 ( .A(n4105), .Y(n4104) );
  INVX2TS U2288 ( .A(n4099), .Y(n4098) );
  INVX2TS U2289 ( .A(n4096), .Y(n4095) );
  INVX2TS U2290 ( .A(n4093), .Y(n4092) );
  INVX2TS U2291 ( .A(n4102), .Y(n4101) );
  INVX2TS U2292 ( .A(n4087), .Y(n4086) );
  INVX2TS U2293 ( .A(n4084), .Y(n4083) );
  INVX2TS U2294 ( .A(n4081), .Y(n4080) );
  INVX2TS U2295 ( .A(n4078), .Y(n4077) );
  INVX2TS U2296 ( .A(n4075), .Y(n4074) );
  INVX2TS U2297 ( .A(n4072), .Y(n4071) );
  INVX2TS U2298 ( .A(n3925), .Y(n3924) );
  INVX2TS U2299 ( .A(n3922), .Y(n3921) );
  INVX2TS U2300 ( .A(n3919), .Y(n3918) );
  INVX2TS U2301 ( .A(n3916), .Y(n3915) );
  INVX2TS U2302 ( .A(n3931), .Y(n3930) );
  INVX2TS U2303 ( .A(n3928), .Y(n3927) );
  INVX2TS U2304 ( .A(n3817), .Y(n3816) );
  INVX2TS U2305 ( .A(n3804), .Y(n3802) );
  INVX2TS U2306 ( .A(n4261), .Y(n4259) );
  INVX2TS U2307 ( .A(n4255), .Y(n4253) );
  INVX2TS U2308 ( .A(n4249), .Y(n4247) );
  INVX2TS U2309 ( .A(n4246), .Y(n4244) );
  INVX2TS U2310 ( .A(n4252), .Y(n4250) );
  INVX2TS U2311 ( .A(n4171), .Y(n4169) );
  INVX2TS U2312 ( .A(n4219), .Y(n4217) );
  INVX2TS U2313 ( .A(n4195), .Y(n4193) );
  INVX2TS U2314 ( .A(n4168), .Y(n4166) );
  INVX2TS U2315 ( .A(n4162), .Y(n4160) );
  INVX2TS U2316 ( .A(n4150), .Y(n4148) );
  INVX2TS U2317 ( .A(n4225), .Y(n4223) );
  INVX2TS U2318 ( .A(n4222), .Y(n4220) );
  INVX2TS U2319 ( .A(n4210), .Y(n4208) );
  INVX2TS U2320 ( .A(n4204), .Y(n4202) );
  INVX2TS U2321 ( .A(n4198), .Y(n4196) );
  INVX2TS U2322 ( .A(n4189), .Y(n4187) );
  INVX2TS U2323 ( .A(n4180), .Y(n4178) );
  INVX2TS U2324 ( .A(n4165), .Y(n4163) );
  INVX2TS U2325 ( .A(n4156), .Y(n4154) );
  INVX2TS U2326 ( .A(n4216), .Y(n4214) );
  INVX2TS U2327 ( .A(n4213), .Y(n4211) );
  INVX2TS U2328 ( .A(n4201), .Y(n4199) );
  INVX2TS U2329 ( .A(n4192), .Y(n4190) );
  INVX2TS U2330 ( .A(n4159), .Y(n4157) );
  INVX2TS U2331 ( .A(n4147), .Y(n4145) );
  INVX2TS U2332 ( .A(n4138), .Y(n4136) );
  INVX2TS U2333 ( .A(n4135), .Y(n4133) );
  INVX2TS U2334 ( .A(n4132), .Y(n4130) );
  INVX2TS U2335 ( .A(n4153), .Y(n4151) );
  INVX2TS U2336 ( .A(n4183), .Y(n4181) );
  INVX2TS U2337 ( .A(n4177), .Y(n4175) );
  INVX2TS U2338 ( .A(n4174), .Y(n4172) );
  INVX2TS U2339 ( .A(n4141), .Y(n4139) );
  INVX2TS U2340 ( .A(n4258), .Y(n4256) );
  INVX2TS U2341 ( .A(n4207), .Y(n4205) );
  INVX2TS U2342 ( .A(n4186), .Y(n4184) );
  INVX2TS U2343 ( .A(n4144), .Y(n4142) );
  INVX2TS U2344 ( .A(n4844), .Y(n6323) );
  INVX2TS U2345 ( .A(n4841), .Y(n6322) );
  CLKBUFX2TS U2346 ( .A(n659), .Y(n612) );
  CLKBUFX2TS U2347 ( .A(n659), .Y(n613) );
  CLKBUFX2TS U2348 ( .A(n624), .Y(n614) );
  CLKBUFX2TS U2349 ( .A(n624), .Y(n622) );
  CLKBUFX2TS U2350 ( .A(n624), .Y(n623) );
  CLKBUFX2TS U2351 ( .A(n245), .Y(n3617) );
  CLKBUFX2TS U2352 ( .A(n8), .Y(n3694) );
  CLKBUFX2TS U2353 ( .A(n8), .Y(n3695) );
  CLKBUFX2TS U2354 ( .A(n245), .Y(n3618) );
  CLKBUFX2TS U2355 ( .A(n1), .Y(n3665) );
  CLKBUFX2TS U2356 ( .A(n6318), .Y(n3633) );
  CLKBUFX2TS U2357 ( .A(n6317), .Y(n3602) );
  INVX2TS U2358 ( .A(n5282), .Y(n6320) );
  CLKBUFX2TS U2359 ( .A(n3634), .Y(n3628) );
  CLKBUFX2TS U2360 ( .A(n6318), .Y(n3634) );
  CLKBUFX2TS U2361 ( .A(n3603), .Y(n3597) );
  CLKBUFX2TS U2362 ( .A(n6317), .Y(n3603) );
  INVX2TS U2363 ( .A(n5294), .Y(n6319) );
  CLKBUFX2TS U2364 ( .A(n611), .Y(n609) );
  CLKBUFX2TS U2365 ( .A(n611), .Y(n610) );
  NOR2X1TS U2366 ( .A(n6331), .B(n5483), .Y(n5559) );
  NOR2X1TS U2367 ( .A(n5521), .B(n5483), .Y(n5552) );
  AOI21X1TS U2368 ( .A0(n6246), .A1(n481), .B0(n5344), .Y(n5311) );
  XNOR2X1TS U2369 ( .A(n4854), .B(n4858), .Y(n6226) );
  XNOR2X1TS U2370 ( .A(n4857), .B(n5323), .Y(n4854) );
  XNOR2X1TS U2371 ( .A(n164), .B(n6226), .Y(n4855) );
  NOR3X1TS U2372 ( .A(n6324), .B(n300), .C(n6245), .Y(n4857) );
  OAI211X1TS U2373 ( .A0(n4849), .A1(n4848), .B0(n4847), .C0(n4846), .Y(n4852)
         );
  NAND3BX1TS U2374 ( .AN(n6222), .B(n6220), .C(n4844), .Y(n4847) );
  OAI21X1TS U2375 ( .A0(n188), .A1(n4861), .B0(n4845), .Y(n4846) );
  OAI32X1TS U2376 ( .A0(n4845), .A1(n188), .A2(n4861), .B0(n6222), .B1(n4853), 
        .Y(n4848) );
  XOR2X1TS U2377 ( .A(n4863), .B(n4862), .Y(n6225) );
  NOR3X1TS U2378 ( .A(n4861), .B(n6324), .C(n188), .Y(n4862) );
  XNOR2X1TS U2379 ( .A(n5326), .B(n4860), .Y(n4863) );
  AOI22X1TS U2380 ( .A0(n4859), .A1(n219), .B0(n4858), .B1(n4857), .Y(n4860)
         );
  INVX2TS U2381 ( .A(n4839), .Y(n6244) );
  INVX2TS U2382 ( .A(n4850), .Y(n6245) );
  OAI221XLTS U2383 ( .A0(n5576), .A1(n264), .B0(n3409), .B1(n17), .C0(n5575), 
        .Y(n2576) );
  OAI221XLTS U2384 ( .A0(n5580), .A1(n263), .B0(n3540), .B1(n6315), .C0(n5579), 
        .Y(n2578) );
  AOI222XLTS U2385 ( .A0(n3799), .A1(n3482), .B0(n3813), .B1(n3494), .C0(n3806), .C1(n3530), .Y(n5579) );
  AOI211X1TS U2386 ( .A0(n6222), .A1(n4853), .B0(n6323), .C0(n6245), .Y(n4849)
         );
  NOR2X1TS U2387 ( .A(n6330), .B(n5326), .Y(n5551) );
  OAI33XLTS U2388 ( .A0(n6233), .A1(n6329), .A2(n5536), .B0(n3811), .B1(n6340), 
        .B2(n5535), .Y(n5537) );
  XOR2X1TS U2389 ( .A(n4851), .B(n9), .Y(n6229) );
  NAND2X1TS U2390 ( .A(n4850), .B(n4852), .Y(n4851) );
  NAND2X1TS U2391 ( .A(n3802), .B(n6339), .Y(n5519) );
  INVX2TS U2392 ( .A(n3810), .Y(n3809) );
  NAND2X1TS U2393 ( .A(n3802), .B(n6336), .Y(n5547) );
  INVX2TS U2394 ( .A(n5309), .Y(n677) );
  NAND4X1TS U2395 ( .A(n5303), .B(n5301), .C(n5299), .D(n4869), .Y(n5309) );
  AND3X2TS U2396 ( .A(n5291), .B(n5302), .C(n5300), .Y(n4869) );
  NOR2X1TS U2397 ( .A(n5302), .B(n6247), .Y(n5278) );
  NOR2X1TS U2398 ( .A(n5303), .B(n6247), .Y(n5277) );
  OAI2BB2XLTS U2399 ( .B0(n238), .B1(n6233), .A0N(n5515), .A1N(n3815), .Y(
        n5542) );
  OAI222X1TS U2400 ( .A0(n3804), .A1(n5303), .B0(n3810), .B1(n5302), .C0(n215), 
        .C1(n5301), .Y(n5304) );
  OR2X2TS U2401 ( .A(n5300), .B(n6247), .Y(n479) );
  OAI211X1TS U2402 ( .A0(n3817), .A1(n5300), .B0(n5299), .C0(n6248), .Y(n5305)
         );
  INVX2TS U2403 ( .A(n5291), .Y(n6247) );
  NOR2X1TS U2404 ( .A(n6248), .B(reset), .Y(n6217) );
  NOR2X1TS U2405 ( .A(n5299), .B(n395), .Y(n5214) );
  INVX2TS U2406 ( .A(readIn_NORTH), .Y(n3817) );
  INVX2TS U2407 ( .A(writeIn_SOUTH), .Y(n3814) );
  INVX2TS U2408 ( .A(writeIn_WEST), .Y(n3801) );
  OAI221XLTS U2409 ( .A0(n263), .A1(n5300), .B0(n3807), .B1(n5302), .C0(n6248), 
        .Y(n5290) );
  INVX2TS U2410 ( .A(readIn_WEST), .Y(n3804) );
  INVX2TS U2411 ( .A(requesterAddressIn_WEST[4]), .Y(n3928) );
  INVX2TS U2412 ( .A(requesterAddressIn_WEST[1]), .Y(n3919) );
  INVX2TS U2413 ( .A(requesterAddressIn_WEST[0]), .Y(n3916) );
  INVX2TS U2414 ( .A(requesterAddressIn_WEST[5]), .Y(n3931) );
  INVX2TS U2415 ( .A(requesterAddressIn_WEST[3]), .Y(n3925) );
  INVX2TS U2416 ( .A(requesterAddressIn_WEST[2]), .Y(n3922) );
  INVX2TS U2417 ( .A(requesterAddressIn_EAST[5]), .Y(n4087) );
  INVX2TS U2418 ( .A(requesterAddressIn_EAST[3]), .Y(n4081) );
  INVX2TS U2419 ( .A(requesterAddressIn_EAST[4]), .Y(n4084) );
  INVX2TS U2420 ( .A(requesterAddressIn_EAST[2]), .Y(n4078) );
  INVX2TS U2421 ( .A(requesterAddressIn_EAST[1]), .Y(n4075) );
  INVX2TS U2422 ( .A(requesterAddressIn_EAST[0]), .Y(n4072) );
  INVX2TS U2423 ( .A(dataIn_EAST[31]), .Y(n4069) );
  INVX2TS U2424 ( .A(dataIn_EAST[30]), .Y(n4066) );
  INVX2TS U2425 ( .A(dataIn_EAST[29]), .Y(n4063) );
  INVX2TS U2426 ( .A(dataIn_EAST[26]), .Y(n4054) );
  INVX2TS U2427 ( .A(dataIn_EAST[24]), .Y(n4048) );
  INVX2TS U2428 ( .A(dataIn_EAST[22]), .Y(n4042) );
  INVX2TS U2429 ( .A(dataIn_EAST[21]), .Y(n4039) );
  INVX2TS U2430 ( .A(dataIn_EAST[19]), .Y(n4033) );
  INVX2TS U2431 ( .A(dataIn_EAST[17]), .Y(n4027) );
  INVX2TS U2432 ( .A(dataIn_EAST[16]), .Y(n4024) );
  INVX2TS U2433 ( .A(dataIn_EAST[14]), .Y(n4018) );
  INVX2TS U2434 ( .A(dataIn_EAST[12]), .Y(n4012) );
  INVX2TS U2435 ( .A(dataIn_EAST[11]), .Y(n4009) );
  INVX2TS U2436 ( .A(dataIn_EAST[10]), .Y(n4006) );
  INVX2TS U2437 ( .A(dataIn_EAST[8]), .Y(n4000) );
  INVX2TS U2438 ( .A(dataIn_EAST[6]), .Y(n3994) );
  INVX2TS U2439 ( .A(dataIn_EAST[3]), .Y(n3985) );
  INVX2TS U2440 ( .A(dataIn_EAST[25]), .Y(n4051) );
  INVX2TS U2441 ( .A(dataIn_EAST[18]), .Y(n4030) );
  INVX2TS U2442 ( .A(dataIn_EAST[15]), .Y(n4021) );
  INVX2TS U2443 ( .A(dataIn_EAST[13]), .Y(n4015) );
  INVX2TS U2444 ( .A(dataIn_EAST[4]), .Y(n3988) );
  INVX2TS U2445 ( .A(dataIn_EAST[28]), .Y(n4060) );
  INVX2TS U2446 ( .A(dataIn_EAST[27]), .Y(n4057) );
  INVX2TS U2447 ( .A(dataIn_EAST[23]), .Y(n4045) );
  INVX2TS U2448 ( .A(dataIn_EAST[20]), .Y(n4036) );
  INVX2TS U2449 ( .A(dataIn_EAST[9]), .Y(n4003) );
  INVX2TS U2450 ( .A(dataIn_EAST[5]), .Y(n3991) );
  INVX2TS U2451 ( .A(dataIn_EAST[2]), .Y(n3982) );
  INVX2TS U2452 ( .A(dataIn_EAST[1]), .Y(n3979) );
  INVX2TS U2453 ( .A(dataIn_EAST[0]), .Y(n3976) );
  INVX2TS U2454 ( .A(dataIn_EAST[7]), .Y(n3997) );
  INVX2TS U2455 ( .A(destinationAddressIn_EAST[5]), .Y(n4105) );
  INVX2TS U2456 ( .A(destinationAddressIn_EAST[3]), .Y(n4099) );
  INVX2TS U2457 ( .A(destinationAddressIn_EAST[1]), .Y(n4093) );
  INVX2TS U2458 ( .A(destinationAddressIn_EAST[4]), .Y(n4102) );
  INVX2TS U2459 ( .A(destinationAddressIn_EAST[0]), .Y(n4090) );
  INVX2TS U2460 ( .A(destinationAddressIn_EAST[2]), .Y(n4096) );
  INVX2TS U2461 ( .A(writeIn_EAST), .Y(n3807) );
  INVX2TS U2462 ( .A(destinationAddressIn_SOUTH[0]), .Y(n4246) );
  INVX2TS U2463 ( .A(requesterAddressIn_SOUTH[5]), .Y(n4243) );
  INVX2TS U2464 ( .A(requesterAddressIn_SOUTH[4]), .Y(n4240) );
  INVX2TS U2465 ( .A(requesterAddressIn_SOUTH[2]), .Y(n4234) );
  INVX2TS U2466 ( .A(destinationAddressIn_SOUTH[5]), .Y(n4261) );
  INVX2TS U2467 ( .A(destinationAddressIn_SOUTH[3]), .Y(n4255) );
  INVX2TS U2468 ( .A(destinationAddressIn_SOUTH[2]), .Y(n4252) );
  INVX2TS U2469 ( .A(destinationAddressIn_SOUTH[1]), .Y(n4249) );
  INVX2TS U2470 ( .A(dataIn_SOUTH[30]), .Y(n4222) );
  INVX2TS U2471 ( .A(dataIn_SOUTH[29]), .Y(n4219) );
  INVX2TS U2472 ( .A(dataIn_SOUTH[26]), .Y(n4210) );
  INVX2TS U2473 ( .A(dataIn_SOUTH[21]), .Y(n4195) );
  INVX2TS U2474 ( .A(dataIn_SOUTH[19]), .Y(n4189) );
  INVX2TS U2475 ( .A(dataIn_SOUTH[13]), .Y(n4171) );
  INVX2TS U2476 ( .A(dataIn_SOUTH[12]), .Y(n4168) );
  INVX2TS U2477 ( .A(dataIn_SOUTH[11]), .Y(n4165) );
  INVX2TS U2478 ( .A(dataIn_SOUTH[10]), .Y(n4162) );
  INVX2TS U2479 ( .A(dataIn_SOUTH[8]), .Y(n4156) );
  INVX2TS U2480 ( .A(requesterAddressIn_SOUTH[3]), .Y(n4237) );
  INVX2TS U2481 ( .A(requesterAddressIn_SOUTH[1]), .Y(n4231) );
  INVX2TS U2482 ( .A(requesterAddressIn_SOUTH[0]), .Y(n4228) );
  INVX2TS U2483 ( .A(dataIn_SOUTH[28]), .Y(n4216) );
  INVX2TS U2484 ( .A(dataIn_SOUTH[27]), .Y(n4213) );
  INVX2TS U2485 ( .A(dataIn_SOUTH[23]), .Y(n4201) );
  INVX2TS U2486 ( .A(dataIn_SOUTH[20]), .Y(n4192) );
  INVX2TS U2487 ( .A(dataIn_SOUTH[9]), .Y(n4159) );
  INVX2TS U2488 ( .A(dataIn_SOUTH[5]), .Y(n4147) );
  INVX2TS U2489 ( .A(dataIn_SOUTH[1]), .Y(n4135) );
  INVX2TS U2490 ( .A(dataIn_SOUTH[31]), .Y(n4225) );
  INVX2TS U2491 ( .A(dataIn_SOUTH[24]), .Y(n4204) );
  INVX2TS U2492 ( .A(dataIn_SOUTH[22]), .Y(n4198) );
  INVX2TS U2493 ( .A(dataIn_SOUTH[16]), .Y(n4180) );
  INVX2TS U2494 ( .A(dataIn_SOUTH[6]), .Y(n4150) );
  INVX2TS U2495 ( .A(dataIn_SOUTH[2]), .Y(n4138) );
  INVX2TS U2496 ( .A(dataIn_SOUTH[0]), .Y(n4132) );
  INVX2TS U2497 ( .A(dataIn_SOUTH[7]), .Y(n4153) );
  INVX2TS U2498 ( .A(dataIn_SOUTH[17]), .Y(n4183) );
  INVX2TS U2499 ( .A(dataIn_SOUTH[15]), .Y(n4177) );
  INVX2TS U2500 ( .A(dataIn_SOUTH[14]), .Y(n4174) );
  INVX2TS U2501 ( .A(dataIn_SOUTH[3]), .Y(n4141) );
  INVX2TS U2502 ( .A(destinationAddressIn_SOUTH[4]), .Y(n4258) );
  INVX2TS U2503 ( .A(dataIn_SOUTH[25]), .Y(n4207) );
  INVX2TS U2504 ( .A(dataIn_SOUTH[18]), .Y(n4186) );
  INVX2TS U2505 ( .A(dataIn_SOUTH[4]), .Y(n4144) );
  INVX2TS U2506 ( .A(dataIn_WEST[31]), .Y(n3913) );
  INVX2TS U2507 ( .A(dataIn_WEST[30]), .Y(n3910) );
  INVX2TS U2508 ( .A(dataIn_WEST[29]), .Y(n3907) );
  INVX2TS U2509 ( .A(dataIn_WEST[26]), .Y(n3898) );
  INVX2TS U2510 ( .A(dataIn_WEST[24]), .Y(n3892) );
  INVX2TS U2511 ( .A(dataIn_WEST[22]), .Y(n3886) );
  INVX2TS U2512 ( .A(dataIn_WEST[21]), .Y(n3883) );
  INVX2TS U2513 ( .A(dataIn_WEST[19]), .Y(n3877) );
  INVX2TS U2514 ( .A(dataIn_WEST[16]), .Y(n3868) );
  INVX2TS U2515 ( .A(dataIn_WEST[13]), .Y(n3859) );
  INVX2TS U2516 ( .A(dataIn_WEST[12]), .Y(n3856) );
  INVX2TS U2517 ( .A(dataIn_WEST[11]), .Y(n3853) );
  INVX2TS U2518 ( .A(dataIn_WEST[10]), .Y(n3850) );
  INVX2TS U2519 ( .A(dataIn_WEST[8]), .Y(n3844) );
  INVX2TS U2520 ( .A(dataIn_WEST[6]), .Y(n3838) );
  INVX2TS U2521 ( .A(dataIn_WEST[28]), .Y(n3904) );
  INVX2TS U2522 ( .A(dataIn_WEST[27]), .Y(n3901) );
  INVX2TS U2523 ( .A(dataIn_WEST[23]), .Y(n3889) );
  INVX2TS U2524 ( .A(dataIn_WEST[20]), .Y(n3880) );
  INVX2TS U2525 ( .A(dataIn_WEST[9]), .Y(n3847) );
  INVX2TS U2526 ( .A(dataIn_WEST[5]), .Y(n3835) );
  INVX2TS U2527 ( .A(dataIn_WEST[2]), .Y(n3826) );
  INVX2TS U2528 ( .A(dataIn_WEST[1]), .Y(n3823) );
  INVX2TS U2529 ( .A(dataIn_WEST[0]), .Y(n3820) );
  INVX2TS U2530 ( .A(dataIn_WEST[7]), .Y(n3841) );
  INVX2TS U2531 ( .A(dataIn_WEST[17]), .Y(n3871) );
  INVX2TS U2532 ( .A(dataIn_WEST[15]), .Y(n3865) );
  INVX2TS U2533 ( .A(dataIn_WEST[14]), .Y(n3862) );
  INVX2TS U2534 ( .A(dataIn_WEST[3]), .Y(n3829) );
  INVX2TS U2535 ( .A(dataIn_WEST[25]), .Y(n3895) );
  INVX2TS U2536 ( .A(dataIn_WEST[18]), .Y(n3874) );
  INVX2TS U2537 ( .A(dataIn_WEST[4]), .Y(n3832) );
  INVX2TS U2538 ( .A(destinationAddressIn_WEST[0]), .Y(n3934) );
  INVX2TS U2539 ( .A(destinationAddressIn_WEST[5]), .Y(n3949) );
  INVX2TS U2540 ( .A(destinationAddressIn_WEST[3]), .Y(n3943) );
  INVX2TS U2541 ( .A(destinationAddressIn_WEST[2]), .Y(n3940) );
  INVX2TS U2542 ( .A(destinationAddressIn_WEST[1]), .Y(n3937) );
  INVX2TS U2543 ( .A(destinationAddressIn_WEST[4]), .Y(n3946) );
  NOR2BX1TS U2544 ( .AN(n6228), .B(n6224), .Y(n2885) );
  AOI31X1TS U2545 ( .A0(n6223), .A1(n6323), .A2(n6222), .B0(n3585), .Y(n6224)
         );
  XNOR2X1TS U2546 ( .A(n6221), .B(n6220), .Y(n6223) );
  CLKBUFX2TS U2547 ( .A(destinationAddressIn_EAST[12]), .Y(n4124) );
  CLKBUFX2TS U2548 ( .A(destinationAddressIn_EAST[6]), .Y(n4106) );
  CLKBUFX2TS U2549 ( .A(destinationAddressIn_WEST[12]), .Y(n3968) );
  CLKBUFX2TS U2550 ( .A(destinationAddressIn_SOUTH[12]), .Y(n4280) );
  CLKBUFX2TS U2551 ( .A(destinationAddressIn_WEST[6]), .Y(n3950) );
  CLKBUFX2TS U2552 ( .A(destinationAddressIn_EAST[10]), .Y(n4118) );
  CLKBUFX2TS U2553 ( .A(destinationAddressIn_SOUTH[10]), .Y(n4274) );
  CLKBUFX2TS U2554 ( .A(destinationAddressIn_WEST[10]), .Y(n3962) );
  CLKBUFX2TS U2555 ( .A(destinationAddressIn_EAST[9]), .Y(n4115) );
  CLKBUFX2TS U2556 ( .A(destinationAddressIn_WEST[9]), .Y(n3959) );
  CLKBUFX2TS U2557 ( .A(destinationAddressIn_SOUTH[9]), .Y(n4271) );
  CLKBUFX2TS U2558 ( .A(destinationAddressIn_WEST[13]), .Y(n3971) );
  CLKBUFX2TS U2559 ( .A(destinationAddressIn_EAST[13]), .Y(n4127) );
  CLKBUFX2TS U2560 ( .A(destinationAddressIn_SOUTH[13]), .Y(n4283) );
  CLKBUFX2TS U2561 ( .A(destinationAddressIn_WEST[11]), .Y(n3965) );
  CLKBUFX2TS U2562 ( .A(destinationAddressIn_EAST[11]), .Y(n4121) );
  CLKBUFX2TS U2563 ( .A(destinationAddressIn_SOUTH[11]), .Y(n4277) );
  CLKBUFX2TS U2564 ( .A(destinationAddressIn_WEST[8]), .Y(n3956) );
  CLKBUFX2TS U2565 ( .A(destinationAddressIn_EAST[8]), .Y(n4112) );
  CLKBUFX2TS U2566 ( .A(destinationAddressIn_SOUTH[8]), .Y(n4268) );
  CLKBUFX2TS U2567 ( .A(destinationAddressIn_WEST[7]), .Y(n3953) );
  CLKBUFX2TS U2568 ( .A(destinationAddressIn_EAST[7]), .Y(n4109) );
  CLKBUFX2TS U2569 ( .A(destinationAddressIn_NORTH[0]), .Y(n4400) );
  CLKBUFX2TS U2570 ( .A(requesterAddressIn_NORTH[5]), .Y(n4397) );
  CLKBUFX2TS U2571 ( .A(requesterAddressIn_NORTH[4]), .Y(n4394) );
  CLKBUFX2TS U2572 ( .A(requesterAddressIn_NORTH[2]), .Y(n4388) );
  CLKBUFX2TS U2573 ( .A(destinationAddressIn_NORTH[5]), .Y(n4415) );
  CLKBUFX2TS U2574 ( .A(destinationAddressIn_NORTH[3]), .Y(n4409) );
  CLKBUFX2TS U2575 ( .A(destinationAddressIn_NORTH[2]), .Y(n4406) );
  CLKBUFX2TS U2576 ( .A(destinationAddressIn_NORTH[1]), .Y(n4403) );
  CLKBUFX2TS U2577 ( .A(dataIn_NORTH[30]), .Y(n4376) );
  CLKBUFX2TS U2578 ( .A(dataIn_NORTH[29]), .Y(n4373) );
  CLKBUFX2TS U2579 ( .A(dataIn_NORTH[26]), .Y(n4364) );
  CLKBUFX2TS U2580 ( .A(dataIn_NORTH[21]), .Y(n4349) );
  CLKBUFX2TS U2581 ( .A(dataIn_NORTH[19]), .Y(n4343) );
  CLKBUFX2TS U2582 ( .A(dataIn_NORTH[13]), .Y(n4325) );
  CLKBUFX2TS U2583 ( .A(dataIn_NORTH[12]), .Y(n4322) );
  CLKBUFX2TS U2584 ( .A(dataIn_NORTH[11]), .Y(n4319) );
  CLKBUFX2TS U2585 ( .A(dataIn_NORTH[10]), .Y(n4316) );
  CLKBUFX2TS U2586 ( .A(dataIn_NORTH[8]), .Y(n4310) );
  CLKBUFX2TS U2587 ( .A(requesterAddressIn_NORTH[3]), .Y(n4391) );
  CLKBUFX2TS U2588 ( .A(requesterAddressIn_NORTH[1]), .Y(n4385) );
  CLKBUFX2TS U2589 ( .A(requesterAddressIn_NORTH[0]), .Y(n4382) );
  CLKBUFX2TS U2590 ( .A(dataIn_NORTH[28]), .Y(n4370) );
  CLKBUFX2TS U2591 ( .A(dataIn_NORTH[27]), .Y(n4367) );
  CLKBUFX2TS U2592 ( .A(dataIn_NORTH[23]), .Y(n4355) );
  CLKBUFX2TS U2593 ( .A(dataIn_NORTH[20]), .Y(n4346) );
  CLKBUFX2TS U2594 ( .A(dataIn_NORTH[9]), .Y(n4313) );
  CLKBUFX2TS U2595 ( .A(dataIn_NORTH[5]), .Y(n4301) );
  CLKBUFX2TS U2596 ( .A(dataIn_NORTH[1]), .Y(n4289) );
  CLKBUFX2TS U2597 ( .A(dataIn_NORTH[31]), .Y(n4379) );
  CLKBUFX2TS U2598 ( .A(dataIn_NORTH[24]), .Y(n4358) );
  CLKBUFX2TS U2599 ( .A(dataIn_NORTH[22]), .Y(n4352) );
  CLKBUFX2TS U2600 ( .A(dataIn_NORTH[16]), .Y(n4334) );
  CLKBUFX2TS U2601 ( .A(dataIn_NORTH[6]), .Y(n4304) );
  CLKBUFX2TS U2602 ( .A(dataIn_NORTH[2]), .Y(n4292) );
  CLKBUFX2TS U2603 ( .A(dataIn_NORTH[0]), .Y(n4286) );
  CLKBUFX2TS U2604 ( .A(dataIn_NORTH[7]), .Y(n4307) );
  CLKBUFX2TS U2605 ( .A(dataIn_NORTH[17]), .Y(n4337) );
  CLKBUFX2TS U2606 ( .A(dataIn_NORTH[15]), .Y(n4331) );
  CLKBUFX2TS U2607 ( .A(dataIn_NORTH[14]), .Y(n4328) );
  CLKBUFX2TS U2608 ( .A(dataIn_NORTH[3]), .Y(n4295) );
  CLKBUFX2TS U2609 ( .A(destinationAddressIn_NORTH[4]), .Y(n4412) );
  CLKBUFX2TS U2610 ( .A(dataIn_NORTH[25]), .Y(n4361) );
  CLKBUFX2TS U2611 ( .A(dataIn_NORTH[18]), .Y(n4340) );
  CLKBUFX2TS U2612 ( .A(dataIn_NORTH[4]), .Y(n4298) );
  INVX2TS U2613 ( .A(readIn_EAST), .Y(n3811) );
  OAI21X1TS U2614 ( .A0(n6248), .A1(n6221), .B0(n4418), .Y(n6219) );
  OAI22X1TS U2615 ( .A0(n3572), .A1(n3653), .B0(n163), .B1(n6219), .Y(n2884)
         );
  XNOR2X1TS U2616 ( .A(n5326), .B(n163), .Y(n6220) );
  AOI21X1TS U2617 ( .A0(n4), .A1(n5327), .B0(n4841), .Y(n4844) );
  XNOR2X1TS U2618 ( .A(n6220), .B(n4843), .Y(n4845) );
  AOI21X1TS U2619 ( .A0(n5323), .A1(n6322), .B0(n4842), .Y(n4843) );
  AOI21X1TS U2620 ( .A0(n4841), .A1(n219), .B0(n164), .Y(n4842) );
  OAI22X1TS U2621 ( .A0(n6303), .A1(n594), .B0(n6281), .B1(n3638), .Y(n5127)
         );
  OAI22X1TS U2622 ( .A0(n6304), .A1(n584), .B0(n6282), .B1(n3637), .Y(n5135)
         );
  OAI22X1TS U2623 ( .A0(n6306), .A1(n584), .B0(n6283), .B1(n3637), .Y(n5151)
         );
  OAI22X1TS U2624 ( .A0(n6307), .A1(n584), .B0(n6310), .B1(n3637), .Y(n5159)
         );
  OAI22X1TS U2625 ( .A0(n6305), .A1(n584), .B0(n6309), .B1(n3637), .Y(n5143)
         );
  OAI22X1TS U2626 ( .A0(n6308), .A1(n582), .B0(n6311), .B1(n3636), .Y(n5167)
         );
  CLKBUFX2TS U2627 ( .A(n5297), .Y(n659) );
  CLKBUFX2TS U2628 ( .A(n5297), .Y(n624) );
  INVX2TS U2629 ( .A(n5295), .Y(n6318) );
  INVX2TS U2630 ( .A(n5285), .Y(n6317) );
  NOR2X1TS U2631 ( .A(n6221), .B(n163), .Y(n5294) );
  INVX2TS U2632 ( .A(n301), .Y(n6316) );
  CLKBUFX2TS U2633 ( .A(n660), .Y(n611) );
  CLKBUFX2TS U2634 ( .A(n5297), .Y(n660) );
  AOI222XLTS U2635 ( .A0(n3969), .A1(n111), .B0(n4282), .B1(n706), .C0(n4125), 
        .C1(n468), .Y(n5321) );
  AOI222XLTS U2636 ( .A0(n3957), .A1(n119), .B0(n4270), .B1(n705), .C0(n4113), 
        .C1(n468), .Y(n5328) );
  AOI222XLTS U2637 ( .A0(n4284), .A1(n860), .B0(destinationAddressIn_EAST[13]), 
        .B1(n843), .C0(n3973), .C1(n1822), .Y(n5367) );
  AOI222XLTS U2638 ( .A0(n3972), .A1(n123), .B0(n4285), .B1(n714), .C0(n4128), 
        .C1(n469), .Y(n5320) );
  AOI222XLTS U2639 ( .A0(n3963), .A1(n114), .B0(n4276), .B1(n706), .C0(n4119), 
        .C1(n468), .Y(n5324) );
  AOI222XLTS U2640 ( .A0(n3951), .A1(n124), .B0(n4264), .B1(n705), .C0(n4107), 
        .C1(n468), .Y(n5330) );
  AOI222XLTS U2641 ( .A0(n3799), .A1(n113), .B0(n3812), .B1(n705), .C0(n3805), 
        .C1(n469), .Y(n5564) );
  AOI222XLTS U2642 ( .A0(n4278), .A1(n860), .B0(destinationAddressIn_EAST[11]), 
        .B1(n845), .C0(n3967), .C1(n1822), .Y(n5369) );
  AOI222XLTS U2643 ( .A0(n4272), .A1(n861), .B0(destinationAddressIn_EAST[9]), 
        .B1(n845), .C0(n3961), .C1(n1894), .Y(n5371) );
  AOI222XLTS U2644 ( .A0(n4266), .A1(n861), .B0(destinationAddressIn_EAST[7]), 
        .B1(n836), .C0(n3955), .C1(n3192), .Y(n5373) );
  AOI222XLTS U2645 ( .A0(n3812), .A1(n862), .B0(n3806), .B1(n836), .C0(n3800), 
        .C1(n3192), .Y(n5569) );
  AOI222XLTS U2646 ( .A0(n3966), .A1(n117), .B0(n4279), .B1(n706), .C0(n4122), 
        .C1(n5563), .Y(n5322) );
  AOI222XLTS U2647 ( .A0(n3960), .A1(n112), .B0(n4273), .B1(n712), .C0(n4116), 
        .C1(n469), .Y(n5325) );
  AOI222XLTS U2648 ( .A0(n3954), .A1(n118), .B0(n4267), .B1(n705), .C0(n4110), 
        .C1(n469), .Y(n5329) );
  AOI222XLTS U2649 ( .A0(n4281), .A1(n860), .B0(destinationAddressIn_EAST[12]), 
        .B1(n845), .C0(n3970), .C1(n1822), .Y(n5368) );
  AOI222XLTS U2650 ( .A0(n4275), .A1(n860), .B0(destinationAddressIn_EAST[10]), 
        .B1(n845), .C0(n3964), .C1(n1894), .Y(n5370) );
  AOI222XLTS U2651 ( .A0(n4269), .A1(n861), .B0(destinationAddressIn_EAST[8]), 
        .B1(n836), .C0(n3958), .C1(n1894), .Y(n5372) );
  AOI222XLTS U2652 ( .A0(n4263), .A1(n861), .B0(destinationAddressIn_EAST[6]), 
        .B1(n836), .C0(n3952), .C1(n3192), .Y(n5374) );
  NOR2X1TS U2653 ( .A(selectBit_SOUTH), .B(selectBit_NORTH), .Y(n4868) );
  INVX2TS U2654 ( .A(selectBit_EAST), .Y(n6232) );
  INVX2TS U2655 ( .A(readReady), .Y(n6230) );
  NOR2X1TS U2656 ( .A(selectBit_WEST), .B(readReady), .Y(n4867) );
  OAI32X1TS U2657 ( .A0(n4865), .A1(n6228), .A2(n4864), .B0(n395), .B1(n96), 
        .Y(N4718) );
  NAND2X1TS U2658 ( .A(n4856), .B(n4855), .Y(n4865) );
  XNOR2X1TS U2659 ( .A(n216), .B(n6225), .Y(n4864) );
  OAI221XLTS U2660 ( .A0(n291), .A1(n272), .B0(n4777), .B1(n678), .C0(n5462), 
        .Y(n2536) );
  OAI221XLTS U2661 ( .A0(n292), .A1(n275), .B0(n4789), .B1(n679), .C0(n5464), 
        .Y(n2538) );
  OAI221XLTS U2662 ( .A0(n290), .A1(n279), .B0(n4797), .B1(n679), .C0(n5465), 
        .Y(n2539) );
  AOI222XLTS U2663 ( .A0(n4272), .A1(n3466), .B0(n4117), .B1(n3441), .C0(n3961), .C1(n3718), .Y(n5465) );
  OAI221XLTS U2664 ( .A0(n291), .A1(n267), .B0(n4821), .B1(n680), .C0(n5468), 
        .Y(n2542) );
  AOI222XLTS U2665 ( .A0(n4263), .A1(n3466), .B0(n4108), .B1(n3437), .C0(n3952), .C1(n3722), .Y(n5468) );
  OAI221XLTS U2666 ( .A0(n379), .A1(n282), .B0(n4766), .B1(n812), .C0(n5345), 
        .Y(n2465) );
  AOI222XLTS U2667 ( .A0(n4128), .A1(n758), .B0(destinationAddressIn_SOUTH[13]), .B1(n761), .C0(n3973), .C1(n808), .Y(n5345) );
  OAI221XLTS U2668 ( .A0(n378), .A1(n272), .B0(n4774), .B1(n811), .C0(n5346), 
        .Y(n2466) );
  AOI222XLTS U2669 ( .A0(n4125), .A1(n751), .B0(destinationAddressIn_SOUTH[12]), .B1(n761), .C0(n3970), .C1(n809), .Y(n5346) );
  OAI221XLTS U2670 ( .A0(n379), .A1(n285), .B0(n4784), .B1(n812), .C0(n5347), 
        .Y(n2467) );
  AOI222XLTS U2671 ( .A0(n4122), .A1(n751), .B0(destinationAddressIn_SOUTH[11]), .B1(n761), .C0(n3967), .C1(n802), .Y(n5347) );
  OAI221XLTS U2672 ( .A0(n378), .A1(n275), .B0(n4790), .B1(n812), .C0(n5348), 
        .Y(n2468) );
  AOI222XLTS U2673 ( .A0(n4119), .A1(n751), .B0(destinationAddressIn_SOUTH[10]), .B1(n761), .C0(n3964), .C1(n802), .Y(n5348) );
  OAI221XLTS U2674 ( .A0(n377), .A1(n278), .B0(n4802), .B1(n813), .C0(n5349), 
        .Y(n2469) );
  AOI222XLTS U2675 ( .A0(n4116), .A1(n751), .B0(destinationAddressIn_SOUTH[9]), 
        .B1(n762), .C0(n3961), .C1(n809), .Y(n5349) );
  OAI221XLTS U2676 ( .A0(n377), .A1(n288), .B0(n4806), .B1(n813), .C0(n5350), 
        .Y(n2470) );
  AOI222XLTS U2677 ( .A0(n4113), .A1(n750), .B0(destinationAddressIn_SOUTH[8]), 
        .B1(n762), .C0(n3958), .C1(n808), .Y(n5350) );
  OAI221XLTS U2678 ( .A0(n377), .A1(n270), .B0(n4814), .B1(n813), .C0(n5351), 
        .Y(n2471) );
  AOI222XLTS U2679 ( .A0(n4110), .A1(n750), .B0(n4265), .B1(n762), .C0(n3955), 
        .C1(n808), .Y(n5351) );
  OAI221XLTS U2680 ( .A0(n379), .A1(n266), .B0(n4826), .B1(n812), .C0(n5352), 
        .Y(n2472) );
  AOI222XLTS U2681 ( .A0(n4107), .A1(n750), .B0(n4262), .B1(n762), .C0(n3952), 
        .C1(n803), .Y(n5352) );
  OAI221XLTS U2682 ( .A0(n377), .A1(n6235), .B0(n810), .B1(n6284), .C0(n5567), 
        .Y(n2572) );
  AOI222XLTS U2683 ( .A0(n3805), .A1(n750), .B0(n3813), .B1(n763), .C0(n3800), 
        .C1(n802), .Y(n5567) );
  OAI221XLTS U2684 ( .A0(n292), .A1(n284), .B0(n4787), .B1(n678), .C0(n5463), 
        .Y(n2537) );
  OAI221XLTS U2685 ( .A0(n290), .A1(n287), .B0(n4811), .B1(n679), .C0(n5466), 
        .Y(n2540) );
  AOI222XLTS U2686 ( .A0(n4269), .A1(n3466), .B0(n4114), .B1(n3427), .C0(n3958), .C1(n3718), .Y(n5466) );
  OAI221XLTS U2687 ( .A0(n291), .A1(n269), .B0(n4817), .B1(n679), .C0(n5467), 
        .Y(n2541) );
  AOI222XLTS U2688 ( .A0(n4266), .A1(n3466), .B0(n4111), .B1(n3427), .C0(n3955), .C1(n3718), .Y(n5467) );
  OAI221XLTS U2689 ( .A0(n292), .A1(n281), .B0(n4767), .B1(n678), .C0(n5461), 
        .Y(n2535) );
  OAI221XLTS U2690 ( .A0(n290), .A1(n264), .B0(n678), .B1(n6314), .C0(n5577), 
        .Y(n2577) );
  AOI222XLTS U2691 ( .A0(n3812), .A1(n3465), .B0(n3806), .B1(n3427), .C0(n3800), .C1(n3719), .Y(n5577) );
  OAI221XLTS U2692 ( .A0(n3240), .A1(n264), .B0(n3272), .B1(n102), .C0(n5573), 
        .Y(n2574) );
  AOI222XLTS U2693 ( .A0(n3799), .A1(n3246), .B0(n3813), .B1(n3210), .C0(n3806), .C1(n463), .Y(n5573) );
  OAI221XLTS U2694 ( .A0(n313), .A1(n263), .B0(n3343), .B1(n100), .C0(n5574), 
        .Y(n2575) );
  AOI222XLTS U2695 ( .A0(n3812), .A1(n3286), .B0(n3800), .B1(n3297), .C0(n3805), .C1(n3336), .Y(n5574) );
  OAI221XLTS U2696 ( .A0(n3238), .A1(n284), .B0(n4783), .B1(n3276), .C0(n5395), 
        .Y(n2495) );
  AOI222XLTS U2697 ( .A0(n3966), .A1(n3244), .B0(n4279), .B1(n3205), .C0(n4123), .C1(n463), .Y(n5395) );
  OAI221XLTS U2698 ( .A0(n3240), .A1(n266), .B0(n4823), .B1(n3276), .C0(n5400), 
        .Y(n2500) );
  AOI222XLTS U2699 ( .A0(n3951), .A1(n3245), .B0(n4264), .B1(n3212), .C0(n4108), .C1(n463), .Y(n5400) );
  OAI221XLTS U2700 ( .A0(n381), .A1(n272), .B0(n4775), .B1(n3344), .C0(n5416), 
        .Y(n2508) );
  AOI222XLTS U2701 ( .A0(n4281), .A1(n3294), .B0(n3970), .B1(n3295), .C0(n4126), .C1(n3335), .Y(n5416) );
  OAI221XLTS U2702 ( .A0(n382), .A1(n284), .B0(n4781), .B1(n3345), .C0(n5417), 
        .Y(n2509) );
  AOI222XLTS U2703 ( .A0(n4278), .A1(n3294), .B0(n3967), .B1(n3295), .C0(n4123), .C1(n3335), .Y(n5417) );
  OAI221XLTS U2704 ( .A0(n382), .A1(n275), .B0(n4791), .B1(n3345), .C0(n5418), 
        .Y(n2510) );
  AOI222XLTS U2705 ( .A0(n4275), .A1(n3285), .B0(n3964), .B1(n3295), .C0(n4120), .C1(n3335), .Y(n5418) );
  OAI221XLTS U2706 ( .A0(n381), .A1(n287), .B0(n4809), .B1(n3346), .C0(n5420), 
        .Y(n2512) );
  AOI222XLTS U2707 ( .A0(n4269), .A1(n3286), .B0(n3958), .B1(n3296), .C0(n4114), .C1(n3336), .Y(n5420) );
  OAI221XLTS U2708 ( .A0(n381), .A1(n269), .B0(n4813), .B1(n3346), .C0(n5421), 
        .Y(n2513) );
  AOI222XLTS U2709 ( .A0(n4266), .A1(n3286), .B0(n3955), .B1(n3296), .C0(n4111), .C1(n3336), .Y(n5421) );
  OAI221XLTS U2710 ( .A0(n381), .A1(n266), .B0(n4825), .B1(n3345), .C0(n5422), 
        .Y(n2514) );
  AOI222XLTS U2711 ( .A0(n4263), .A1(n3294), .B0(n3952), .B1(n3296), .C0(n4108), .C1(n3338), .Y(n5422) );
  OAI221XLTS U2712 ( .A0(n3238), .A1(n273), .B0(n4776), .B1(n3273), .C0(n5394), 
        .Y(n2494) );
  AOI222XLTS U2713 ( .A0(n3969), .A1(n3244), .B0(n4282), .B1(n3205), .C0(n4126), .C1(n463), .Y(n5394) );
  OAI221XLTS U2714 ( .A0(n3239), .A1(n278), .B0(n4798), .B1(n3274), .C0(n5397), 
        .Y(n2497) );
  AOI222XLTS U2715 ( .A0(n3960), .A1(n3245), .B0(n4273), .B1(n3205), .C0(n4117), .C1(n5572), .Y(n5397) );
  OAI221XLTS U2716 ( .A0(n3239), .A1(n287), .B0(n4812), .B1(n3275), .C0(n5398), 
        .Y(n2498) );
  AOI222XLTS U2717 ( .A0(n3957), .A1(n3245), .B0(n4270), .B1(n3209), .C0(n4114), .C1(n464), .Y(n5398) );
  OAI221XLTS U2718 ( .A0(n374), .A1(n281), .B0(n4770), .B1(n3411), .C0(n5438), 
        .Y(n2521) );
  OAI221XLTS U2719 ( .A0(n374), .A1(n272), .B0(n4780), .B1(n3410), .C0(n5439), 
        .Y(n2522) );
  AOI222XLTS U2720 ( .A0(n3969), .A1(n3371), .B0(n4282), .B1(n331), .C0(n4125), 
        .C1(n3403), .Y(n5439) );
  OAI221XLTS U2721 ( .A0(n375), .A1(n285), .B0(n4786), .B1(n3411), .C0(n5440), 
        .Y(n2523) );
  AOI222XLTS U2722 ( .A0(n3966), .A1(n3371), .B0(n4279), .B1(n303), .C0(n4122), 
        .C1(n3403), .Y(n5440) );
  OAI221XLTS U2723 ( .A0(n374), .A1(n276), .B0(n4796), .B1(n3411), .C0(n5441), 
        .Y(n2524) );
  AOI222XLTS U2724 ( .A0(n3963), .A1(n3371), .B0(n4276), .B1(n303), .C0(n4119), 
        .C1(n3403), .Y(n5441) );
  OAI221XLTS U2725 ( .A0(n375), .A1(n278), .B0(n4800), .B1(n3412), .C0(n5442), 
        .Y(n2525) );
  AOI222XLTS U2726 ( .A0(n3960), .A1(n3370), .B0(n4273), .B1(n331), .C0(n4116), 
        .C1(n3403), .Y(n5442) );
  OAI221XLTS U2727 ( .A0(n375), .A1(n288), .B0(n4810), .B1(n3412), .C0(n5443), 
        .Y(n2526) );
  AOI222XLTS U2728 ( .A0(n3957), .A1(n3369), .B0(n4270), .B1(n331), .C0(n4113), 
        .C1(n3404), .Y(n5443) );
  OAI221XLTS U2729 ( .A0(n374), .A1(n269), .B0(n4816), .B1(n3412), .C0(n5444), 
        .Y(n2527) );
  AOI222XLTS U2730 ( .A0(n3954), .A1(n3369), .B0(n4267), .B1(n303), .C0(n4110), 
        .C1(n3404), .Y(n5444) );
  OAI221XLTS U2731 ( .A0(n375), .A1(n267), .B0(n4822), .B1(n3411), .C0(n5445), 
        .Y(n2528) );
  AOI222XLTS U2732 ( .A0(n3951), .A1(n3369), .B0(n4264), .B1(n303), .C0(n4107), 
        .C1(n3405), .Y(n5445) );
  OAI221XLTS U2733 ( .A0(n3238), .A1(n6243), .B0(n4769), .B1(n3273), .C0(n5393), .Y(n2493) );
  AOI222XLTS U2734 ( .A0(n3972), .A1(n3244), .B0(n4285), .B1(n3211), .C0(n4129), .C1(n464), .Y(n5393) );
  OAI221XLTS U2735 ( .A0(n3239), .A1(n275), .B0(n4795), .B1(n3274), .C0(n5396), 
        .Y(n2496) );
  AOI222XLTS U2736 ( .A0(n3963), .A1(n3244), .B0(n4276), .B1(n3205), .C0(n4120), .C1(n464), .Y(n5396) );
  OAI221XLTS U2737 ( .A0(n3240), .A1(n270), .B0(n4819), .B1(n3275), .C0(n5399), 
        .Y(n2499) );
  AOI222XLTS U2738 ( .A0(n3954), .A1(n3245), .B0(n4267), .B1(n3212), .C0(n4111), .C1(n464), .Y(n5399) );
  OAI221XLTS U2739 ( .A0(n382), .A1(n282), .B0(n4771), .B1(n3345), .C0(n5415), 
        .Y(n2507) );
  AOI222XLTS U2740 ( .A0(n4284), .A1(n3292), .B0(n3973), .B1(n3295), .C0(n4129), .C1(n3339), .Y(n5415) );
  OAI221XLTS U2741 ( .A0(n382), .A1(n279), .B0(n4803), .B1(n3346), .C0(n5419), 
        .Y(n2511) );
  AOI222XLTS U2742 ( .A0(n4272), .A1(n3285), .B0(n3961), .B1(n3296), .C0(n4117), .C1(n3335), .Y(n5419) );
  OAI221XLTS U2743 ( .A0(n372), .A1(n6239), .B0(n4801), .B1(n3543), .C0(n5490), 
        .Y(n2553) );
  AOI222XLTS U2744 ( .A0(n3960), .A1(n3483), .B0(n4273), .B1(n3493), .C0(n4117), .C1(n3531), .Y(n5490) );
  OAI221XLTS U2745 ( .A0(n371), .A1(n6243), .B0(n4768), .B1(n3542), .C0(n5486), 
        .Y(n2549) );
  AOI222XLTS U2746 ( .A0(n3972), .A1(n3489), .B0(n4285), .B1(n3492), .C0(n4129), .C1(n3535), .Y(n5486) );
  OAI221XLTS U2747 ( .A0(n372), .A1(n6242), .B0(n4778), .B1(n3541), .C0(n5487), 
        .Y(n2550) );
  AOI222XLTS U2748 ( .A0(n3969), .A1(n3483), .B0(n4282), .B1(n3492), .C0(n4126), .C1(n3531), .Y(n5487) );
  OAI221XLTS U2749 ( .A0(n371), .A1(n6241), .B0(n4782), .B1(n3542), .C0(n5488), 
        .Y(n2551) );
  AOI222XLTS U2750 ( .A0(n3966), .A1(n3483), .B0(n4279), .B1(n3492), .C0(n4123), .C1(n3531), .Y(n5488) );
  OAI221XLTS U2751 ( .A0(n372), .A1(n6240), .B0(n4792), .B1(n3542), .C0(n5489), 
        .Y(n2552) );
  AOI222XLTS U2752 ( .A0(n3963), .A1(n3483), .B0(n4276), .B1(n3492), .C0(n4120), .C1(n3531), .Y(n5489) );
  OAI221XLTS U2753 ( .A0(n371), .A1(n6238), .B0(n4808), .B1(n3543), .C0(n5491), 
        .Y(n2554) );
  AOI222XLTS U2754 ( .A0(n3957), .A1(n3482), .B0(n4270), .B1(n3493), .C0(n4114), .C1(n3530), .Y(n5491) );
  OAI221XLTS U2755 ( .A0(n372), .A1(n6237), .B0(n4818), .B1(n3543), .C0(n5492), 
        .Y(n2555) );
  AOI222XLTS U2756 ( .A0(n3954), .A1(n3482), .B0(n4267), .B1(n3493), .C0(n4111), .C1(n3530), .Y(n5492) );
  OAI221XLTS U2757 ( .A0(n371), .A1(n6236), .B0(n4824), .B1(n3542), .C0(n5493), 
        .Y(n2556) );
  AOI222XLTS U2758 ( .A0(n3951), .A1(n3482), .B0(n4264), .B1(n3493), .C0(n4108), .C1(n3530), .Y(n5493) );
  AOI22X1TS U2759 ( .A0(n3278), .A1(n4235), .B0(n311), .B1(n4392), .Y(n6158)
         );
  AOI222XLTS U2760 ( .A0(n3326), .A1(n4080), .B0(n3318), .B1(n150), .C0(n3297), 
        .C1(n3924), .Y(n6157) );
  AOI22X1TS U2761 ( .A0(n3278), .A1(n4232), .B0(n315), .B1(n4389), .Y(n6160)
         );
  AOI222XLTS U2762 ( .A0(n3326), .A1(n4077), .B0(n3318), .B1(n145), .C0(n3297), 
        .C1(n3921), .Y(n6159) );
  AOI22X1TS U2763 ( .A0(n3278), .A1(n4229), .B0(n307), .B1(n4386), .Y(n6162)
         );
  AOI222XLTS U2764 ( .A0(n3326), .A1(n4074), .B0(n3318), .B1(n140), .C0(n3297), 
        .C1(n3918), .Y(n6161) );
  AOI22X1TS U2765 ( .A0(n3279), .A1(n4226), .B0(n310), .B1(n4383), .Y(n6168)
         );
  AOI222XLTS U2766 ( .A0(n3327), .A1(n4071), .B0(n3319), .B1(n135), .C0(n3298), 
        .C1(n3915), .Y(n6167) );
  AOI22X1TS U2767 ( .A0(n3279), .A1(n4241), .B0(n314), .B1(n4398), .Y(n6154)
         );
  AOI222XLTS U2768 ( .A0(n3327), .A1(n4086), .B0(n3319), .B1(n162), .C0(n3298), 
        .C1(n3930), .Y(n6153) );
  AOI22X1TS U2769 ( .A0(n3278), .A1(n4238), .B0(n306), .B1(n4395), .Y(n6156)
         );
  AOI222XLTS U2770 ( .A0(n3326), .A1(n4083), .B0(n3319), .B1(n155), .C0(n3298), 
        .C1(n3927), .Y(n6155) );
  AOI22X1TS U2771 ( .A0(n3362), .A1(n3929), .B0(n3726), .B1(n4398), .Y(n6170)
         );
  AOI222XLTS U2772 ( .A0(n3393), .A1(n4086), .B0(n3385), .B1(n161), .C0(n332), 
        .C1(n4242), .Y(n6169) );
  AOI22X1TS U2773 ( .A0(n3361), .A1(n3926), .B0(n3726), .B1(n4395), .Y(n6172)
         );
  AOI222XLTS U2774 ( .A0(n3392), .A1(n4083), .B0(n3385), .B1(n156), .C0(n333), 
        .C1(n4239), .Y(n6171) );
  AOI22X1TS U2775 ( .A0(n3361), .A1(n3923), .B0(n3725), .B1(n4392), .Y(n6174)
         );
  AOI222XLTS U2776 ( .A0(n3392), .A1(n4080), .B0(n3384), .B1(n151), .C0(n334), 
        .C1(n4236), .Y(n6173) );
  AOI22X1TS U2777 ( .A0(n3361), .A1(n3920), .B0(n3725), .B1(n4389), .Y(n6176)
         );
  AOI222XLTS U2778 ( .A0(n3392), .A1(n4077), .B0(n3384), .B1(n146), .C0(n304), 
        .C1(n4233), .Y(n6175) );
  AOI22X1TS U2779 ( .A0(n3361), .A1(n3917), .B0(n3725), .B1(n4386), .Y(n6178)
         );
  AOI222XLTS U2780 ( .A0(n3392), .A1(n4074), .B0(n3384), .B1(n141), .C0(n305), 
        .C1(n4230), .Y(n6177) );
  AOI22X1TS U2781 ( .A0(n3362), .A1(n3914), .B0(n3725), .B1(n4383), .Y(n6184)
         );
  AOI222XLTS U2782 ( .A0(n3393), .A1(n4071), .B0(n3385), .B1(n136), .C0(n247), 
        .C1(n4227), .Y(n6183) );
  AOI22X1TS U2783 ( .A0(n3215), .A1(readRequesterAddress[5]), .B0(n3197), .B1(
        n4241), .Y(n6139) );
  AOI222XLTS U2784 ( .A0(\requesterAddressbuffer[3][5] ), .A1(n3270), .B0(
        n6150), .B1(n3930), .C0(n3228), .C1(n4399), .Y(n6138) );
  AOI22X1TS U2785 ( .A0(n3215), .A1(readRequesterAddress[4]), .B0(n3196), .B1(
        n4238), .Y(n6141) );
  AOI222XLTS U2786 ( .A0(\requesterAddressbuffer[3][4] ), .A1(n3270), .B0(
        n3258), .B1(n3927), .C0(n3228), .C1(n4396), .Y(n6140) );
  AOI22X1TS U2787 ( .A0(n3215), .A1(readRequesterAddress[3]), .B0(n3196), .B1(
        n4235), .Y(n6143) );
  AOI222XLTS U2788 ( .A0(\requesterAddressbuffer[3][3] ), .A1(n3271), .B0(
        n3254), .B1(n3924), .C0(n3227), .C1(n4393), .Y(n6142) );
  AOI22X1TS U2789 ( .A0(n3214), .A1(readRequesterAddress[2]), .B0(n3196), .B1(
        n4232), .Y(n6145) );
  AOI222XLTS U2790 ( .A0(\requesterAddressbuffer[3][2] ), .A1(n3271), .B0(
        n3255), .B1(n3921), .C0(n3227), .C1(n4390), .Y(n6144) );
  AOI22X1TS U2791 ( .A0(n3213), .A1(readRequesterAddress[1]), .B0(n3196), .B1(
        n4229), .Y(n6147) );
  AOI222XLTS U2792 ( .A0(\requesterAddressbuffer[3][1] ), .A1(n3271), .B0(
        n3256), .B1(n3918), .C0(n3227), .C1(n4387), .Y(n6146) );
  AOI22X1TS U2793 ( .A0(n3215), .A1(n136), .B0(n3197), .B1(n4226), .Y(n6152)
         );
  AOI222XLTS U2794 ( .A0(\requesterAddressbuffer[3][0] ), .A1(n3271), .B0(
        n3258), .B1(n3915), .C0(n3227), .C1(n4384), .Y(n6151) );
  AOI22X1TS U2795 ( .A0(n753), .A1(n4085), .B0(n185), .B1(n4398), .Y(n6108) );
  AOI22X1TS U2796 ( .A0(n759), .A1(n4082), .B0(n186), .B1(n4395), .Y(n6110) );
  AOI222XLTS U2797 ( .A0(n793), .A1(n3926), .B0(n787), .B1(n157), .C0(n774), 
        .C1(n4239), .Y(n6109) );
  AOI22X1TS U2798 ( .A0(n760), .A1(n4079), .B0(n179), .B1(n4392), .Y(n6112) );
  AOI222XLTS U2799 ( .A0(n793), .A1(n3923), .B0(n787), .B1(n152), .C0(n763), 
        .C1(n4236), .Y(n6111) );
  AOI22X1TS U2800 ( .A0(n757), .A1(n4076), .B0(n181), .B1(n4389), .Y(n6114) );
  AOI222XLTS U2801 ( .A0(n793), .A1(n3920), .B0(n6119), .B1(n147), .C0(n763), 
        .C1(n4233), .Y(n6113) );
  AOI22X1TS U2802 ( .A0(n752), .A1(n4073), .B0(n179), .B1(n4386), .Y(n6116) );
  AOI222XLTS U2803 ( .A0(n793), .A1(n3917), .B0(n788), .B1(n142), .C0(n763), 
        .C1(n4230), .Y(n6115) );
  AOI22X1TS U2804 ( .A0(n6117), .A1(n4070), .B0(n180), .B1(n4383), .Y(n6122)
         );
  AOI222XLTS U2805 ( .A0(n794), .A1(n3914), .B0(n791), .B1(n137), .C0(n770), 
        .C1(n4227), .Y(n6121) );
  AOI222XLTS U2806 ( .A0(\requesterAddressbuffer[6][5] ), .A1(n691), .B0(n3467), .B1(n4241), .C0(n252), .C1(n4399), .Y(n6185) );
  AOI22X1TS U2807 ( .A0(n3445), .A1(n156), .B0(n3441), .B1(n4082), .Y(n6188)
         );
  AOI222XLTS U2808 ( .A0(\requesterAddressbuffer[6][4] ), .A1(n690), .B0(n3468), .B1(n4238), .C0(n252), .C1(n4396), .Y(n6187) );
  AOI22X1TS U2809 ( .A0(n3444), .A1(n146), .B0(n3439), .B1(n4076), .Y(n6192)
         );
  AOI222XLTS U2810 ( .A0(\requesterAddressbuffer[6][2] ), .A1(n693), .B0(n3468), .B1(n4232), .C0(n252), .C1(n4390), .Y(n6191) );
  AOI22X1TS U2811 ( .A0(n4259), .A1(n6163), .B0(n4417), .B1(n315), .Y(n5424)
         );
  AOI22X1TS U2812 ( .A0(n4253), .A1(n3291), .B0(n4411), .B1(n307), .Y(n5428)
         );
  AOI222XLTS U2813 ( .A0(n4097), .A1(n3336), .B0(n3320), .B1(n150), .C0(n3942), 
        .C1(n3306), .Y(n5427) );
  AOI22X1TS U2814 ( .A0(n4250), .A1(n3293), .B0(n4408), .B1(n311), .Y(n5430)
         );
  AOI222XLTS U2815 ( .A0(n4094), .A1(n3337), .B0(n3320), .B1(n145), .C0(n3939), 
        .C1(n3306), .Y(n5429) );
  AOI22X1TS U2816 ( .A0(n4247), .A1(n3290), .B0(n4405), .B1(n316), .Y(n5432)
         );
  AOI222XLTS U2817 ( .A0(n4091), .A1(n3340), .B0(n3320), .B1(n140), .C0(n3936), 
        .C1(n3305), .Y(n5431) );
  AOI22X1TS U2818 ( .A0(n4244), .A1(n3288), .B0(n4402), .B1(n308), .Y(n5434)
         );
  AOI222XLTS U2819 ( .A0(n4088), .A1(n3337), .B0(n3319), .B1(n135), .C0(n3933), 
        .C1(n3311), .Y(n5433) );
  AOI22X1TS U2820 ( .A0(n4220), .A1(n3287), .B0(n4377), .B1(n3739), .Y(n5776)
         );
  AOI222XLTS U2821 ( .A0(n4064), .A1(n3342), .B0(cacheDataOut[30]), .B1(n3324), 
        .C0(n3909), .C1(n3311), .Y(n5775) );
  AOI22X1TS U2822 ( .A0(n4214), .A1(n3289), .B0(n4371), .B1(n3739), .Y(n5780)
         );
  AOI222XLTS U2823 ( .A0(n4058), .A1(n3334), .B0(cacheDataOut[28]), .B1(n3324), 
        .C0(n3903), .C1(n3311), .Y(n5779) );
  AOI22X1TS U2824 ( .A0(n4211), .A1(n3290), .B0(n4368), .B1(n343), .Y(n5782)
         );
  AOI222XLTS U2825 ( .A0(n4055), .A1(n3334), .B0(cacheDataOut[27]), .B1(n3323), 
        .C0(n3900), .C1(n6164), .Y(n5781) );
  AOI22X1TS U2826 ( .A0(n4208), .A1(n3289), .B0(n4365), .B1(n312), .Y(n5784)
         );
  AOI222XLTS U2827 ( .A0(n4052), .A1(n3334), .B0(cacheDataOut[26]), .B1(n3313), 
        .C0(n3897), .C1(n3307), .Y(n5783) );
  AOI22X1TS U2828 ( .A0(n4205), .A1(n3288), .B0(n4362), .B1(n308), .Y(n5786)
         );
  AOI222XLTS U2829 ( .A0(n4049), .A1(n3333), .B0(cacheDataOut[25]), .B1(n3313), 
        .C0(n3894), .C1(n3309), .Y(n5785) );
  AOI22X1TS U2830 ( .A0(n4202), .A1(n3288), .B0(n4359), .B1(n343), .Y(n5788)
         );
  AOI222XLTS U2831 ( .A0(n4046), .A1(n3333), .B0(cacheDataOut[24]), .B1(n3312), 
        .C0(n3891), .C1(n3308), .Y(n5787) );
  AOI22X1TS U2832 ( .A0(n4199), .A1(n3287), .B0(n4356), .B1(n316), .Y(n5790)
         );
  AOI222XLTS U2833 ( .A0(n4043), .A1(n3333), .B0(cacheDataOut[23]), .B1(n3314), 
        .C0(n3888), .C1(n3304), .Y(n5789) );
  AOI22X1TS U2834 ( .A0(n4184), .A1(n3283), .B0(n4341), .B1(n314), .Y(n5800)
         );
  AOI222XLTS U2835 ( .A0(n4028), .A1(n3331), .B0(cacheDataOut[18]), .B1(n3313), 
        .C0(n3873), .C1(n3303), .Y(n5799) );
  AOI22X1TS U2836 ( .A0(n4169), .A1(n3282), .B0(n4326), .B1(n306), .Y(n5810)
         );
  AOI222XLTS U2837 ( .A0(n4013), .A1(n3330), .B0(cacheDataOut[13]), .B1(n3316), 
        .C0(n3858), .C1(n3302), .Y(n5809) );
  AOI22X1TS U2838 ( .A0(n4157), .A1(n3284), .B0(n4314), .B1(n315), .Y(n5818)
         );
  AOI222XLTS U2839 ( .A0(n4001), .A1(n3332), .B0(cacheDataOut[9]), .B1(n3316), 
        .C0(n3846), .C1(n3301), .Y(n5817) );
  AOI22X1TS U2840 ( .A0(n4151), .A1(n3281), .B0(n4308), .B1(n307), .Y(n5822)
         );
  AOI222XLTS U2841 ( .A0(n3995), .A1(n3329), .B0(cacheDataOut[7]), .B1(n3316), 
        .C0(n3840), .C1(n3300), .Y(n5821) );
  AOI22X1TS U2842 ( .A0(n4145), .A1(n3280), .B0(n4302), .B1(n310), .Y(n5826)
         );
  AOI222XLTS U2843 ( .A0(n3989), .A1(n3328), .B0(cacheDataOut[5]), .B1(n3323), 
        .C0(n3834), .C1(n3300), .Y(n5825) );
  AOI22X1TS U2844 ( .A0(n4142), .A1(n3280), .B0(n4299), .B1(n316), .Y(n5828)
         );
  AOI222XLTS U2845 ( .A0(n3986), .A1(n3328), .B0(cacheDataOut[4]), .B1(n3321), 
        .C0(n3831), .C1(n3300), .Y(n5827) );
  AOI22X1TS U2846 ( .A0(n4136), .A1(n3280), .B0(n4293), .B1(n308), .Y(n5832)
         );
  AOI222XLTS U2847 ( .A0(n3980), .A1(n3328), .B0(cacheDataOut[2]), .B1(n3322), 
        .C0(n3825), .C1(n3299), .Y(n5831) );
  AOI22X1TS U2848 ( .A0(n4223), .A1(n3287), .B0(n4380), .B1(n343), .Y(n5774)
         );
  AOI222XLTS U2849 ( .A0(n4067), .A1(n3338), .B0(cacheDataOut[31]), .B1(n3312), 
        .C0(n3912), .C1(n3309), .Y(n5773) );
  AOI22X1TS U2850 ( .A0(n4217), .A1(n3291), .B0(n4374), .B1(n344), .Y(n5778)
         );
  AOI222XLTS U2851 ( .A0(n4061), .A1(n3334), .B0(cacheDataOut[29]), .B1(n3312), 
        .C0(n3906), .C1(n3308), .Y(n5777) );
  AOI22X1TS U2852 ( .A0(n4196), .A1(n3287), .B0(n4353), .B1(n344), .Y(n5792)
         );
  AOI222XLTS U2853 ( .A0(n4040), .A1(n3333), .B0(cacheDataOut[22]), .B1(n3314), 
        .C0(n3885), .C1(n3304), .Y(n5791) );
  AOI22X1TS U2854 ( .A0(n4193), .A1(n3284), .B0(n4350), .B1(n306), .Y(n5794)
         );
  AOI222XLTS U2855 ( .A0(n4037), .A1(n3332), .B0(cacheDataOut[21]), .B1(n3312), 
        .C0(n3882), .C1(n3304), .Y(n5793) );
  AOI22X1TS U2856 ( .A0(n4190), .A1(n3284), .B0(n4347), .B1(n310), .Y(n5796)
         );
  AOI222XLTS U2857 ( .A0(n4034), .A1(n3332), .B0(cacheDataOut[20]), .B1(n3314), 
        .C0(n3879), .C1(n3304), .Y(n5795) );
  AOI22X1TS U2858 ( .A0(n4187), .A1(n3284), .B0(n4344), .B1(n344), .Y(n5798)
         );
  AOI222XLTS U2859 ( .A0(n4031), .A1(n3332), .B0(cacheDataOut[19]), .B1(n3315), 
        .C0(n3876), .C1(n3303), .Y(n5797) );
  AOI22X1TS U2860 ( .A0(n4178), .A1(n3283), .B0(n4335), .B1(n312), .Y(n5804)
         );
  AOI222XLTS U2861 ( .A0(n4022), .A1(n3331), .B0(cacheDataOut[16]), .B1(n3324), 
        .C0(n3867), .C1(n3303), .Y(n5803) );
  AOI22X1TS U2862 ( .A0(n4166), .A1(n3282), .B0(n4323), .B1(n310), .Y(n5812)
         );
  AOI222XLTS U2863 ( .A0(n4010), .A1(n3330), .B0(cacheDataOut[12]), .B1(n3315), 
        .C0(n3855), .C1(n3301), .Y(n5811) );
  AOI22X1TS U2864 ( .A0(n4163), .A1(n3282), .B0(n4320), .B1(n316), .Y(n5814)
         );
  AOI222XLTS U2865 ( .A0(n4007), .A1(n3330), .B0(cacheDataOut[11]), .B1(n3317), 
        .C0(n3852), .C1(n3301), .Y(n5813) );
  AOI22X1TS U2866 ( .A0(n4160), .A1(n3281), .B0(n4317), .B1(n308), .Y(n5816)
         );
  AOI222XLTS U2867 ( .A0(n4004), .A1(n3329), .B0(cacheDataOut[10]), .B1(n3317), 
        .C0(n3849), .C1(n3301), .Y(n5815) );
  AOI22X1TS U2868 ( .A0(n4154), .A1(n3281), .B0(n4311), .B1(n311), .Y(n5820)
         );
  AOI222XLTS U2869 ( .A0(n3998), .A1(n3329), .B0(cacheDataOut[8]), .B1(n3317), 
        .C0(n3843), .C1(n3300), .Y(n5819) );
  AOI22X1TS U2870 ( .A0(n4148), .A1(n3281), .B0(n4305), .B1(n314), .Y(n5824)
         );
  AOI222XLTS U2871 ( .A0(n3992), .A1(n3329), .B0(cacheDataOut[6]), .B1(n3316), 
        .C0(n3837), .C1(n3302), .Y(n5823) );
  AOI22X1TS U2872 ( .A0(n4133), .A1(n3279), .B0(n4290), .B1(n314), .Y(n5834)
         );
  AOI222XLTS U2873 ( .A0(n3977), .A1(n3327), .B0(cacheDataOut[1]), .B1(n3325), 
        .C0(n3822), .C1(n3299), .Y(n5833) );
  AOI22X1TS U2874 ( .A0(n4130), .A1(n3279), .B0(n4287), .B1(n306), .Y(n5836)
         );
  AOI222XLTS U2875 ( .A0(n3974), .A1(n3327), .B0(cacheDataOut[0]), .B1(n3315), 
        .C0(n3819), .C1(n3299), .Y(n5835) );
  AOI22X1TS U2876 ( .A0(n4181), .A1(n3283), .B0(n4338), .B1(n315), .Y(n5802)
         );
  AOI222XLTS U2877 ( .A0(n4025), .A1(n3331), .B0(cacheDataOut[17]), .B1(n3315), 
        .C0(n3870), .C1(n3303), .Y(n5801) );
  AOI22X1TS U2878 ( .A0(n4175), .A1(n3283), .B0(n4332), .B1(n307), .Y(n5806)
         );
  AOI222XLTS U2879 ( .A0(n4019), .A1(n3331), .B0(cacheDataOut[15]), .B1(n3314), 
        .C0(n3864), .C1(n3302), .Y(n5805) );
  AOI22X1TS U2880 ( .A0(n4172), .A1(n3282), .B0(n4329), .B1(n311), .Y(n5808)
         );
  AOI222XLTS U2881 ( .A0(n4016), .A1(n3330), .B0(cacheDataOut[14]), .B1(n3313), 
        .C0(n3861), .C1(n3302), .Y(n5807) );
  AOI22X1TS U2882 ( .A0(n4139), .A1(n3280), .B0(n4296), .B1(n312), .Y(n5830)
         );
  AOI222XLTS U2883 ( .A0(n3983), .A1(n3328), .B0(cacheDataOut[3]), .B1(n3317), 
        .C0(n3828), .C1(n3299), .Y(n5829) );
  AOI22X1TS U2884 ( .A0(n4055), .A1(n747), .B0(n4368), .B1(n176), .Y(n5974) );
  AOI22X1TS U2885 ( .A0(n4040), .A1(n746), .B0(n4353), .B1(n183), .Y(n5984) );
  AOI22X1TS U2886 ( .A0(n4034), .A1(n745), .B0(n4347), .B1(n178), .Y(n5988) );
  AOI22X1TS U2887 ( .A0(n4031), .A1(n745), .B0(n4344), .B1(n184), .Y(n5990) );
  AOI22X1TS U2888 ( .A0(n4004), .A1(n743), .B0(n4317), .B1(n185), .Y(n6008) );
  AOI22X1TS U2889 ( .A0(n3998), .A1(n743), .B0(n4311), .B1(n183), .Y(n6012) );
  AOI22X1TS U2890 ( .A0(n3989), .A1(n755), .B0(n4302), .B1(n180), .Y(n6018) );
  AOI22X1TS U2891 ( .A0(n3980), .A1(n755), .B0(n4293), .B1(n177), .Y(n6024) );
  AOI22X1TS U2892 ( .A0(n4256), .A1(n3286), .B0(n4414), .B1(n312), .Y(n5426)
         );
  AOI222XLTS U2893 ( .A0(n4100), .A1(n3340), .B0(n3320), .B1(
        readRequesterAddress[4]), .C0(n3945), .C1(n3311), .Y(n5425) );
  AOI22X1TS U2894 ( .A0(n3911), .A1(n3373), .B0(n4380), .B1(n3737), .Y(n5710)
         );
  AOI22X1TS U2895 ( .A0(n3866), .A1(n3366), .B0(n4335), .B1(n3730), .Y(n5740)
         );
  AOI22X1TS U2896 ( .A0(n3863), .A1(n3366), .B0(n4332), .B1(n3730), .Y(n5742)
         );
  AOI22X1TS U2897 ( .A0(n3851), .A1(n3365), .B0(n4320), .B1(n3729), .Y(n5750)
         );
  AOI22X1TS U2898 ( .A0(n3821), .A1(n3362), .B0(n4290), .B1(n3726), .Y(n5770)
         );
  AOI22X1TS U2899 ( .A0(n4259), .A1(n3471), .B0(n4416), .B1(n317), .Y(n5471)
         );
  AOI222XLTS U2900 ( .A0(n3947), .A1(n3722), .B0(n3452), .B1(n130), .C0(n4104), 
        .C1(n3427), .Y(n5470) );
  AOI22X1TS U2901 ( .A0(n4253), .A1(n3465), .B0(n4410), .B1(n317), .Y(n5475)
         );
  AOI222XLTS U2902 ( .A0(n3941), .A1(n3718), .B0(n3452), .B1(
        readRequesterAddress[3]), .C0(n4098), .C1(n3436), .Y(n5474) );
  AOI22X1TS U2903 ( .A0(n4250), .A1(n3464), .B0(n4407), .B1(n317), .Y(n5477)
         );
  AOI222XLTS U2904 ( .A0(n3938), .A1(n3721), .B0(n3452), .B1(
        readRequesterAddress[2]), .C0(n4095), .C1(n3436), .Y(n5476) );
  AOI22X1TS U2905 ( .A0(n4247), .A1(n3464), .B0(n4404), .B1(n329), .Y(n5479)
         );
  AOI222XLTS U2906 ( .A0(n3935), .A1(n3720), .B0(n3451), .B1(
        readRequesterAddress[1]), .C0(n4092), .C1(n3436), .Y(n5478) );
  AOI22X1TS U2907 ( .A0(n4244), .A1(n3464), .B0(n4401), .B1(n317), .Y(n5481)
         );
  AOI222XLTS U2908 ( .A0(n3932), .A1(n3723), .B0(n3451), .B1(
        readRequesterAddress[0]), .C0(n4089), .C1(n3436), .Y(n5480) );
  AOI22X1TS U2909 ( .A0(n4217), .A1(n3470), .B0(n4374), .B1(n6344), .Y(n5650)
         );
  AOI22X1TS U2910 ( .A0(n4199), .A1(n3463), .B0(n4356), .B1(n240), .Y(n5662)
         );
  AOI22X1TS U2911 ( .A0(n4193), .A1(n3463), .B0(n4350), .B1(n241), .Y(n5666)
         );
  AOI22X1TS U2912 ( .A0(n4190), .A1(n3463), .B0(n4347), .B1(n241), .Y(n5668)
         );
  AOI22X1TS U2913 ( .A0(n4169), .A1(n3461), .B0(n4326), .B1(n328), .Y(n5682)
         );
  AOI22X1TS U2914 ( .A0(n4166), .A1(n3461), .B0(n4323), .B1(n327), .Y(n5684)
         );
  AOI22X1TS U2915 ( .A0(n4160), .A1(n3460), .B0(n4317), .B1(n319), .Y(n5688)
         );
  AOI22X1TS U2916 ( .A0(n4148), .A1(n3459), .B0(n4305), .B1(n328), .Y(n5696)
         );
  AOI22X1TS U2917 ( .A0(n3944), .A1(n3481), .B0(n4413), .B1(n3696), .Y(n5499)
         );
  AOI222XLTS U2918 ( .A0(n4101), .A1(n3529), .B0(n155), .B1(n3517), .C0(n4257), 
        .C1(n3501), .Y(n5498) );
  AOI22X1TS U2919 ( .A0(n3932), .A1(n3491), .B0(n4401), .B1(n3697), .Y(n5507)
         );
  AOI222XLTS U2920 ( .A0(n4089), .A1(n3528), .B0(n138), .B1(n3509), .C0(n4245), 
        .C1(n3500), .Y(n5506) );
  AOI22X1TS U2921 ( .A0(n4103), .A1(n749), .B0(n4416), .B1(n380), .Y(n5355) );
  OAI211X1TS U2922 ( .A0(n4722), .A1(n823), .B0(n5357), .C0(n5356), .Y(n2474)
         );
  INVX2TS U2923 ( .A(n827), .Y(n823) );
  AOI22X1TS U2924 ( .A0(n4100), .A1(n749), .B0(n4413), .B1(n380), .Y(n5357) );
  AOI222XLTS U2925 ( .A0(n3945), .A1(n801), .B0(n6119), .B1(n155), .C0(n4257), 
        .C1(n775), .Y(n5356) );
  AOI22X1TS U2926 ( .A0(n4097), .A1(n749), .B0(n4410), .B1(n183), .Y(n5359) );
  AOI222XLTS U2927 ( .A0(n3942), .A1(n801), .B0(n790), .B1(n152), .C0(n4254), 
        .C1(n777), .Y(n5358) );
  AOI22X1TS U2928 ( .A0(n4094), .A1(n749), .B0(n4407), .B1(n175), .Y(n5361) );
  AOI222XLTS U2929 ( .A0(n3939), .A1(n801), .B0(n789), .B1(n147), .C0(n4251), 
        .C1(n770), .Y(n5360) );
  AOI22X1TS U2930 ( .A0(n4091), .A1(n748), .B0(n4404), .B1(n175), .Y(n5363) );
  AOI222XLTS U2931 ( .A0(n3936), .A1(n807), .B0(n788), .B1(n142), .C0(n4248), 
        .C1(n770), .Y(n5362) );
  AOI22X1TS U2932 ( .A0(n4088), .A1(n748), .B0(n4401), .B1(n184), .Y(n5365) );
  AOI222XLTS U2933 ( .A0(n3933), .A1(n809), .B0(n791), .B1(n137), .C0(n4245), 
        .C1(n777), .Y(n5364) );
  AOI22X1TS U2934 ( .A0(n4067), .A1(n748), .B0(n4380), .B1(n175), .Y(n5966) );
  AOI22X1TS U2935 ( .A0(n4064), .A1(n748), .B0(n4377), .B1(n176), .Y(n5968) );
  AOI22X1TS U2936 ( .A0(n4061), .A1(n747), .B0(n4374), .B1(n181), .Y(n5970) );
  AOI22X1TS U2937 ( .A0(n4058), .A1(n747), .B0(n4371), .B1(n3768), .Y(n5972)
         );
  AOI22X1TS U2938 ( .A0(n4052), .A1(n747), .B0(n4365), .B1(n183), .Y(n5976) );
  AOI22X1TS U2939 ( .A0(n4049), .A1(n746), .B0(n4362), .B1(n186), .Y(n5978) );
  AOI22X1TS U2940 ( .A0(n4046), .A1(n746), .B0(n4359), .B1(n176), .Y(n5980) );
  AOI22X1TS U2941 ( .A0(n4043), .A1(n746), .B0(n4356), .B1(n175), .Y(n5982) );
  AOI22X1TS U2942 ( .A0(n4037), .A1(n745), .B0(n4350), .B1(n176), .Y(n5986) );
  AOI22X1TS U2943 ( .A0(n4028), .A1(n757), .B0(n4341), .B1(n180), .Y(n5992) );
  AOI22X1TS U2944 ( .A0(n4025), .A1(n753), .B0(n4338), .B1(n184), .Y(n5994) );
  AOI22X1TS U2945 ( .A0(n4022), .A1(n756), .B0(n4335), .B1(n177), .Y(n5996) );
  AOI22X1TS U2946 ( .A0(n4019), .A1(n756), .B0(n4332), .B1(n178), .Y(n5998) );
  AOI22X1TS U2947 ( .A0(n4016), .A1(n754), .B0(n4329), .B1(n3768), .Y(n6000)
         );
  AOI22X1TS U2948 ( .A0(n4013), .A1(n757), .B0(n4326), .B1(n178), .Y(n6002) );
  AOI22X1TS U2949 ( .A0(n4010), .A1(n756), .B0(n4323), .B1(n185), .Y(n6004) );
  AOI22X1TS U2950 ( .A0(n4007), .A1(n756), .B0(n4320), .B1(n181), .Y(n6006) );
  AOI22X1TS U2951 ( .A0(n4001), .A1(n745), .B0(n4314), .B1(n177), .Y(n6010) );
  AOI22X1TS U2952 ( .A0(n3995), .A1(n743), .B0(n4308), .B1(n184), .Y(n6014) );
  AOI22X1TS U2953 ( .A0(n3992), .A1(n743), .B0(n4305), .B1(n185), .Y(n6016) );
  AOI22X1TS U2954 ( .A0(n3986), .A1(n760), .B0(n4299), .B1(n178), .Y(n6020) );
  AOI22X1TS U2955 ( .A0(n3983), .A1(n754), .B0(n4296), .B1(n180), .Y(n6022) );
  AOI22X1TS U2956 ( .A0(n3977), .A1(n760), .B0(n4290), .B1(n177), .Y(n6026) );
  AOI22X1TS U2957 ( .A0(n3947), .A1(n3368), .B0(n4416), .B1(n3735), .Y(n5448)
         );
  AOI222XLTS U2958 ( .A0(n4103), .A1(n3402), .B0(n3384), .B1(n130), .C0(n4260), 
        .C1(n333), .Y(n5447) );
  AOI22X1TS U2959 ( .A0(n3944), .A1(n3368), .B0(n4413), .B1(n3734), .Y(n5450)
         );
  AOI222XLTS U2960 ( .A0(n4100), .A1(n3402), .B0(n3386), .B1(n157), .C0(n4257), 
        .C1(n305), .Y(n5449) );
  AOI22X1TS U2961 ( .A0(n3941), .A1(n3368), .B0(n4410), .B1(n3737), .Y(n5452)
         );
  AOI222XLTS U2962 ( .A0(n4097), .A1(n3402), .B0(n3386), .B1(n153), .C0(n4254), 
        .C1(n304), .Y(n5451) );
  AOI22X1TS U2963 ( .A0(n3938), .A1(n3368), .B0(n4407), .B1(n3735), .Y(n5454)
         );
  AOI222XLTS U2964 ( .A0(n4094), .A1(n3402), .B0(n3386), .B1(n148), .C0(n4251), 
        .C1(n304), .Y(n5453) );
  AOI22X1TS U2965 ( .A0(n3935), .A1(n3377), .B0(n4404), .B1(n3737), .Y(n5456)
         );
  AOI222XLTS U2966 ( .A0(n4091), .A1(n3401), .B0(n3386), .B1(n143), .C0(n4248), 
        .C1(n334), .Y(n5455) );
  AOI22X1TS U2967 ( .A0(n3932), .A1(n6179), .B0(n4401), .B1(n6345), .Y(n5458)
         );
  AOI222XLTS U2968 ( .A0(n4088), .A1(n3401), .B0(n3385), .B1(n138), .C0(n4245), 
        .C1(n332), .Y(n5457) );
  AOI22X1TS U2969 ( .A0(n3908), .A1(n3371), .B0(n4377), .B1(n3736), .Y(n5712)
         );
  AOI22X1TS U2970 ( .A0(n3905), .A1(n3374), .B0(n4374), .B1(n3733), .Y(n5714)
         );
  AOI22X1TS U2971 ( .A0(n3902), .A1(n3375), .B0(n4371), .B1(n3733), .Y(n5716)
         );
  AOI22X1TS U2972 ( .A0(n3899), .A1(n3374), .B0(n4368), .B1(n3733), .Y(n5718)
         );
  AOI22X1TS U2973 ( .A0(n3896), .A1(n3375), .B0(n4365), .B1(n3733), .Y(n5720)
         );
  AOI22X1TS U2974 ( .A0(n3893), .A1(n3372), .B0(n4362), .B1(n3732), .Y(n5722)
         );
  AOI22X1TS U2975 ( .A0(n3890), .A1(n3372), .B0(n4359), .B1(n3732), .Y(n5724)
         );
  AOI22X1TS U2976 ( .A0(n3887), .A1(n3372), .B0(n4356), .B1(n3732), .Y(n5726)
         );
  AOI22X1TS U2977 ( .A0(n3884), .A1(n3373), .B0(n4353), .B1(n3732), .Y(n5728)
         );
  AOI22X1TS U2978 ( .A0(n3881), .A1(n3367), .B0(n4350), .B1(n3731), .Y(n5730)
         );
  AOI22X1TS U2979 ( .A0(n3878), .A1(n3367), .B0(n4347), .B1(n3731), .Y(n5732)
         );
  AOI22X1TS U2980 ( .A0(n3875), .A1(n3367), .B0(n4344), .B1(n3731), .Y(n5734)
         );
  AOI22X1TS U2981 ( .A0(n3872), .A1(n3366), .B0(n4341), .B1(n3731), .Y(n5736)
         );
  AOI22X1TS U2982 ( .A0(n3869), .A1(n3366), .B0(n4338), .B1(n3730), .Y(n5738)
         );
  AOI22X1TS U2983 ( .A0(n3860), .A1(n3365), .B0(n4329), .B1(n3730), .Y(n5744)
         );
  AOI22X1TS U2984 ( .A0(n3857), .A1(n3365), .B0(n4326), .B1(n3729), .Y(n5746)
         );
  AOI22X1TS U2985 ( .A0(n3854), .A1(n3365), .B0(n4323), .B1(n3729), .Y(n5748)
         );
  AOI22X1TS U2986 ( .A0(n3848), .A1(n3364), .B0(n4317), .B1(n3729), .Y(n5752)
         );
  AOI22X1TS U2987 ( .A0(n3845), .A1(n3367), .B0(n4314), .B1(n3728), .Y(n5754)
         );
  AOI22X1TS U2988 ( .A0(n3842), .A1(n3364), .B0(n4311), .B1(n3728), .Y(n5756)
         );
  AOI22X1TS U2989 ( .A0(n3839), .A1(n3364), .B0(n4308), .B1(n3728), .Y(n5758)
         );
  AOI22X1TS U2990 ( .A0(n3836), .A1(n3364), .B0(n4305), .B1(n3728), .Y(n5760)
         );
  AOI22X1TS U2991 ( .A0(n3833), .A1(n3363), .B0(n4302), .B1(n3727), .Y(n5762)
         );
  AOI22X1TS U2992 ( .A0(n3830), .A1(n3363), .B0(n4299), .B1(n3727), .Y(n5764)
         );
  AOI22X1TS U2993 ( .A0(n3827), .A1(n3363), .B0(n4296), .B1(n3727), .Y(n5766)
         );
  AOI22X1TS U2994 ( .A0(n3824), .A1(n3363), .B0(n4293), .B1(n3727), .Y(n5768)
         );
  AOI22X1TS U2995 ( .A0(n3818), .A1(n3362), .B0(n4287), .B1(n3726), .Y(n5772)
         );
  AOI22X1TS U2996 ( .A0(n4223), .A1(n3464), .B0(n4380), .B1(n241), .Y(n5646)
         );
  AOI22X1TS U2997 ( .A0(n4220), .A1(n3470), .B0(n4377), .B1(n319), .Y(n5648)
         );
  AOI22X1TS U2998 ( .A0(n4214), .A1(n3473), .B0(n4371), .B1(n318), .Y(n5652)
         );
  AOI22X1TS U2999 ( .A0(n4211), .A1(n3473), .B0(n4368), .B1(n319), .Y(n5654)
         );
  AOI22X1TS U3000 ( .A0(n4208), .A1(n3472), .B0(n4365), .B1(n6344), .Y(n5656)
         );
  AOI22X1TS U3001 ( .A0(n4202), .A1(n3472), .B0(n4359), .B1(n240), .Y(n5660)
         );
  AOI22X1TS U3002 ( .A0(n4196), .A1(n3463), .B0(n4353), .B1(n240), .Y(n5664)
         );
  AOI22X1TS U3003 ( .A0(n4187), .A1(n3462), .B0(n4344), .B1(n240), .Y(n5670)
         );
  AOI22X1TS U3004 ( .A0(n4181), .A1(n3462), .B0(n4338), .B1(n325), .Y(n5674)
         );
  AOI22X1TS U3005 ( .A0(n4178), .A1(n3462), .B0(n4335), .B1(n325), .Y(n5676)
         );
  AOI22X1TS U3006 ( .A0(n4175), .A1(n3461), .B0(n4332), .B1(n325), .Y(n5678)
         );
  AOI22X1TS U3007 ( .A0(n4172), .A1(n3461), .B0(n4329), .B1(n318), .Y(n5680)
         );
  AOI22X1TS U3008 ( .A0(n4163), .A1(n3460), .B0(n4320), .B1(n326), .Y(n5686)
         );
  AOI22X1TS U3009 ( .A0(n4157), .A1(n3460), .B0(n4314), .B1(n318), .Y(n5690)
         );
  AOI22X1TS U3010 ( .A0(n4154), .A1(n3460), .B0(n4311), .B1(n327), .Y(n5692)
         );
  AOI22X1TS U3011 ( .A0(n4151), .A1(n3459), .B0(n4308), .B1(n326), .Y(n5694)
         );
  AOI22X1TS U3012 ( .A0(n4145), .A1(n3459), .B0(n4302), .B1(n328), .Y(n5698)
         );
  AOI22X1TS U3013 ( .A0(n4139), .A1(n3458), .B0(n4296), .B1(n327), .Y(n5702)
         );
  AOI22X1TS U3014 ( .A0(n4136), .A1(n3458), .B0(n4293), .B1(n326), .Y(n5704)
         );
  AOI22X1TS U3015 ( .A0(n3947), .A1(n3481), .B0(n4416), .B1(n3696), .Y(n5497)
         );
  AOI222XLTS U3016 ( .A0(n4104), .A1(n3529), .B0(n161), .B1(n3517), .C0(n4260), 
        .C1(n3494), .Y(n5496) );
  AOI22X1TS U3017 ( .A0(n3941), .A1(n3481), .B0(n4410), .B1(n3696), .Y(n5501)
         );
  AOI222XLTS U3018 ( .A0(n4098), .A1(n3529), .B0(n153), .B1(n3519), .C0(n4254), 
        .C1(n3500), .Y(n5500) );
  AOI22X1TS U3019 ( .A0(n3938), .A1(n3481), .B0(n4407), .B1(n3696), .Y(n5503)
         );
  AOI222XLTS U3020 ( .A0(n4095), .A1(n3529), .B0(n148), .B1(n3519), .C0(n4251), 
        .C1(n3500), .Y(n5502) );
  AOI22X1TS U3021 ( .A0(n3935), .A1(n3488), .B0(n4404), .B1(n3697), .Y(n5505)
         );
  AOI222XLTS U3022 ( .A0(n4092), .A1(n3528), .B0(n143), .B1(n3509), .C0(n4248), 
        .C1(n3500), .Y(n5504) );
  AOI22X1TS U3023 ( .A0(n3911), .A1(n3491), .B0(n4381), .B1(n3697), .Y(n5582)
         );
  AOI22X1TS U3024 ( .A0(n3908), .A1(n3491), .B0(n4378), .B1(n3697), .Y(n5584)
         );
  AOI22X1TS U3025 ( .A0(n3905), .A1(n3484), .B0(n4375), .B1(n3698), .Y(n5586)
         );
  AOI22X1TS U3026 ( .A0(n3902), .A1(n3485), .B0(n4372), .B1(n3698), .Y(n5588)
         );
  AOI22X1TS U3027 ( .A0(n3899), .A1(n3487), .B0(n4369), .B1(n3698), .Y(n5590)
         );
  AOI22X1TS U3028 ( .A0(n3896), .A1(n3486), .B0(n4366), .B1(n3698), .Y(n5592)
         );
  AOI22X1TS U3029 ( .A0(n3893), .A1(n3490), .B0(n4363), .B1(n3707), .Y(n5594)
         );
  AOI22X1TS U3030 ( .A0(n3890), .A1(n3487), .B0(n4360), .B1(n3706), .Y(n5596)
         );
  AOI22X1TS U3031 ( .A0(n3887), .A1(n3486), .B0(n4357), .B1(n6342), .Y(n5598)
         );
  AOI22X1TS U3032 ( .A0(n3884), .A1(n3488), .B0(n4354), .B1(n3709), .Y(n5600)
         );
  AOI22X1TS U3033 ( .A0(n3881), .A1(n6211), .B0(n4351), .B1(n3707), .Y(n5602)
         );
  AOI22X1TS U3034 ( .A0(n3878), .A1(n3490), .B0(n4348), .B1(n3708), .Y(n5604)
         );
  AOI22X1TS U3035 ( .A0(n3875), .A1(n3490), .B0(n4345), .B1(n3707), .Y(n5606)
         );
  AOI22X1TS U3036 ( .A0(n3872), .A1(n3480), .B0(n4342), .B1(n3708), .Y(n5608)
         );
  AOI22X1TS U3037 ( .A0(n3869), .A1(n3480), .B0(n4339), .B1(n3699), .Y(n5610)
         );
  AOI22X1TS U3038 ( .A0(n3866), .A1(n3480), .B0(n4336), .B1(n3699), .Y(n5612)
         );
  AOI22X1TS U3039 ( .A0(n3863), .A1(n3480), .B0(n4333), .B1(n3699), .Y(n5614)
         );
  AOI22X1TS U3040 ( .A0(n3860), .A1(n3479), .B0(n4330), .B1(n3699), .Y(n5616)
         );
  AOI22X1TS U3041 ( .A0(n3857), .A1(n3479), .B0(n4327), .B1(n3700), .Y(n5618)
         );
  AOI22X1TS U3042 ( .A0(n3854), .A1(n3479), .B0(n4324), .B1(n3700), .Y(n5620)
         );
  AOI22X1TS U3043 ( .A0(n3851), .A1(n3479), .B0(n4321), .B1(n3700), .Y(n5622)
         );
  AOI22X1TS U3044 ( .A0(n3848), .A1(n3478), .B0(n4318), .B1(n3700), .Y(n5624)
         );
  AOI22X1TS U3045 ( .A0(n3845), .A1(n3478), .B0(n4315), .B1(n3701), .Y(n5626)
         );
  AOI22X1TS U3046 ( .A0(n3842), .A1(n3478), .B0(n4312), .B1(n3701), .Y(n5628)
         );
  AOI22X1TS U3047 ( .A0(n3839), .A1(n3478), .B0(n4309), .B1(n3701), .Y(n5630)
         );
  AOI22X1TS U3048 ( .A0(n3836), .A1(n3477), .B0(n4306), .B1(n3701), .Y(n5632)
         );
  AOI22X1TS U3049 ( .A0(n3833), .A1(n3477), .B0(n4303), .B1(n3702), .Y(n5634)
         );
  AOI22X1TS U3050 ( .A0(n3830), .A1(n3477), .B0(n4300), .B1(n3702), .Y(n5636)
         );
  AOI22X1TS U3051 ( .A0(n3827), .A1(n3477), .B0(n4297), .B1(n3702), .Y(n5638)
         );
  AOI22X1TS U3052 ( .A0(n3824), .A1(n3476), .B0(n4294), .B1(n3702), .Y(n5640)
         );
  AOI22X1TS U3053 ( .A0(n3821), .A1(n3476), .B0(n4291), .B1(n3703), .Y(n5642)
         );
  AOI22X1TS U3054 ( .A0(n3818), .A1(n3476), .B0(n4288), .B1(n3703), .Y(n5644)
         );
  AOI22X1TS U3055 ( .A0(n3974), .A1(n757), .B0(n4287), .B1(n179), .Y(n6028) );
  AOI22X1TS U3056 ( .A0(n4256), .A1(n3465), .B0(n4413), .B1(n318), .Y(n5473)
         );
  AOI222XLTS U3057 ( .A0(n3944), .A1(n3721), .B0(n3452), .B1(n158), .C0(n4101), 
        .C1(n3441), .Y(n5472) );
  AOI22X1TS U3058 ( .A0(n4205), .A1(n3471), .B0(n4362), .B1(n241), .Y(n5658)
         );
  AOI22X1TS U3059 ( .A0(n4184), .A1(n3462), .B0(n4341), .B1(n319), .Y(n5672)
         );
  AOI22X1TS U3060 ( .A0(n4142), .A1(n3459), .B0(n4299), .B1(n325), .Y(n5700)
         );
  AOI22X1TS U3061 ( .A0(n6134), .A1(n142), .B0(n829), .B1(n4073), .Y(n6132) );
  AOI222XLTS U3062 ( .A0(\requesterAddressbuffer[2][1] ), .A1(n299), .B0(n957), 
        .B1(n4230), .C0(n3754), .C1(n4387), .Y(n6131) );
  AOI22X1TS U3063 ( .A0(n857), .A1(n137), .B0(n830), .B1(n4070), .Y(n6137) );
  AOI222XLTS U3064 ( .A0(\requesterAddressbuffer[2][0] ), .A1(n297), .B0(n957), 
        .B1(n4227), .C0(n3754), .C1(n4384), .Y(n6136) );
  AOI22X1TS U3065 ( .A0(n856), .A1(n152), .B0(n829), .B1(n4079), .Y(n6128) );
  AOI222XLTS U3066 ( .A0(\requesterAddressbuffer[2][3] ), .A1(n298), .B0(n957), 
        .B1(n4236), .C0(n3754), .C1(n4393), .Y(n6127) );
  AOI22X1TS U3067 ( .A0(n858), .A1(n147), .B0(n829), .B1(n4076), .Y(n6130) );
  AOI222XLTS U3068 ( .A0(\requesterAddressbuffer[2][2] ), .A1(n297), .B0(n871), 
        .B1(n4233), .C0(n3754), .C1(n4390), .Y(n6129) );
  AOI22X1TS U3069 ( .A0(n857), .A1(n157), .B0(n829), .B1(n4082), .Y(n6126) );
  AOI222XLTS U3070 ( .A0(\requesterAddressbuffer[2][4] ), .A1(n299), .B0(n870), 
        .B1(n4239), .C0(n3755), .C1(n4396), .Y(n6125) );
  AOI22X1TS U3071 ( .A0(n855), .A1(n160), .B0(n830), .B1(n4085), .Y(n6124) );
  AOI222XLTS U3072 ( .A0(\requesterAddressbuffer[2][5] ), .A1(n298), .B0(n936), 
        .B1(n4242), .C0(n3755), .C1(n4399), .Y(n6123) );
  AOI22X1TS U3073 ( .A0(n3444), .A1(n151), .B0(n3437), .B1(n4079), .Y(n6190)
         );
  AOI222XLTS U3074 ( .A0(\requesterAddressbuffer[6][3] ), .A1(n692), .B0(n3468), .B1(n4235), .C0(n6344), .C1(n4393), .Y(n6189) );
  AOI22X1TS U3075 ( .A0(n3444), .A1(n141), .B0(n3438), .B1(n4073), .Y(n6194)
         );
  AOI222XLTS U3076 ( .A0(\requesterAddressbuffer[6][1] ), .A1(n692), .B0(n3468), .B1(n4229), .C0(n6344), .C1(n4387), .Y(n6193) );
  AOI222XLTS U3077 ( .A0(\requesterAddressbuffer[6][0] ), .A1(n692), .B0(n3474), .B1(n4226), .C0(n252), .C1(n4384), .Y(n6198) );
  AOI22X1TS U3078 ( .A0(n740), .A1(n130), .B0(n697), .B1(n4241), .Y(n6094) );
  AOI222XLTS U3079 ( .A0(\requesterAddressbuffer[0][5] ), .A1(n230), .B0(n118), 
        .B1(n3930), .C0(n3793), .C1(n4399), .Y(n6093) );
  AOI22X1TS U3080 ( .A0(n739), .A1(n151), .B0(n696), .B1(n4235), .Y(n6098) );
  AOI222XLTS U3081 ( .A0(\requesterAddressbuffer[0][3] ), .A1(n337), .B0(n117), 
        .B1(n3924), .C0(n3795), .C1(n4393), .Y(n6097) );
  AOI22X1TS U3082 ( .A0(n740), .A1(n156), .B0(n696), .B1(n4238), .Y(n6096) );
  AOI222XLTS U3083 ( .A0(\requesterAddressbuffer[0][4] ), .A1(n229), .B0(n124), 
        .B1(n3927), .C0(n3794), .C1(n4396), .Y(n6095) );
  AOI22X1TS U3084 ( .A0(n741), .A1(n146), .B0(n696), .B1(n4232), .Y(n6100) );
  AOI222XLTS U3085 ( .A0(\requesterAddressbuffer[0][2] ), .A1(n228), .B0(n114), 
        .B1(n3921), .C0(n254), .C1(n4390), .Y(n6099) );
  AOI22X1TS U3086 ( .A0(n6104), .A1(n141), .B0(n696), .B1(n4229), .Y(n6102) );
  AOI222XLTS U3087 ( .A0(\requesterAddressbuffer[0][1] ), .A1(n230), .B0(n113), 
        .B1(n3918), .C0(n254), .C1(n4387), .Y(n6101) );
  AOI22X1TS U3088 ( .A0(n736), .A1(n138), .B0(n697), .B1(n4226), .Y(n6106) );
  AOI222XLTS U3089 ( .A0(\requesterAddressbuffer[0][0] ), .A1(n337), .B0(n123), 
        .B1(n3915), .C0(n3797), .C1(n4384), .Y(n6105) );
  AOI22X1TS U3090 ( .A0(n740), .A1(n160), .B0(n4259), .B1(n708), .Y(n5332) );
  AOI222XLTS U3091 ( .A0(n209), .A1(n20), .B0(n3948), .B1(n123), .C0(n4417), 
        .C1(n3791), .Y(n5331) );
  AOI22X1TS U3092 ( .A0(n716), .A1(n153), .B0(n4253), .B1(n711), .Y(n5336) );
  AOI222XLTS U3093 ( .A0(n230), .A1(n21), .B0(n3942), .B1(n112), .C0(n4411), 
        .C1(n3791), .Y(n5335) );
  AOI22X1TS U3094 ( .A0(n716), .A1(n148), .B0(n4250), .B1(n712), .Y(n5338) );
  AOI222XLTS U3095 ( .A0(n337), .A1(n22), .B0(n3939), .B1(n112), .C0(n4408), 
        .C1(n3791), .Y(n5337) );
  AOI22X1TS U3096 ( .A0(n736), .A1(n143), .B0(n4247), .B1(n707), .Y(n5340) );
  AOI222XLTS U3097 ( .A0(n208), .A1(n23), .B0(n3936), .B1(n113), .C0(n4405), 
        .C1(n3790), .Y(n5339) );
  AOI22X1TS U3098 ( .A0(n397), .A1(n735), .B0(n4223), .B1(n707), .Y(n6030) );
  AOI222XLTS U3099 ( .A0(n338), .A1(n24), .B0(n3912), .B1(n121), .C0(n4381), 
        .C1(n3790), .Y(n6029) );
  AOI22X1TS U3100 ( .A0(n399), .A1(n739), .B0(n4220), .B1(n708), .Y(n6032) );
  AOI222XLTS U3101 ( .A0(n208), .A1(n25), .B0(n3909), .B1(n118), .C0(n4378), 
        .C1(n3790), .Y(n6031) );
  AOI22X1TS U3102 ( .A0(n401), .A1(n739), .B0(n4217), .B1(n704), .Y(n6034) );
  AOI222XLTS U3103 ( .A0(n208), .A1(n26), .B0(n3906), .B1(n116), .C0(n4375), 
        .C1(n3789), .Y(n6033) );
  AOI22X1TS U3104 ( .A0(n407), .A1(n732), .B0(n4208), .B1(n704), .Y(n6040) );
  AOI222XLTS U3105 ( .A0(n228), .A1(n27), .B0(n3897), .B1(n122), .C0(n4366), 
        .C1(n3789), .Y(n6039) );
  AOI22X1TS U3106 ( .A0(n409), .A1(n738), .B0(n4205), .B1(n703), .Y(n6042) );
  AOI222XLTS U3107 ( .A0(n233), .A1(n28), .B0(n3894), .B1(n125), .C0(n4363), 
        .C1(n3788), .Y(n6041) );
  AOI22X1TS U3108 ( .A0(n411), .A1(n742), .B0(n4202), .B1(n703), .Y(n6044) );
  AOI222XLTS U3109 ( .A0(n231), .A1(n29), .B0(n3891), .B1(n121), .C0(n4360), 
        .C1(n3788), .Y(n6043) );
  AOI22X1TS U3110 ( .A0(n415), .A1(n6104), .B0(n4196), .B1(n703), .Y(n6048) );
  AOI222XLTS U3111 ( .A0(n208), .A1(n30), .B0(n3885), .B1(n125), .C0(n4354), 
        .C1(n3788), .Y(n6047) );
  AOI22X1TS U3112 ( .A0(n417), .A1(n717), .B0(n4193), .B1(n702), .Y(n6050) );
  AOI222XLTS U3113 ( .A0(n338), .A1(n31), .B0(n3882), .B1(n124), .C0(n4351), 
        .C1(n3787), .Y(n6049) );
  AOI22X1TS U3114 ( .A0(n421), .A1(n717), .B0(n4187), .B1(n702), .Y(n6054) );
  AOI222XLTS U3115 ( .A0(n231), .A1(n32), .B0(n3876), .B1(n116), .C0(n4345), 
        .C1(n3787), .Y(n6053) );
  AOI22X1TS U3116 ( .A0(n423), .A1(n729), .B0(n4184), .B1(n701), .Y(n6056) );
  AOI222XLTS U3117 ( .A0(n229), .A1(n33), .B0(n3873), .B1(n122), .C0(n4342), 
        .C1(n3787), .Y(n6055) );
  AOI22X1TS U3118 ( .A0(n425), .A1(n717), .B0(n4181), .B1(n701), .Y(n6058) );
  AOI222XLTS U3119 ( .A0(n190), .A1(n34), .B0(n3870), .B1(n120), .C0(n4339), 
        .C1(n3786), .Y(n6057) );
  AOI22X1TS U3120 ( .A0(n427), .A1(n729), .B0(n4178), .B1(n701), .Y(n6060) );
  AOI222XLTS U3121 ( .A0(n209), .A1(n35), .B0(n3867), .B1(n112), .C0(n4336), 
        .C1(n3786), .Y(n6059) );
  AOI22X1TS U3122 ( .A0(n429), .A1(n732), .B0(n4175), .B1(n701), .Y(n6062) );
  AOI222XLTS U3123 ( .A0(n233), .A1(n36), .B0(n3864), .B1(n116), .C0(n4333), 
        .C1(n3786), .Y(n6061) );
  AOI22X1TS U3124 ( .A0(n431), .A1(n729), .B0(n4172), .B1(n700), .Y(n6064) );
  AOI222XLTS U3125 ( .A0(n209), .A1(n37), .B0(n3861), .B1(n113), .C0(n4330), 
        .C1(n3786), .Y(n6063) );
  AOI22X1TS U3126 ( .A0(n433), .A1(n729), .B0(n4169), .B1(n700), .Y(n6066) );
  AOI222XLTS U3127 ( .A0(n210), .A1(n38), .B0(n3858), .B1(n122), .C0(n4327), 
        .C1(n3785), .Y(n6065) );
  AOI22X1TS U3128 ( .A0(n435), .A1(n732), .B0(n4166), .B1(n700), .Y(n6068) );
  AOI222XLTS U3129 ( .A0(n231), .A1(n39), .B0(n3855), .B1(n120), .C0(n4324), 
        .C1(n3785), .Y(n6067) );
  AOI22X1TS U3130 ( .A0(n437), .A1(n732), .B0(n4163), .B1(n700), .Y(n6070) );
  AOI222XLTS U3131 ( .A0(n338), .A1(n40), .B0(n3852), .B1(n121), .C0(n4321), 
        .C1(n3785), .Y(n6069) );
  AOI22X1TS U3132 ( .A0(n439), .A1(n735), .B0(n4160), .B1(n699), .Y(n6072) );
  AOI222XLTS U3133 ( .A0(n228), .A1(n41), .B0(n3849), .B1(n120), .C0(n4318), 
        .C1(n3785), .Y(n6071) );
  AOI22X1TS U3134 ( .A0(n443), .A1(n733), .B0(n4154), .B1(n699), .Y(n6076) );
  AOI222XLTS U3135 ( .A0(n231), .A1(n42), .B0(n3843), .B1(n121), .C0(n4312), 
        .C1(n3784), .Y(n6075) );
  AOI22X1TS U3136 ( .A0(n445), .A1(n733), .B0(n4151), .B1(n699), .Y(n6078) );
  AOI222XLTS U3137 ( .A0(n233), .A1(n43), .B0(n3840), .B1(n117), .C0(n4309), 
        .C1(n3784), .Y(n6077) );
  AOI22X1TS U3138 ( .A0(n447), .A1(n734), .B0(n4148), .B1(n699), .Y(n6080) );
  AOI222XLTS U3139 ( .A0(n229), .A1(n44), .B0(n3837), .B1(n118), .C0(n4306), 
        .C1(n3784), .Y(n6079) );
  AOI22X1TS U3140 ( .A0(n451), .A1(n734), .B0(n4142), .B1(n698), .Y(n6084) );
  AOI222XLTS U3141 ( .A0(n209), .A1(n45), .B0(n3831), .B1(n123), .C0(n4300), 
        .C1(n3798), .Y(n6083) );
  AOI22X1TS U3142 ( .A0(n453), .A1(n735), .B0(n4139), .B1(n698), .Y(n6086) );
  AOI222XLTS U3143 ( .A0(n233), .A1(n46), .B0(n3828), .B1(n114), .C0(n4297), 
        .C1(n3796), .Y(n6085) );
  AOI22X1TS U3144 ( .A0(n716), .A1(n158), .B0(n4256), .B1(n6103), .Y(n5334) );
  AOI222XLTS U3145 ( .A0(n229), .A1(n47), .B0(n3945), .B1(n119), .C0(n4414), 
        .C1(n3791), .Y(n5333) );
  AOI22X1TS U3146 ( .A0(n716), .A1(n135), .B0(n4244), .B1(n711), .Y(n5342) );
  AOI222XLTS U3147 ( .A0(n228), .A1(n48), .B0(n3933), .B1(n114), .C0(n4402), 
        .C1(n3790), .Y(n5341) );
  AOI22X1TS U3148 ( .A0(n403), .A1(n737), .B0(n4214), .B1(n704), .Y(n6036) );
  AOI222XLTS U3149 ( .A0(n6347), .A1(n49), .B0(n3903), .B1(n124), .C0(n4372), 
        .C1(n3789), .Y(n6035) );
  AOI22X1TS U3150 ( .A0(n405), .A1(n739), .B0(n4211), .B1(n704), .Y(n6038) );
  AOI222XLTS U3151 ( .A0(n3769), .A1(n50), .B0(n3900), .B1(n120), .C0(n4369), 
        .C1(n3789), .Y(n6037) );
  AOI22X1TS U3152 ( .A0(n413), .A1(n741), .B0(n4199), .B1(n703), .Y(n6046) );
  AOI222XLTS U3153 ( .A0(n230), .A1(n51), .B0(n3888), .B1(n119), .C0(n4357), 
        .C1(n3788), .Y(n6045) );
  AOI22X1TS U3154 ( .A0(n419), .A1(n717), .B0(n4190), .B1(n702), .Y(n6052) );
  AOI222XLTS U3155 ( .A0(n210), .A1(n52), .B0(n3879), .B1(n111), .C0(n4348), 
        .C1(n3787), .Y(n6051) );
  AOI22X1TS U3156 ( .A0(n441), .A1(n733), .B0(n4157), .B1(n702), .Y(n6074) );
  AOI222XLTS U3157 ( .A0(n3769), .A1(n53), .B0(n3846), .B1(n116), .C0(n4315), 
        .C1(n3784), .Y(n6073) );
  AOI22X1TS U3158 ( .A0(n449), .A1(n733), .B0(n4145), .B1(n698), .Y(n6082) );
  AOI222XLTS U3159 ( .A0(n338), .A1(n54), .B0(n3834), .B1(n119), .C0(n4303), 
        .C1(n3796), .Y(n6081) );
  AOI22X1TS U3160 ( .A0(n455), .A1(n734), .B0(n4136), .B1(n698), .Y(n6088) );
  AOI222XLTS U3161 ( .A0(n210), .A1(n55), .B0(n3825), .B1(n111), .C0(n4294), 
        .C1(n3796), .Y(n6087) );
  AOI22X1TS U3162 ( .A0(n457), .A1(n734), .B0(n4133), .B1(n697), .Y(n6090) );
  AOI222XLTS U3163 ( .A0(n3769), .A1(n56), .B0(n3822), .B1(n111), .C0(n4291), 
        .C1(n3792), .Y(n6089) );
  AOI22X1TS U3164 ( .A0(n459), .A1(n735), .B0(n4130), .B1(n697), .Y(n6092) );
  AOI222XLTS U3165 ( .A0(n210), .A1(n57), .B0(n3819), .B1(n117), .C0(n4288), 
        .C1(n3796), .Y(n6091) );
  AOI22X1TS U3166 ( .A0(n3213), .A1(n161), .B0(n4259), .B1(n3204), .Y(n5402)
         );
  AOI222XLTS U3167 ( .A0(n3261), .A1(n6250), .B0(n3948), .B1(n3246), .C0(n4417), .C1(n3237), .Y(n5401) );
  AOI22X1TS U3168 ( .A0(n3213), .A1(n158), .B0(n4256), .B1(n3204), .Y(n5404)
         );
  AOI222XLTS U3169 ( .A0(n3261), .A1(n6251), .B0(n3945), .B1(n3253), .C0(n4414), .C1(n3237), .Y(n5403) );
  AOI22X1TS U3170 ( .A0(n3213), .A1(n153), .B0(n4253), .B1(n3204), .Y(n5406)
         );
  AOI222XLTS U3171 ( .A0(n3261), .A1(n6252), .B0(n3942), .B1(n3256), .C0(n4411), .C1(n3237), .Y(n5405) );
  AOI22X1TS U3172 ( .A0(n3214), .A1(n143), .B0(n4247), .B1(n3206), .Y(n5410)
         );
  AOI222XLTS U3173 ( .A0(n3262), .A1(n6253), .B0(n3936), .B1(n3252), .C0(n4405), .C1(n3236), .Y(n5409) );
  AOI22X1TS U3174 ( .A0(n3214), .A1(readRequesterAddress[0]), .B0(n4244), .B1(
        n3206), .Y(n5412) );
  AOI222XLTS U3175 ( .A0(n3262), .A1(n6254), .B0(n3933), .B1(n3252), .C0(n4402), .C1(n3236), .Y(n5411) );
  AOI22X1TS U3176 ( .A0(n397), .A1(n3220), .B0(n4223), .B1(n3210), .Y(n5838)
         );
  AOI222XLTS U3177 ( .A0(n3262), .A1(n6255), .B0(n3912), .B1(n3252), .C0(n4381), .C1(n3236), .Y(n5837) );
  AOI22X1TS U3178 ( .A0(n399), .A1(n3220), .B0(n4220), .B1(n3209), .Y(n5840)
         );
  AOI222XLTS U3179 ( .A0(n3262), .A1(n6256), .B0(n3909), .B1(n3252), .C0(n4378), .C1(n3236), .Y(n5839) );
  AOI22X1TS U3180 ( .A0(n401), .A1(n3220), .B0(n4217), .B1(n3207), .Y(n5842)
         );
  AOI222XLTS U3181 ( .A0(n3263), .A1(n6257), .B0(n3906), .B1(n3251), .C0(n4375), .C1(n3235), .Y(n5841) );
  AOI22X1TS U3182 ( .A0(n403), .A1(n3225), .B0(n4214), .B1(n3207), .Y(n5844)
         );
  AOI222XLTS U3183 ( .A0(n3263), .A1(n6258), .B0(n3903), .B1(n3251), .C0(n4372), .C1(n3235), .Y(n5843) );
  AOI22X1TS U3184 ( .A0(n405), .A1(n3220), .B0(n4211), .B1(n3206), .Y(n5846)
         );
  AOI222XLTS U3185 ( .A0(n3263), .A1(n6259), .B0(n3900), .B1(n3251), .C0(n4369), .C1(n3235), .Y(n5845) );
  AOI22X1TS U3186 ( .A0(n407), .A1(n3219), .B0(n4208), .B1(n3206), .Y(n5848)
         );
  AOI222XLTS U3187 ( .A0(n3263), .A1(n6260), .B0(n3897), .B1(n3251), .C0(n4366), .C1(n3235), .Y(n5847) );
  AOI22X1TS U3188 ( .A0(n411), .A1(n3219), .B0(n4202), .B1(n3203), .Y(n5852)
         );
  AOI222XLTS U3189 ( .A0(n3264), .A1(n6261), .B0(n3891), .B1(n3250), .C0(n4360), .C1(n3234), .Y(n5851) );
  AOI22X1TS U3190 ( .A0(n415), .A1(n3222), .B0(n4196), .B1(n3203), .Y(n5856)
         );
  AOI222XLTS U3191 ( .A0(n3264), .A1(n6262), .B0(n3885), .B1(n3250), .C0(n4354), .C1(n3234), .Y(n5855) );
  AOI22X1TS U3192 ( .A0(n417), .A1(n6149), .B0(n4193), .B1(n3202), .Y(n5858)
         );
  AOI222XLTS U3193 ( .A0(n3265), .A1(n6263), .B0(n3882), .B1(n3255), .C0(n4351), .C1(n3233), .Y(n5857) );
  AOI22X1TS U3194 ( .A0(n421), .A1(n6149), .B0(n4187), .B1(n3202), .Y(n5862)
         );
  AOI222XLTS U3195 ( .A0(n3265), .A1(n6264), .B0(n3876), .B1(n3255), .C0(n4345), .C1(n3233), .Y(n5861) );
  AOI22X1TS U3196 ( .A0(n425), .A1(n3224), .B0(n4181), .B1(n3201), .Y(n5866)
         );
  AOI222XLTS U3197 ( .A0(n3266), .A1(n6265), .B0(n3870), .B1(n3257), .C0(n4339), .C1(n3232), .Y(n5865) );
  AOI22X1TS U3198 ( .A0(n427), .A1(n3224), .B0(n4178), .B1(n3201), .Y(n5868)
         );
  AOI222XLTS U3199 ( .A0(n3266), .A1(n6266), .B0(n3867), .B1(n3253), .C0(n4336), .C1(n3232), .Y(n5867) );
  AOI22X1TS U3200 ( .A0(n431), .A1(n3222), .B0(n4172), .B1(n3200), .Y(n5872)
         );
  AOI222XLTS U3201 ( .A0(n3266), .A1(n6267), .B0(n3861), .B1(n3249), .C0(n4330), .C1(n3232), .Y(n5871) );
  AOI22X1TS U3202 ( .A0(n435), .A1(n3223), .B0(n4166), .B1(n3200), .Y(n5876)
         );
  AOI222XLTS U3203 ( .A0(n3267), .A1(n6268), .B0(n3855), .B1(n3249), .C0(n4324), .C1(n3231), .Y(n5875) );
  AOI22X1TS U3204 ( .A0(n437), .A1(n3218), .B0(n4163), .B1(n3200), .Y(n5878)
         );
  AOI222XLTS U3205 ( .A0(n3267), .A1(n6269), .B0(n3852), .B1(n3249), .C0(n4321), .C1(n3231), .Y(n5877) );
  AOI22X1TS U3206 ( .A0(n439), .A1(n3218), .B0(n4160), .B1(n3199), .Y(n5880)
         );
  AOI222XLTS U3207 ( .A0(n3267), .A1(n6270), .B0(n3849), .B1(n3248), .C0(n4318), .C1(n3231), .Y(n5879) );
  AOI22X1TS U3208 ( .A0(n441), .A1(n3218), .B0(n4157), .B1(n3202), .Y(n5882)
         );
  AOI222XLTS U3209 ( .A0(n3268), .A1(n6271), .B0(n3846), .B1(n3248), .C0(n4315), .C1(n3230), .Y(n5881) );
  AOI22X1TS U3210 ( .A0(n443), .A1(n3218), .B0(n4154), .B1(n3199), .Y(n5884)
         );
  AOI222XLTS U3211 ( .A0(n3268), .A1(n6272), .B0(n3843), .B1(n3248), .C0(n4312), .C1(n3230), .Y(n5883) );
  AOI22X1TS U3212 ( .A0(n447), .A1(n3217), .B0(n4148), .B1(n3199), .Y(n5888)
         );
  AOI222XLTS U3213 ( .A0(n3268), .A1(n6273), .B0(n3837), .B1(n3253), .C0(n4306), .C1(n3230), .Y(n5887) );
  AOI22X1TS U3214 ( .A0(n453), .A1(n3216), .B0(n4139), .B1(n3198), .Y(n5894)
         );
  AOI222XLTS U3215 ( .A0(n3269), .A1(n6274), .B0(n3828), .B1(n3247), .C0(n4297), .C1(n3229), .Y(n5893) );
  AOI22X1TS U3216 ( .A0(n457), .A1(n3216), .B0(n4133), .B1(n3197), .Y(n5898)
         );
  AOI222XLTS U3217 ( .A0(n3270), .A1(n6275), .B0(n3822), .B1(n3246), .C0(n4291), .C1(n3228), .Y(n5897) );
  AOI22X1TS U3218 ( .A0(n459), .A1(n3216), .B0(n4130), .B1(n3197), .Y(n5900)
         );
  AOI222XLTS U3219 ( .A0(n3270), .A1(n6276), .B0(n3819), .B1(n3246), .C0(n4288), .C1(n3228), .Y(n5899) );
  AOI22X1TS U3220 ( .A0(n3214), .A1(n148), .B0(n4250), .B1(n3204), .Y(n5408)
         );
  AOI222XLTS U3221 ( .A0(n3261), .A1(n6291), .B0(n3939), .B1(n3259), .C0(n4408), .C1(n3237), .Y(n5407) );
  AOI22X1TS U3222 ( .A0(n409), .A1(n3219), .B0(n4205), .B1(n3203), .Y(n5850)
         );
  AOI222XLTS U3223 ( .A0(n3264), .A1(n6292), .B0(n3894), .B1(n3250), .C0(n4363), .C1(n3234), .Y(n5849) );
  AOI22X1TS U3224 ( .A0(n413), .A1(n3219), .B0(n4199), .B1(n3203), .Y(n5854)
         );
  AOI222XLTS U3225 ( .A0(n3264), .A1(n6293), .B0(n3888), .B1(n3250), .C0(n4357), .C1(n3234), .Y(n5853) );
  AOI22X1TS U3226 ( .A0(n419), .A1(n3221), .B0(n4190), .B1(n3202), .Y(n5860)
         );
  AOI222XLTS U3227 ( .A0(n3265), .A1(n6294), .B0(n3879), .B1(n3254), .C0(n4348), .C1(n3233), .Y(n5859) );
  AOI22X1TS U3228 ( .A0(n423), .A1(n3222), .B0(n4184), .B1(n3201), .Y(n5864)
         );
  AOI222XLTS U3229 ( .A0(n3265), .A1(n6295), .B0(n3873), .B1(n3255), .C0(n4342), .C1(n3233), .Y(n5863) );
  AOI22X1TS U3230 ( .A0(n429), .A1(n3223), .B0(n4175), .B1(n3201), .Y(n5870)
         );
  AOI222XLTS U3231 ( .A0(n3266), .A1(n6296), .B0(n3864), .B1(n3257), .C0(n4333), .C1(n3232), .Y(n5869) );
  AOI22X1TS U3232 ( .A0(n433), .A1(n3225), .B0(n4169), .B1(n3200), .Y(n5874)
         );
  AOI222XLTS U3233 ( .A0(n3267), .A1(n6297), .B0(n3858), .B1(n3249), .C0(n4327), .C1(n3231), .Y(n5873) );
  AOI22X1TS U3234 ( .A0(n449), .A1(n3217), .B0(n4145), .B1(n3198), .Y(n5890)
         );
  AOI222XLTS U3235 ( .A0(n3269), .A1(n6298), .B0(n3834), .B1(n3247), .C0(n4303), .C1(n3229), .Y(n5889) );
  AOI22X1TS U3236 ( .A0(n451), .A1(n3217), .B0(n4142), .B1(n3198), .Y(n5892)
         );
  AOI222XLTS U3237 ( .A0(n3269), .A1(n6299), .B0(n3831), .B1(n3247), .C0(n4300), .C1(n3229), .Y(n5891) );
  AOI22X1TS U3238 ( .A0(n455), .A1(n3216), .B0(n4136), .B1(n3198), .Y(n5896)
         );
  AOI222XLTS U3239 ( .A0(n3269), .A1(n6300), .B0(n3825), .B1(n3247), .C0(n4294), .C1(n3229), .Y(n5895) );
  AOI22X1TS U3240 ( .A0(n445), .A1(n3217), .B0(n4151), .B1(n3199), .Y(n5886)
         );
  AOI222XLTS U3241 ( .A0(n3268), .A1(n6313), .B0(n3840), .B1(n3248), .C0(n4309), .C1(n3230), .Y(n5885) );
  AOI22X1TS U3242 ( .A0(n846), .A1(n145), .B0(n4094), .B1(n835), .Y(n5382) );
  AOI222XLTS U3243 ( .A0(n250), .A1(n58), .B0(n4251), .B1(n957), .C0(n4408), 
        .C1(n3760), .Y(n5381) );
  AOI22X1TS U3244 ( .A0(n400), .A1(n856), .B0(n4064), .B1(n838), .Y(n5904) );
  AOI222XLTS U3245 ( .A0(n257), .A1(n59), .B0(n4221), .B1(n919), .C0(n4378), 
        .C1(n3759), .Y(n5903) );
  AOI22X1TS U3246 ( .A0(n402), .A1(n856), .B0(n4061), .B1(n838), .Y(n5906) );
  AOI222XLTS U3247 ( .A0(n339), .A1(n60), .B0(n4218), .B1(n869), .C0(n4375), 
        .C1(n3762), .Y(n5905) );
  AOI22X1TS U3248 ( .A0(n404), .A1(n853), .B0(n4058), .B1(n842), .Y(n5908) );
  AOI222XLTS U3249 ( .A0(n339), .A1(n61), .B0(n4215), .B1(n869), .C0(n4372), 
        .C1(n3762), .Y(n5907) );
  AOI22X1TS U3250 ( .A0(n408), .A1(n849), .B0(n4052), .B1(n844), .Y(n5912) );
  AOI222XLTS U3251 ( .A0(n250), .A1(n62), .B0(n4209), .B1(n869), .C0(n4366), 
        .C1(n3762), .Y(n5911) );
  AOI22X1TS U3252 ( .A0(n410), .A1(n854), .B0(n4049), .B1(n839), .Y(n5914) );
  AOI222XLTS U3253 ( .A0(n259), .A1(n63), .B0(n4206), .B1(n868), .C0(n4363), 
        .C1(n3763), .Y(n5913) );
  AOI22X1TS U3254 ( .A0(n414), .A1(n859), .B0(n4043), .B1(n839), .Y(n5918) );
  AOI222XLTS U3255 ( .A0(n261), .A1(n64), .B0(n4200), .B1(n868), .C0(n4357), 
        .C1(n3762), .Y(n5917) );
  AOI22X1TS U3256 ( .A0(n418), .A1(n847), .B0(n4037), .B1(n839), .Y(n5922) );
  AOI222XLTS U3257 ( .A0(n257), .A1(n65), .B0(n4194), .B1(n867), .C0(n4351), 
        .C1(n3765), .Y(n5921) );
  AOI22X1TS U3258 ( .A0(n420), .A1(n847), .B0(n4034), .B1(n841), .Y(n5924) );
  AOI222XLTS U3259 ( .A0(n259), .A1(n66), .B0(n4191), .B1(n867), .C0(n4348), 
        .C1(n3765), .Y(n5923) );
  AOI22X1TS U3260 ( .A0(n422), .A1(n847), .B0(n4031), .B1(n840), .Y(n5926) );
  AOI222XLTS U3261 ( .A0(n251), .A1(n67), .B0(n4188), .B1(n867), .C0(n4345), 
        .C1(n3765), .Y(n5925) );
  AOI22X1TS U3262 ( .A0(n424), .A1(n848), .B0(n4028), .B1(n834), .Y(n5928) );
  AOI222XLTS U3263 ( .A0(n261), .A1(n68), .B0(n4185), .B1(n866), .C0(n4342), 
        .C1(n3767), .Y(n5927) );
  AOI22X1TS U3264 ( .A0(n426), .A1(n847), .B0(n4025), .B1(n834), .Y(n5930) );
  AOI222XLTS U3265 ( .A0(n341), .A1(n69), .B0(n4182), .B1(n866), .C0(n4339), 
        .C1(n3758), .Y(n5929) );
  AOI22X1TS U3266 ( .A0(n430), .A1(n849), .B0(n4019), .B1(n834), .Y(n5934) );
  AOI222XLTS U3267 ( .A0(n250), .A1(n70), .B0(n4176), .B1(n866), .C0(n4333), 
        .C1(n3758), .Y(n5933) );
  AOI22X1TS U3268 ( .A0(n432), .A1(n848), .B0(n4016), .B1(n833), .Y(n5936) );
  AOI222XLTS U3269 ( .A0(n260), .A1(n71), .B0(n4173), .B1(n865), .C0(n4330), 
        .C1(n3758), .Y(n5935) );
  AOI22X1TS U3270 ( .A0(n434), .A1(n848), .B0(n4013), .B1(n833), .Y(n5938) );
  AOI222XLTS U3271 ( .A0(n250), .A1(n72), .B0(n4170), .B1(n865), .C0(n4327), 
        .C1(n3763), .Y(n5937) );
  AOI22X1TS U3272 ( .A0(n436), .A1(n849), .B0(n4010), .B1(n833), .Y(n5940) );
  AOI222XLTS U3273 ( .A0(n261), .A1(n73), .B0(n4167), .B1(n865), .C0(n4324), 
        .C1(n3763), .Y(n5939) );
  AOI22X1TS U3274 ( .A0(n438), .A1(n849), .B0(n4007), .B1(n833), .Y(n5942) );
  AOI222XLTS U3275 ( .A0(n257), .A1(n74), .B0(n4164), .B1(n865), .C0(n4321), 
        .C1(n3761), .Y(n5941) );
  AOI22X1TS U3276 ( .A0(n442), .A1(n850), .B0(n4001), .B1(n842), .Y(n5946) );
  AOI222XLTS U3277 ( .A0(n299), .A1(n75), .B0(n4158), .B1(n864), .C0(n4315), 
        .C1(n3757), .Y(n5945) );
  AOI22X1TS U3278 ( .A0(n444), .A1(n850), .B0(n3998), .B1(n832), .Y(n5948) );
  AOI222XLTS U3279 ( .A0(n260), .A1(n76), .B0(n4155), .B1(n864), .C0(n4312), 
        .C1(n3757), .Y(n5947) );
  AOI22X1TS U3280 ( .A0(n446), .A1(n850), .B0(n3995), .B1(n832), .Y(n5950) );
  AOI222XLTS U3281 ( .A0(n340), .A1(n77), .B0(n4152), .B1(n864), .C0(n4309), 
        .C1(n3757), .Y(n5949) );
  AOI22X1TS U3282 ( .A0(n450), .A1(n850), .B0(n3989), .B1(n831), .Y(n5954) );
  AOI222XLTS U3283 ( .A0(n339), .A1(n78), .B0(n4146), .B1(n863), .C0(n4303), 
        .C1(n3756), .Y(n5953) );
  AOI22X1TS U3284 ( .A0(n452), .A1(n851), .B0(n3986), .B1(n831), .Y(n5956) );
  AOI222XLTS U3285 ( .A0(n341), .A1(n79), .B0(n4143), .B1(n863), .C0(n4300), 
        .C1(n3756), .Y(n5955) );
  AOI22X1TS U3286 ( .A0(n454), .A1(n852), .B0(n3983), .B1(n831), .Y(n5958) );
  AOI222XLTS U3287 ( .A0(n259), .A1(n80), .B0(n4140), .B1(n863), .C0(n4297), 
        .C1(n3756), .Y(n5957) );
  AOI22X1TS U3288 ( .A0(n857), .A1(readRequesterAddress[5]), .B0(n4103), .B1(
        n835), .Y(n5376) );
  AOI222XLTS U3289 ( .A0(n297), .A1(n81), .B0(n4260), .B1(n862), .C0(n4417), 
        .C1(n3760), .Y(n5375) );
  AOI22X1TS U3290 ( .A0(n846), .A1(n155), .B0(n4100), .B1(n835), .Y(n5378) );
  AOI222XLTS U3291 ( .A0(n297), .A1(n82), .B0(n4257), .B1(n870), .C0(n4414), 
        .C1(n3760), .Y(n5377) );
  AOI22X1TS U3292 ( .A0(n846), .A1(n150), .B0(n4097), .B1(n835), .Y(n5380) );
  AOI222XLTS U3293 ( .A0(n298), .A1(n83), .B0(n4254), .B1(n936), .C0(n4411), 
        .C1(n3760), .Y(n5379) );
  AOI22X1TS U3294 ( .A0(n855), .A1(n140), .B0(n4091), .B1(n838), .Y(n5384) );
  AOI222XLTS U3295 ( .A0(n261), .A1(n84), .B0(n4248), .B1(n919), .C0(n4405), 
        .C1(n3759), .Y(n5383) );
  AOI22X1TS U3296 ( .A0(n846), .A1(n136), .B0(n4088), .B1(n841), .Y(n5386) );
  AOI222XLTS U3297 ( .A0(n251), .A1(n85), .B0(n4245), .B1(n886), .C0(n4402), 
        .C1(n3759), .Y(n5385) );
  AOI22X1TS U3298 ( .A0(n406), .A1(n6134), .B0(n4055), .B1(n6133), .Y(n5910)
         );
  AOI222XLTS U3299 ( .A0(n341), .A1(n86), .B0(n4212), .B1(n869), .C0(n4369), 
        .C1(n3761), .Y(n5909) );
  AOI22X1TS U3300 ( .A0(n440), .A1(n852), .B0(n4004), .B1(n832), .Y(n5944) );
  AOI222XLTS U3301 ( .A0(n257), .A1(n87), .B0(n4161), .B1(n864), .C0(n4318), 
        .C1(n3764), .Y(n5943) );
  AOI22X1TS U3302 ( .A0(n458), .A1(n851), .B0(n3977), .B1(n830), .Y(n5962) );
  AOI222XLTS U3303 ( .A0(n299), .A1(n88), .B0(n4134), .B1(n862), .C0(n4291), 
        .C1(n3755), .Y(n5961) );
  AOI22X1TS U3304 ( .A0(n398), .A1(n852), .B0(n4067), .B1(n840), .Y(n5902) );
  AOI222XLTS U3305 ( .A0(n260), .A1(n89), .B0(n4224), .B1(n6135), .C0(n4381), 
        .C1(n3759), .Y(n5901) );
  AOI22X1TS U3306 ( .A0(n412), .A1(n856), .B0(n4046), .B1(n838), .Y(n5916) );
  AOI222XLTS U3307 ( .A0(n260), .A1(n90), .B0(n4203), .B1(n868), .C0(n4360), 
        .C1(n3764), .Y(n5915) );
  AOI22X1TS U3308 ( .A0(n416), .A1(n858), .B0(n4040), .B1(n839), .Y(n5920) );
  AOI222XLTS U3309 ( .A0(n340), .A1(n91), .B0(n4197), .B1(n868), .C0(n4354), 
        .C1(n3766), .Y(n5919) );
  AOI22X1TS U3310 ( .A0(n428), .A1(n848), .B0(n4022), .B1(n834), .Y(n5932) );
  AOI222XLTS U3311 ( .A0(n341), .A1(n92), .B0(n4179), .B1(n866), .C0(n4336), 
        .C1(n3758), .Y(n5931) );
  AOI22X1TS U3312 ( .A0(n448), .A1(n851), .B0(n3992), .B1(n832), .Y(n5952) );
  AOI222XLTS U3313 ( .A0(n340), .A1(n93), .B0(n4149), .B1(n867), .C0(n4306), 
        .C1(n3757), .Y(n5951) );
  AOI22X1TS U3314 ( .A0(n456), .A1(n851), .B0(n3980), .B1(n831), .Y(n5960) );
  AOI222XLTS U3315 ( .A0(n298), .A1(n94), .B0(n4137), .B1(n863), .C0(n4294), 
        .C1(n3756), .Y(n5959) );
  AOI22X1TS U3316 ( .A0(n460), .A1(n852), .B0(n3974), .B1(n830), .Y(n5964) );
  AOI222XLTS U3317 ( .A0(n251), .A1(n95), .B0(n4131), .B1(n862), .C0(n4288), 
        .C1(n3755), .Y(n5963) );
  AOI22X1TS U3318 ( .A0(n3929), .A1(n3476), .B0(n4398), .B1(n3703), .Y(n6202)
         );
  AOI222XLTS U3319 ( .A0(n4085), .A1(n3524), .B0(n160), .B1(n3514), .C0(n4242), 
        .C1(n3495), .Y(n6201) );
  AOI22X1TS U3320 ( .A0(n3926), .A1(n3475), .B0(n4395), .B1(n3703), .Y(n6204)
         );
  AOI222XLTS U3321 ( .A0(n4082), .A1(n3523), .B0(n158), .B1(n3514), .C0(n4239), 
        .C1(n3495), .Y(n6203) );
  AOI22X1TS U3322 ( .A0(n3920), .A1(n3475), .B0(n4389), .B1(n3704), .Y(n6208)
         );
  AOI222XLTS U3323 ( .A0(n4076), .A1(n3523), .B0(n145), .B1(n3515), .C0(n4233), 
        .C1(n3495), .Y(n6207) );
  AOI22X1TS U3324 ( .A0(n3923), .A1(n3475), .B0(n4392), .B1(n3704), .Y(n6206)
         );
  AOI222XLTS U3325 ( .A0(n4079), .A1(n3523), .B0(n150), .B1(n3515), .C0(n4236), 
        .C1(n3494), .Y(n6205) );
  AOI22X1TS U3326 ( .A0(n3917), .A1(n3475), .B0(n4386), .B1(n3704), .Y(n6210)
         );
  AOI222XLTS U3327 ( .A0(n4073), .A1(n3523), .B0(n140), .B1(n3515), .C0(n4230), 
        .C1(n3494), .Y(n6209) );
  AOI22X1TS U3328 ( .A0(n3914), .A1(n3485), .B0(n4383), .B1(n3704), .Y(n6216)
         );
  AOI222XLTS U3329 ( .A0(n4070), .A1(n3525), .B0(n135), .B1(n3515), .C0(n4227), 
        .C1(n3499), .Y(n6215) );
  NAND2X1TS U3330 ( .A(n3802), .B(n6340), .Y(n5540) );
  AOI2BB2X1TS U3331 ( .B0(n5534), .B1(n5533), .A0N(n3272), .A1N(
        readOutbuffer[3]), .Y(n2566) );
  OAI22X1TS U3332 ( .A0(n387), .A1(n6226), .B0(n173), .B1(n6227), .Y(n2887) );
  OAI22X1TS U3333 ( .A0(n6225), .A1(n6228), .B0(n5326), .B1(n6227), .Y(n2886)
         );
  OAI22X1TS U3334 ( .A0(n6229), .A1(n387), .B0(n5327), .B1(n6227), .Y(n2888)
         );
  OAI221XLTS U3335 ( .A0(readIn_SOUTH), .A1(n6326), .B0(n3816), .B1(n5557), 
        .C0(n5556), .Y(n5561) );
  AOI222XLTS U3336 ( .A0(n3808), .A1(n5552), .B0(readIn_SOUTH), .B1(n5551), 
        .C0(n3816), .C1(n5550), .Y(n5553) );
  OAI22X1TS U3337 ( .A0(n662), .A1(n4707), .B0(n5130), .B1(n3575), .Y(n5131)
         );
  NOR4XLTS U3338 ( .A(n5129), .B(n5128), .C(n5127), .D(n5126), .Y(n5130) );
  AO22X1TS U3339 ( .A0(n207), .A1(\requesterAddressbuffer[3][5] ), .B0(
        \requesterAddressbuffer[6][5] ), .B1(n5282), .Y(n5128) );
  OAI2BB2XLTS U3340 ( .B0(n6301), .B1(n3632), .A0N(
        \requesterAddressbuffer[0][5] ), .A1N(n246), .Y(n5129) );
  OAI22X1TS U3341 ( .A0(n662), .A1(n4708), .B0(n5138), .B1(n3575), .Y(n5139)
         );
  NOR4XLTS U3342 ( .A(n5137), .B(n5136), .C(n5135), .D(n5134), .Y(n5138) );
  AO22X1TS U3343 ( .A0(n253), .A1(\requesterAddressbuffer[3][4] ), .B0(
        \requesterAddressbuffer[6][4] ), .B1(n5282), .Y(n5136) );
  OAI2BB2XLTS U3344 ( .B0(n6302), .B1(n3632), .A0N(
        \requesterAddressbuffer[0][4] ), .A1N(n5283), .Y(n5137) );
  OAI22X1TS U3345 ( .A0(n661), .A1(n4709), .B0(n5154), .B1(n3574), .Y(n5155)
         );
  NOR4XLTS U3346 ( .A(n5153), .B(n5152), .C(n5151), .D(n5150), .Y(n5154) );
  AO22X1TS U3347 ( .A0(n207), .A1(\requesterAddressbuffer[3][2] ), .B0(
        \requesterAddressbuffer[6][2] ), .B1(n5282), .Y(n5152) );
  OAI2BB2XLTS U3348 ( .B0(n6278), .B1(n3619), .A0N(
        \requesterAddressbuffer[0][2] ), .A1N(n246), .Y(n5153) );
  OAI22X1TS U3349 ( .A0(n661), .A1(n4710), .B0(n5162), .B1(n3574), .Y(n5163)
         );
  NOR4XLTS U3350 ( .A(n5161), .B(n5160), .C(n5159), .D(n5158), .Y(n5162) );
  AO22X1TS U3351 ( .A0(n253), .A1(\requesterAddressbuffer[3][1] ), .B0(
        \requesterAddressbuffer[6][1] ), .B1(n396), .Y(n5160) );
  OAI2BB2XLTS U3352 ( .B0(n6279), .B1(n3619), .A0N(
        \requesterAddressbuffer[0][1] ), .A1N(n5283), .Y(n5161) );
  OAI22X1TS U3353 ( .A0(n661), .A1(n4834), .B0(n5146), .B1(n3574), .Y(n5147)
         );
  NOR4XLTS U3354 ( .A(n5145), .B(n5144), .C(n5143), .D(n5142), .Y(n5146) );
  AO22X1TS U3355 ( .A0(n207), .A1(\requesterAddressbuffer[3][3] ), .B0(
        \requesterAddressbuffer[6][3] ), .B1(n396), .Y(n5144) );
  OAI2BB2XLTS U3356 ( .B0(n6277), .B1(n3619), .A0N(
        \requesterAddressbuffer[0][3] ), .A1N(n246), .Y(n5145) );
  OAI22X1TS U3357 ( .A0(n661), .A1(n4833), .B0(n5170), .B1(n3574), .Y(n5171)
         );
  NOR4XLTS U3358 ( .A(n5169), .B(n5168), .C(n5167), .D(n5166), .Y(n5170) );
  AO22X1TS U3359 ( .A0(n253), .A1(\requesterAddressbuffer[3][0] ), .B0(
        \requesterAddressbuffer[6][0] ), .B1(n396), .Y(n5168) );
  OAI2BB2XLTS U3360 ( .B0(n6280), .B1(n3619), .A0N(
        \requesterAddressbuffer[0][0] ), .A1N(n5283), .Y(n5169) );
  OAI22X1TS U3361 ( .A0(n4419), .A1(n662), .B0(n4874), .B1(n3572), .Y(n4875)
         );
  NOR4XLTS U3362 ( .A(n4873), .B(n4872), .C(n4871), .D(n4870), .Y(n4874) );
  OAI22X1TS U3363 ( .A0(n4420), .A1(n3616), .B0(n4421), .B1(n3620), .Y(n4873)
         );
  OAI22X1TS U3364 ( .A0(n4422), .A1(n3664), .B0(n4423), .B1(n3666), .Y(n4872)
         );
  OAI22X1TS U3365 ( .A0(n4428), .A1(n671), .B0(n4882), .B1(n3586), .Y(n4883)
         );
  NOR4XLTS U3366 ( .A(n4881), .B(n4880), .C(n4879), .D(n4878), .Y(n4882) );
  OAI22X1TS U3367 ( .A0(n4433), .A1(n3616), .B0(n4429), .B1(n3625), .Y(n4881)
         );
  OAI22X1TS U3368 ( .A0(n4435), .A1(n3657), .B0(n4434), .B1(n3666), .Y(n4880)
         );
  OAI22X1TS U3369 ( .A0(n4437), .A1(n671), .B0(n4890), .B1(n3584), .Y(n4891)
         );
  NOR4XLTS U3370 ( .A(n4889), .B(n4888), .C(n4887), .D(n4886), .Y(n4890) );
  OAI22X1TS U3371 ( .A0(n4444), .A1(n3614), .B0(n4445), .B1(n3625), .Y(n4889)
         );
  OAI22X1TS U3372 ( .A0(n4440), .A1(n3657), .B0(n4442), .B1(n3666), .Y(n4888)
         );
  OAI22X1TS U3373 ( .A0(n4446), .A1(n671), .B0(n4898), .B1(n3581), .Y(n4899)
         );
  NOR4XLTS U3374 ( .A(n4897), .B(n4896), .C(n4895), .D(n4894), .Y(n4898) );
  OAI22X1TS U3375 ( .A0(n4453), .A1(n3615), .B0(n4447), .B1(n3625), .Y(n4897)
         );
  OAI22X1TS U3376 ( .A0(n4451), .A1(n3657), .B0(n4450), .B1(n3666), .Y(n4896)
         );
  OAI22X1TS U3377 ( .A0(n4455), .A1(n671), .B0(n4906), .B1(n3586), .Y(n4907)
         );
  NOR4XLTS U3378 ( .A(n4905), .B(n4904), .C(n4903), .D(n4902), .Y(n4906) );
  OAI22X1TS U3379 ( .A0(n4462), .A1(n3615), .B0(n4458), .B1(n3625), .Y(n4905)
         );
  OAI22X1TS U3380 ( .A0(n4460), .A1(n3656), .B0(n4459), .B1(n3667), .Y(n4904)
         );
  OAI22X1TS U3381 ( .A0(n4464), .A1(n670), .B0(n4914), .B1(n3582), .Y(n4915)
         );
  NOR4XLTS U3382 ( .A(n4913), .B(n4912), .C(n4911), .D(n4910), .Y(n4914) );
  OAI22X1TS U3383 ( .A0(n4469), .A1(n3611), .B0(n4465), .B1(n3624), .Y(n4913)
         );
  OAI22X1TS U3384 ( .A0(n4471), .A1(n3656), .B0(n4470), .B1(n3667), .Y(n4912)
         );
  OAI22X1TS U3385 ( .A0(n4473), .A1(n670), .B0(n4922), .B1(n3581), .Y(n4923)
         );
  NOR4XLTS U3386 ( .A(n4921), .B(n4920), .C(n4919), .D(n4918), .Y(n4922) );
  OAI22X1TS U3387 ( .A0(n4476), .A1(n3616), .B0(n4478), .B1(n3624), .Y(n4921)
         );
  OAI22X1TS U3388 ( .A0(n4475), .A1(n3656), .B0(n4480), .B1(n3667), .Y(n4920)
         );
  OAI22X1TS U3389 ( .A0(n4482), .A1(n670), .B0(n4930), .B1(n3583), .Y(n4931)
         );
  NOR4XLTS U3390 ( .A(n4929), .B(n4928), .C(n4927), .D(n4926), .Y(n4930) );
  OAI22X1TS U3391 ( .A0(n4485), .A1(n3613), .B0(n4483), .B1(n3624), .Y(n4929)
         );
  OAI22X1TS U3392 ( .A0(n4487), .A1(n3656), .B0(n4490), .B1(n3667), .Y(n4928)
         );
  OAI22X1TS U3393 ( .A0(n4491), .A1(n670), .B0(n4938), .B1(n3583), .Y(n4939)
         );
  NOR4XLTS U3394 ( .A(n4937), .B(n4936), .C(n4935), .D(n4934), .Y(n4938) );
  OAI22X1TS U3395 ( .A0(n4498), .A1(n3617), .B0(n4494), .B1(n3624), .Y(n4937)
         );
  OAI22X1TS U3396 ( .A0(n4499), .A1(n3655), .B0(n4492), .B1(n3679), .Y(n4936)
         );
  OAI22X1TS U3397 ( .A0(n4500), .A1(n669), .B0(n4946), .B1(n3586), .Y(n4947)
         );
  NOR4XLTS U3398 ( .A(n4945), .B(n4944), .C(n4943), .D(n4942), .Y(n4946) );
  OAI22X1TS U3399 ( .A0(n4501), .A1(n3613), .B0(n4504), .B1(n3623), .Y(n4945)
         );
  OAI22X1TS U3400 ( .A0(n4503), .A1(n3655), .B0(n4508), .B1(n3676), .Y(n4944)
         );
  OAI22X1TS U3401 ( .A0(n4509), .A1(n669), .B0(n4954), .B1(n3582), .Y(n4955)
         );
  NOR4XLTS U3402 ( .A(n4953), .B(n4952), .C(n4951), .D(n4950), .Y(n4954) );
  OAI22X1TS U3403 ( .A0(n4516), .A1(n3614), .B0(n4515), .B1(n3623), .Y(n4953)
         );
  OAI22X1TS U3404 ( .A0(n4514), .A1(n3655), .B0(n4512), .B1(n3678), .Y(n4952)
         );
  OAI22X1TS U3405 ( .A0(n4518), .A1(n669), .B0(n4962), .B1(n3580), .Y(n4963)
         );
  NOR4XLTS U3406 ( .A(n4961), .B(n4960), .C(n4959), .D(n4958), .Y(n4962) );
  OAI22X1TS U3407 ( .A0(n4525), .A1(n3617), .B0(n4524), .B1(n3623), .Y(n4961)
         );
  OAI22X1TS U3408 ( .A0(n4526), .A1(n3655), .B0(n4519), .B1(n3674), .Y(n4960)
         );
  OAI22X1TS U3409 ( .A0(n4527), .A1(n669), .B0(n4970), .B1(n3580), .Y(n4971)
         );
  NOR4XLTS U3410 ( .A(n4969), .B(n4968), .C(n4967), .D(n4966), .Y(n4970) );
  OAI22X1TS U3411 ( .A0(n4530), .A1(n3612), .B0(n4529), .B1(n3623), .Y(n4969)
         );
  OAI22X1TS U3412 ( .A0(n4534), .A1(n3654), .B0(n4531), .B1(n3677), .Y(n4968)
         );
  OAI22X1TS U3413 ( .A0(n4536), .A1(n668), .B0(n4978), .B1(n3580), .Y(n4979)
         );
  NOR4XLTS U3414 ( .A(n4977), .B(n4976), .C(n4975), .D(n4974), .Y(n4978) );
  OAI22X1TS U3415 ( .A0(n4539), .A1(n3612), .B0(n4537), .B1(n3622), .Y(n4977)
         );
  OAI22X1TS U3416 ( .A0(n4542), .A1(n3654), .B0(n4543), .B1(n6320), .Y(n4976)
         );
  OAI22X1TS U3417 ( .A0(n4545), .A1(n668), .B0(n4986), .B1(n3580), .Y(n4987)
         );
  NOR4XLTS U3418 ( .A(n4985), .B(n4984), .C(n4983), .D(n4982), .Y(n4986) );
  OAI22X1TS U3419 ( .A0(n4548), .A1(n3616), .B0(n4552), .B1(n3622), .Y(n4985)
         );
  OAI22X1TS U3420 ( .A0(n4546), .A1(n3654), .B0(n4553), .B1(n3676), .Y(n4984)
         );
  OAI22X1TS U3421 ( .A0(n4554), .A1(n668), .B0(n4994), .B1(n3579), .Y(n4995)
         );
  NOR4XLTS U3422 ( .A(n4993), .B(n4992), .C(n4991), .D(n4990), .Y(n4994) );
  OAI22X1TS U3423 ( .A0(n4557), .A1(n3618), .B0(n4556), .B1(n3622), .Y(n4993)
         );
  OAI22X1TS U3424 ( .A0(n4555), .A1(n3654), .B0(n4558), .B1(n3677), .Y(n4992)
         );
  OAI22X1TS U3425 ( .A0(n4563), .A1(n668), .B0(n5002), .B1(n3579), .Y(n5003)
         );
  NOR4XLTS U3426 ( .A(n5001), .B(n5000), .C(n4999), .D(n4998), .Y(n5002) );
  OAI22X1TS U3427 ( .A0(n4568), .A1(n3604), .B0(n4570), .B1(n3622), .Y(n5001)
         );
  OAI22X1TS U3428 ( .A0(n4567), .A1(n3660), .B0(n4571), .B1(n3675), .Y(n5000)
         );
  OAI22X1TS U3429 ( .A0(n4572), .A1(n667), .B0(n5010), .B1(n3579), .Y(n5011)
         );
  NOR4XLTS U3430 ( .A(n5009), .B(n5008), .C(n5007), .D(n5006), .Y(n5010) );
  OAI22X1TS U3431 ( .A0(n4575), .A1(n3604), .B0(n4579), .B1(n3621), .Y(n5009)
         );
  OAI22X1TS U3432 ( .A0(n4577), .A1(n3660), .B0(n4578), .B1(n3675), .Y(n5008)
         );
  OAI22X1TS U3433 ( .A0(n4581), .A1(n667), .B0(n5018), .B1(n3579), .Y(n5019)
         );
  NOR4XLTS U3434 ( .A(n5017), .B(n5016), .C(n5015), .D(n5014), .Y(n5018) );
  OAI22X1TS U3435 ( .A0(n4588), .A1(n3604), .B0(n4582), .B1(n3621), .Y(n5017)
         );
  OAI22X1TS U3436 ( .A0(n4585), .A1(n3659), .B0(n4586), .B1(n3678), .Y(n5016)
         );
  OAI22X1TS U3437 ( .A0(n4590), .A1(n667), .B0(n5026), .B1(n3578), .Y(n5027)
         );
  NOR4XLTS U3438 ( .A(n5025), .B(n5024), .C(n5023), .D(n5022), .Y(n5026) );
  OAI22X1TS U3439 ( .A0(n4595), .A1(n3604), .B0(n4594), .B1(n3621), .Y(n5025)
         );
  OAI22X1TS U3440 ( .A0(n4593), .A1(n3662), .B0(n4597), .B1(n3679), .Y(n5024)
         );
  OAI22X1TS U3441 ( .A0(n4599), .A1(n667), .B0(n5034), .B1(n3578), .Y(n5035)
         );
  NOR4XLTS U3442 ( .A(n5033), .B(n5032), .C(n5031), .D(n5030), .Y(n5034) );
  OAI22X1TS U3443 ( .A0(n4600), .A1(n3605), .B0(n4605), .B1(n3621), .Y(n5033)
         );
  OAI22X1TS U3444 ( .A0(n4604), .A1(n3653), .B0(n4607), .B1(n3668), .Y(n5032)
         );
  OAI22X1TS U3445 ( .A0(n4608), .A1(n666), .B0(n5042), .B1(n3578), .Y(n5043)
         );
  NOR4XLTS U3446 ( .A(n5041), .B(n5040), .C(n5039), .D(n5038), .Y(n5042) );
  OAI22X1TS U3447 ( .A0(n4613), .A1(n3605), .B0(n4612), .B1(n3620), .Y(n5041)
         );
  OAI22X1TS U3448 ( .A0(n4611), .A1(n3653), .B0(n4609), .B1(n3668), .Y(n5040)
         );
  OAI22X1TS U3449 ( .A0(n4617), .A1(n666), .B0(n5050), .B1(n3578), .Y(n5051)
         );
  NOR4XLTS U3450 ( .A(n5049), .B(n5048), .C(n5047), .D(n5046), .Y(n5050) );
  OAI22X1TS U3451 ( .A0(n4624), .A1(n3605), .B0(n4622), .B1(n3620), .Y(n5049)
         );
  OAI22X1TS U3452 ( .A0(n4620), .A1(n3653), .B0(n4623), .B1(n3668), .Y(n5048)
         );
  OAI22X1TS U3453 ( .A0(n4626), .A1(n666), .B0(n5058), .B1(n3577), .Y(n5059)
         );
  NOR4XLTS U3454 ( .A(n5057), .B(n5056), .C(n5055), .D(n5054), .Y(n5058) );
  OAI22X1TS U3455 ( .A0(n4633), .A1(n3605), .B0(n4628), .B1(n3620), .Y(n5057)
         );
  OAI22X1TS U3456 ( .A0(n4627), .A1(n3652), .B0(n4634), .B1(n3668), .Y(n5056)
         );
  OAI22X1TS U3457 ( .A0(n4635), .A1(n665), .B0(n5066), .B1(n3577), .Y(n5067)
         );
  NOR4XLTS U3458 ( .A(n5065), .B(n5064), .C(n5063), .D(n5062), .Y(n5066) );
  OAI22X1TS U3459 ( .A0(n4638), .A1(n3606), .B0(n4640), .B1(n3629), .Y(n5065)
         );
  OAI22X1TS U3460 ( .A0(n4642), .A1(n3652), .B0(n4639), .B1(n3669), .Y(n5064)
         );
  OAI22X1TS U3461 ( .A0(n4644), .A1(n665), .B0(n5074), .B1(n3577), .Y(n5075)
         );
  NOR4XLTS U3462 ( .A(n5073), .B(n5072), .C(n5071), .D(n5070), .Y(n5074) );
  OAI22X1TS U3463 ( .A0(n4647), .A1(n3606), .B0(n4650), .B1(n3629), .Y(n5073)
         );
  OAI22X1TS U3464 ( .A0(n4649), .A1(n3652), .B0(n4645), .B1(n3669), .Y(n5072)
         );
  OAI22X1TS U3465 ( .A0(n4653), .A1(n665), .B0(n5082), .B1(n3576), .Y(n5083)
         );
  NOR4XLTS U3466 ( .A(n5081), .B(n5080), .C(n5079), .D(n5078), .Y(n5082) );
  OAI22X1TS U3467 ( .A0(n4660), .A1(n3606), .B0(n4656), .B1(n3633), .Y(n5081)
         );
  OAI22X1TS U3468 ( .A0(n4659), .A1(n3652), .B0(n4657), .B1(n3669), .Y(n5080)
         );
  OAI22X1TS U3469 ( .A0(n4662), .A1(n665), .B0(n5090), .B1(n3576), .Y(n5091)
         );
  NOR4XLTS U3470 ( .A(n5089), .B(n5088), .C(n5087), .D(n5086), .Y(n5090) );
  OAI22X1TS U3471 ( .A0(n4663), .A1(n3606), .B0(n4667), .B1(n3630), .Y(n5089)
         );
  OAI22X1TS U3472 ( .A0(n4666), .A1(n3651), .B0(n4669), .B1(n3669), .Y(n5088)
         );
  OAI22X1TS U3473 ( .A0(n4671), .A1(n664), .B0(n5098), .B1(n3576), .Y(n5099)
         );
  NOR4XLTS U3474 ( .A(n5097), .B(n5096), .C(n5095), .D(n5094), .Y(n5098) );
  OAI22X1TS U3475 ( .A0(n4674), .A1(n3607), .B0(n4678), .B1(n3630), .Y(n5097)
         );
  OAI22X1TS U3476 ( .A0(n4676), .A1(n3651), .B0(n4673), .B1(n3670), .Y(n5096)
         );
  OAI22X1TS U3477 ( .A0(n4680), .A1(n664), .B0(n5106), .B1(n3576), .Y(n5107)
         );
  NOR4XLTS U3478 ( .A(n5105), .B(n5104), .C(n5103), .D(n5102), .Y(n5106) );
  OAI22X1TS U3479 ( .A0(n4687), .A1(n3607), .B0(n4683), .B1(n3631), .Y(n5105)
         );
  OAI22X1TS U3480 ( .A0(n4686), .A1(n3651), .B0(n4688), .B1(n3670), .Y(n5104)
         );
  OAI22X1TS U3481 ( .A0(n4689), .A1(n664), .B0(n5114), .B1(n3575), .Y(n5115)
         );
  NOR4XLTS U3482 ( .A(n5113), .B(n5112), .C(n5111), .D(n5110), .Y(n5114) );
  OAI22X1TS U3483 ( .A0(n4696), .A1(n3607), .B0(n4691), .B1(n3631), .Y(n5113)
         );
  OAI22X1TS U3484 ( .A0(n4690), .A1(n3651), .B0(n4692), .B1(n3670), .Y(n5112)
         );
  OAI22X1TS U3485 ( .A0(n4698), .A1(n664), .B0(n5122), .B1(n3575), .Y(n5123)
         );
  NOR4XLTS U3486 ( .A(n5121), .B(n5120), .C(n5119), .D(n5118), .Y(n5122) );
  OAI22X1TS U3487 ( .A0(n4703), .A1(n3607), .B0(n4702), .B1(n6318), .Y(n5121)
         );
  OAI22X1TS U3488 ( .A0(n4699), .A1(n3664), .B0(n4704), .B1(n3670), .Y(n5120)
         );
  OAI22X1TS U3489 ( .A0(n4711), .A1(n663), .B0(n5178), .B1(n3573), .Y(n5179)
         );
  NOR4XLTS U3490 ( .A(n5177), .B(n5176), .C(n5175), .D(n5174), .Y(n5178) );
  OAI22X1TS U3491 ( .A0(n4712), .A1(n3608), .B0(n4714), .B1(n3634), .Y(n5177)
         );
  OAI22X1TS U3492 ( .A0(n4718), .A1(n3664), .B0(n4716), .B1(n3671), .Y(n5176)
         );
  OAI22X1TS U3493 ( .A0(n4720), .A1(n663), .B0(n5186), .B1(n3573), .Y(n5187)
         );
  NOR4XLTS U3494 ( .A(n5185), .B(n5184), .C(n5183), .D(n5182), .Y(n5186) );
  OAI22X1TS U3495 ( .A0(n4724), .A1(n3608), .B0(n4725), .B1(n3634), .Y(n5185)
         );
  OAI22X1TS U3496 ( .A0(n4723), .A1(n3661), .B0(n4727), .B1(n3671), .Y(n5184)
         );
  OAI22X1TS U3497 ( .A0(n4729), .A1(n666), .B0(n5194), .B1(n3573), .Y(n5195)
         );
  NOR4XLTS U3498 ( .A(n5193), .B(n5192), .C(n5191), .D(n5190), .Y(n5194) );
  OAI22X1TS U3499 ( .A0(n4732), .A1(n3608), .B0(n4734), .B1(n3634), .Y(n5193)
         );
  OAI22X1TS U3500 ( .A0(n4736), .A1(n3662), .B0(n4730), .B1(n3671), .Y(n5192)
         );
  OAI22X1TS U3501 ( .A0(n4738), .A1(n663), .B0(n5202), .B1(n3573), .Y(n5203)
         );
  NOR4XLTS U3502 ( .A(n5201), .B(n5200), .C(n5199), .D(n5198), .Y(n5202) );
  OAI22X1TS U3503 ( .A0(n4743), .A1(n3608), .B0(n4739), .B1(n3628), .Y(n5201)
         );
  OAI22X1TS U3504 ( .A0(n4740), .A1(n3663), .B0(n4741), .B1(n3671), .Y(n5200)
         );
  OAI22X1TS U3505 ( .A0(n4747), .A1(n662), .B0(n5210), .B1(n3572), .Y(n5211)
         );
  NOR4XLTS U3506 ( .A(n5209), .B(n5208), .C(n5207), .D(n5206), .Y(n5210) );
  OAI22X1TS U3507 ( .A0(n4748), .A1(n3609), .B0(n4752), .B1(n3628), .Y(n5209)
         );
  OAI22X1TS U3508 ( .A0(n4754), .A1(n3664), .B0(n4750), .B1(n3672), .Y(n5208)
         );
  OAI22X1TS U3509 ( .A0(n4756), .A1(n663), .B0(n5219), .B1(n3572), .Y(n5220)
         );
  NOR4XLTS U3510 ( .A(n5218), .B(n5217), .C(n5216), .D(n5215), .Y(n5219) );
  OAI22X1TS U3511 ( .A0(n4762), .A1(n3609), .B0(n4757), .B1(n3632), .Y(n5218)
         );
  OAI22X1TS U3512 ( .A0(n4761), .A1(n3663), .B0(n4759), .B1(n3672), .Y(n5217)
         );
  OAI221XLTS U3513 ( .A0(n5307), .A1(n5306), .B0(n5305), .B1(n5304), .C0(n4418), .Y(n5308) );
  OAI211X1TS U3514 ( .A0(n3603), .A1(n16), .B0(n4830), .C0(n5298), .Y(n5306)
         );
  OAI221XLTS U3515 ( .A0(n3611), .A1(n6312), .B0(n3674), .B1(n18), .C0(n5296), 
        .Y(n5307) );
  OAI211X1TS U3516 ( .A0(n282), .A1(n514), .B0(n5229), .C0(n5228), .Y(n2441)
         );
  AOI22X1TS U3517 ( .A0(n461), .A1(n5227), .B0(n673), .B1(
        destinationAddressOut[13]), .Y(n5229) );
  AOI222XLTS U3518 ( .A0(n391), .A1(n4284), .B0(n566), .B1(n4128), .C0(n554), 
        .C1(destinationAddressIn_WEST[13]), .Y(n5228) );
  NAND4X1TS U3519 ( .A(n5226), .B(n5225), .C(n5224), .D(n5223), .Y(n5227) );
  OAI211X1TS U3520 ( .A0(n273), .A1(n514), .B0(n5236), .C0(n5235), .Y(n2442)
         );
  AOI22X1TS U3521 ( .A0(n462), .A1(n5234), .B0(n673), .B1(
        destinationAddressOut[12]), .Y(n5236) );
  AOI222XLTS U3522 ( .A0(n390), .A1(n4281), .B0(n566), .B1(n4125), .C0(n561), 
        .C1(destinationAddressIn_WEST[12]), .Y(n5235) );
  NAND4X1TS U3523 ( .A(n5233), .B(n5232), .C(n5231), .D(n5230), .Y(n5234) );
  OAI211X1TS U3524 ( .A0(n285), .A1(n514), .B0(n5243), .C0(n5242), .Y(n2443)
         );
  AOI22X1TS U3525 ( .A0(n462), .A1(n5241), .B0(n673), .B1(
        destinationAddressOut[11]), .Y(n5243) );
  AOI222XLTS U3526 ( .A0(n391), .A1(n4278), .B0(n566), .B1(n4122), .C0(n557), 
        .C1(destinationAddressIn_WEST[11]), .Y(n5242) );
  NAND4X1TS U3527 ( .A(n5240), .B(n5239), .C(n5238), .D(n5237), .Y(n5241) );
  OAI211X1TS U3528 ( .A0(n276), .A1(n516), .B0(n5250), .C0(n5249), .Y(n2444)
         );
  AOI22X1TS U3529 ( .A0(n461), .A1(n5248), .B0(n673), .B1(
        destinationAddressOut[10]), .Y(n5250) );
  AOI222XLTS U3530 ( .A0(n390), .A1(n4275), .B0(n566), .B1(n4119), .C0(n556), 
        .C1(destinationAddressIn_WEST[10]), .Y(n5249) );
  NAND4X1TS U3531 ( .A(n5247), .B(n5246), .C(n5245), .D(n5244), .Y(n5248) );
  OAI211X1TS U3532 ( .A0(n279), .A1(n516), .B0(n5257), .C0(n5256), .Y(n2445)
         );
  AOI22X1TS U3533 ( .A0(n462), .A1(n5255), .B0(n674), .B1(
        destinationAddressOut[9]), .Y(n5257) );
  AOI222XLTS U3534 ( .A0(n391), .A1(n4272), .B0(n565), .B1(n4116), .C0(n564), 
        .C1(destinationAddressIn_WEST[9]), .Y(n5256) );
  NAND4X1TS U3535 ( .A(n5254), .B(n5253), .C(n5252), .D(n5251), .Y(n5255) );
  OAI211X1TS U3536 ( .A0(n288), .A1(n516), .B0(n5264), .C0(n5263), .Y(n2446)
         );
  AOI22X1TS U3537 ( .A0(n461), .A1(n5262), .B0(n674), .B1(
        destinationAddressOut[8]), .Y(n5264) );
  AOI222XLTS U3538 ( .A0(n390), .A1(n4269), .B0(n565), .B1(n4113), .C0(n563), 
        .C1(destinationAddressIn_WEST[8]), .Y(n5263) );
  NAND4X1TS U3539 ( .A(n5261), .B(n5260), .C(n5259), .D(n5258), .Y(n5262) );
  OAI211X1TS U3540 ( .A0(n270), .A1(n517), .B0(n5271), .C0(n5270), .Y(n2447)
         );
  AOI22X1TS U3541 ( .A0(n461), .A1(n5269), .B0(n674), .B1(
        destinationAddressOut[7]), .Y(n5271) );
  AOI222XLTS U3542 ( .A0(n391), .A1(n4266), .B0(n565), .B1(n4110), .C0(n562), 
        .C1(destinationAddressIn_WEST[7]), .Y(n5270) );
  NAND4X1TS U3543 ( .A(n5268), .B(n5267), .C(n5266), .D(n5265), .Y(n5269) );
  OAI211X1TS U3544 ( .A0(n267), .A1(n517), .B0(n5281), .C0(n5280), .Y(n2448)
         );
  AOI22X1TS U3545 ( .A0(n462), .A1(n5276), .B0(n674), .B1(
        destinationAddressOut[6]), .Y(n5281) );
  AOI222XLTS U3546 ( .A0(n390), .A1(n4263), .B0(n565), .B1(n4107), .C0(n555), 
        .C1(destinationAddressIn_WEST[6]), .Y(n5280) );
  NAND4X1TS U3547 ( .A(n5275), .B(n5274), .C(n5273), .D(n5272), .Y(n5276) );
  OAI211X1TS U3548 ( .A0(n4225), .A1(n3569), .B0(n4877), .C0(n4876), .Y(n2397)
         );
  AOI22X1TS U3549 ( .A0(n494), .A1(n398), .B0(n562), .B1(n3911), .Y(n4877) );
  AOI221X1TS U3550 ( .A0(n496), .A1(n4379), .B0(n579), .B1(n4068), .C0(n4875), 
        .Y(n4876) );
  OAI211X1TS U3551 ( .A0(n4222), .A1(n3568), .B0(n4885), .C0(n4884), .Y(n2398)
         );
  AOI22X1TS U3552 ( .A0(n493), .A1(n400), .B0(n562), .B1(n3908), .Y(n4885) );
  AOI221X1TS U3553 ( .A0(n496), .A1(n4376), .B0(n577), .B1(n4065), .C0(n4883), 
        .Y(n4884) );
  OAI211X1TS U3554 ( .A0(n4219), .A1(n3570), .B0(n4893), .C0(n4892), .Y(n2399)
         );
  AOI22X1TS U3555 ( .A0(n494), .A1(n402), .B0(n562), .B1(n3905), .Y(n4893) );
  AOI221X1TS U3556 ( .A0(n496), .A1(n4373), .B0(n577), .B1(n4062), .C0(n4891), 
        .Y(n4892) );
  OAI211X1TS U3557 ( .A0(n4216), .A1(n3571), .B0(n4901), .C0(n4900), .Y(n2400)
         );
  AOI22X1TS U3558 ( .A0(n493), .A1(n404), .B0(n5277), .B1(n3902), .Y(n4901) );
  AOI221X1TS U3559 ( .A0(n496), .A1(n4370), .B0(n5278), .B1(n4059), .C0(n4899), 
        .Y(n4900) );
  OAI211X1TS U3560 ( .A0(n4213), .A1(n3558), .B0(n4909), .C0(n4908), .Y(n2401)
         );
  AOI22X1TS U3561 ( .A0(n482), .A1(n406), .B0(n537), .B1(n3899), .Y(n4909) );
  AOI221X1TS U3562 ( .A0(n500), .A1(n4367), .B0(n5278), .B1(n4056), .C0(n4907), 
        .Y(n4908) );
  OAI211X1TS U3563 ( .A0(n4210), .A1(n3558), .B0(n4917), .C0(n4916), .Y(n2402)
         );
  AOI22X1TS U3564 ( .A0(n482), .A1(n408), .B0(n537), .B1(n3896), .Y(n4917) );
  AOI221X1TS U3565 ( .A0(n500), .A1(n4364), .B0(n578), .B1(n4053), .C0(n4915), 
        .Y(n4916) );
  OAI211X1TS U3566 ( .A0(n4207), .A1(n3558), .B0(n4925), .C0(n4924), .Y(n2403)
         );
  AOI22X1TS U3567 ( .A0(n482), .A1(n410), .B0(n537), .B1(n3893), .Y(n4925) );
  AOI221X1TS U3568 ( .A0(n500), .A1(n4361), .B0(n579), .B1(n4050), .C0(n4923), 
        .Y(n4924) );
  OAI211X1TS U3569 ( .A0(n4204), .A1(n3558), .B0(n4933), .C0(n4932), .Y(n2404)
         );
  AOI22X1TS U3570 ( .A0(n482), .A1(n412), .B0(n537), .B1(n3890), .Y(n4933) );
  AOI221X1TS U3571 ( .A0(n500), .A1(n4358), .B0(n580), .B1(n4047), .C0(n4931), 
        .Y(n4932) );
  OAI211X1TS U3572 ( .A0(n4201), .A1(n3567), .B0(n4941), .C0(n4940), .Y(n2405)
         );
  AOI22X1TS U3573 ( .A0(n483), .A1(n414), .B0(n541), .B1(n3887), .Y(n4941) );
  AOI221X1TS U3574 ( .A0(n501), .A1(n4355), .B0(n575), .B1(n4044), .C0(n4939), 
        .Y(n4940) );
  OAI211X1TS U3575 ( .A0(n4198), .A1(n3566), .B0(n4949), .C0(n4948), .Y(n2406)
         );
  AOI22X1TS U3576 ( .A0(n483), .A1(n416), .B0(n541), .B1(n3884), .Y(n4949) );
  AOI221X1TS U3577 ( .A0(n501), .A1(n4352), .B0(n576), .B1(n4041), .C0(n4947), 
        .Y(n4948) );
  OAI211X1TS U3578 ( .A0(n4195), .A1(n3565), .B0(n4957), .C0(n4956), .Y(n2407)
         );
  AOI22X1TS U3579 ( .A0(n483), .A1(n418), .B0(n541), .B1(n3881), .Y(n4957) );
  AOI221X1TS U3580 ( .A0(n501), .A1(n4349), .B0(n579), .B1(n4038), .C0(n4955), 
        .Y(n4956) );
  OAI211X1TS U3581 ( .A0(n4192), .A1(n3569), .B0(n4965), .C0(n4964), .Y(n2408)
         );
  AOI22X1TS U3582 ( .A0(n483), .A1(n420), .B0(n541), .B1(n3878), .Y(n4965) );
  AOI221X1TS U3583 ( .A0(n501), .A1(n4346), .B0(n575), .B1(n4035), .C0(n4963), 
        .Y(n4964) );
  OAI211X1TS U3584 ( .A0(n4189), .A1(n3568), .B0(n4973), .C0(n4972), .Y(n2409)
         );
  AOI22X1TS U3585 ( .A0(n484), .A1(n422), .B0(n561), .B1(n3875), .Y(n4973) );
  AOI221X1TS U3586 ( .A0(n502), .A1(n4343), .B0(n574), .B1(n4032), .C0(n4971), 
        .Y(n4972) );
  OAI211X1TS U3587 ( .A0(n4186), .A1(n3568), .B0(n4981), .C0(n4980), .Y(n2410)
         );
  AOI22X1TS U3588 ( .A0(n484), .A1(n424), .B0(n556), .B1(n3872), .Y(n4981) );
  AOI221X1TS U3589 ( .A0(n502), .A1(n4340), .B0(n574), .B1(n4029), .C0(n4979), 
        .Y(n4980) );
  OAI211X1TS U3590 ( .A0(n4183), .A1(n3569), .B0(n4989), .C0(n4988), .Y(n2411)
         );
  AOI22X1TS U3591 ( .A0(n484), .A1(n426), .B0(n557), .B1(n3869), .Y(n4989) );
  AOI221X1TS U3592 ( .A0(n502), .A1(n4337), .B0(n574), .B1(n4026), .C0(n4987), 
        .Y(n4988) );
  OAI211X1TS U3593 ( .A0(n4180), .A1(n3570), .B0(n4997), .C0(n4996), .Y(n2412)
         );
  AOI22X1TS U3594 ( .A0(n484), .A1(n428), .B0(n5277), .B1(n3866), .Y(n4997) );
  AOI221X1TS U3595 ( .A0(n502), .A1(n4334), .B0(n574), .B1(n4023), .C0(n4995), 
        .Y(n4996) );
  OAI211X1TS U3596 ( .A0(n4177), .A1(n3568), .B0(n5005), .C0(n5004), .Y(n2413)
         );
  AOI22X1TS U3597 ( .A0(n485), .A1(n430), .B0(n557), .B1(n3863), .Y(n5005) );
  AOI221X1TS U3598 ( .A0(n503), .A1(n4331), .B0(n573), .B1(n4020), .C0(n5003), 
        .Y(n5004) );
  OAI211X1TS U3599 ( .A0(n4174), .A1(n3567), .B0(n5013), .C0(n5012), .Y(n2414)
         );
  AOI22X1TS U3600 ( .A0(n485), .A1(n432), .B0(n557), .B1(n3860), .Y(n5013) );
  AOI221X1TS U3601 ( .A0(n503), .A1(n4328), .B0(n573), .B1(n4017), .C0(n5011), 
        .Y(n5012) );
  OAI211X1TS U3602 ( .A0(n4171), .A1(n3566), .B0(n5021), .C0(n5020), .Y(n2415)
         );
  AOI22X1TS U3603 ( .A0(n485), .A1(n434), .B0(n555), .B1(n3857), .Y(n5021) );
  AOI221X1TS U3604 ( .A0(n503), .A1(n4325), .B0(n573), .B1(n4014), .C0(n5019), 
        .Y(n5020) );
  OAI211X1TS U3605 ( .A0(n4168), .A1(n3565), .B0(n5029), .C0(n5028), .Y(n2416)
         );
  AOI22X1TS U3606 ( .A0(n485), .A1(n436), .B0(n554), .B1(n3854), .Y(n5029) );
  AOI221X1TS U3607 ( .A0(n503), .A1(n4322), .B0(n573), .B1(n4011), .C0(n5027), 
        .Y(n5028) );
  OAI211X1TS U3608 ( .A0(n4165), .A1(n3559), .B0(n5037), .C0(n5036), .Y(n2417)
         );
  AOI22X1TS U3609 ( .A0(n494), .A1(n438), .B0(n543), .B1(n3851), .Y(n5037) );
  AOI221X1TS U3610 ( .A0(n504), .A1(n4319), .B0(n572), .B1(n4008), .C0(n5035), 
        .Y(n5036) );
  OAI211X1TS U3611 ( .A0(n4162), .A1(n3559), .B0(n5045), .C0(n5044), .Y(n2418)
         );
  AOI22X1TS U3612 ( .A0(n491), .A1(n440), .B0(n543), .B1(n3848), .Y(n5045) );
  AOI221X1TS U3613 ( .A0(n504), .A1(n4316), .B0(n572), .B1(n4005), .C0(n5043), 
        .Y(n5044) );
  OAI211X1TS U3614 ( .A0(n4159), .A1(n3559), .B0(n5053), .C0(n5052), .Y(n2419)
         );
  AOI22X1TS U3615 ( .A0(n495), .A1(n442), .B0(n543), .B1(n3845), .Y(n5053) );
  AOI221X1TS U3616 ( .A0(n504), .A1(n4313), .B0(n572), .B1(n4002), .C0(n5051), 
        .Y(n5052) );
  OAI211X1TS U3617 ( .A0(n4156), .A1(n3559), .B0(n5061), .C0(n5060), .Y(n2420)
         );
  AOI22X1TS U3618 ( .A0(n492), .A1(n444), .B0(n543), .B1(n3842), .Y(n5061) );
  AOI221X1TS U3619 ( .A0(n504), .A1(n4310), .B0(n572), .B1(n3999), .C0(n5059), 
        .Y(n5060) );
  OAI211X1TS U3620 ( .A0(n4153), .A1(n3560), .B0(n5069), .C0(n5068), .Y(n2421)
         );
  AOI22X1TS U3621 ( .A0(n486), .A1(n446), .B0(n544), .B1(n3839), .Y(n5069) );
  AOI221X1TS U3622 ( .A0(n505), .A1(n4307), .B0(n571), .B1(n3996), .C0(n5067), 
        .Y(n5068) );
  OAI211X1TS U3623 ( .A0(n4150), .A1(n3560), .B0(n5077), .C0(n5076), .Y(n2422)
         );
  AOI22X1TS U3624 ( .A0(n486), .A1(n448), .B0(n544), .B1(n3836), .Y(n5077) );
  AOI221X1TS U3625 ( .A0(n505), .A1(n4304), .B0(n571), .B1(n3993), .C0(n5075), 
        .Y(n5076) );
  OAI211X1TS U3626 ( .A0(n4147), .A1(n3560), .B0(n5085), .C0(n5084), .Y(n2423)
         );
  AOI22X1TS U3627 ( .A0(n486), .A1(n450), .B0(n544), .B1(n3833), .Y(n5085) );
  AOI221X1TS U3628 ( .A0(n505), .A1(n4301), .B0(n571), .B1(n3990), .C0(n5083), 
        .Y(n5084) );
  OAI211X1TS U3629 ( .A0(n4144), .A1(n3560), .B0(n5093), .C0(n5092), .Y(n2424)
         );
  AOI22X1TS U3630 ( .A0(n486), .A1(n452), .B0(n544), .B1(n3830), .Y(n5093) );
  AOI221X1TS U3631 ( .A0(n505), .A1(n4298), .B0(n571), .B1(n3987), .C0(n5091), 
        .Y(n5092) );
  OAI211X1TS U3632 ( .A0(n4141), .A1(n3561), .B0(n5101), .C0(n5100), .Y(n2425)
         );
  AOI22X1TS U3633 ( .A0(n487), .A1(n454), .B0(n545), .B1(n3827), .Y(n5101) );
  AOI221X1TS U3634 ( .A0(n507), .A1(n4295), .B0(n570), .B1(n3984), .C0(n5099), 
        .Y(n5100) );
  OAI211X1TS U3635 ( .A0(n4138), .A1(n3561), .B0(n5109), .C0(n5108), .Y(n2426)
         );
  AOI22X1TS U3636 ( .A0(n487), .A1(n456), .B0(n545), .B1(n3824), .Y(n5109) );
  AOI221X1TS U3637 ( .A0(n507), .A1(n4292), .B0(n570), .B1(n3981), .C0(n5107), 
        .Y(n5108) );
  OAI211X1TS U3638 ( .A0(n4135), .A1(n3561), .B0(n5117), .C0(n5116), .Y(n2427)
         );
  AOI22X1TS U3639 ( .A0(n487), .A1(n458), .B0(n545), .B1(n3821), .Y(n5117) );
  AOI221X1TS U3640 ( .A0(n507), .A1(n4289), .B0(n570), .B1(n3978), .C0(n5115), 
        .Y(n5116) );
  OAI211X1TS U3641 ( .A0(n4132), .A1(n3561), .B0(n5125), .C0(n5124), .Y(n2428)
         );
  AOI22X1TS U3642 ( .A0(n487), .A1(n460), .B0(n545), .B1(n3818), .Y(n5125) );
  AOI221X1TS U3643 ( .A0(n507), .A1(n4286), .B0(n570), .B1(n3975), .C0(n5123), 
        .Y(n5124) );
  OAI211X1TS U3644 ( .A0(n4243), .A1(n3562), .B0(n5133), .C0(n5132), .Y(n2429)
         );
  AOI22X1TS U3645 ( .A0(n488), .A1(n162), .B0(n546), .B1(n3929), .Y(n5133) );
  AOI221X1TS U3646 ( .A0(n508), .A1(n4397), .B0(n569), .B1(n4086), .C0(n5131), 
        .Y(n5132) );
  OAI211X1TS U3647 ( .A0(n4240), .A1(n3562), .B0(n5141), .C0(n5140), .Y(n2430)
         );
  AOI22X1TS U3648 ( .A0(n488), .A1(n156), .B0(n546), .B1(n3926), .Y(n5141) );
  AOI221X1TS U3649 ( .A0(n508), .A1(n4394), .B0(n569), .B1(n4083), .C0(n5139), 
        .Y(n5140) );
  OAI211X1TS U3650 ( .A0(n4234), .A1(n3562), .B0(n5157), .C0(n5156), .Y(n2432)
         );
  AOI22X1TS U3651 ( .A0(n488), .A1(n146), .B0(n546), .B1(n3920), .Y(n5157) );
  AOI221X1TS U3652 ( .A0(n508), .A1(n4388), .B0(n569), .B1(n4077), .C0(n5155), 
        .Y(n5156) );
  OAI211X1TS U3653 ( .A0(n4231), .A1(n3563), .B0(n5165), .C0(n5164), .Y(n2433)
         );
  AOI22X1TS U3654 ( .A0(n489), .A1(n141), .B0(n548), .B1(n3917), .Y(n5165) );
  AOI221X1TS U3655 ( .A0(n509), .A1(n4385), .B0(n568), .B1(n4074), .C0(n5163), 
        .Y(n5164) );
  OAI211X1TS U3656 ( .A0(n4261), .A1(n3563), .B0(n5181), .C0(n5180), .Y(n2435)
         );
  AOI22X1TS U3657 ( .A0(n489), .A1(n161), .B0(n548), .B1(n3947), .Y(n5181) );
  AOI221X1TS U3658 ( .A0(n509), .A1(n4415), .B0(n568), .B1(n4104), .C0(n5179), 
        .Y(n5180) );
  OAI211X1TS U3659 ( .A0(n4258), .A1(n3563), .B0(n5189), .C0(n5188), .Y(n2436)
         );
  AOI22X1TS U3660 ( .A0(n489), .A1(n157), .B0(n548), .B1(n3944), .Y(n5189) );
  AOI221X1TS U3661 ( .A0(n509), .A1(n4412), .B0(n568), .B1(n4101), .C0(n5187), 
        .Y(n5188) );
  OAI211X1TS U3662 ( .A0(n4255), .A1(n3564), .B0(n5197), .C0(n5196), .Y(n2437)
         );
  AOI22X1TS U3663 ( .A0(n490), .A1(n151), .B0(n551), .B1(n3941), .Y(n5197) );
  AOI221X1TS U3664 ( .A0(n511), .A1(n4409), .B0(n567), .B1(n4098), .C0(n5195), 
        .Y(n5196) );
  OAI211X1TS U3665 ( .A0(n4252), .A1(n3564), .B0(n5205), .C0(n5204), .Y(n2438)
         );
  AOI22X1TS U3666 ( .A0(n490), .A1(n147), .B0(n551), .B1(n3938), .Y(n5205) );
  AOI221X1TS U3667 ( .A0(n511), .A1(n4406), .B0(n567), .B1(n4095), .C0(n5203), 
        .Y(n5204) );
  OAI211X1TS U3668 ( .A0(n4249), .A1(n3564), .B0(n5213), .C0(n5212), .Y(n2439)
         );
  AOI22X1TS U3669 ( .A0(n490), .A1(n142), .B0(n551), .B1(n3935), .Y(n5213) );
  AOI221X1TS U3670 ( .A0(n511), .A1(n4403), .B0(n567), .B1(n4092), .C0(n5211), 
        .Y(n5212) );
  OAI211X1TS U3671 ( .A0(n4246), .A1(n3564), .B0(n5222), .C0(n5221), .Y(n2440)
         );
  AOI22X1TS U3672 ( .A0(n490), .A1(n137), .B0(n551), .B1(n3932), .Y(n5222) );
  AOI221X1TS U3673 ( .A0(n511), .A1(n4400), .B0(n567), .B1(n4089), .C0(n5220), 
        .Y(n5221) );
  OAI211X1TS U3674 ( .A0(n4237), .A1(n3562), .B0(n5149), .C0(n5148), .Y(n2431)
         );
  AOI22X1TS U3675 ( .A0(n488), .A1(n152), .B0(n546), .B1(n3923), .Y(n5149) );
  AOI221X1TS U3676 ( .A0(n508), .A1(n4391), .B0(n569), .B1(n4080), .C0(n5147), 
        .Y(n5148) );
  OAI211X1TS U3677 ( .A0(n4228), .A1(n3563), .B0(n5173), .C0(n5172), .Y(n2434)
         );
  AOI22X1TS U3678 ( .A0(n489), .A1(n138), .B0(n548), .B1(n3914), .Y(n5173) );
  AOI221X1TS U3679 ( .A0(n509), .A1(n4382), .B0(n568), .B1(n4071), .C0(n5171), 
        .Y(n5172) );
  NOR2X1TS U3680 ( .A(reset), .B(n4830), .Y(n5291) );
  INVX2TS U3681 ( .A(readIn_SOUTH), .Y(n6233) );
  INVX2TS U3682 ( .A(writeIn_NORTH), .Y(n6235) );
  OAI22X1TS U3683 ( .A0(n5292), .A1(n5291), .B0(n5290), .B1(n5289), .Y(n5293)
         );
  AOI31X1TS U3684 ( .A0(n5288), .A1(n5287), .A2(n5286), .B0(reset), .Y(n5292)
         );
  OAI22X1TS U3685 ( .A0(n3814), .A1(n5301), .B0(n3801), .B1(n5303), .Y(n5289)
         );
  OAI22X1TS U3686 ( .A0(n395), .A1(n6316), .B0(n4), .B1(n3577), .Y(n2889) );
  INVX2TS U3687 ( .A(destinationAddressIn_NORTH[6]), .Y(n6236) );
  INVX2TS U3688 ( .A(destinationAddressIn_NORTH[7]), .Y(n6237) );
  INVX2TS U3689 ( .A(destinationAddressIn_NORTH[12]), .Y(n6242) );
  INVX2TS U3690 ( .A(destinationAddressIn_NORTH[10]), .Y(n6240) );
  INVX2TS U3691 ( .A(destinationAddressIn_NORTH[9]), .Y(n6239) );
  INVX2TS U3692 ( .A(destinationAddressIn_NORTH[13]), .Y(n6243) );
  INVX2TS U3693 ( .A(destinationAddressIn_NORTH[11]), .Y(n6241) );
  INVX2TS U3694 ( .A(destinationAddressIn_NORTH[8]), .Y(n6238) );
  NOR2X1TS U3695 ( .A(n6218), .B(n6219), .Y(n2883) );
  AOI21X1TS U3696 ( .A0(n301), .A1(n6217), .B0(n5), .Y(n6218) );
  XNOR2X1TS U3697 ( .A(n4840), .B(n6322), .Y(n6222) );
  XNOR2X1TS U3698 ( .A(n217), .B(n218), .Y(n4840) );
  OAI22X1TS U3699 ( .A0(n4426), .A1(n3694), .B0(n4427), .B1(n3592), .Y(n4870)
         );
  OAI22X1TS U3700 ( .A0(n4431), .A1(n3689), .B0(n4436), .B1(n3601), .Y(n4878)
         );
  OAI22X1TS U3701 ( .A0(n4438), .A1(n3693), .B0(n4441), .B1(n3599), .Y(n4886)
         );
  OAI22X1TS U3702 ( .A0(n4449), .A1(n3691), .B0(n4448), .B1(n6317), .Y(n4894)
         );
  OAI22X1TS U3703 ( .A0(n4463), .A1(n3691), .B0(n4456), .B1(n3600), .Y(n4902)
         );
  OAI22X1TS U3704 ( .A0(n4467), .A1(n3693), .B0(n4472), .B1(n3595), .Y(n4910)
         );
  OAI22X1TS U3705 ( .A0(n4474), .A1(n3692), .B0(n4479), .B1(n3595), .Y(n4918)
         );
  OAI22X1TS U3706 ( .A0(n4489), .A1(n3689), .B0(n4484), .B1(n3595), .Y(n4926)
         );
  OAI22X1TS U3707 ( .A0(n4496), .A1(n3690), .B0(n4493), .B1(n3595), .Y(n4934)
         );
  OAI22X1TS U3708 ( .A0(n4507), .A1(n3690), .B0(n4505), .B1(n3598), .Y(n4942)
         );
  OAI22X1TS U3709 ( .A0(n4510), .A1(n3692), .B0(n4511), .B1(n3598), .Y(n4950)
         );
  OAI22X1TS U3710 ( .A0(n4523), .A1(n3695), .B0(n4521), .B1(n3603), .Y(n4958)
         );
  OAI22X1TS U3711 ( .A0(n4528), .A1(n3681), .B0(n4532), .B1(n3601), .Y(n4966)
         );
  OAI22X1TS U3712 ( .A0(n4541), .A1(n3681), .B0(n4544), .B1(n3594), .Y(n4974)
         );
  OAI22X1TS U3713 ( .A0(n4550), .A1(n3681), .B0(n4547), .B1(n3594), .Y(n4982)
         );
  OAI22X1TS U3714 ( .A0(n4561), .A1(n3681), .B0(n4562), .B1(n3594), .Y(n4990)
         );
  OAI22X1TS U3715 ( .A0(n4566), .A1(n3682), .B0(n4569), .B1(n3594), .Y(n4998)
         );
  OAI22X1TS U3716 ( .A0(n4573), .A1(n3682), .B0(n4576), .B1(n3593), .Y(n5006)
         );
  OAI22X1TS U3717 ( .A0(n4584), .A1(n3682), .B0(n4589), .B1(n3593), .Y(n5014)
         );
  OAI22X1TS U3718 ( .A0(n4591), .A1(n3682), .B0(n4598), .B1(n3593), .Y(n5022)
         );
  OAI22X1TS U3719 ( .A0(n4606), .A1(n3683), .B0(n4601), .B1(n3593), .Y(n5030)
         );
  OAI22X1TS U3720 ( .A0(n4614), .A1(n3683), .B0(n4615), .B1(n3592), .Y(n5038)
         );
  OAI22X1TS U3721 ( .A0(n4618), .A1(n3683), .B0(n4619), .B1(n3592), .Y(n5046)
         );
  OAI22X1TS U3722 ( .A0(n4631), .A1(n3683), .B0(n4629), .B1(n3592), .Y(n5054)
         );
  OAI22X1TS U3723 ( .A0(n4636), .A1(n3684), .B0(n4643), .B1(n3591), .Y(n5062)
         );
  OAI22X1TS U3724 ( .A0(n4651), .A1(n3684), .B0(n4646), .B1(n3591), .Y(n5070)
         );
  OAI22X1TS U3725 ( .A0(n4658), .A1(n3684), .B0(n4654), .B1(n3591), .Y(n5078)
         );
  OAI22X1TS U3726 ( .A0(n4665), .A1(n3684), .B0(n4670), .B1(n3591), .Y(n5086)
         );
  OAI22X1TS U3727 ( .A0(n4672), .A1(n3685), .B0(n4675), .B1(n3590), .Y(n5094)
         );
  OAI22X1TS U3728 ( .A0(n4685), .A1(n3685), .B0(n4681), .B1(n3590), .Y(n5102)
         );
  OAI22X1TS U3729 ( .A0(n4697), .A1(n3685), .B0(n4693), .B1(n3590), .Y(n5110)
         );
  OAI22X1TS U3730 ( .A0(n4701), .A1(n3685), .B0(n4705), .B1(n3590), .Y(n5118)
         );
  OAI22X1TS U3731 ( .A0(n4715), .A1(n3686), .B0(n4713), .B1(n3589), .Y(n5174)
         );
  OAI22X1TS U3732 ( .A0(n4728), .A1(n3686), .B0(n4722), .B1(n3589), .Y(n5182)
         );
  OAI22X1TS U3733 ( .A0(n4737), .A1(n3686), .B0(n4733), .B1(n3589), .Y(n5190)
         );
  OAI22X1TS U3734 ( .A0(n4745), .A1(n3686), .B0(n4746), .B1(n3588), .Y(n5198)
         );
  OAI22X1TS U3735 ( .A0(n4751), .A1(n3687), .B0(n4755), .B1(n3589), .Y(n5206)
         );
  OAI22X1TS U3736 ( .A0(n4758), .A1(n3687), .B0(n4764), .B1(n3588), .Y(n5215)
         );
  OAI22X1TS U3737 ( .A0(n4424), .A1(n608), .B0(n4425), .B1(n3635), .Y(n4871)
         );
  OAI22X1TS U3738 ( .A0(n4432), .A1(n610), .B0(n4430), .B1(n3647), .Y(n4879)
         );
  OAI22X1TS U3739 ( .A0(n4443), .A1(n612), .B0(n4439), .B1(n3650), .Y(n4887)
         );
  OAI22X1TS U3740 ( .A0(n4454), .A1(n612), .B0(n4452), .B1(n3646), .Y(n4895)
         );
  OAI22X1TS U3741 ( .A0(n4457), .A1(n622), .B0(n4461), .B1(n3648), .Y(n4903)
         );
  OAI22X1TS U3742 ( .A0(n4466), .A1(n610), .B0(n4468), .B1(n3645), .Y(n4911)
         );
  OAI22X1TS U3743 ( .A0(n4481), .A1(n613), .B0(n4477), .B1(n3646), .Y(n4919)
         );
  OAI22X1TS U3744 ( .A0(n4488), .A1(n613), .B0(n4486), .B1(n6319), .Y(n4927)
         );
  OAI22X1TS U3745 ( .A0(n4495), .A1(n613), .B0(n4497), .B1(n3649), .Y(n4935)
         );
  OAI22X1TS U3746 ( .A0(n4506), .A1(n612), .B0(n4502), .B1(n3650), .Y(n4943)
         );
  OAI22X1TS U3747 ( .A0(n4513), .A1(n613), .B0(n4517), .B1(n3643), .Y(n4951)
         );
  OAI22X1TS U3748 ( .A0(n4520), .A1(n623), .B0(n4522), .B1(n3643), .Y(n4959)
         );
  OAI22X1TS U3749 ( .A0(n4533), .A1(n614), .B0(n4535), .B1(n3643), .Y(n4967)
         );
  OAI22X1TS U3750 ( .A0(n4540), .A1(n622), .B0(n4538), .B1(n3643), .Y(n4975)
         );
  OAI22X1TS U3751 ( .A0(n4551), .A1(n611), .B0(n4549), .B1(n3642), .Y(n4983)
         );
  OAI22X1TS U3752 ( .A0(n4559), .A1(n659), .B0(n4560), .B1(n3642), .Y(n4991)
         );
  OAI22X1TS U3753 ( .A0(n4564), .A1(n624), .B0(n4565), .B1(n3642), .Y(n4999)
         );
  OAI22X1TS U3754 ( .A0(n4574), .A1(n659), .B0(n4580), .B1(n3642), .Y(n5007)
         );
  OAI22X1TS U3755 ( .A0(n4587), .A1(n660), .B0(n4583), .B1(n3641), .Y(n5015)
         );
  OAI22X1TS U3756 ( .A0(n4596), .A1(n660), .B0(n4592), .B1(n3641), .Y(n5023)
         );
  OAI22X1TS U3757 ( .A0(n4602), .A1(n660), .B0(n4603), .B1(n3641), .Y(n5031)
         );
  OAI22X1TS U3758 ( .A0(n4610), .A1(n611), .B0(n4616), .B1(n3641), .Y(n5039)
         );
  OAI22X1TS U3759 ( .A0(n4621), .A1(n608), .B0(n4625), .B1(n3640), .Y(n5047)
         );
  OAI22X1TS U3760 ( .A0(n4632), .A1(n608), .B0(n4630), .B1(n3640), .Y(n5055)
         );
  OAI22X1TS U3761 ( .A0(n4641), .A1(n608), .B0(n4637), .B1(n3640), .Y(n5063)
         );
  OAI22X1TS U3762 ( .A0(n4648), .A1(n607), .B0(n4652), .B1(n3639), .Y(n5071)
         );
  OAI22X1TS U3763 ( .A0(n4661), .A1(n607), .B0(n4655), .B1(n3639), .Y(n5079)
         );
  OAI22X1TS U3764 ( .A0(n4668), .A1(n607), .B0(n4664), .B1(n3639), .Y(n5087)
         );
  OAI22X1TS U3765 ( .A0(n4679), .A1(n607), .B0(n4677), .B1(n3639), .Y(n5095)
         );
  OAI22X1TS U3766 ( .A0(n4684), .A1(n594), .B0(n4682), .B1(n3638), .Y(n5103)
         );
  OAI22X1TS U3767 ( .A0(n4694), .A1(n594), .B0(n4695), .B1(n3638), .Y(n5111)
         );
  OAI22X1TS U3768 ( .A0(n4706), .A1(n594), .B0(n4700), .B1(n3638), .Y(n5119)
         );
  OAI22X1TS U3769 ( .A0(n4717), .A1(n582), .B0(n4719), .B1(n3636), .Y(n5175)
         );
  OAI22X1TS U3770 ( .A0(n4726), .A1(n582), .B0(n4721), .B1(n3636), .Y(n5183)
         );
  OAI22X1TS U3771 ( .A0(n4735), .A1(n582), .B0(n4731), .B1(n3636), .Y(n5191)
         );
  OAI22X1TS U3772 ( .A0(n4744), .A1(n581), .B0(n4742), .B1(n3635), .Y(n5199)
         );
  OAI22X1TS U3773 ( .A0(n4753), .A1(n581), .B0(n4749), .B1(n3635), .Y(n5207)
         );
  OAI22X1TS U3774 ( .A0(n4760), .A1(n581), .B0(n4763), .B1(n3635), .Y(n5216)
         );
  NOR3X1TS U3775 ( .A(n4), .B(n217), .C(n163), .Y(n5295) );
  NOR3X1TS U3776 ( .A(n5), .B(n216), .C(n6316), .Y(n5285) );
  NAND3X1TS U3777 ( .A(n302), .B(n388), .C(n3), .Y(n5297) );
  AOI2BB2X1TS U3778 ( .B0(readOutbuffer[3]), .B1(n253), .A0N(n19), .A1N(n612), 
        .Y(n5298) );
  AOI222XLTS U3779 ( .A0(readOutbuffer[4]), .A1(n5295), .B0(readOutbuffer[7]), 
        .B1(n5294), .C0(readOutbuffer[2]), .C1(n205), .Y(n5296) );
  AOI221X1TS U3780 ( .A0(n5285), .A1(writeOutbuffer[1]), .B0(n205), .B1(
        writeOutbuffer[2]), .C0(n5284), .Y(n5286) );
  OAI22X1TS U3781 ( .A0(n17), .A1(n581), .B0(n6315), .B1(n3640), .Y(n5284) );
  OA22X1TS U3782 ( .A0(n3597), .A1(n4766), .B0(n3687), .B1(n4765), .Y(n5226)
         );
  OA22X1TS U3783 ( .A0(n3597), .A1(n4774), .B0(n3687), .B1(n4779), .Y(n5233)
         );
  OA22X1TS U3784 ( .A0(n3597), .A1(n4784), .B0(n3688), .B1(n4788), .Y(n5240)
         );
  OA22X1TS U3785 ( .A0(n3602), .A1(n4790), .B0(n3688), .B1(n4793), .Y(n5247)
         );
  OA22X1TS U3786 ( .A0(n3596), .A1(n4802), .B0(n3688), .B1(n4804), .Y(n5254)
         );
  OA22X1TS U3787 ( .A0(n3596), .A1(n4806), .B0(n3688), .B1(n4807), .Y(n5261)
         );
  OA22X1TS U3788 ( .A0(n3596), .A1(n4814), .B0(n3689), .B1(n4820), .Y(n5268)
         );
  OA22X1TS U3789 ( .A0(n3596), .A1(n4826), .B0(n3689), .B1(n4827), .Y(n5275)
         );
  OA22X1TS U3790 ( .A0(n3626), .A1(n4771), .B0(n3609), .B1(n4772), .Y(n5223)
         );
  OA22X1TS U3791 ( .A0(n3626), .A1(n4775), .B0(n3609), .B1(n4773), .Y(n5230)
         );
  OA22X1TS U3792 ( .A0(n3626), .A1(n4781), .B0(n3610), .B1(n4785), .Y(n5237)
         );
  OA22X1TS U3793 ( .A0(n3626), .A1(n4791), .B0(n3610), .B1(n4794), .Y(n5244)
         );
  OA22X1TS U3794 ( .A0(n3627), .A1(n4803), .B0(n3610), .B1(n4799), .Y(n5251)
         );
  OA22X1TS U3795 ( .A0(n3627), .A1(n4809), .B0(n3610), .B1(n4805), .Y(n5258)
         );
  OA22X1TS U3796 ( .A0(n3627), .A1(n4813), .B0(n3611), .B1(n4815), .Y(n5265)
         );
  OA22X1TS U3797 ( .A0(n3627), .A1(n4825), .B0(n3611), .B1(n4828), .Y(n5272)
         );
  OA22X1TS U3798 ( .A0(n3648), .A1(n4768), .B0(n623), .B1(n4770), .Y(n5225) );
  OA22X1TS U3799 ( .A0(n3645), .A1(n4778), .B0(n609), .B1(n4780), .Y(n5232) );
  OA22X1TS U3800 ( .A0(n3647), .A1(n4782), .B0(n614), .B1(n4786), .Y(n5239) );
  AOI2BB2X1TS U3801 ( .B0(n5294), .B1(n480), .A0N(n610), .A1N(n4796), .Y(n5246) );
  OA22X1TS U3802 ( .A0(n3644), .A1(n4801), .B0(n609), .B1(n4800), .Y(n5253) );
  OA22X1TS U3803 ( .A0(n3644), .A1(n4808), .B0(n609), .B1(n4810), .Y(n5260) );
  OA22X1TS U3804 ( .A0(n3644), .A1(n4818), .B0(n609), .B1(n4816), .Y(n5267) );
  OA22X1TS U3805 ( .A0(n3644), .A1(n4824), .B0(n610), .B1(n4822), .Y(n5274) );
  OA22X1TS U3806 ( .A0(n3672), .A1(n4767), .B0(n3657), .B1(n4769), .Y(n5224)
         );
  OA22X1TS U3807 ( .A0(n3672), .A1(n4777), .B0(n3658), .B1(n4776), .Y(n5231)
         );
  OA22X1TS U3808 ( .A0(n3673), .A1(n4787), .B0(n3658), .B1(n4783), .Y(n5238)
         );
  OA22X1TS U3809 ( .A0(n3673), .A1(n4789), .B0(n3659), .B1(n4795), .Y(n5245)
         );
  OA22X1TS U3810 ( .A0(n3673), .A1(n4797), .B0(n3658), .B1(n4798), .Y(n5252)
         );
  OA22X1TS U3811 ( .A0(n3673), .A1(n4811), .B0(n3658), .B1(n4812), .Y(n5259)
         );
  OA22X1TS U3812 ( .A0(n3674), .A1(n4817), .B0(n3659), .B1(n4819), .Y(n5266)
         );
  OA22X1TS U3813 ( .A0(n3674), .A1(n4821), .B0(n3659), .B1(n4823), .Y(n5273)
         );
  AOI22X1TS U3814 ( .A0(n396), .A1(writeOutbuffer[6]), .B0(writeOutbuffer[3]), 
        .B1(n207), .Y(n5288) );
  AOI22X1TS U3815 ( .A0(n5295), .A1(writeOutbuffer[4]), .B0(n246), .B1(
        writeOutbuffer[0]), .Y(n5287) );
  AOI32XLTS U3816 ( .A0(n109), .A1(n5540), .A2(n5539), .B0(n3357), .B1(n97), 
        .Y(n2567) );
  AOI32XLTS U3817 ( .A0(n193), .A1(n5526), .A2(n5525), .B0(n259), .B1(n99), 
        .Y(n2565) );
  AOI21XLTS U3818 ( .A0(n3803), .A1(n6337), .B0(n203), .Y(n5534) );
  AOI32XLTS U3819 ( .A0(n5532), .A1(n5531), .A2(n3808), .B0(n5530), .B1(n5529), 
        .Y(n5533) );
  AOI21XLTS U3820 ( .A0(n3815), .A1(n197), .B0(n6348), .Y(n5514) );
  OAI221XLTS U3821 ( .A0(n256), .A1(n264), .B0(n191), .B1(n103), .C0(n5564), 
        .Y(n2571) );
  OAI221XLTS U3822 ( .A0(n255), .A1(n266), .B0(n4828), .B1(n383), .C0(n5330), 
        .Y(n2458) );
  OAI221XLTS U3823 ( .A0(n5566), .A1(n269), .B0(n4815), .B1(n191), .C0(n5329), 
        .Y(n2457) );
  OAI221XLTS U3824 ( .A0(n256), .A1(n287), .B0(n4805), .B1(n383), .C0(n5328), 
        .Y(n2456) );
  OAI221XLTS U3825 ( .A0(n255), .A1(n278), .B0(n4799), .B1(n191), .C0(n5325), 
        .Y(n2455) );
  OAI221XLTS U3826 ( .A0(n5566), .A1(n6240), .B0(n4794), .B1(n232), .C0(n5324), 
        .Y(n2454) );
  OAI221XLTS U3827 ( .A0(n256), .A1(n284), .B0(n4785), .B1(n191), .C0(n5322), 
        .Y(n2453) );
  OAI221XLTS U3828 ( .A0(n255), .A1(n6242), .B0(n4773), .B1(n383), .C0(n5321), 
        .Y(n2452) );
  OAI221XLTS U3829 ( .A0(n5566), .A1(n281), .B0(n4772), .B1(n383), .C0(n5320), 
        .Y(n2451) );
  AND3X2TS U3830 ( .A(n5512), .B(n5511), .C(n5319), .Y(n6103) );
  OAI221XLTS U3831 ( .A0(n295), .A1(n6235), .B0(n222), .B1(n101), .C0(n5569), 
        .Y(n2573) );
  OAI221XLTS U3832 ( .A0(n5571), .A1(n6236), .B0(n4827), .B1(n5570), .C0(n5374), .Y(n2486) );
  OAI221XLTS U3833 ( .A0(n295), .A1(n6237), .B0(n4820), .B1(n221), .C0(n5373), 
        .Y(n2485) );
  OAI221XLTS U3834 ( .A0(n5571), .A1(n6238), .B0(n4807), .B1(n5570), .C0(n5372), .Y(n2484) );
  OAI221XLTS U3835 ( .A0(n295), .A1(n6239), .B0(n4804), .B1(n221), .C0(n5371), 
        .Y(n2483) );
  OAI221XLTS U3836 ( .A0(n294), .A1(n276), .B0(n4793), .B1(n5570), .C0(n5370), 
        .Y(n2482) );
  OAI221XLTS U3837 ( .A0(n295), .A1(n6241), .B0(n4788), .B1(n222), .C0(n5369), 
        .Y(n2481) );
  OAI221XLTS U3838 ( .A0(n5571), .A1(n273), .B0(n4779), .B1(n221), .C0(n5368), 
        .Y(n2480) );
  OAI221XLTS U3839 ( .A0(n294), .A1(n281), .B0(n4765), .B1(n222), .C0(n5367), 
        .Y(n2479) );
endmodule


module outputPortArbiter_3 ( clk, reset, selectBit_NORTH, 
        destinationAddressIn_NORTH, requesterAddressIn_NORTH, readIn_NORTH, 
        writeIn_NORTH, dataIn_NORTH, selectBit_SOUTH, 
        destinationAddressIn_SOUTH, requesterAddressIn_SOUTH, readIn_SOUTH, 
        writeIn_SOUTH, dataIn_SOUTH, selectBit_EAST, destinationAddressIn_EAST, 
        requesterAddressIn_EAST, readIn_EAST, writeIn_EAST, dataIn_EAST, 
        selectBit_WEST, destinationAddressIn_WEST, requesterAddressIn_WEST, 
        readIn_WEST, writeIn_WEST, dataIn_WEST, readReady, 
        readRequesterAddress, cacheDataOut, destinationAddressOut, 
        requesterAddressOut, readOut, writeOut, dataOut );
  input [13:0] destinationAddressIn_NORTH;
  input [5:0] requesterAddressIn_NORTH;
  input [31:0] dataIn_NORTH;
  input [13:0] destinationAddressIn_SOUTH;
  input [5:0] requesterAddressIn_SOUTH;
  input [31:0] dataIn_SOUTH;
  input [13:0] destinationAddressIn_EAST;
  input [5:0] requesterAddressIn_EAST;
  input [31:0] dataIn_EAST;
  input [13:0] destinationAddressIn_WEST;
  input [5:0] requesterAddressIn_WEST;
  input [31:0] dataIn_WEST;
  input [5:0] readRequesterAddress;
  input [31:0] cacheDataOut;
  output [13:0] destinationAddressOut;
  output [5:0] requesterAddressOut;
  output [31:0] dataOut;
  input clk, reset, selectBit_NORTH, readIn_NORTH, writeIn_NORTH,
         selectBit_SOUTH, readIn_SOUTH, writeIn_SOUTH, selectBit_EAST,
         readIn_EAST, writeIn_EAST, selectBit_WEST, readIn_WEST, writeIn_WEST,
         readReady;
  output readOut, writeOut;
  wire   N4718, n2888, n5327, n2886, n5326, n2889, n2883, n2887, n5323, n2569,
         n2567, n2566, n2578, n2638, n2624, n2617, n2577, n2544, n2541, n2540,
         n2537, n2535, n2703, n2692, n2691, n2689, n2511, n2507, n2731, n2574,
         n2499, n2496, n2493, n2770, n2768, n2764, n2754, n2748, n2746, n2739,
         n2486, n2484, n2482, n2480, n2802, n2834, n2833, n2832, n2829, n2825,
         n2814, n2811, n2807, n2806, n2457, n2455, n2453, n2570, n2565, n2573,
         n2568, n2564, n2563, n2575, n2882, n2881, n2879, n2610, n2609, n2608,
         n2607, n2606, n2605, n2604, n2603, n2602, n2601, n2600, n2599, n2598,
         n2597, n2596, n2595, n2594, n2593, n2592, n2591, n2590, n2589, n2588,
         n2587, n2586, n2585, n2584, n2583, n2582, n2581, n2580, n2579, n2561,
         n2560, n2559, n2557, n2556, n2555, n2554, n2552, n2551, n2550, n2549,
         n2642, n2640, n2639, n2637, n2635, n2634, n2633, n2631, n2628, n2627,
         n2626, n2625, n2623, n2620, n2618, n2616, n2615, n2614, n2612, n2611,
         n2870, n2869, n2868, n2867, n2866, n2865, n2674, n2672, n2671, n2670,
         n2669, n2668, n2667, n2666, n2665, n2664, n2662, n2661, n2660, n2657,
         n2656, n2655, n2654, n2653, n2652, n2651, n2650, n2649, n2648, n2647,
         n2646, n2645, n2644, n2576, n2534, n2533, n2532, n2531, n2530, n2529,
         n2528, n2527, n2526, n2525, n2524, n2523, n2522, n2521, n2860, n2859,
         n2706, n2705, n2700, n2698, n2696, n2695, n2694, n2690, n2687, n2686,
         n2685, n2684, n2677, n2675, n2736, n2734, n2733, n2725, n2723, n2720,
         n2718, n2715, n2713, n2504, n2498, n2497, n2494, n2850,
         \requesterAddressbuffer[2][2] , n2849, \requesterAddressbuffer[2][3] ,
         n2847, \requesterAddressbuffer[2][5] , n2769, n2760, n2743, n2492,
         n2491, n2489, n2488, n2487, n2485, n2483, n2481, n2846, n2845, n2844,
         n2843, n2842, n2841, n2801, n2799, n2798, n2796, n2795, n2793, n2791,
         n2790, n2789, n2788, n2787, n2786, n2785, n2784, n2781, n2779, n2778,
         n2777, n2776, n2774, n2773, n2772, n2771, n2572, n2478, n2477, n2476,
         n2475, n2474, n2473, n2472, n2471, n2470, n2469, n2468, n2467, n2466,
         n2465, n2840, \requesterAddressbuffer[0][0] , n2839,
         \requesterAddressbuffer[0][1] , n2838, \requesterAddressbuffer[0][2] ,
         n2836, \requesterAddressbuffer[0][4] , n2571, n2464, n2460, n2458,
         n2454, n2451, n2880, n2878, n2877, n2562, n2558, n2553, n2876,
         \requesterAddressbuffer[6][0] , n2875, \requesterAddressbuffer[6][1] ,
         n2874, \requesterAddressbuffer[6][2] , n2873,
         \requesterAddressbuffer[6][3] , n2872, \requesterAddressbuffer[6][4] ,
         n2871, \requesterAddressbuffer[6][5] , n2641, n2636, n2632, n2630,
         n2629, n2622, n2621, n2619, n2613, n2548, n2547, n2546, n2545, n2543,
         n2542, n2539, n2538, n2536, n2673, n2663, n2659, n2658, n2643, n2864,
         n2863, n2862, n2861, n2704, n2702, n2701, n2699, n2697, n2693, n2688,
         n2683, n2682, n2681, n2680, n2679, n2678, n2676, n2520, n2519, n2518,
         n2517, n2516, n2515, n2514, n2513, n2512, n2510, n2509, n2508, n2858,
         \requesterAddressbuffer[3][0] , n2857, \requesterAddressbuffer[3][1] ,
         n2856, \requesterAddressbuffer[3][2] , n2855,
         \requesterAddressbuffer[3][3] , n2854, \requesterAddressbuffer[3][4] ,
         n2853, \requesterAddressbuffer[3][5] , n2738, n2737, n2735, n2732,
         n2730, n2729, n2728, n2727, n2726, n2724, n2722, n2721, n2719, n2717,
         n2716, n2714, n2712, n2711, n2710, n2709, n2708, n2707, n2506, n2505,
         n2503, n2502, n2501, n2500, n2495, n2852,
         \requesterAddressbuffer[2][0] , n2851, \requesterAddressbuffer[2][1] ,
         n2848, \requesterAddressbuffer[2][4] , n2767, n2766, n2765, n2763,
         n2762, n2761, n2759, n2758, n2757, n2756, n2755, n2753, n2752, n2751,
         n2750, n2749, n2747, n2745, n2744, n2742, n2741, n2740, n2490, n2479,
         n2800, n2797, n2794, n2792, n2783, n2782, n2780, n2775, n2837,
         \requesterAddressbuffer[0][3] , n2835, \requesterAddressbuffer[0][5] ,
         n2831, n2830, n2828, n2827, n2826, n2824, n2823, n2822, n2821, n2820,
         n2819, n2818, n2817, n2816, n2815, n2813, n2812, n2810, n2809, n2808,
         n2805, n2804, n2803, n2463, n2462, n2461, n2459, n2456, n2452, n2885,
         n2449, n2434, n2431, n2450, n2448, n2447, n2446, n2445, n2444, n2443,
         n2442, n2441, n2440, n2439, n2438, n2437, n2436, n2435, n2433, n2432,
         n2430, n2429, n2428, n2427, n2426, n2425, n2424, n2423, n2422, n2421,
         n2420, n2419, n2418, n2417, n2416, n2415, n2414, n2413, n2412, n2411,
         n2410, n2409, n2408, n2407, n2406, n2405, n2404, n2403, n2402, n2401,
         n2400, n2399, n2398, n2397, n2884, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n496, n499, n500, n501, n502, n503,
         n505, n507, n508, n509, n511, n514, n516, n517, n526, n536, n537,
         n541, n543, n544, n545, n546, n548, n551, n554, n555, n556, n557,
         n558, n559, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n581,
         n582, n583, n584, n585, n586, n587, n594, n607, n608, n609, n610,
         n611, n612, n613, n614, n622, n623, n624, n625, n626, n627, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n711, n712, n714, n715, n716, n729,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n886, n919, n936, n955, n957,
         n959, n970, n986, n1402, n1602, n1654, n1728, n1764, n1797, n1817,
         n1822, n1894, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5324, n5325, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347;
  wire   [0:7] readOutbuffer;
  wire   [0:7] writeOutbuffer;

  DFFNSRX2TS \destinationAddressbuffer_reg[0][7]  ( .D(n2457), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4819) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][6]  ( .D(n2458), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4832) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][8]  ( .D(n2456), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4809) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][7]  ( .D(n2499), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4823) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][10]  ( .D(n2496), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4799) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][13]  ( .D(n2493), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4773) );
  DFFNSRX2TS \destinationAddressbuffer_reg[5][6]  ( .D(n2528), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4826) );
  DFFNSRX2TS \destinationAddressbuffer_reg[5][7]  ( .D(n2527), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4820) );
  DFFNSRX2TS \destinationAddressbuffer_reg[5][8]  ( .D(n2526), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4814) );
  DFFNSRX2TS \destinationAddressbuffer_reg[5][9]  ( .D(n2525), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4804) );
  DFFNSRX2TS \destinationAddressbuffer_reg[5][10]  ( .D(n2524), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4800) );
  DFFNSRX2TS \destinationAddressbuffer_reg[5][11]  ( .D(n2523), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4790) );
  DFFNSRX2TS \destinationAddressbuffer_reg[5][12]  ( .D(n2522), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4784) );
  DFFNSRX2TS \destinationAddressbuffer_reg[5][13]  ( .D(n2521), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4774) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][8]  ( .D(n2498), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4816) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][9]  ( .D(n2497), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4802) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][12]  ( .D(n2494), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4780) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][6]  ( .D(n2500), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4827) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][11]  ( .D(n2495), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4787) );
  DFFNSRX2TS \destinationAddressbuffer_reg[6][7]  ( .D(n2541), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4821) );
  DFFNSRX2TS \destinationAddressbuffer_reg[6][8]  ( .D(n2540), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4815) );
  DFFNSRX2TS \destinationAddressbuffer_reg[6][11]  ( .D(n2537), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4791) );
  DFFNSRX2TS \destinationAddressbuffer_reg[6][13]  ( .D(n2535), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4771) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][9]  ( .D(n2511), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4807) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][13]  ( .D(n2507), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4775) );
  DFFNSRX2TS \destinationAddressbuffer_reg[7][6]  ( .D(n2556), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4828) );
  DFFNSRX2TS \destinationAddressbuffer_reg[7][7]  ( .D(n2555), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4822) );
  DFFNSRX2TS \destinationAddressbuffer_reg[7][8]  ( .D(n2554), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4812) );
  DFFNSRX2TS \destinationAddressbuffer_reg[7][10]  ( .D(n2552), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n431), .QN(n4796) );
  DFFNSRX2TS \destinationAddressbuffer_reg[7][11]  ( .D(n2551), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4786) );
  DFFNSRX2TS \destinationAddressbuffer_reg[7][12]  ( .D(n2550), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4782) );
  DFFNSRX2TS \destinationAddressbuffer_reg[7][13]  ( .D(n2549), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4772) );
  DFFNSRX2TS \destinationAddressbuffer_reg[7][9]  ( .D(n2553), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4805) );
  DFFNSRX2TS \destinationAddressbuffer_reg[6][6]  ( .D(n2542), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4825) );
  DFFNSRX2TS \destinationAddressbuffer_reg[6][9]  ( .D(n2539), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4801) );
  DFFNSRX2TS \destinationAddressbuffer_reg[6][10]  ( .D(n2538), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4793) );
  DFFNSRX2TS \destinationAddressbuffer_reg[6][12]  ( .D(n2536), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4781) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][6]  ( .D(n2514), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4829) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][7]  ( .D(n2513), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4817) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][8]  ( .D(n2512), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4813) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][10]  ( .D(n2510), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4795) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][11]  ( .D(n2509), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4785) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][12]  ( .D(n2508), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4779) );
  DFFNSRX2TS \dataoutbuffer_reg[6][4]  ( .D(n2638), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4673) );
  DFFNSRX2TS \destinationAddressbuffer_reg[6][4]  ( .D(n2544), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4731) );
  DFFNSRX2TS \dataoutbuffer_reg[7][1]  ( .D(n2609), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4699) );
  DFFNSRX2TS \dataoutbuffer_reg[7][2]  ( .D(n2608), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4686) );
  DFFNSRX2TS \dataoutbuffer_reg[7][3]  ( .D(n2607), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4681) );
  DFFNSRX2TS \dataoutbuffer_reg[7][4]  ( .D(n2606), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4668) );
  DFFNSRX2TS \dataoutbuffer_reg[7][5]  ( .D(n2605), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4659) );
  DFFNSRX2TS \dataoutbuffer_reg[7][6]  ( .D(n2604), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4656) );
  DFFNSRX2TS \dataoutbuffer_reg[7][7]  ( .D(n2603), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4641) );
  DFFNSRX2TS \dataoutbuffer_reg[7][8]  ( .D(n2602), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4634) );
  DFFNSRX2TS \dataoutbuffer_reg[7][9]  ( .D(n2601), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4629) );
  DFFNSRX2TS \dataoutbuffer_reg[7][10]  ( .D(n2600), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4620) );
  DFFNSRX2TS \dataoutbuffer_reg[7][11]  ( .D(n2599), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4607) );
  DFFNSRX2TS \dataoutbuffer_reg[7][12]  ( .D(n2598), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4596) );
  DFFNSRX2TS \dataoutbuffer_reg[7][16]  ( .D(n2594), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4564) );
  DFFNSRX2TS \dataoutbuffer_reg[7][17]  ( .D(n2593), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4553) );
  DFFNSRX2TS \dataoutbuffer_reg[7][18]  ( .D(n2592), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4542) );
  DFFNSRX2TS \dataoutbuffer_reg[7][19]  ( .D(n2591), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4539) );
  DFFNSRX2TS \dataoutbuffer_reg[7][20]  ( .D(n2590), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4526) );
  DFFNSRX2TS \dataoutbuffer_reg[7][21]  ( .D(n2589), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4521) );
  DFFNSRX2TS \dataoutbuffer_reg[7][22]  ( .D(n2588), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4506) );
  DFFNSRX2TS \dataoutbuffer_reg[7][23]  ( .D(n2587), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4501) );
  DFFNSRX2TS \dataoutbuffer_reg[7][24]  ( .D(n2586), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4490) );
  DFFNSRX2TS \dataoutbuffer_reg[7][25]  ( .D(n2585), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4481) );
  DFFNSRX2TS \dataoutbuffer_reg[7][26]  ( .D(n2584), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4472) );
  DFFNSRX2TS \dataoutbuffer_reg[7][27]  ( .D(n2583), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4465) );
  DFFNSRX2TS \dataoutbuffer_reg[7][28]  ( .D(n2582), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4456) );
  DFFNSRX2TS \dataoutbuffer_reg[7][29]  ( .D(n2581), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4443) );
  DFFNSRX2TS \dataoutbuffer_reg[7][30]  ( .D(n2580), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4434) );
  DFFNSRX2TS \dataoutbuffer_reg[7][31]  ( .D(n2579), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4429) );
  DFFNSRX2TS \destinationAddressbuffer_reg[7][1]  ( .D(n2561), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4753) );
  DFFNSRX2TS \destinationAddressbuffer_reg[7][2]  ( .D(n2560), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4746) );
  DFFNSRX2TS \destinationAddressbuffer_reg[7][3]  ( .D(n2559), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4735) );
  DFFNSRX2TS \destinationAddressbuffer_reg[7][5]  ( .D(n2557), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4723) );
  DFFNSRX2TS \dataoutbuffer_reg[6][0]  ( .D(n2642), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4708) );
  DFFNSRX2TS \dataoutbuffer_reg[6][2]  ( .D(n2640), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4692) );
  DFFNSRX2TS \dataoutbuffer_reg[6][3]  ( .D(n2639), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4677) );
  DFFNSRX2TS \dataoutbuffer_reg[6][5]  ( .D(n2637), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4661) );
  DFFNSRX2TS \dataoutbuffer_reg[6][7]  ( .D(n2635), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4643) );
  DFFNSRX2TS \dataoutbuffer_reg[6][8]  ( .D(n2634), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4638) );
  DFFNSRX2TS \dataoutbuffer_reg[6][9]  ( .D(n2633), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4627) );
  DFFNSRX2TS \dataoutbuffer_reg[6][11]  ( .D(n2631), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4611) );
  DFFNSRX2TS \dataoutbuffer_reg[6][30]  ( .D(n2612), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4438) );
  DFFNSRX2TS \dataoutbuffer_reg[6][31]  ( .D(n2611), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4427) );
  DFFNSRX2TS \destinationAddressbuffer_reg[7][0]  ( .D(n2562), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4767) );
  DFFNSRX2TS \destinationAddressbuffer_reg[7][4]  ( .D(n2558), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4725) );
  DFFNSRX2TS \dataoutbuffer_reg[6][1]  ( .D(n2641), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4696) );
  DFFNSRX2TS \dataoutbuffer_reg[6][6]  ( .D(n2636), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4649) );
  DFFNSRX2TS \dataoutbuffer_reg[6][10]  ( .D(n2632), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4613) );
  DFFNSRX2TS \destinationAddressbuffer_reg[6][0]  ( .D(n2548), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4763) );
  DFFNSRX2TS \destinationAddressbuffer_reg[6][1]  ( .D(n2547), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4754) );
  DFFNSRX2TS \destinationAddressbuffer_reg[6][2]  ( .D(n2546), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4745) );
  DFFNSRX2TS \destinationAddressbuffer_reg[6][3]  ( .D(n2545), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4734) );
  DFFNSRX2TS \destinationAddressbuffer_reg[6][5]  ( .D(n2543), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4720) );
  DFFNSRX2TS \requesterAddressbuffer_reg[6][0]  ( .D(n2876), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][0] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[6][1]  ( .D(n2875), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][1] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[6][2]  ( .D(n2874), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][2] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[6][3]  ( .D(n2873), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][3] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[6][4]  ( .D(n2872), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][4] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[6][5]  ( .D(n2871), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][5] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[2][2]  ( .D(n2850), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][2] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[2][3]  ( .D(n2849), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][3] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[2][5]  ( .D(n2847), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][5] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[0][0]  ( .D(n2840), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][0] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[0][1]  ( .D(n2839), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][1] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[0][2]  ( .D(n2838), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][2] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[0][4]  ( .D(n2836), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][4] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[2][0]  ( .D(n2852), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][0] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[2][1]  ( .D(n2851), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][1] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[2][4]  ( .D(n2848), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][4] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[0][3]  ( .D(n2837), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][3] ) );
  DFFNSRX2TS \requesterAddressbuffer_reg[0][5]  ( .D(n2835), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][5] ) );
  DFFNSRX2TS \readOutbuffer_reg[3]  ( .D(n2566), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[3]) );
  DFFNSRX2TS \readOutbuffer_reg[6]  ( .D(n2569), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n11) );
  DFFNSRX2TS \writeOutbuffer_reg[7]  ( .D(n2578), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n10) );
  DFFNSRX2TS \readOutbuffer_reg[5]  ( .D(n2568), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n25) );
  DFFNSRX2TS \readOutbuffer_reg[1]  ( .D(n2564), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n17) );
  DFFNSRX2TS \readOutbuffer_reg[0]  ( .D(n2563), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n26) );
  DFFNSRX2TS \requesterAddressbuffer_reg[7][0]  ( .D(n2882), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n24) );
  DFFNSRX2TS \requesterAddressbuffer_reg[7][1]  ( .D(n2881), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n22) );
  DFFNSRX2TS \requesterAddressbuffer_reg[7][3]  ( .D(n2879), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n23) );
  DFFNSRX2TS \writeOutbuffer_reg[5]  ( .D(n2576), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n18) );
  DFFNSRX2TS \requesterAddressbuffer_reg[7][2]  ( .D(n2880), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n21) );
  DFFNSRX2TS \requesterAddressbuffer_reg[7][4]  ( .D(n2878), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n20) );
  DFFNSRX2TS \requesterAddressbuffer_reg[7][5]  ( .D(n2877), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n19) );
  DFFNSRX2TS \dataoutbuffer_reg[2][0]  ( .D(n2770), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n102), .QN(n4705) );
  DFFNSRX2TS \dataoutbuffer_reg[2][2]  ( .D(n2768), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n101), .QN(n4689) );
  DFFNSRX2TS \dataoutbuffer_reg[2][6]  ( .D(n2764), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n100), .QN(n4655) );
  DFFNSRX2TS \dataoutbuffer_reg[2][16]  ( .D(n2754), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n99), .QN(n4565) );
  DFFNSRX2TS \dataoutbuffer_reg[2][22]  ( .D(n2748), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n98), .QN(n4511) );
  DFFNSRX2TS \dataoutbuffer_reg[2][24]  ( .D(n2746), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n97), .QN(n4493) );
  DFFNSRX2TS \dataoutbuffer_reg[2][31]  ( .D(n2739), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n96), .QN(n4430) );
  DFFNSRX2TS \dataoutbuffer_reg[0][0]  ( .D(n2834), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n64), .QN(n4707) );
  DFFNSRX2TS \dataoutbuffer_reg[0][1]  ( .D(n2833), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n63), .QN(n4700) );
  DFFNSRX2TS \dataoutbuffer_reg[0][2]  ( .D(n2832), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n62), .QN(n4691) );
  DFFNSRX2TS \dataoutbuffer_reg[0][5]  ( .D(n2829), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n61), .QN(n4664) );
  DFFNSRX2TS \dataoutbuffer_reg[0][9]  ( .D(n2825), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n60), .QN(n4628) );
  DFFNSRX2TS \dataoutbuffer_reg[0][20]  ( .D(n2814), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n59), .QN(n4529) );
  DFFNSRX2TS \dataoutbuffer_reg[0][23]  ( .D(n2811), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n58), .QN(n4502) );
  DFFNSRX2TS \dataoutbuffer_reg[0][27]  ( .D(n2807), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n57), .QN(n4466) );
  DFFNSRX2TS \dataoutbuffer_reg[0][28]  ( .D(n2806), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n56), .QN(n4457) );
  DFFNSRX2TS \dataoutbuffer_reg[2][1]  ( .D(n2769), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n95), .QN(n4701) );
  DFFNSRX2TS \dataoutbuffer_reg[2][10]  ( .D(n2760), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n94), .QN(n4618) );
  DFFNSRX2TS \dataoutbuffer_reg[2][27]  ( .D(n2743), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n93), .QN(n4467) );
  DFFNSRX2TS \destinationAddressbuffer_reg[2][0]  ( .D(n2492), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n92), .QN(n4762) );
  DFFNSRX2TS \destinationAddressbuffer_reg[2][1]  ( .D(n2491), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n91), .QN(n4755) );
  DFFNSRX2TS \destinationAddressbuffer_reg[2][3]  ( .D(n2489), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n90), .QN(n4741) );
  DFFNSRX2TS \destinationAddressbuffer_reg[2][4]  ( .D(n2488), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n89), .QN(n4732) );
  DFFNSRX2TS \destinationAddressbuffer_reg[2][5]  ( .D(n2487), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n88), .QN(n4719) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][0]  ( .D(n2464), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n55), .QN(n4766) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][4]  ( .D(n2460), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n54), .QN(n4728) );
  DFFNSRX2TS \dataoutbuffer_reg[2][3]  ( .D(n2767), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n87), .QN(n4676) );
  DFFNSRX2TS \dataoutbuffer_reg[2][4]  ( .D(n2766), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n86), .QN(n4669) );
  DFFNSRX2TS \dataoutbuffer_reg[2][5]  ( .D(n2765), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n85), .QN(n4662) );
  DFFNSRX2TS \dataoutbuffer_reg[2][7]  ( .D(n2763), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n84), .QN(n4640) );
  DFFNSRX2TS \dataoutbuffer_reg[2][8]  ( .D(n2762), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n83), .QN(n4635) );
  DFFNSRX2TS \dataoutbuffer_reg[2][9]  ( .D(n2761), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n82), .QN(n4622) );
  DFFNSRX2TS \dataoutbuffer_reg[2][11]  ( .D(n2759), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n81), .QN(n4610) );
  DFFNSRX2TS \dataoutbuffer_reg[2][12]  ( .D(n2758), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n80), .QN(n4595) );
  DFFNSRX2TS \dataoutbuffer_reg[2][13]  ( .D(n2757), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n79), .QN(n4588) );
  DFFNSRX2TS \dataoutbuffer_reg[2][14]  ( .D(n2756), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n78), .QN(n4577) );
  DFFNSRX2TS \dataoutbuffer_reg[2][15]  ( .D(n2755), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n77), .QN(n4570) );
  DFFNSRX2TS \dataoutbuffer_reg[2][17]  ( .D(n2753), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n76), .QN(n4554) );
  DFFNSRX2TS \dataoutbuffer_reg[2][18]  ( .D(n2752), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n75), .QN(n4545) );
  DFFNSRX2TS \dataoutbuffer_reg[2][19]  ( .D(n2751), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n74), .QN(n4532) );
  DFFNSRX2TS \dataoutbuffer_reg[2][20]  ( .D(n2750), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n73), .QN(n4527) );
  DFFNSRX2TS \dataoutbuffer_reg[2][21]  ( .D(n2749), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n72), .QN(n4514) );
  DFFNSRX2TS \dataoutbuffer_reg[2][23]  ( .D(n2747), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n71), .QN(n4500) );
  DFFNSRX2TS \dataoutbuffer_reg[2][25]  ( .D(n2745), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n70), .QN(n4478) );
  DFFNSRX2TS \dataoutbuffer_reg[2][26]  ( .D(n2744), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n69), .QN(n4471) );
  DFFNSRX2TS \dataoutbuffer_reg[2][28]  ( .D(n2742), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n68), .QN(n4453) );
  DFFNSRX2TS \dataoutbuffer_reg[2][29]  ( .D(n2741), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n67), .QN(n4442) );
  DFFNSRX2TS \dataoutbuffer_reg[2][30]  ( .D(n2740), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n66), .QN(n4435) );
  DFFNSRX2TS \destinationAddressbuffer_reg[2][2]  ( .D(n2490), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n65), .QN(n4749) );
  DFFNSRX2TS \dataoutbuffer_reg[0][3]  ( .D(n2831), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n53), .QN(n4678) );
  DFFNSRX2TS \dataoutbuffer_reg[0][4]  ( .D(n2830), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n52), .QN(n4667) );
  DFFNSRX2TS \dataoutbuffer_reg[0][6]  ( .D(n2828), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n51), .QN(n4651) );
  DFFNSRX2TS \dataoutbuffer_reg[0][7]  ( .D(n2827), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n50), .QN(n4642) );
  DFFNSRX2TS \dataoutbuffer_reg[0][8]  ( .D(n2826), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n49), .QN(n4637) );
  DFFNSRX2TS \dataoutbuffer_reg[0][10]  ( .D(n2824), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n48), .QN(n4617) );
  DFFNSRX2TS \dataoutbuffer_reg[0][11]  ( .D(n2823), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n47), .QN(n4604) );
  DFFNSRX2TS \dataoutbuffer_reg[0][12]  ( .D(n2822), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n46), .QN(n4599) );
  DFFNSRX2TS \dataoutbuffer_reg[0][13]  ( .D(n2821), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n45), .QN(n4592) );
  DFFNSRX2TS \dataoutbuffer_reg[0][14]  ( .D(n2820), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n44), .QN(n4579) );
  DFFNSRX2TS \dataoutbuffer_reg[0][15]  ( .D(n2819), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n43), .QN(n4572) );
  DFFNSRX2TS \dataoutbuffer_reg[0][16]  ( .D(n2818), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n42), .QN(n4561) );
  DFFNSRX2TS \dataoutbuffer_reg[0][17]  ( .D(n2817), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n41), .QN(n4552) );
  DFFNSRX2TS \dataoutbuffer_reg[0][18]  ( .D(n2816), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n40), .QN(n4543) );
  DFFNSRX2TS \dataoutbuffer_reg[0][19]  ( .D(n2815), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n39), .QN(n4534) );
  DFFNSRX2TS \dataoutbuffer_reg[0][21]  ( .D(n2813), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n38), .QN(n4520) );
  DFFNSRX2TS \dataoutbuffer_reg[0][22]  ( .D(n2812), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n37), .QN(n4505) );
  DFFNSRX2TS \dataoutbuffer_reg[0][24]  ( .D(n2810), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n36), .QN(n4489) );
  DFFNSRX2TS \dataoutbuffer_reg[0][25]  ( .D(n2809), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n35), .QN(n4480) );
  DFFNSRX2TS \dataoutbuffer_reg[0][26]  ( .D(n2808), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n34), .QN(n4473) );
  DFFNSRX2TS \dataoutbuffer_reg[0][29]  ( .D(n2805), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n33), .QN(n4448) );
  DFFNSRX2TS \dataoutbuffer_reg[0][30]  ( .D(n2804), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n32), .QN(n4437) );
  DFFNSRX2TS \dataoutbuffer_reg[0][31]  ( .D(n2803), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n31), .QN(n4424) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][1]  ( .D(n2463), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n30), .QN(n4752) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][2]  ( .D(n2462), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n29), .QN(n4747) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][3]  ( .D(n2461), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n28), .QN(n4736) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][5]  ( .D(n2459), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n27), .QN(n4716) );
  DFFNSRX2TS \writeOutbuffer_reg[0]  ( .D(n2571), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[0]), .QN(n109) );
  DFFNSRX2TS \writeOutbuffer_reg[3]  ( .D(n2574), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[3]), .QN(n108) );
  DFFNSRX2TS \writeOutbuffer_reg[6]  ( .D(n2577), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[6]), .QN(n106) );
  DFFNSRX2TS \writeOutbuffer_reg[4]  ( .D(n2575), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[4]), .QN(n107) );
  DFFNSRX2TS \readOutbuffer_reg[7]  ( .D(n2570), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[7]), .QN(n104) );
  DFFNSRX2TS \readOutbuffer_reg[2]  ( .D(n2565), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[2]), .QN(n105) );
  DFFNSRX2TS \readOutbuffer_reg[4]  ( .D(n2567), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[4]), .QN(n103) );
  DFFNSRX2TS \read_reg_reg[0]  ( .D(n2889), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n4), .QN(n8) );
  DFFNSRX2TS \write_reg_reg[1]  ( .D(n2887), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n343), .QN(n5323) );
  DFFNSRX2TS writeOut_reg ( .D(n2449), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        writeOut), .QN(n4833) );
  DFFNSRX2TS \requesterAddressOut_reg[0]  ( .D(n2434), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[0]), .QN(n4837) );
  DFFNSRX2TS \requesterAddressOut_reg[3]  ( .D(n2431), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[3]), .QN(n4838) );
  DFFNSRX2TS readOut_reg ( .D(n2450), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        readOut), .QN(n4835) );
  DFFNSRX2TS \destinationAddressOut_reg[0]  ( .D(n2440), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[0]), .QN(n4760) );
  DFFNSRX2TS \destinationAddressOut_reg[1]  ( .D(n2439), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[1]), .QN(n4751) );
  DFFNSRX2TS \destinationAddressOut_reg[2]  ( .D(n2438), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[2]), .QN(n4742) );
  DFFNSRX2TS \destinationAddressOut_reg[3]  ( .D(n2437), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[3]), .QN(n4733) );
  DFFNSRX2TS \destinationAddressOut_reg[4]  ( .D(n2436), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[4]), .QN(n4724) );
  DFFNSRX2TS \destinationAddressOut_reg[5]  ( .D(n2435), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[5]), .QN(n4715) );
  DFFNSRX2TS \requesterAddressOut_reg[1]  ( .D(n2433), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[1]), .QN(n4714) );
  DFFNSRX2TS \requesterAddressOut_reg[2]  ( .D(n2432), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[2]), .QN(n4713) );
  DFFNSRX2TS \requesterAddressOut_reg[4]  ( .D(n2430), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[4]), .QN(n4712) );
  DFFNSRX2TS \requesterAddressOut_reg[5]  ( .D(n2429), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[5]), .QN(n4711) );
  DFFNSRX2TS \dataOut_reg[0]  ( .D(n2428), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[0]), .QN(n4702) );
  DFFNSRX2TS \dataOut_reg[1]  ( .D(n2427), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[1]), .QN(n4693) );
  DFFNSRX2TS \dataOut_reg[2]  ( .D(n2426), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[2]), .QN(n4684) );
  DFFNSRX2TS \dataOut_reg[3]  ( .D(n2425), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[3]), .QN(n4675) );
  DFFNSRX2TS \dataOut_reg[4]  ( .D(n2424), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[4]), .QN(n4666) );
  DFFNSRX2TS \dataOut_reg[5]  ( .D(n2423), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[5]), .QN(n4657) );
  DFFNSRX2TS \dataOut_reg[6]  ( .D(n2422), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[6]), .QN(n4648) );
  DFFNSRX2TS \dataOut_reg[7]  ( .D(n2421), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[7]), .QN(n4639) );
  DFFNSRX2TS \dataOut_reg[8]  ( .D(n2420), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[8]), .QN(n4630) );
  DFFNSRX2TS \dataOut_reg[9]  ( .D(n2419), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[9]), .QN(n4621) );
  DFFNSRX2TS \dataOut_reg[10]  ( .D(n2418), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[10]), .QN(n4612) );
  DFFNSRX2TS \dataOut_reg[11]  ( .D(n2417), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[11]), .QN(n4603) );
  DFFNSRX2TS \dataOut_reg[12]  ( .D(n2416), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[12]), .QN(n4594) );
  DFFNSRX2TS \dataOut_reg[13]  ( .D(n2415), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[13]), .QN(n4585) );
  DFFNSRX2TS \dataOut_reg[14]  ( .D(n2414), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[14]), .QN(n4576) );
  DFFNSRX2TS \dataOut_reg[15]  ( .D(n2413), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[15]), .QN(n4567) );
  DFFNSRX2TS \dataOut_reg[16]  ( .D(n2412), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[16]), .QN(n4558) );
  DFFNSRX2TS \dataOut_reg[17]  ( .D(n2411), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[17]), .QN(n4549) );
  DFFNSRX2TS \dataOut_reg[18]  ( .D(n2410), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[18]), .QN(n4540) );
  DFFNSRX2TS \dataOut_reg[19]  ( .D(n2409), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[19]), .QN(n4531) );
  DFFNSRX2TS \dataOut_reg[20]  ( .D(n2408), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[20]), .QN(n4522) );
  DFFNSRX2TS \dataOut_reg[21]  ( .D(n2407), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[21]), .QN(n4513) );
  DFFNSRX2TS \dataOut_reg[22]  ( .D(n2406), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[22]), .QN(n4504) );
  DFFNSRX2TS \dataOut_reg[23]  ( .D(n2405), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[23]), .QN(n4495) );
  DFFNSRX2TS \dataOut_reg[24]  ( .D(n2404), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[24]), .QN(n4486) );
  DFFNSRX2TS \dataOut_reg[25]  ( .D(n2403), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[25]), .QN(n4477) );
  DFFNSRX2TS \dataOut_reg[26]  ( .D(n2402), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[26]), .QN(n4468) );
  DFFNSRX2TS \dataOut_reg[27]  ( .D(n2401), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[27]), .QN(n4459) );
  DFFNSRX2TS \dataOut_reg[28]  ( .D(n2400), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[28]), .QN(n4450) );
  DFFNSRX2TS \dataOut_reg[29]  ( .D(n2399), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[29]), .QN(n4441) );
  DFFNSRX2TS \dataOut_reg[30]  ( .D(n2398), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[30]), .QN(n4432) );
  DFFNSRX2TS \dataOut_reg[31]  ( .D(n2397), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[31]), .QN(n4423) );
  DFFNSRX2TS \destinationAddressOut_reg[6]  ( .D(n2448), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[6]) );
  DFFNSRX2TS \destinationAddressOut_reg[7]  ( .D(n2447), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[7]) );
  DFFNSRX2TS \destinationAddressOut_reg[8]  ( .D(n2446), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[8]) );
  DFFNSRX2TS \destinationAddressOut_reg[9]  ( .D(n2445), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[9]) );
  DFFNSRX2TS \destinationAddressOut_reg[10]  ( .D(n2444), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[10]) );
  DFFNSRX2TS \destinationAddressOut_reg[11]  ( .D(n2443), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[11]) );
  DFFNSRX2TS \destinationAddressOut_reg[12]  ( .D(n2442), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[12]) );
  DFFNSRX2TS \destinationAddressOut_reg[13]  ( .D(n2441), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[13]) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][6]  ( .D(n2486), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4831) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][8]  ( .D(n2484), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4811) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][7]  ( .D(n2485), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4824) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][6]  ( .D(n2472), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4830) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][7]  ( .D(n2471), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4818) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][8]  ( .D(n2470), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4810) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][9]  ( .D(n2469), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4806) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][10]  ( .D(n2468), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4794) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][11]  ( .D(n2467), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4788) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][12]  ( .D(n2466), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4778) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][13]  ( .D(n2465), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4770) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][4]  ( .D(n2530), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4730) );
  DFFNSRXLTS \dataoutbuffer_reg[5][0]  ( .D(n2674), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4710) );
  DFFNSRXLTS \dataoutbuffer_reg[5][2]  ( .D(n2672), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4688) );
  DFFNSRXLTS \dataoutbuffer_reg[5][3]  ( .D(n2671), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4683) );
  DFFNSRXLTS \dataoutbuffer_reg[5][4]  ( .D(n2670), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4672) );
  DFFNSRXLTS \dataoutbuffer_reg[5][5]  ( .D(n2669), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4665) );
  DFFNSRXLTS \dataoutbuffer_reg[5][6]  ( .D(n2668), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4652) );
  DFFNSRXLTS \dataoutbuffer_reg[5][7]  ( .D(n2667), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4645) );
  DFFNSRXLTS \dataoutbuffer_reg[5][8]  ( .D(n2666), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4636) );
  DFFNSRXLTS \dataoutbuffer_reg[5][9]  ( .D(n2665), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4625) );
  DFFNSRXLTS \dataoutbuffer_reg[5][10]  ( .D(n2664), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4614) );
  DFFNSRXLTS \dataoutbuffer_reg[5][12]  ( .D(n2662), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4600) );
  DFFNSRXLTS \dataoutbuffer_reg[5][13]  ( .D(n2661), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4591) );
  DFFNSRXLTS \dataoutbuffer_reg[5][14]  ( .D(n2660), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4578) );
  DFFNSRXLTS \dataoutbuffer_reg[5][17]  ( .D(n2657), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4555) );
  DFFNSRXLTS \dataoutbuffer_reg[5][18]  ( .D(n2656), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4544) );
  DFFNSRXLTS \dataoutbuffer_reg[5][19]  ( .D(n2655), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4537) );
  DFFNSRXLTS \dataoutbuffer_reg[5][20]  ( .D(n2654), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4524) );
  DFFNSRXLTS \dataoutbuffer_reg[5][21]  ( .D(n2653), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4517) );
  DFFNSRXLTS \dataoutbuffer_reg[5][22]  ( .D(n2652), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4510) );
  DFFNSRXLTS \dataoutbuffer_reg[5][23]  ( .D(n2651), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4499) );
  DFFNSRXLTS \dataoutbuffer_reg[5][24]  ( .D(n2650), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4492) );
  DFFNSRXLTS \dataoutbuffer_reg[5][25]  ( .D(n2649), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4485) );
  DFFNSRXLTS \dataoutbuffer_reg[5][26]  ( .D(n2648), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4470) );
  DFFNSRXLTS \dataoutbuffer_reg[5][27]  ( .D(n2647), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4461) );
  DFFNSRXLTS \dataoutbuffer_reg[5][28]  ( .D(n2646), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4458) );
  DFFNSRXLTS \dataoutbuffer_reg[5][29]  ( .D(n2645), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4447) );
  DFFNSRXLTS \dataoutbuffer_reg[5][30]  ( .D(n2644), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4436) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][0]  ( .D(n2534), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4764) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][1]  ( .D(n2533), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4757) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][2]  ( .D(n2532), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4748) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][3]  ( .D(n2531), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4739) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][5]  ( .D(n2529), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4721) );
  DFFNSRXLTS \dataoutbuffer_reg[5][1]  ( .D(n2673), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4698) );
  DFFNSRXLTS \dataoutbuffer_reg[5][11]  ( .D(n2663), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4606) );
  DFFNSRXLTS \dataoutbuffer_reg[5][15]  ( .D(n2659), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4568) );
  DFFNSRXLTS \dataoutbuffer_reg[5][16]  ( .D(n2658), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4563) );
  DFFNSRXLTS \dataoutbuffer_reg[5][31]  ( .D(n2643), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4428) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][4]  ( .D(n2516), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4729) );
  DFFNSRXLTS \dataoutbuffer_reg[4][3]  ( .D(n2703), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4682) );
  DFFNSRXLTS \dataoutbuffer_reg[4][14]  ( .D(n2692), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4583) );
  DFFNSRXLTS \dataoutbuffer_reg[4][15]  ( .D(n2691), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4574) );
  DFFNSRXLTS \dataoutbuffer_reg[4][17]  ( .D(n2689), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4556) );
  DFFNSRXLTS \dataoutbuffer_reg[1][0]  ( .D(n2802), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4709) );
  DFFNSRXLTS \dataoutbuffer_reg[4][0]  ( .D(n2706), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4706) );
  DFFNSRXLTS \dataoutbuffer_reg[4][1]  ( .D(n2705), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4695) );
  DFFNSRXLTS \dataoutbuffer_reg[4][6]  ( .D(n2700), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4654) );
  DFFNSRXLTS \dataoutbuffer_reg[4][8]  ( .D(n2698), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4632) );
  DFFNSRXLTS \dataoutbuffer_reg[4][10]  ( .D(n2696), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4616) );
  DFFNSRXLTS \dataoutbuffer_reg[4][11]  ( .D(n2695), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4609) );
  DFFNSRXLTS \dataoutbuffer_reg[4][12]  ( .D(n2694), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4598) );
  DFFNSRXLTS \dataoutbuffer_reg[4][16]  ( .D(n2690), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4560) );
  DFFNSRXLTS \dataoutbuffer_reg[4][19]  ( .D(n2687), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4533) );
  DFFNSRXLTS \dataoutbuffer_reg[4][20]  ( .D(n2686), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4528) );
  DFFNSRXLTS \dataoutbuffer_reg[4][21]  ( .D(n2685), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4519) );
  DFFNSRXLTS \dataoutbuffer_reg[4][22]  ( .D(n2684), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4508) );
  DFFNSRXLTS \dataoutbuffer_reg[4][29]  ( .D(n2677), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4449) );
  DFFNSRXLTS \dataoutbuffer_reg[4][31]  ( .D(n2675), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4425) );
  DFFNSRXLTS \dataoutbuffer_reg[1][1]  ( .D(n2801), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4697) );
  DFFNSRXLTS \dataoutbuffer_reg[1][3]  ( .D(n2799), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4679) );
  DFFNSRXLTS \dataoutbuffer_reg[1][4]  ( .D(n2798), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4674) );
  DFFNSRXLTS \dataoutbuffer_reg[1][6]  ( .D(n2796), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4650) );
  DFFNSRXLTS \dataoutbuffer_reg[1][7]  ( .D(n2795), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4647) );
  DFFNSRXLTS \dataoutbuffer_reg[1][9]  ( .D(n2793), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4623) );
  DFFNSRXLTS \dataoutbuffer_reg[1][11]  ( .D(n2791), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4605) );
  DFFNSRXLTS \dataoutbuffer_reg[1][12]  ( .D(n2790), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4602) );
  DFFNSRXLTS \dataoutbuffer_reg[1][13]  ( .D(n2789), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4593) );
  DFFNSRXLTS \dataoutbuffer_reg[1][14]  ( .D(n2788), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4580) );
  DFFNSRXLTS \dataoutbuffer_reg[1][15]  ( .D(n2787), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4573) );
  DFFNSRXLTS \dataoutbuffer_reg[1][16]  ( .D(n2786), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4566) );
  DFFNSRXLTS \dataoutbuffer_reg[1][17]  ( .D(n2785), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4551) );
  DFFNSRXLTS \dataoutbuffer_reg[1][18]  ( .D(n2784), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4548) );
  DFFNSRXLTS \dataoutbuffer_reg[1][21]  ( .D(n2781), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4515) );
  DFFNSRXLTS \dataoutbuffer_reg[1][23]  ( .D(n2779), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4497) );
  DFFNSRXLTS \dataoutbuffer_reg[1][24]  ( .D(n2778), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4488) );
  DFFNSRXLTS \dataoutbuffer_reg[1][25]  ( .D(n2777), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4483) );
  DFFNSRXLTS \dataoutbuffer_reg[1][26]  ( .D(n2776), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4476) );
  DFFNSRXLTS \dataoutbuffer_reg[1][28]  ( .D(n2774), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4452) );
  DFFNSRXLTS \dataoutbuffer_reg[1][29]  ( .D(n2773), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4445) );
  DFFNSRXLTS \dataoutbuffer_reg[1][30]  ( .D(n2772), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4440) );
  DFFNSRXLTS \dataoutbuffer_reg[1][31]  ( .D(n2771), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4431) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][0]  ( .D(n2478), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4768) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][1]  ( .D(n2477), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4759) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][2]  ( .D(n2476), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4750) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][3]  ( .D(n2475), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4737) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][5]  ( .D(n2473), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4717) );
  DFFNSRXLTS \dataoutbuffer_reg[4][2]  ( .D(n2704), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4687) );
  DFFNSRXLTS \dataoutbuffer_reg[4][4]  ( .D(n2702), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4671) );
  DFFNSRXLTS \dataoutbuffer_reg[4][5]  ( .D(n2701), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4660) );
  DFFNSRXLTS \dataoutbuffer_reg[4][7]  ( .D(n2699), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4644) );
  DFFNSRXLTS \dataoutbuffer_reg[4][9]  ( .D(n2697), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4626) );
  DFFNSRXLTS \dataoutbuffer_reg[4][13]  ( .D(n2693), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4586) );
  DFFNSRXLTS \dataoutbuffer_reg[4][18]  ( .D(n2688), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4541) );
  DFFNSRXLTS \dataoutbuffer_reg[4][23]  ( .D(n2683), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4498) );
  DFFNSRXLTS \dataoutbuffer_reg[4][24]  ( .D(n2682), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4487) );
  DFFNSRXLTS \dataoutbuffer_reg[4][25]  ( .D(n2681), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4482) );
  DFFNSRXLTS \dataoutbuffer_reg[4][26]  ( .D(n2680), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4469) );
  DFFNSRXLTS \dataoutbuffer_reg[4][27]  ( .D(n2679), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4462) );
  DFFNSRXLTS \dataoutbuffer_reg[4][28]  ( .D(n2678), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4451) );
  DFFNSRXLTS \dataoutbuffer_reg[4][30]  ( .D(n2676), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4433) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][0]  ( .D(n2520), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4761) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][1]  ( .D(n2519), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4756) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][2]  ( .D(n2518), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4743) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][3]  ( .D(n2517), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4738) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][5]  ( .D(n2515), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4718) );
  DFFNSRXLTS \dataoutbuffer_reg[1][2]  ( .D(n2800), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4685) );
  DFFNSRXLTS \dataoutbuffer_reg[1][5]  ( .D(n2797), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4658) );
  DFFNSRXLTS \dataoutbuffer_reg[1][8]  ( .D(n2794), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4633) );
  DFFNSRXLTS \dataoutbuffer_reg[1][10]  ( .D(n2792), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4619) );
  DFFNSRXLTS \dataoutbuffer_reg[1][19]  ( .D(n2783), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4536) );
  DFFNSRXLTS \dataoutbuffer_reg[1][20]  ( .D(n2782), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4525) );
  DFFNSRXLTS \dataoutbuffer_reg[1][22]  ( .D(n2780), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4509) );
  DFFNSRXLTS \dataoutbuffer_reg[1][27]  ( .D(n2775), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4460) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][4]  ( .D(n2474), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4726) );
  DFFNSRXLTS \dataoutbuffer_reg[3][7]  ( .D(n2731), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n6312), .QN(n4646) );
  DFFNSRXLTS \dataoutbuffer_reg[3][2]  ( .D(n2736), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n6302), .QN(n4690) );
  DFFNSRXLTS \dataoutbuffer_reg[3][4]  ( .D(n2734), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n6301), .QN(n4670) );
  DFFNSRXLTS \dataoutbuffer_reg[3][5]  ( .D(n2733), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n6300), .QN(n4663) );
  DFFNSRXLTS \dataoutbuffer_reg[3][13]  ( .D(n2725), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6299), .QN(n4589) );
  DFFNSRXLTS \dataoutbuffer_reg[3][15]  ( .D(n2723), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6298), .QN(n4571) );
  DFFNSRXLTS \dataoutbuffer_reg[3][18]  ( .D(n2720), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6297), .QN(n4546) );
  DFFNSRXLTS \dataoutbuffer_reg[3][20]  ( .D(n2718), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6296), .QN(n4530) );
  DFFNSRXLTS \dataoutbuffer_reg[3][23]  ( .D(n2715), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6295), .QN(n4503) );
  DFFNSRXLTS \dataoutbuffer_reg[3][25]  ( .D(n2713), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6294), .QN(n4479) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][2]  ( .D(n2504), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n6293), .QN(n4744) );
  DFFNSRXLTS \dataoutbuffer_reg[3][0]  ( .D(n2738), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n6281), .QN(n4703) );
  DFFNSRXLTS \dataoutbuffer_reg[3][1]  ( .D(n2737), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n6280), .QN(n4694) );
  DFFNSRXLTS \dataoutbuffer_reg[3][3]  ( .D(n2735), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n6279), .QN(n4680) );
  DFFNSRXLTS \dataoutbuffer_reg[3][6]  ( .D(n2732), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n6278), .QN(n4653) );
  DFFNSRXLTS \dataoutbuffer_reg[3][8]  ( .D(n2730), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n6277), .QN(n4631) );
  DFFNSRXLTS \dataoutbuffer_reg[3][9]  ( .D(n2729), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n6276), .QN(n4624) );
  DFFNSRXLTS \dataoutbuffer_reg[3][10]  ( .D(n2728), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6275), .QN(n4615) );
  DFFNSRXLTS \dataoutbuffer_reg[3][11]  ( .D(n2727), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6274), .QN(n4608) );
  DFFNSRXLTS \dataoutbuffer_reg[3][12]  ( .D(n2726), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6273), .QN(n4597) );
  DFFNSRXLTS \dataoutbuffer_reg[3][14]  ( .D(n2724), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6272), .QN(n4581) );
  DFFNSRXLTS \dataoutbuffer_reg[3][16]  ( .D(n2722), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6271), .QN(n4559) );
  DFFNSRXLTS \dataoutbuffer_reg[3][17]  ( .D(n2721), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6270), .QN(n4550) );
  DFFNSRXLTS \dataoutbuffer_reg[3][19]  ( .D(n2719), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6269), .QN(n4538) );
  DFFNSRXLTS \dataoutbuffer_reg[3][21]  ( .D(n2717), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6268), .QN(n4518) );
  DFFNSRXLTS \dataoutbuffer_reg[3][22]  ( .D(n2716), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6267), .QN(n4507) );
  DFFNSRXLTS \dataoutbuffer_reg[3][24]  ( .D(n2714), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6266), .QN(n4491) );
  DFFNSRXLTS \dataoutbuffer_reg[3][26]  ( .D(n2712), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6265), .QN(n4475) );
  DFFNSRXLTS \dataoutbuffer_reg[3][27]  ( .D(n2711), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6264), .QN(n4464) );
  DFFNSRXLTS \dataoutbuffer_reg[3][28]  ( .D(n2710), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6263), .QN(n4455) );
  DFFNSRXLTS \dataoutbuffer_reg[3][29]  ( .D(n2709), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6262), .QN(n4444) );
  DFFNSRXLTS \dataoutbuffer_reg[3][30]  ( .D(n2708), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6261), .QN(n4439) );
  DFFNSRXLTS \dataoutbuffer_reg[3][31]  ( .D(n2707), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6260), .QN(n4426) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][0]  ( .D(n2506), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n6259), .QN(n4765) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][1]  ( .D(n2505), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n6258), .QN(n4758) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][3]  ( .D(n2503), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n6257), .QN(n4740) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][4]  ( .D(n2502), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n6256), .QN(n4727) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][5]  ( .D(n2501), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n6255), .QN(n4722) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][0]  ( .D(n2858), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][0] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][1]  ( .D(n2857), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][1] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][2]  ( .D(n2856), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][2] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][3]  ( .D(n2855), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][3] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][5]  ( .D(n2853), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][5] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][4]  ( .D(n2854), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][4] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[5][0]  ( .D(n2870), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6310) );
  DFFNSRXLTS \requesterAddressbuffer_reg[5][1]  ( .D(n2869), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6309) );
  DFFNSRXLTS \requesterAddressbuffer_reg[5][2]  ( .D(n2868), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6308) );
  DFFNSRXLTS \requesterAddressbuffer_reg[5][3]  ( .D(n2867), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6307) );
  DFFNSRXLTS \requesterAddressbuffer_reg[5][4]  ( .D(n2866), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6306) );
  DFFNSRXLTS \requesterAddressbuffer_reg[5][5]  ( .D(n2865), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6305) );
  DFFNSRXLTS \requesterAddressbuffer_reg[4][4]  ( .D(n2860), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6304) );
  DFFNSRXLTS \requesterAddressbuffer_reg[4][5]  ( .D(n2859), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6303) );
  DFFNSRXLTS \requesterAddressbuffer_reg[4][0]  ( .D(n2864), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6285) );
  DFFNSRXLTS \requesterAddressbuffer_reg[4][1]  ( .D(n2863), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6284) );
  DFFNSRXLTS \requesterAddressbuffer_reg[4][2]  ( .D(n2862), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6283) );
  DFFNSRXLTS \requesterAddressbuffer_reg[4][3]  ( .D(n2861), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6282) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][0]  ( .D(n2846), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6292) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][1]  ( .D(n2845), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6291) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][2]  ( .D(n2844), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6290) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][3]  ( .D(n2843), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6289) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][4]  ( .D(n2842), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6288) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][5]  ( .D(n2841), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n6287) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][9]  ( .D(n2455), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4803) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][11]  ( .D(n2453), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4789) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][10]  ( .D(n2454), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4798) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][12]  ( .D(n2452), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4777) );
  DFFNSRXLTS \writeOutbuffer_reg[2]  ( .D(n2573), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[2]), .QN(n6311) );
  DFFNSRXLTS \writeOutbuffer_reg[1]  ( .D(n2572), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[1]), .QN(n6286) );
  DFFNSRX2TS \read_reg_reg[1]  ( .D(n2883), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n5), .QN(n335) );
  DFFNSRX2TS \read_reg_reg[2]  ( .D(n2884), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n3), .QN(n333) );
  DFFNSRXLTS full_reg_reg ( .D(N4718), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        n4836), .QN(n6347) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][13]  ( .D(n2479), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4769) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][13]  ( .D(n2451), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4776) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][12]  ( .D(n2480), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4783) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][11]  ( .D(n2481), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4792) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][10]  ( .D(n2482), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4797) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][9]  ( .D(n2483), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n4808) );
  DFFNSRXLTS empty_reg_reg ( .D(n2885), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        n6253), .QN(n4834) );
  DFFNSRXLTS \write_reg_reg[0]  ( .D(n2888), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n16), .QN(n5327) );
  DFFNSRXLTS \write_reg_reg[2]  ( .D(n2886), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n7), .QN(n5326) );
  DFFNSRXLTS \dataoutbuffer_reg[7][0]  ( .D(n2610), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n4704) );
  DFFNSRXLTS \dataoutbuffer_reg[7][15]  ( .D(n2595), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4569) );
  DFFNSRXLTS \dataoutbuffer_reg[7][14]  ( .D(n2596), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4584) );
  DFFNSRXLTS \dataoutbuffer_reg[7][13]  ( .D(n2597), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4587) );
  DFFNSRXLTS \dataoutbuffer_reg[6][29]  ( .D(n2613), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4446) );
  DFFNSRXLTS \dataoutbuffer_reg[6][28]  ( .D(n2614), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4454) );
  DFFNSRXLTS \dataoutbuffer_reg[6][27]  ( .D(n2615), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4463) );
  DFFNSRXLTS \dataoutbuffer_reg[6][26]  ( .D(n2616), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4474) );
  DFFNSRXLTS \dataoutbuffer_reg[6][25]  ( .D(n2617), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4484) );
  DFFNSRXLTS \dataoutbuffer_reg[6][24]  ( .D(n2618), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4494) );
  DFFNSRXLTS \dataoutbuffer_reg[6][23]  ( .D(n2619), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4496) );
  DFFNSRXLTS \dataoutbuffer_reg[6][22]  ( .D(n2620), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4512) );
  DFFNSRXLTS \dataoutbuffer_reg[6][21]  ( .D(n2621), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4516) );
  DFFNSRXLTS \dataoutbuffer_reg[6][20]  ( .D(n2622), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4523) );
  DFFNSRXLTS \dataoutbuffer_reg[6][19]  ( .D(n2623), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4535) );
  DFFNSRXLTS \dataoutbuffer_reg[6][18]  ( .D(n2624), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4547) );
  DFFNSRXLTS \dataoutbuffer_reg[6][17]  ( .D(n2625), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4557) );
  DFFNSRXLTS \dataoutbuffer_reg[6][16]  ( .D(n2626), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4562) );
  DFFNSRXLTS \dataoutbuffer_reg[6][15]  ( .D(n2627), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4575) );
  DFFNSRXLTS \dataoutbuffer_reg[6][14]  ( .D(n2628), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4582) );
  DFFNSRXLTS \dataoutbuffer_reg[6][13]  ( .D(n2629), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4590) );
  DFFNSRXLTS \dataoutbuffer_reg[6][12]  ( .D(n2630), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n4601) );
  INVX2TS U2 ( .A(selectBit_SOUTH), .Y(n189) );
  INVX2TS U3 ( .A(n278), .Y(n205) );
  INVXLTS U4 ( .A(n5438), .Y(n334) );
  NAND3XLTS U5 ( .A(n5486), .B(n5438), .C(n6332), .Y(n5548) );
  INVX4TS U6 ( .A(n5438), .Y(n6331) );
  XOR2X4TS U7 ( .A(n5321), .B(n7), .Y(n5438) );
  BUFX2TS U8 ( .A(n684), .Y(n673) );
  BUFX4TS U9 ( .A(n611), .Y(n610) );
  CLKBUFX2TS U10 ( .A(n680), .Y(n678) );
  XOR2X1TS U11 ( .A(n121), .B(n6248), .Y(n5346) );
  AND2X2TS U12 ( .A(n5523), .B(n6336), .Y(n6126) );
  AND3X2TS U13 ( .A(n172), .B(n5520), .C(n113), .Y(n6123) );
  AOI21X1TS U14 ( .A0(n342), .A1(n5356), .B0(n429), .Y(n5523) );
  INVX2TS U15 ( .A(n5391), .Y(n6332) );
  NOR2BX1TS U16 ( .AN(n5346), .B(n6236), .Y(n5486) );
  NAND3X1TS U17 ( .A(n5463), .B(n5438), .C(n6332), .Y(n5417) );
  OA21X2TS U18 ( .A0(n157), .A1(n5416), .B0(n5515), .Y(n5512) );
  NOR2BX1TS U19 ( .AN(n5523), .B(n5518), .Y(n6124) );
  CLKBUFX2TS U20 ( .A(n6187), .Y(n3372) );
  NOR3X1TS U21 ( .A(n6323), .B(n196), .C(n5316), .Y(n5561) );
  CLKBUFX2TS U22 ( .A(n3338), .Y(n3327) );
  CLKBUFX2TS U23 ( .A(n5523), .Y(n113) );
  NOR3X1TS U24 ( .A(n5555), .B(n5556), .C(n5553), .Y(n5554) );
  CLKBUFX2TS U25 ( .A(n3282), .Y(n3281) );
  CLKBUFX2TS U26 ( .A(n3236), .Y(n3235) );
  CLKBUFX2TS U27 ( .A(n3432), .Y(n3430) );
  AOI222XLTS U28 ( .A0(n206), .A1(n54), .B0(n3949), .B1(n678), .C0(n4418), 
        .C1(n3797), .Y(n5336) );
  AOI222XLTS U29 ( .A0(n3973), .A1(n1894), .B0(n4286), .B1(n221), .C0(n4130), 
        .C1(n414), .Y(n5397) );
  NOR2X1TS U30 ( .A(n215), .B(n6325), .Y(n5392) );
  AND2X2TS U31 ( .A(n5555), .B(n165), .Y(n6202) );
  OA22X1TS U32 ( .A0(n5542), .A1(n188), .B0(n204), .B1(n153), .Y(n426) );
  OA22X1TS U33 ( .A0(n5547), .A1(n188), .B0(n5488), .B1(n153), .Y(n425) );
  OR2X2TS U34 ( .A(n6226), .B(n194), .Y(n1) );
  AND2X2TS U35 ( .A(n5556), .B(n5559), .Y(n6200) );
  AND2X2TS U36 ( .A(n5566), .B(n5561), .Y(n6217) );
  OA21XLTS U37 ( .A0(n5440), .A1(n5439), .B0(n5548), .Y(n5547) );
  INVX2TS U38 ( .A(n171), .Y(n172) );
  AND3XLTS U39 ( .A(n5463), .B(n5391), .C(n6331), .Y(n5525) );
  INVXLTS U40 ( .A(n5548), .Y(n6333) );
  INVXLTS U41 ( .A(n5532), .Y(n156) );
  INVX1TS U42 ( .A(n5532), .Y(n6323) );
  OAI22X2TS U43 ( .A0(n5512), .A1(n187), .B0(n203), .B1(n6318), .Y(n5569) );
  INVX1TS U44 ( .A(n205), .Y(n206) );
  NAND3XLTS U45 ( .A(n5523), .B(n217), .C(n5519), .Y(n5572) );
  INVXLTS U46 ( .A(n5520), .Y(n6336) );
  OA21XLTS U47 ( .A0(n6325), .A1(n5439), .B0(n5520), .Y(n5519) );
  NAND3X1TS U48 ( .A(n337), .B(n5486), .C(n334), .Y(n5520) );
  INVX1TS U49 ( .A(n5440), .Y(n6325) );
  CLKBUFX2TS U50 ( .A(n3289), .Y(n3282) );
  CLKBUFX2TS U51 ( .A(n6184), .Y(n3324) );
  CLKBUFX2TS U52 ( .A(n6340), .Y(n3688) );
  OA22X1TS U53 ( .A0(n5554), .A1(n418), .B0(n201), .B1(n203), .Y(n427) );
  CLKBUFX2TS U54 ( .A(n6108), .Y(n625) );
  OA22X1TS U55 ( .A0(n5519), .A1(n188), .B0(n5488), .B1(n6318), .Y(n429) );
  NOR2BX1TS U56 ( .AN(n5552), .B(n5518), .Y(n6185) );
  CLKBUFX2TS U57 ( .A(n6126), .Y(n769) );
  CLKBUFX2TS U58 ( .A(n805), .Y(n798) );
  OAI21X1TS U59 ( .A0(n5317), .A1(n157), .B0(n6324), .Y(n5440) );
  AOI21X1TS U60 ( .A0(n342), .A1(n154), .B0(n425), .Y(n5552) );
  OA22X1TS U61 ( .A0(n5560), .A1(n187), .B0(n201), .B1(n5488), .Y(n428) );
  CLKBUFX2TS U62 ( .A(n6219), .Y(n3498) );
  CLKBUFX2TS U63 ( .A(n3455), .Y(n3449) );
  AOI21X1TS U64 ( .A0(n176), .A1(n5449), .B0(n426), .Y(n5545) );
  CLKBUFX2TS U65 ( .A(n3438), .Y(n3432) );
  AOI21X1TS U66 ( .A0(n176), .A1(n200), .B0(n158), .Y(n5322) );
  NAND2X1TS U67 ( .A(n5527), .B(n5530), .Y(n5575) );
  OAI21X1TS U68 ( .A0(n5487), .A1(n5539), .B0(n5417), .Y(n5540) );
  NOR3BX1TS U69 ( .AN(n5463), .B(n6331), .C(n6332), .Y(n5553) );
  CLKBUFX2TS U70 ( .A(n5559), .Y(n165) );
  AOI21X2TS U71 ( .A0(n5536), .A1(n5392), .B0(n6334), .Y(n5534) );
  CLKBUFX2TS U72 ( .A(n837), .Y(n831) );
  CLKBUFX2TS U73 ( .A(n3407), .Y(n3401) );
  CLKBUFX2TS U74 ( .A(n3466), .Y(n3465) );
  CLKBUFX2TS U75 ( .A(n3406), .Y(n3392) );
  CLKBUFX2TS U76 ( .A(n3500), .Y(n3497) );
  CLKBUFX2TS U77 ( .A(n3371), .Y(n3364) );
  CLKBUFX2TS U78 ( .A(n3365), .Y(n3363) );
  AOI222XLTS U79 ( .A0(n3859), .A1(n3676), .B0(n385), .B1(n3412), .C0(n4015), 
        .C1(n3395), .Y(n5688) );
  AOI222XLTS U80 ( .A0(n3862), .A1(n3677), .B0(n383), .B1(n3412), .C0(n4018), 
        .C1(n3396), .Y(n5686) );
  AOI222XLTS U81 ( .A0(n3865), .A1(n3677), .B0(n381), .B1(n3413), .C0(n4021), 
        .C1(n3396), .Y(n5684) );
  AOI222XLTS U82 ( .A0(n3868), .A1(n3677), .B0(n379), .B1(n3413), .C0(n4024), 
        .C1(n3396), .Y(n5682) );
  AOI222XLTS U83 ( .A0(n3871), .A1(n3677), .B0(n377), .B1(n3413), .C0(n4027), 
        .C1(n3397), .Y(n5680) );
  AOI222XLTS U84 ( .A0(n3874), .A1(n3678), .B0(n375), .B1(n3413), .C0(n4030), 
        .C1(n3397), .Y(n5678) );
  AOI222XLTS U85 ( .A0(n3877), .A1(n3678), .B0(n374), .B1(n3414), .C0(n4033), 
        .C1(n3397), .Y(n5676) );
  AOI222XLTS U86 ( .A0(n3880), .A1(n3678), .B0(n371), .B1(n3414), .C0(n4036), 
        .C1(n3397), .Y(n5674) );
  AOI222XLTS U87 ( .A0(n3883), .A1(n3678), .B0(n369), .B1(n3414), .C0(n4039), 
        .C1(n3398), .Y(n5672) );
  AOI222XLTS U88 ( .A0(n3886), .A1(n3679), .B0(n367), .B1(n3414), .C0(n4042), 
        .C1(n3398), .Y(n5670) );
  AOI222XLTS U89 ( .A0(n3889), .A1(n3679), .B0(n365), .B1(n3415), .C0(n4045), 
        .C1(n3398), .Y(n5668) );
  AOI222XLTS U90 ( .A0(n3892), .A1(n3679), .B0(n363), .B1(n3415), .C0(n4048), 
        .C1(n3398), .Y(n5666) );
  AOI222XLTS U91 ( .A0(n3895), .A1(n3680), .B0(n361), .B1(n3415), .C0(n4051), 
        .C1(n3399), .Y(n5664) );
  AOI222XLTS U92 ( .A0(n3898), .A1(n3680), .B0(n360), .B1(n3415), .C0(n4054), 
        .C1(n3399), .Y(n5662) );
  AOI222XLTS U93 ( .A0(n3901), .A1(n3680), .B0(n357), .B1(n3419), .C0(n4057), 
        .C1(n3399), .Y(n5660) );
  AOI222XLTS U94 ( .A0(n3904), .A1(n3680), .B0(n355), .B1(n3419), .C0(n4060), 
        .C1(n3399), .Y(n5658) );
  AOI222XLTS U95 ( .A0(n3907), .A1(n3681), .B0(n353), .B1(n3419), .C0(n4063), 
        .C1(n3400), .Y(n5656) );
  AOI222XLTS U96 ( .A0(n3910), .A1(n3681), .B0(n351), .B1(n3420), .C0(n4066), 
        .C1(n3400), .Y(n5654) );
  AOI222XLTS U97 ( .A0(n4018), .A1(n3491), .B0(n384), .B1(n3478), .C0(n4174), 
        .C1(n3463), .Y(n5622) );
  AOI222XLTS U98 ( .A0(n4021), .A1(n3491), .B0(n382), .B1(n3477), .C0(n4177), 
        .C1(n3463), .Y(n5620) );
  AOI222XLTS U99 ( .A0(n4024), .A1(n3492), .B0(n380), .B1(n3477), .C0(n4180), 
        .C1(n3463), .Y(n5618) );
  AOI222XLTS U100 ( .A0(n3979), .A1(n3488), .B0(n410), .B1(n3481), .C0(n4135), 
        .C1(n3459), .Y(n5648) );
  AOI222XLTS U101 ( .A0(n3903), .A1(n761), .B0(n355), .B1(n738), .C0(n4216), 
        .C1(n715), .Y(n5978) );
  AOI222XLTS U102 ( .A0(n3888), .A1(n760), .B0(n365), .B1(n741), .C0(n4201), 
        .C1(n714), .Y(n5988) );
  AOI222XLTS U103 ( .A0(n3882), .A1(n759), .B0(n369), .B1(n741), .C0(n4195), 
        .C1(n714), .Y(n5992) );
  AOI222XLTS U104 ( .A0(n3879), .A1(n759), .B0(n371), .B1(n742), .C0(n4192), 
        .C1(n712), .Y(n5994) );
  AOI222XLTS U105 ( .A0(n3852), .A1(n756), .B0(n389), .B1(n747), .C0(n4165), 
        .C1(n732), .Y(n6012) );
  AOI222XLTS U106 ( .A0(n3846), .A1(n756), .B0(n393), .B1(n750), .C0(n4159), 
        .C1(n711), .Y(n6016) );
  AOI222XLTS U107 ( .A0(n3837), .A1(n755), .B0(n399), .B1(n746), .C0(n4150), 
        .C1(n711), .Y(n6022) );
  AOI222XLTS U108 ( .A0(n3828), .A1(n755), .B0(n405), .B1(n746), .C0(n4141), 
        .C1(n708), .Y(n6028) );
  AOI222XLTS U109 ( .A0(n3915), .A1(n769), .B0(n348), .B1(n739), .C0(n4228), 
        .C1(n716), .Y(n5970) );
  AOI222XLTS U110 ( .A0(n3912), .A1(n765), .B0(n349), .B1(n738), .C0(n4225), 
        .C1(n716), .Y(n5972) );
  AOI222XLTS U111 ( .A0(n3909), .A1(n761), .B0(n351), .B1(n739), .C0(n4222), 
        .C1(n716), .Y(n5974) );
  AOI222XLTS U112 ( .A0(n3906), .A1(n761), .B0(n353), .B1(n738), .C0(n4219), 
        .C1(n716), .Y(n5976) );
  AOI222XLTS U113 ( .A0(n3900), .A1(n761), .B0(n357), .B1(n740), .C0(n4213), 
        .C1(n715), .Y(n5980) );
  AOI222XLTS U114 ( .A0(n3897), .A1(n760), .B0(n359), .B1(n740), .C0(n4210), 
        .C1(n715), .Y(n5982) );
  AOI222XLTS U115 ( .A0(n3894), .A1(n760), .B0(n361), .B1(n739), .C0(n4207), 
        .C1(n715), .Y(n5984) );
  AOI222XLTS U116 ( .A0(n3891), .A1(n760), .B0(n363), .B1(n741), .C0(n4204), 
        .C1(n714), .Y(n5986) );
  AOI222XLTS U117 ( .A0(n3885), .A1(n759), .B0(n367), .B1(n739), .C0(n4198), 
        .C1(n714), .Y(n5990) );
  AOI222XLTS U118 ( .A0(n3876), .A1(n758), .B0(n373), .B1(n740), .C0(n4189), 
        .C1(n712), .Y(n5996) );
  AOI222XLTS U119 ( .A0(n3873), .A1(n758), .B0(n375), .B1(n742), .C0(n4186), 
        .C1(n712), .Y(n5998) );
  AOI222XLTS U120 ( .A0(n3870), .A1(n758), .B0(n378), .B1(n738), .C0(n4183), 
        .C1(n712), .Y(n6000) );
  AOI222XLTS U121 ( .A0(n3867), .A1(n758), .B0(n380), .B1(n741), .C0(n4180), 
        .C1(n735), .Y(n6002) );
  AOI222XLTS U122 ( .A0(n3864), .A1(n757), .B0(n381), .B1(n740), .C0(n4177), 
        .C1(n735), .Y(n6004) );
  AOI222XLTS U123 ( .A0(n3861), .A1(n757), .B0(n383), .B1(n743), .C0(n4174), 
        .C1(n732), .Y(n6006) );
  AOI222XLTS U124 ( .A0(n3858), .A1(n757), .B0(n385), .B1(n742), .C0(n4171), 
        .C1(n732), .Y(n6008) );
  AOI222XLTS U125 ( .A0(n3855), .A1(n757), .B0(n388), .B1(n747), .C0(n4168), 
        .C1(n732), .Y(n6010) );
  AOI222XLTS U126 ( .A0(n3849), .A1(n759), .B0(n391), .B1(n743), .C0(n4162), 
        .C1(n6124), .Y(n6014) );
  AOI222XLTS U127 ( .A0(n3843), .A1(n756), .B0(n395), .B1(n743), .C0(n4156), 
        .C1(n711), .Y(n6018) );
  AOI222XLTS U128 ( .A0(n3840), .A1(n756), .B0(n397), .B1(n743), .C0(n4153), 
        .C1(n734), .Y(n6020) );
  AOI222XLTS U129 ( .A0(n3834), .A1(n755), .B0(n401), .B1(n749), .C0(n4147), 
        .C1(n711), .Y(n6024) );
  AOI222XLTS U130 ( .A0(n3831), .A1(n755), .B0(n403), .B1(n6125), .C0(n4144), 
        .C1(n708), .Y(n6026) );
  AOI222XLTS U131 ( .A0(n3825), .A1(n754), .B0(n408), .B1(n747), .C0(n4138), 
        .C1(n708), .Y(n6030) );
  AOI222XLTS U132 ( .A0(n3822), .A1(n754), .B0(n410), .B1(n742), .C0(n4135), 
        .C1(n708), .Y(n6032) );
  AOI222XLTS U133 ( .A0(n4071), .A1(n3366), .B0(n347), .B1(n3342), .C0(n4228), 
        .C1(n3332), .Y(n5714) );
  AOI222XLTS U134 ( .A0(n4026), .A1(n3361), .B0(n377), .B1(n3349), .C0(n4183), 
        .C1(n3335), .Y(n5744) );
  AOI222XLTS U135 ( .A0(n4023), .A1(n3361), .B0(n379), .B1(n3352), .C0(n4180), 
        .C1(n3336), .Y(n5746) );
  AOI222XLTS U136 ( .A0(n4011), .A1(n3360), .B0(n387), .B1(n3344), .C0(n4168), 
        .C1(n3336), .Y(n5754) );
  AOI222XLTS U137 ( .A0(n3981), .A1(n3357), .B0(n407), .B1(n3345), .C0(n4138), 
        .C1(n3328), .Y(n5774) );
  AOI222XLTS U138 ( .A0(n4068), .A1(n3372), .B0(n350), .B1(n3349), .C0(n4225), 
        .C1(n3332), .Y(n5716) );
  AOI222XLTS U139 ( .A0(n4065), .A1(n3366), .B0(n352), .B1(n3342), .C0(n4222), 
        .C1(n3332), .Y(n5718) );
  AOI222XLTS U140 ( .A0(n4062), .A1(n3368), .B0(n354), .B1(n3353), .C0(n4219), 
        .C1(n3332), .Y(n5720) );
  AOI222XLTS U141 ( .A0(n4059), .A1(n3369), .B0(n356), .B1(n3352), .C0(n4216), 
        .C1(n3331), .Y(n5722) );
  AOI222XLTS U142 ( .A0(n4056), .A1(n3370), .B0(n358), .B1(n3353), .C0(n4213), 
        .C1(n3331), .Y(n5724) );
  AOI222XLTS U143 ( .A0(n4053), .A1(n3367), .B0(n360), .B1(n3354), .C0(n4210), 
        .C1(n3331), .Y(n5726) );
  AOI222XLTS U144 ( .A0(n4050), .A1(n3368), .B0(n362), .B1(n3342), .C0(n4207), 
        .C1(n3331), .Y(n5728) );
  AOI222XLTS U145 ( .A0(n4047), .A1(n3369), .B0(n364), .B1(n3353), .C0(n4204), 
        .C1(n3330), .Y(n5730) );
  AOI222XLTS U146 ( .A0(n4044), .A1(n3370), .B0(n366), .B1(n3351), .C0(n4201), 
        .C1(n3330), .Y(n5732) );
  AOI222XLTS U147 ( .A0(n4041), .A1(n3366), .B0(n368), .B1(n3342), .C0(n4198), 
        .C1(n3330), .Y(n5734) );
  AOI222XLTS U148 ( .A0(n4038), .A1(n3367), .B0(n370), .B1(n3350), .C0(n4195), 
        .C1(n3330), .Y(n5736) );
  AOI222XLTS U149 ( .A0(n4035), .A1(n3366), .B0(n372), .B1(n3352), .C0(n4192), 
        .C1(n3335), .Y(n5738) );
  AOI222XLTS U150 ( .A0(n4032), .A1(n3361), .B0(n374), .B1(n3354), .C0(n4189), 
        .C1(n3334), .Y(n5740) );
  AOI222XLTS U151 ( .A0(n4029), .A1(n3361), .B0(n376), .B1(n3352), .C0(n4186), 
        .C1(n3339), .Y(n5742) );
  AOI222XLTS U152 ( .A0(n4020), .A1(n3360), .B0(n382), .B1(n3355), .C0(n4177), 
        .C1(n3338), .Y(n5748) );
  AOI222XLTS U153 ( .A0(n4017), .A1(n3360), .B0(n384), .B1(n3343), .C0(n4174), 
        .C1(n3336), .Y(n5750) );
  AOI222XLTS U154 ( .A0(n4014), .A1(n3360), .B0(n386), .B1(n6186), .C0(n4171), 
        .C1(n3336), .Y(n5752) );
  AOI222XLTS U155 ( .A0(n4008), .A1(n3359), .B0(n390), .B1(n3344), .C0(n4165), 
        .C1(n3334), .Y(n5756) );
  AOI222XLTS U156 ( .A0(n4005), .A1(n3367), .B0(n392), .B1(n3343), .C0(n4162), 
        .C1(n3335), .Y(n5758) );
  AOI222XLTS U157 ( .A0(n4002), .A1(n3359), .B0(n394), .B1(n3344), .C0(n4159), 
        .C1(n3329), .Y(n5760) );
  AOI222XLTS U158 ( .A0(n3999), .A1(n3359), .B0(n396), .B1(n3343), .C0(n4156), 
        .C1(n3329), .Y(n5762) );
  AOI222XLTS U159 ( .A0(n3996), .A1(n3359), .B0(n398), .B1(n3343), .C0(n4153), 
        .C1(n3337), .Y(n5764) );
  AOI222XLTS U160 ( .A0(n3993), .A1(n3358), .B0(n400), .B1(n3345), .C0(n4150), 
        .C1(n3329), .Y(n5766) );
  AOI222XLTS U161 ( .A0(n3990), .A1(n3358), .B0(n402), .B1(n3345), .C0(n4147), 
        .C1(n3329), .Y(n5768) );
  AOI222XLTS U162 ( .A0(n3987), .A1(n3358), .B0(n404), .B1(n3344), .C0(n4144), 
        .C1(n3328), .Y(n5770) );
  AOI222XLTS U163 ( .A0(n3984), .A1(n3358), .B0(n406), .B1(n3345), .C0(n4141), 
        .C1(n3328), .Y(n5772) );
  AOI222XLTS U164 ( .A0(n3978), .A1(n3357), .B0(n409), .B1(n6186), .C0(n4135), 
        .C1(n3328), .Y(n5776) );
  AOI222XLTS U165 ( .A0(n3816), .A1(n3235), .B0(n3804), .B1(n3256), .C0(n3809), 
        .C1(n3281), .Y(n5578) );
  AOI222XLTS U166 ( .A0(n3853), .A1(n3676), .B0(n389), .B1(n3412), .C0(n4009), 
        .C1(n3395), .Y(n5692) );
  AOI222XLTS U167 ( .A0(n3841), .A1(n3675), .B0(n397), .B1(n3411), .C0(n3997), 
        .C1(n3396), .Y(n5700) );
  AOI222XLTS U168 ( .A0(n3826), .A1(n3674), .B0(n407), .B1(n3409), .C0(n3982), 
        .C1(n3393), .Y(n5710) );
  AOI222XLTS U169 ( .A0(n3916), .A1(n3681), .B0(n347), .B1(n3421), .C0(n4072), 
        .C1(n3400), .Y(n5650) );
  AOI222XLTS U170 ( .A0(n3913), .A1(n3681), .B0(n349), .B1(n3421), .C0(n4069), 
        .C1(n3400), .Y(n5652) );
  AOI222XLTS U171 ( .A0(n3856), .A1(n3676), .B0(n387), .B1(n3412), .C0(n4012), 
        .C1(n3395), .Y(n5690) );
  AOI222XLTS U172 ( .A0(n3850), .A1(n3676), .B0(n391), .B1(n3411), .C0(n4006), 
        .C1(n3395), .Y(n5694) );
  AOI222XLTS U173 ( .A0(n3847), .A1(n3675), .B0(n393), .B1(n3411), .C0(n4003), 
        .C1(n3394), .Y(n5696) );
  AOI222XLTS U174 ( .A0(n3844), .A1(n3675), .B0(n395), .B1(n3411), .C0(n4000), 
        .C1(n3394), .Y(n5698) );
  AOI222XLTS U175 ( .A0(n3838), .A1(n3675), .B0(n399), .B1(n3410), .C0(n3994), 
        .C1(n3394), .Y(n5702) );
  AOI222XLTS U176 ( .A0(n3832), .A1(n3674), .B0(n403), .B1(n3410), .C0(n3988), 
        .C1(n3393), .Y(n5706) );
  AOI222XLTS U177 ( .A0(n3829), .A1(n3674), .B0(n405), .B1(n3410), .C0(n3985), 
        .C1(n3393), .Y(n5708) );
  AOI222XLTS U178 ( .A0(n3823), .A1(n3679), .B0(n409), .B1(n3409), .C0(n3979), 
        .C1(n3393), .Y(n5712) );
  AOI222XLTS U179 ( .A0(n4072), .A1(n3494), .B0(n348), .B1(n3473), .C0(n4228), 
        .C1(n3468), .Y(n5586) );
  AOI222XLTS U180 ( .A0(n4069), .A1(n3494), .B0(n350), .B1(n3473), .C0(n4225), 
        .C1(n3469), .Y(n5588) );
  AOI222XLTS U181 ( .A0(n4066), .A1(n3493), .B0(n352), .B1(n3474), .C0(n4222), 
        .C1(n3470), .Y(n5590) );
  AOI222XLTS U182 ( .A0(n4063), .A1(n3493), .B0(n354), .B1(n3474), .C0(n4219), 
        .C1(n3466), .Y(n5592) );
  AOI222XLTS U183 ( .A0(n4060), .A1(n3493), .B0(n356), .B1(n3474), .C0(n4216), 
        .C1(n3466), .Y(n5594) );
  AOI222XLTS U184 ( .A0(n4057), .A1(n3493), .B0(n358), .B1(n3474), .C0(n4213), 
        .C1(n3467), .Y(n5596) );
  AOI222XLTS U185 ( .A0(n4054), .A1(n3500), .B0(n359), .B1(n3475), .C0(n4210), 
        .C1(n3466), .Y(n5598) );
  AOI222XLTS U186 ( .A0(n4051), .A1(n3498), .B0(n362), .B1(n3475), .C0(n4207), 
        .C1(n3467), .Y(n5600) );
  AOI222XLTS U187 ( .A0(n4048), .A1(n3502), .B0(n364), .B1(n3475), .C0(n4204), 
        .C1(n3471), .Y(n5602) );
  AOI222XLTS U188 ( .A0(n4045), .A1(n3503), .B0(n366), .B1(n3475), .C0(n4201), 
        .C1(n3471), .Y(n5604) );
  AOI222XLTS U189 ( .A0(n4042), .A1(n3501), .B0(n368), .B1(n3476), .C0(n4198), 
        .C1(n3472), .Y(n5606) );
  AOI222XLTS U190 ( .A0(n4039), .A1(n3500), .B0(n370), .B1(n3476), .C0(n4195), 
        .C1(n3468), .Y(n5608) );
  AOI222XLTS U191 ( .A0(n4036), .A1(n3500), .B0(n372), .B1(n3476), .C0(n4192), 
        .C1(n3464), .Y(n5610) );
  AOI222XLTS U192 ( .A0(n4033), .A1(n3492), .B0(n373), .B1(n3476), .C0(n4189), 
        .C1(n3464), .Y(n5612) );
  AOI222XLTS U193 ( .A0(n4030), .A1(n3492), .B0(n376), .B1(n3477), .C0(n4186), 
        .C1(n3464), .Y(n5614) );
  AOI222XLTS U194 ( .A0(n4027), .A1(n3492), .B0(n378), .B1(n3477), .C0(n4183), 
        .C1(n3464), .Y(n5616) );
  AOI222XLTS U195 ( .A0(n4015), .A1(n3491), .B0(n386), .B1(n3478), .C0(n4171), 
        .C1(n3462), .Y(n5624) );
  AOI222XLTS U196 ( .A0(n4012), .A1(n3491), .B0(n388), .B1(n3478), .C0(n4168), 
        .C1(n3462), .Y(n5626) );
  AOI222XLTS U197 ( .A0(n4009), .A1(n3490), .B0(n390), .B1(n3478), .C0(n4165), 
        .C1(n3462), .Y(n5628) );
  AOI222XLTS U198 ( .A0(n4006), .A1(n3490), .B0(n392), .B1(n3479), .C0(n4162), 
        .C1(n3462), .Y(n5630) );
  AOI222XLTS U199 ( .A0(n4003), .A1(n3490), .B0(n394), .B1(n3479), .C0(n4159), 
        .C1(n3461), .Y(n5632) );
  AOI222XLTS U200 ( .A0(n4000), .A1(n3490), .B0(n396), .B1(n3479), .C0(n4156), 
        .C1(n3461), .Y(n5634) );
  AOI222XLTS U201 ( .A0(n3997), .A1(n3489), .B0(n398), .B1(n3479), .C0(n4153), 
        .C1(n3461), .Y(n5636) );
  AOI222XLTS U202 ( .A0(n3994), .A1(n3489), .B0(n400), .B1(n3480), .C0(n4150), 
        .C1(n3461), .Y(n5638) );
  AOI222XLTS U203 ( .A0(n3991), .A1(n3489), .B0(n401), .B1(n3480), .C0(n4147), 
        .C1(n3460), .Y(n5640) );
  AOI222XLTS U204 ( .A0(n3988), .A1(n3489), .B0(n404), .B1(n3480), .C0(n4144), 
        .C1(n3460), .Y(n5642) );
  AOI222XLTS U205 ( .A0(n3985), .A1(n3488), .B0(n406), .B1(n3480), .C0(n4141), 
        .C1(n3460), .Y(n5644) );
  AOI222XLTS U206 ( .A0(n3982), .A1(n3488), .B0(n408), .B1(n3481), .C0(n4138), 
        .C1(n3460), .Y(n5646) );
  AOI222XLTS U207 ( .A0(n3835), .A1(n3674), .B0(n402), .B1(n3410), .C0(n3991), 
        .C1(n3394), .Y(n5704) );
  AOI222XLTS U208 ( .A0(n3976), .A1(n3319), .B0(n4289), .B1(n3325), .C0(n4132), 
        .C1(n3367), .Y(n5441) );
  INVX2TS U209 ( .A(n284), .Y(n285) );
  INVX2TS U210 ( .A(n233), .Y(n284) );
  OR3X1TS U211 ( .A(n6335), .B(n157), .C(n5531), .Y(n2) );
  OR2X2TS U212 ( .A(n4836), .B(n5314), .Y(n6) );
  OR3X1TS U213 ( .A(n276), .B(n194), .C(n335), .Y(n9) );
  NAND2BX1TS U214 ( .AN(n5369), .B(n5390), .Y(n5539) );
  AND2X2TS U215 ( .A(n432), .B(n168), .Y(n12) );
  OR2X2TS U216 ( .A(n189), .B(n5315), .Y(n13) );
  XOR2X1TS U217 ( .A(n174), .B(n197), .Y(n14) );
  OA22X2TS U218 ( .A0(n6250), .A1(n190), .B0(n4872), .B1(n331), .Y(n15) );
  AOI221X1TS U219 ( .A0(n202), .A1(n174), .B0(n6322), .B1(n5326), .C0(n200), 
        .Y(n5532) );
  INVX2TS U220 ( .A(n262), .Y(n263) );
  CLKBUFX2TS U221 ( .A(n5525), .Y(n110) );
  INVX2TS U222 ( .A(n5545), .Y(n111) );
  INVXLTS U223 ( .A(n111), .Y(n112) );
  INVXLTS U224 ( .A(n122), .Y(n114) );
  INVXLTS U225 ( .A(n126), .Y(n115) );
  INVXLTS U226 ( .A(n130), .Y(n116) );
  INVXLTS U227 ( .A(n134), .Y(n117) );
  INVXLTS U228 ( .A(n143), .Y(n118) );
  CLKBUFX2TS U229 ( .A(selectBit_NORTH), .Y(n119) );
  INVXLTS U230 ( .A(n6237), .Y(n120) );
  CLKBUFX2TS U231 ( .A(n5327), .Y(n121) );
  INVXLTS U232 ( .A(readRequesterAddress[0]), .Y(n122) );
  INVXLTS U233 ( .A(n122), .Y(n123) );
  INVXLTS U234 ( .A(n122), .Y(n124) );
  INVXLTS U235 ( .A(n122), .Y(n125) );
  INVXLTS U236 ( .A(readRequesterAddress[1]), .Y(n126) );
  INVXLTS U237 ( .A(n126), .Y(n127) );
  INVXLTS U238 ( .A(n126), .Y(n128) );
  INVXLTS U239 ( .A(n126), .Y(n129) );
  INVXLTS U240 ( .A(readRequesterAddress[2]), .Y(n130) );
  INVXLTS U241 ( .A(n130), .Y(n131) );
  INVXLTS U242 ( .A(n130), .Y(n132) );
  INVXLTS U243 ( .A(n130), .Y(n133) );
  INVXLTS U244 ( .A(readRequesterAddress[3]), .Y(n134) );
  INVXLTS U245 ( .A(n134), .Y(n135) );
  INVXLTS U246 ( .A(n134), .Y(n136) );
  INVXLTS U247 ( .A(n134), .Y(n137) );
  INVXLTS U248 ( .A(readRequesterAddress[4]), .Y(n138) );
  INVXLTS U249 ( .A(n138), .Y(n139) );
  INVXLTS U250 ( .A(n138), .Y(n140) );
  INVXLTS U251 ( .A(n138), .Y(n141) );
  INVXLTS U252 ( .A(n138), .Y(n142) );
  INVXLTS U253 ( .A(readRequesterAddress[5]), .Y(n143) );
  INVXLTS U254 ( .A(n143), .Y(n144) );
  INVXLTS U255 ( .A(n143), .Y(n145) );
  INVXLTS U256 ( .A(n143), .Y(n146) );
  INVXLTS U257 ( .A(n3), .Y(n147) );
  INVXLTS U258 ( .A(n5), .Y(n148) );
  INVXLTS U259 ( .A(n14), .Y(n149) );
  INVXLTS U260 ( .A(n14), .Y(n150) );
  INVXLTS U261 ( .A(n5393), .Y(n151) );
  INVXLTS U262 ( .A(n151), .Y(n152) );
  INVXLTS U263 ( .A(n5449), .Y(n153) );
  INVXLTS U264 ( .A(n153), .Y(n154) );
  INVXLTS U265 ( .A(n197), .Y(n155) );
  INVX2TS U266 ( .A(selectBit_NORTH), .Y(n6250) );
  CLKINVX1TS U267 ( .A(n156), .Y(n157) );
  CLKINVX2TS U268 ( .A(n5569), .Y(n158) );
  INVXLTS U269 ( .A(n15), .Y(n159) );
  INVXLTS U270 ( .A(n15), .Y(n160) );
  CLKINVX2TS U271 ( .A(n5530), .Y(n161) );
  INVXLTS U272 ( .A(n161), .Y(n162) );
  CLKBUFX2TS U273 ( .A(n5552), .Y(n163) );
  CLKBUFX2TS U274 ( .A(n5512), .Y(n164) );
  AOI21X1TS U275 ( .A0(n177), .A1(n5392), .B0(n6338), .Y(n5515) );
  AOI21X1TS U276 ( .A0(n202), .A1(n5464), .B0(n427), .Y(n5559) );
  CLKBUFX2TS U277 ( .A(n5566), .Y(n166) );
  AOI21X1TS U278 ( .A0(n5489), .A1(n5498), .B0(n428), .Y(n5566) );
  INVXLTS U279 ( .A(n6), .Y(n167) );
  INVXLTS U280 ( .A(n6), .Y(n168) );
  INVXLTS U281 ( .A(n13), .Y(n169) );
  INVXLTS U282 ( .A(n13), .Y(n170) );
  INVXLTS U283 ( .A(n5549), .Y(n171) );
  CLKBUFX2TS U284 ( .A(n5531), .Y(n173) );
  INVXLTS U285 ( .A(n6322), .Y(n174) );
  INVXLTS U286 ( .A(n5464), .Y(n175) );
  INVXLTS U287 ( .A(n175), .Y(n176) );
  AOI21X1TS U288 ( .A0(n176), .A1(n5393), .B0(n6344), .Y(n5530) );
  INVXLTS U289 ( .A(n5539), .Y(n177) );
  INVXLTS U290 ( .A(n177), .Y(n178) );
  INVXLTS U291 ( .A(n9), .Y(n179) );
  INVXLTS U292 ( .A(n9), .Y(n180) );
  INVXLTS U293 ( .A(n1), .Y(n181) );
  INVXLTS U294 ( .A(n198), .Y(n182) );
  INVXLTS U295 ( .A(n182), .Y(n183) );
  INVXLTS U296 ( .A(n277), .Y(n184) );
  INVXLTS U297 ( .A(n205), .Y(n185) );
  INVXLTS U298 ( .A(n271), .Y(n186) );
  INVXLTS U299 ( .A(n167), .Y(n187) );
  INVXLTS U300 ( .A(n167), .Y(n188) );
  INVXLTS U301 ( .A(n341), .Y(n190) );
  NAND2X1TS U302 ( .A(n6326), .B(n196), .Y(n5518) );
  INVXLTS U303 ( .A(n4843), .Y(n191) );
  INVXLTS U304 ( .A(n6238), .Y(n192) );
  INVXLTS U305 ( .A(n192), .Y(n193) );
  INVXLTS U306 ( .A(n333), .Y(n194) );
  INVXLTS U307 ( .A(n335), .Y(n195) );
  INVXLTS U308 ( .A(n343), .Y(n196) );
  INVXLTS U309 ( .A(n196), .Y(n197) );
  INVXLTS U310 ( .A(n329), .Y(n198) );
  INVXLTS U311 ( .A(n198), .Y(n199) );
  INVXLTS U312 ( .A(n6318), .Y(n200) );
  INVXLTS U313 ( .A(n5498), .Y(n201) );
  INVXLTS U314 ( .A(n201), .Y(n202) );
  INVXLTS U315 ( .A(n12), .Y(n203) );
  INVXLTS U316 ( .A(n12), .Y(n204) );
  INVXLTS U317 ( .A(n281), .Y(n207) );
  INVXLTS U318 ( .A(n205), .Y(n208) );
  INVXLTS U319 ( .A(n284), .Y(n209) );
  INVXLTS U320 ( .A(n285), .Y(n210) );
  INVXLTS U321 ( .A(n210), .Y(n211) );
  INVXLTS U322 ( .A(n285), .Y(n212) );
  INVXLTS U323 ( .A(n212), .Y(n213) );
  INVXLTS U324 ( .A(n212), .Y(n214) );
  INVXLTS U325 ( .A(n212), .Y(n286) );
  CLKBUFX2TS U326 ( .A(n331), .Y(n215) );
  INVX2TS U327 ( .A(n5518), .Y(n216) );
  INVXLTS U328 ( .A(n216), .Y(n217) );
  INVXLTS U329 ( .A(n212), .Y(n218) );
  INVXLTS U330 ( .A(n2), .Y(n219) );
  INVXLTS U331 ( .A(n210), .Y(n220) );
  INVXLTS U332 ( .A(n284), .Y(n221) );
  INVXLTS U333 ( .A(n5287), .Y(n222) );
  INVXLTS U334 ( .A(n222), .Y(n223) );
  INVXLTS U335 ( .A(n7), .Y(n224) );
  INVXLTS U336 ( .A(n3745), .Y(n225) );
  INVXLTS U337 ( .A(n225), .Y(n226) );
  INVXLTS U338 ( .A(n225), .Y(n227) );
  INVXLTS U339 ( .A(n5570), .Y(n228) );
  INVXLTS U340 ( .A(n228), .Y(n229) );
  INVXLTS U341 ( .A(n228), .Y(n230) );
  INVXLTS U342 ( .A(n3629), .Y(n231) );
  INVXLTS U343 ( .A(n2), .Y(n232) );
  INVXLTS U344 ( .A(n2), .Y(n233) );
  INVXLTS U345 ( .A(n199), .Y(n234) );
  INVXLTS U346 ( .A(n6239), .Y(n235) );
  INVXLTS U347 ( .A(n235), .Y(n236) );
  INVXLTS U348 ( .A(n235), .Y(n237) );
  INVXLTS U349 ( .A(n6241), .Y(n238) );
  INVXLTS U350 ( .A(n238), .Y(n239) );
  INVXLTS U351 ( .A(n238), .Y(n240) );
  INVXLTS U352 ( .A(n6240), .Y(n241) );
  INVXLTS U353 ( .A(n241), .Y(n242) );
  INVXLTS U354 ( .A(n241), .Y(n243) );
  INVXLTS U355 ( .A(n6246), .Y(n244) );
  INVXLTS U356 ( .A(n244), .Y(n245) );
  INVXLTS U357 ( .A(n244), .Y(n246) );
  INVXLTS U358 ( .A(n6244), .Y(n247) );
  INVXLTS U359 ( .A(n247), .Y(n248) );
  INVXLTS U360 ( .A(n247), .Y(n249) );
  INVXLTS U361 ( .A(n6243), .Y(n250) );
  INVXLTS U362 ( .A(n250), .Y(n251) );
  INVXLTS U363 ( .A(n250), .Y(n252) );
  INVXLTS U364 ( .A(n6247), .Y(n253) );
  INVXLTS U365 ( .A(n253), .Y(n254) );
  INVXLTS U366 ( .A(n253), .Y(n255) );
  INVXLTS U367 ( .A(n6245), .Y(n256) );
  INVXLTS U368 ( .A(n256), .Y(n257) );
  INVXLTS U369 ( .A(n256), .Y(n258) );
  INVXLTS U370 ( .A(n6242), .Y(n259) );
  INVXLTS U371 ( .A(n259), .Y(n260) );
  INVXLTS U372 ( .A(n259), .Y(n261) );
  INVXLTS U373 ( .A(n5572), .Y(n262) );
  INVXLTS U374 ( .A(n262), .Y(n264) );
  INVXLTS U375 ( .A(n5579), .Y(n265) );
  INVXLTS U376 ( .A(n265), .Y(n266) );
  INVXLTS U377 ( .A(n265), .Y(n267) );
  INVX2TS U378 ( .A(n5575), .Y(n268) );
  INVX2TS U379 ( .A(n268), .Y(n269) );
  INVXLTS U380 ( .A(n268), .Y(n270) );
  INVXLTS U381 ( .A(n183), .Y(n271) );
  INVXLTS U382 ( .A(n271), .Y(n272) );
  INVXLTS U383 ( .A(n271), .Y(n273) );
  INVXLTS U384 ( .A(n271), .Y(n274) );
  INVXLTS U385 ( .A(n8), .Y(n275) );
  INVXLTS U386 ( .A(n8), .Y(n276) );
  INVXLTS U387 ( .A(n3776), .Y(n277) );
  INVXLTS U388 ( .A(n277), .Y(n278) );
  INVXLTS U389 ( .A(n277), .Y(n279) );
  INVXLTS U390 ( .A(n277), .Y(n280) );
  INVXLTS U391 ( .A(n3775), .Y(n281) );
  INVXLTS U392 ( .A(n281), .Y(n282) );
  INVXLTS U393 ( .A(n281), .Y(n283) );
  INVXLTS U394 ( .A(n284), .Y(n287) );
  INVXLTS U395 ( .A(n210), .Y(n288) );
  INVXLTS U396 ( .A(n225), .Y(n289) );
  INVXLTS U397 ( .A(n225), .Y(n290) );
  CLKBUFX2TS U430 ( .A(n5585), .Y(n323) );
  CLKBUFX2TS U431 ( .A(n5585), .Y(n324) );
  CLKBUFX2TS U432 ( .A(n5581), .Y(n325) );
  CLKBUFX2TS U433 ( .A(n5581), .Y(n326) );
  CLKBUFX2TS U434 ( .A(n5583), .Y(n327) );
  CLKBUFX2TS U435 ( .A(n5583), .Y(n328) );
  OAI22X1TS U436 ( .A0(n5527), .A1(n188), .B0(n204), .B1(n151), .Y(n329) );
  OAI22X1TS U437 ( .A0(n5527), .A1(n187), .B0(n204), .B1(n151), .Y(n5574) );
  INVXLTS U438 ( .A(n5417), .Y(n6337) );
  OAI22X1TS U439 ( .A0(n164), .A1(n6), .B0(n203), .B1(n6318), .Y(n330) );
  XNOR2X4TS U440 ( .A(n155), .B(n5320), .Y(n5318) );
  NAND2X1TS U441 ( .A(n6325), .B(selectBit_EAST), .Y(n5487) );
  INVX1TS U442 ( .A(selectBit_EAST), .Y(n6237) );
  AND3XLTS U443 ( .A(n5515), .B(n170), .C(n5322), .Y(n6108) );
  NOR3BX1TS U444 ( .AN(n162), .B(n5524), .C(n5525), .Y(n6139) );
  XNOR2X1TS U445 ( .A(selectBit_NORTH), .B(selectBit_EAST), .Y(n4839) );
  BUFX3TS U446 ( .A(n6237), .Y(n331) );
  NAND2XLTS U447 ( .A(n5553), .B(n5559), .Y(n6205) );
  CLKBUFX2TS U448 ( .A(n6233), .Y(n332) );
  CLKBUFX2TS U449 ( .A(readReady), .Y(n336) );
  INVXLTS U450 ( .A(n5391), .Y(n337) );
  NAND3X1TS U451 ( .A(n6332), .B(n5463), .C(n6331), .Y(n5513) );
  OR2X2TS U452 ( .A(n5305), .B(n6252), .Y(n5283) );
  INVX2TS U453 ( .A(n5283), .Y(n338) );
  INVX2TS U454 ( .A(n5283), .Y(n339) );
  CLKBUFX2TS U455 ( .A(selectBit_WEST), .Y(n340) );
  CLKBUFX2TS U456 ( .A(selectBit_SOUTH), .Y(n341) );
  NOR2X1TS U457 ( .A(selectBit_SOUTH), .B(selectBit_NORTH), .Y(n4872) );
  CLKBUFX2TS U458 ( .A(n5489), .Y(n342) );
  OAI31XLTS U459 ( .A0(n5489), .A1(n6326), .A2(n174), .B0(n167), .Y(n5488) );
  OAI21X1TS U460 ( .A0(n5320), .A1(n159), .B0(n343), .Y(n5319) );
  INVX2TS U461 ( .A(n3684), .Y(n344) );
  INVX1TS U462 ( .A(n6205), .Y(n6340) );
  INVX2TS U463 ( .A(n5295), .Y(n345) );
  OAI32XLTS U464 ( .A0(n4869), .A1(n332), .A2(n4868), .B0(n345), .B1(n6347), 
        .Y(N4718) );
  INVX2TS U465 ( .A(n3644), .Y(n346) );
  CLKBUFX2TS U466 ( .A(cacheDataOut[31]), .Y(n347) );
  CLKBUFX2TS U467 ( .A(cacheDataOut[31]), .Y(n348) );
  CLKBUFX2TS U468 ( .A(cacheDataOut[30]), .Y(n349) );
  CLKBUFX2TS U469 ( .A(cacheDataOut[30]), .Y(n350) );
  CLKBUFX2TS U470 ( .A(cacheDataOut[29]), .Y(n351) );
  CLKBUFX2TS U471 ( .A(cacheDataOut[29]), .Y(n352) );
  CLKBUFX2TS U472 ( .A(cacheDataOut[28]), .Y(n353) );
  CLKBUFX2TS U473 ( .A(cacheDataOut[28]), .Y(n354) );
  CLKBUFX2TS U474 ( .A(cacheDataOut[27]), .Y(n355) );
  CLKBUFX2TS U475 ( .A(cacheDataOut[27]), .Y(n356) );
  CLKBUFX2TS U476 ( .A(cacheDataOut[26]), .Y(n357) );
  CLKBUFX2TS U477 ( .A(cacheDataOut[26]), .Y(n358) );
  CLKBUFX2TS U478 ( .A(cacheDataOut[25]), .Y(n359) );
  CLKBUFX2TS U479 ( .A(cacheDataOut[25]), .Y(n360) );
  CLKBUFX2TS U480 ( .A(cacheDataOut[24]), .Y(n361) );
  CLKBUFX2TS U481 ( .A(cacheDataOut[24]), .Y(n362) );
  CLKBUFX2TS U482 ( .A(cacheDataOut[23]), .Y(n363) );
  CLKBUFX2TS U483 ( .A(cacheDataOut[23]), .Y(n364) );
  CLKBUFX2TS U484 ( .A(cacheDataOut[22]), .Y(n365) );
  CLKBUFX2TS U485 ( .A(cacheDataOut[22]), .Y(n366) );
  CLKBUFX2TS U486 ( .A(cacheDataOut[21]), .Y(n367) );
  CLKBUFX2TS U487 ( .A(cacheDataOut[21]), .Y(n368) );
  CLKBUFX2TS U488 ( .A(cacheDataOut[20]), .Y(n369) );
  CLKBUFX2TS U489 ( .A(cacheDataOut[20]), .Y(n370) );
  CLKBUFX2TS U490 ( .A(cacheDataOut[19]), .Y(n371) );
  CLKBUFX2TS U491 ( .A(cacheDataOut[19]), .Y(n372) );
  CLKBUFX2TS U492 ( .A(cacheDataOut[18]), .Y(n373) );
  CLKBUFX2TS U493 ( .A(cacheDataOut[18]), .Y(n374) );
  CLKBUFX2TS U494 ( .A(cacheDataOut[17]), .Y(n375) );
  CLKBUFX2TS U495 ( .A(cacheDataOut[17]), .Y(n376) );
  CLKBUFX2TS U496 ( .A(cacheDataOut[16]), .Y(n377) );
  CLKBUFX2TS U497 ( .A(cacheDataOut[16]), .Y(n378) );
  CLKBUFX2TS U498 ( .A(cacheDataOut[15]), .Y(n379) );
  CLKBUFX2TS U499 ( .A(cacheDataOut[15]), .Y(n380) );
  CLKBUFX2TS U500 ( .A(cacheDataOut[14]), .Y(n381) );
  CLKBUFX2TS U501 ( .A(cacheDataOut[14]), .Y(n382) );
  CLKBUFX2TS U502 ( .A(cacheDataOut[13]), .Y(n383) );
  CLKBUFX2TS U503 ( .A(cacheDataOut[13]), .Y(n384) );
  CLKBUFX2TS U504 ( .A(cacheDataOut[12]), .Y(n385) );
  CLKBUFX2TS U505 ( .A(cacheDataOut[12]), .Y(n386) );
  CLKBUFX2TS U506 ( .A(cacheDataOut[11]), .Y(n387) );
  CLKBUFX2TS U507 ( .A(cacheDataOut[11]), .Y(n388) );
  CLKBUFX2TS U508 ( .A(cacheDataOut[10]), .Y(n389) );
  CLKBUFX2TS U509 ( .A(cacheDataOut[10]), .Y(n390) );
  CLKBUFX2TS U510 ( .A(cacheDataOut[9]), .Y(n391) );
  CLKBUFX2TS U511 ( .A(cacheDataOut[9]), .Y(n392) );
  CLKBUFX2TS U512 ( .A(cacheDataOut[8]), .Y(n393) );
  CLKBUFX2TS U513 ( .A(cacheDataOut[8]), .Y(n394) );
  CLKBUFX2TS U514 ( .A(cacheDataOut[7]), .Y(n395) );
  CLKBUFX2TS U515 ( .A(cacheDataOut[7]), .Y(n396) );
  CLKBUFX2TS U516 ( .A(cacheDataOut[6]), .Y(n397) );
  CLKBUFX2TS U517 ( .A(cacheDataOut[6]), .Y(n398) );
  CLKBUFX2TS U518 ( .A(cacheDataOut[5]), .Y(n399) );
  CLKBUFX2TS U519 ( .A(cacheDataOut[5]), .Y(n400) );
  CLKBUFX2TS U520 ( .A(cacheDataOut[4]), .Y(n401) );
  CLKBUFX2TS U521 ( .A(cacheDataOut[4]), .Y(n402) );
  CLKBUFX2TS U522 ( .A(cacheDataOut[3]), .Y(n403) );
  CLKBUFX2TS U523 ( .A(cacheDataOut[3]), .Y(n404) );
  CLKBUFX2TS U524 ( .A(cacheDataOut[2]), .Y(n405) );
  CLKBUFX2TS U525 ( .A(cacheDataOut[2]), .Y(n406) );
  CLKBUFX2TS U526 ( .A(cacheDataOut[1]), .Y(n407) );
  CLKBUFX2TS U527 ( .A(cacheDataOut[1]), .Y(n408) );
  CLKBUFX2TS U528 ( .A(cacheDataOut[0]), .Y(n409) );
  CLKBUFX2TS U529 ( .A(cacheDataOut[0]), .Y(n410) );
  CLKBUFX2TS U530 ( .A(n6222), .Y(n411) );
  CLKBUFX2TS U531 ( .A(n6222), .Y(n412) );
  CLKBUFX2TS U532 ( .A(n5576), .Y(n413) );
  CLKBUFX2TS U533 ( .A(n5576), .Y(n414) );
  NOR3XLTS U534 ( .A(n6329), .B(n6334), .C(n173), .Y(n5576) );
  OR3XLTS U535 ( .A(n5539), .B(n6338), .C(n6345), .Y(n5567) );
  INVXLTS U536 ( .A(n5567), .Y(n415) );
  CLKINVX1TS U537 ( .A(n5567), .Y(n416) );
  INVXLTS U538 ( .A(n5567), .Y(n417) );
  INVX1TS U539 ( .A(n5322), .Y(n6345) );
  INVX2TS U540 ( .A(n168), .Y(n418) );
  NAND3XLTS U541 ( .A(n163), .B(n217), .C(n5547), .Y(n5581) );
  INVX2TS U542 ( .A(n4856), .Y(n6321) );
  AOI211X1TS U543 ( .A0(n6227), .A1(n4857), .B0(n6320), .C0(n6249), .Y(n4853)
         );
  AND3X2TS U544 ( .A(n5545), .B(n177), .C(n5417), .Y(n6171) );
  OAI21X1TS U545 ( .A0(n5394), .A1(n418), .B0(n420), .Y(n419) );
  AND2XLTS U546 ( .A(n5563), .B(n5566), .Y(n6219) );
  NAND2XLTS U547 ( .A(n5315), .B(n341), .Y(n5316) );
  CLKBUFX2TS U548 ( .A(n685), .Y(n679) );
  CLKBUFX2TS U549 ( .A(n805), .Y(n797) );
  NOR2XLTS U550 ( .A(n6327), .B(n149), .Y(n5462) );
  NAND2XLTS U551 ( .A(n5512), .B(n5322), .Y(n5570) );
  NAND3XLTS U552 ( .A(n166), .B(n6324), .C(n5560), .Y(n5585) );
  NAND2XLTS U553 ( .A(n5554), .B(n5559), .Y(n5583) );
  AND2XLTS U554 ( .A(n5562), .B(n5566), .Y(n6216) );
  NAND2X1TS U555 ( .A(n5390), .B(n5369), .Y(n5524) );
  NOR2BXLTS U556 ( .AN(n150), .B(n5390), .Y(n5549) );
  NOR2XLTS U557 ( .A(n4857), .B(n6321), .Y(n4862) );
  NAND2XLTS U558 ( .A(n169), .B(n149), .Y(n5416) );
  INVX2TS U559 ( .A(n863), .Y(n420) );
  XNOR2XLTS U560 ( .A(n4861), .B(n5323), .Y(n4858) );
  NOR3XLTS U561 ( .A(n4865), .B(n6321), .C(n6251), .Y(n4866) );
  AOI22XLTS U562 ( .A0(n4863), .A1(n197), .B0(n4862), .B1(n4861), .Y(n4864) );
  NAND2XLTS U563 ( .A(n4854), .B(n4856), .Y(n4855) );
  XOR2X2TS U564 ( .A(n5318), .B(n160), .Y(n5391) );
  OAI211XLTS U565 ( .A0(n5567), .A1(n3983), .B0(n6095), .C0(n6094), .Y(n2833)
         );
  OAI211XLTS U566 ( .A0(n3786), .A1(n3980), .B0(n6097), .C0(n6096), .Y(n2834)
         );
  OAI211XLTS U567 ( .A0(n3777), .A1(n4109), .B0(n5335), .C0(n5334), .Y(n2459)
         );
  OAI211XLTS U568 ( .A0(n3777), .A1(n4103), .B0(n5339), .C0(n5338), .Y(n2461)
         );
  OAI211XLTS U569 ( .A0(n3777), .A1(n4100), .B0(n5341), .C0(n5340), .Y(n2462)
         );
  OAI211XLTS U570 ( .A0(n3778), .A1(n4097), .B0(n5343), .C0(n5342), .Y(n2463)
         );
  OAI22XLTS U571 ( .A0(n6230), .A1(n6233), .B0(n5326), .B1(n6232), .Y(n2886)
         );
  INVXLTS U572 ( .A(n853), .Y(n848) );
  INVXLTS U573 ( .A(n852), .Y(n849) );
  INVXLTS U574 ( .A(n851), .Y(n850) );
  INVXLTS U575 ( .A(n3518), .Y(n3516) );
  INVXLTS U576 ( .A(n428), .Y(n3515) );
  CLKBUFX2TS U577 ( .A(n3307), .Y(n3304) );
  CLKBUFX2TS U578 ( .A(n582), .Y(n578) );
  CLKBUFX2TS U579 ( .A(n582), .Y(n577) );
  CLKBUFX2TS U580 ( .A(n788), .Y(n785) );
  CLKBUFX2TS U581 ( .A(n3390), .Y(n3387) );
  CLKBUFX2TS U582 ( .A(n3521), .Y(n3518) );
  CLKBUFX2TS U583 ( .A(n3307), .Y(n3305) );
  CLKBUFX2TS U584 ( .A(n3390), .Y(n3388) );
  CLKBUFX2TS U585 ( .A(n3521), .Y(n3519) );
  CLKBUFX2TS U586 ( .A(n788), .Y(n786) );
  NOR2XLTS U587 ( .A(n5513), .B(n6345), .Y(n6110) );
  CLKAND2X2TS U588 ( .A(n162), .B(n5462), .Y(n6141) );
  AND2XLTS U589 ( .A(n5525), .B(n162), .Y(n423) );
  NAND2X2TS U590 ( .A(n3223), .B(n5395), .Y(n5531) );
  OR2XLTS U591 ( .A(n5531), .B(n6323), .Y(n424) );
  CLKBUFX2TS U592 ( .A(n564), .Y(n558) );
  CLKBUFX2TS U593 ( .A(n564), .Y(n559) );
  NOR3BXLTS U594 ( .AN(n5486), .B(n334), .C(n337), .Y(n5562) );
  NOR3BX1TS U595 ( .AN(n112), .B(n5540), .C(n6327), .Y(n6168) );
  NAND3XLTS U596 ( .A(n5486), .B(n5391), .C(n6331), .Y(n5535) );
  NOR2X1TS U597 ( .A(n343), .B(n7), .Y(n5356) );
  AOI221X2TS U598 ( .A0(n6330), .A1(n5392), .B0(n5326), .B1(n5462), .C0(n5525), 
        .Y(n5527) );
  NOR2X4TS U599 ( .A(n6248), .B(n121), .Y(n5320) );
  XOR2XLTS U600 ( .A(n4865), .B(n160), .Y(n4857) );
  NOR2X1TS U601 ( .A(n6235), .B(n432), .Y(n5489) );
  NOR2X1TS U602 ( .A(n6250), .B(n5327), .Y(n5347) );
  AOI21X1TS U603 ( .A0(n190), .A1(n5315), .B0(n169), .Y(n5390) );
  AOI32XLTS U604 ( .A0(n163), .A1(n5551), .A2(n5550), .B0(n3389), .B1(n25), 
        .Y(n2568) );
  AOI32XLTS U605 ( .A0(n5549), .A1(n5548), .A2(n3812), .B0(n5547), .B1(n5546), 
        .Y(n5550) );
  AOI32XLTS U606 ( .A0(n113), .A1(n5522), .A2(n5521), .B0(n787), .B1(n17), .Y(
        n2564) );
  AOI32XLTS U607 ( .A0(n172), .A1(n5520), .A2(n3813), .B0(n5519), .B1(n5546), 
        .Y(n5521) );
  INVXLTS U608 ( .A(n5347), .Y(n6322) );
  NOR2X1TS U609 ( .A(n6235), .B(n16), .Y(n5464) );
  OAI32XLTS U610 ( .A0(n3814), .A1(n110), .A2(n5524), .B0(n6328), .B1(n193), 
        .Y(n5526) );
  AND2XLTS U611 ( .A(n342), .B(n168), .Y(n5499) );
  NAND2XLTS U612 ( .A(n167), .B(n4422), .Y(n6233) );
  NOR2X1TS U613 ( .A(n224), .B(n5323), .Y(n5498) );
  NOR2X1TS U614 ( .A(n7), .B(n155), .Y(n5393) );
  NOR2X1TS U615 ( .A(n343), .B(n224), .Y(n5449) );
  NOR2X1TS U616 ( .A(n275), .B(n121), .Y(n4845) );
  NOR3X1TS U617 ( .A(n333), .B(n4), .C(n148), .Y(n5286) );
  OAI211XLTS U618 ( .A0(n849), .A1(n3827), .B0(n5967), .C0(n5966), .Y(n2769)
         );
  OAI211XLTS U619 ( .A0(n849), .A1(n3824), .B0(n5969), .C0(n5968), .Y(n2770)
         );
  OAI211XLTS U620 ( .A0(n840), .A1(n3944), .B0(n5385), .C0(n5384), .Y(n2490)
         );
  OAI211XLTS U621 ( .A0(n841), .A1(n3914), .B0(n5909), .C0(n5908), .Y(n2740)
         );
  OAI211XLTS U622 ( .A0(n842), .A1(n3911), .B0(n5911), .C0(n5910), .Y(n2741)
         );
  OAI211XLTS U623 ( .A0(n842), .A1(n3908), .B0(n5913), .C0(n5912), .Y(n2742)
         );
  OAI211XLTS U624 ( .A0(n842), .A1(n3902), .B0(n5917), .C0(n5916), .Y(n2744)
         );
  OAI211XLTS U625 ( .A0(n843), .A1(n3899), .B0(n5919), .C0(n5918), .Y(n2745)
         );
  OAI211XLTS U626 ( .A0(n843), .A1(n3893), .B0(n5923), .C0(n5922), .Y(n2747)
         );
  OAI211XLTS U627 ( .A0(n844), .A1(n3887), .B0(n5927), .C0(n5926), .Y(n2749)
         );
  OAI211XLTS U628 ( .A0(n844), .A1(n3884), .B0(n5929), .C0(n5928), .Y(n2750)
         );
  OAI211XLTS U629 ( .A0(n844), .A1(n3881), .B0(n5931), .C0(n5930), .Y(n2751)
         );
  OAI211XLTS U630 ( .A0(n844), .A1(n3878), .B0(n5933), .C0(n5932), .Y(n2752)
         );
  OAI211XLTS U631 ( .A0(n845), .A1(n3875), .B0(n5935), .C0(n5934), .Y(n2753)
         );
  OAI211XLTS U632 ( .A0(n845), .A1(n3869), .B0(n5939), .C0(n5938), .Y(n2755)
         );
  OAI211XLTS U633 ( .A0(n845), .A1(n3866), .B0(n5941), .C0(n5940), .Y(n2756)
         );
  OAI211XLTS U634 ( .A0(n846), .A1(n3863), .B0(n5943), .C0(n5942), .Y(n2757)
         );
  OAI211XLTS U635 ( .A0(n846), .A1(n3860), .B0(n5945), .C0(n5944), .Y(n2758)
         );
  OAI211XLTS U636 ( .A0(n846), .A1(n3857), .B0(n5947), .C0(n5946), .Y(n2759)
         );
  OAI211XLTS U637 ( .A0(n847), .A1(n3851), .B0(n5951), .C0(n5950), .Y(n2761)
         );
  OAI211XLTS U638 ( .A0(n847), .A1(n3848), .B0(n5953), .C0(n5952), .Y(n2762)
         );
  OAI211XLTS U639 ( .A0(n847), .A1(n3845), .B0(n5955), .C0(n5954), .Y(n2763)
         );
  OAI211XLTS U640 ( .A0(n848), .A1(n3839), .B0(n5959), .C0(n5958), .Y(n2765)
         );
  OAI211XLTS U641 ( .A0(n848), .A1(n3836), .B0(n5961), .C0(n5960), .Y(n2766)
         );
  OAI211XLTS U642 ( .A0(n848), .A1(n3833), .B0(n5963), .C0(n5962), .Y(n2767)
         );
  OAI211XLTS U643 ( .A0(n840), .A1(n3953), .B0(n5379), .C0(n5378), .Y(n2487)
         );
  OAI211XLTS U644 ( .A0(n840), .A1(n3950), .B0(n5381), .C0(n5380), .Y(n2488)
         );
  OAI211XLTS U645 ( .A0(n840), .A1(n3947), .B0(n5383), .C0(n5382), .Y(n2489)
         );
  OAI211XLTS U646 ( .A0(n841), .A1(n3941), .B0(n5387), .C0(n5386), .Y(n2491)
         );
  OAI211XLTS U647 ( .A0(n841), .A1(n3938), .B0(n5389), .C0(n5388), .Y(n2492)
         );
  OAI211XLTS U648 ( .A0(n842), .A1(n3905), .B0(n5915), .C0(n5914), .Y(n2743)
         );
  OAI211XLTS U649 ( .A0(n846), .A1(n3854), .B0(n5949), .C0(n5948), .Y(n2760)
         );
  OAI211XLTS U650 ( .A0(n841), .A1(n3917), .B0(n5907), .C0(n5906), .Y(n2739)
         );
  OAI211XLTS U651 ( .A0(n843), .A1(n3896), .B0(n5921), .C0(n5920), .Y(n2746)
         );
  OAI211XLTS U652 ( .A0(n843), .A1(n3890), .B0(n5925), .C0(n5924), .Y(n2748)
         );
  OAI211XLTS U653 ( .A0(n845), .A1(n3872), .B0(n5937), .C0(n5936), .Y(n2754)
         );
  OAI211XLTS U654 ( .A0(n847), .A1(n3842), .B0(n5957), .C0(n5956), .Y(n2764)
         );
  OAI211XLTS U655 ( .A0(n848), .A1(n3830), .B0(n5965), .C0(n5964), .Y(n2768)
         );
  OAI211XLTS U656 ( .A0(n4091), .A1(n3787), .B0(n6099), .C0(n6098), .Y(n2835)
         );
  OAI211XLTS U657 ( .A0(n4088), .A1(n3789), .B0(n6101), .C0(n6100), .Y(n2836)
         );
  OAI211XLTS U658 ( .A0(n4085), .A1(n3785), .B0(n6103), .C0(n6102), .Y(n2837)
         );
  OAI211XLTS U659 ( .A0(n4082), .A1(n3788), .B0(n6105), .C0(n6104), .Y(n2838)
         );
  OAI211XLTS U660 ( .A0(n4079), .A1(n3785), .B0(n6107), .C0(n6106), .Y(n2839)
         );
  OAI211XLTS U661 ( .A0(n4076), .A1(n3788), .B0(n6112), .C0(n6111), .Y(n2840)
         );
  OAI211XLTS U662 ( .A0(n3932), .A1(n849), .B0(n6132), .C0(n6131), .Y(n2848)
         );
  OAI211XLTS U663 ( .A0(n3935), .A1(n849), .B0(n6130), .C0(n6129), .Y(n2847)
         );
  OAI211XLTS U664 ( .A0(n3923), .A1(n850), .B0(n6138), .C0(n6137), .Y(n2851)
         );
  OAI211XLTS U665 ( .A0(n3920), .A1(n850), .B0(n6143), .C0(n6142), .Y(n2852)
         );
  OAI211XLTS U666 ( .A0(n3929), .A1(n850), .B0(n6134), .C0(n6133), .Y(n2849)
         );
  OAI211XLTS U667 ( .A0(n3926), .A1(n850), .B0(n6136), .C0(n6135), .Y(n2850)
         );
  OAI211XLTS U668 ( .A0(n3778), .A1(n4073), .B0(n6035), .C0(n6034), .Y(n2803)
         );
  OAI211XLTS U669 ( .A0(n3778), .A1(n4070), .B0(n6037), .C0(n6036), .Y(n2804)
         );
  OAI211XLTS U670 ( .A0(n3779), .A1(n4067), .B0(n6039), .C0(n6038), .Y(n2805)
         );
  OAI211XLTS U671 ( .A0(n3779), .A1(n4058), .B0(n6045), .C0(n6044), .Y(n2808)
         );
  OAI211XLTS U672 ( .A0(n3780), .A1(n4055), .B0(n6047), .C0(n6046), .Y(n2809)
         );
  OAI211XLTS U673 ( .A0(n3780), .A1(n4052), .B0(n6049), .C0(n6048), .Y(n2810)
         );
  OAI211XLTS U674 ( .A0(n3780), .A1(n4046), .B0(n6053), .C0(n6052), .Y(n2812)
         );
  OAI211XLTS U675 ( .A0(n3781), .A1(n4043), .B0(n6055), .C0(n6054), .Y(n2813)
         );
  OAI211XLTS U676 ( .A0(n3781), .A1(n4037), .B0(n6059), .C0(n6058), .Y(n2815)
         );
  OAI211XLTS U677 ( .A0(n3781), .A1(n4034), .B0(n6061), .C0(n6060), .Y(n2816)
         );
  OAI211XLTS U678 ( .A0(n3782), .A1(n4031), .B0(n6063), .C0(n6062), .Y(n2817)
         );
  OAI211XLTS U679 ( .A0(n3782), .A1(n4028), .B0(n6065), .C0(n6064), .Y(n2818)
         );
  OAI211XLTS U680 ( .A0(n3782), .A1(n4025), .B0(n6067), .C0(n6066), .Y(n2819)
         );
  OAI211XLTS U681 ( .A0(n3782), .A1(n4022), .B0(n6069), .C0(n6068), .Y(n2820)
         );
  OAI211XLTS U682 ( .A0(n3783), .A1(n4019), .B0(n6071), .C0(n6070), .Y(n2821)
         );
  OAI211XLTS U683 ( .A0(n3783), .A1(n4016), .B0(n6073), .C0(n6072), .Y(n2822)
         );
  OAI211XLTS U684 ( .A0(n3783), .A1(n4013), .B0(n6075), .C0(n6074), .Y(n2823)
         );
  OAI211XLTS U685 ( .A0(n3783), .A1(n4010), .B0(n6077), .C0(n6076), .Y(n2824)
         );
  OAI211XLTS U686 ( .A0(n3784), .A1(n4004), .B0(n6081), .C0(n6080), .Y(n2826)
         );
  OAI211XLTS U687 ( .A0(n3784), .A1(n4001), .B0(n6083), .C0(n6082), .Y(n2827)
         );
  OAI211XLTS U688 ( .A0(n3784), .A1(n3998), .B0(n6085), .C0(n6084), .Y(n2828)
         );
  OAI211XLTS U689 ( .A0(n3785), .A1(n3992), .B0(n6089), .C0(n6088), .Y(n2830)
         );
  OAI211XLTS U690 ( .A0(n3787), .A1(n3989), .B0(n6091), .C0(n6090), .Y(n2831)
         );
  OAI211XLTS U691 ( .A0(n3777), .A1(n4106), .B0(n5337), .C0(n5336), .Y(n2460)
         );
  OAI211XLTS U692 ( .A0(n3778), .A1(n4094), .B0(n5345), .C0(n5344), .Y(n2464)
         );
  OAI211XLTS U693 ( .A0(n3779), .A1(n4064), .B0(n6041), .C0(n6040), .Y(n2806)
         );
  OAI211XLTS U694 ( .A0(n3779), .A1(n4061), .B0(n6043), .C0(n6042), .Y(n2807)
         );
  OAI211XLTS U695 ( .A0(n3780), .A1(n4049), .B0(n6051), .C0(n6050), .Y(n2811)
         );
  OAI211XLTS U696 ( .A0(n3781), .A1(n4040), .B0(n6057), .C0(n6056), .Y(n2814)
         );
  OAI211XLTS U697 ( .A0(n3784), .A1(n4007), .B0(n6079), .C0(n6078), .Y(n2825)
         );
  OAI211XLTS U698 ( .A0(n3789), .A1(n3995), .B0(n6087), .C0(n6086), .Y(n2829)
         );
  OAI211XLTS U699 ( .A0(n3789), .A1(n3986), .B0(n6093), .C0(n6092), .Y(n2832)
         );
  AOI21XLTS U700 ( .A0(n3819), .A1(n5527), .B0(n5526), .Y(n5528) );
  NAND2XLTS U701 ( .A(n3807), .B(n110), .Y(n5529) );
  AOI2BB2XLTS U702 ( .B0(readReady), .B1(selectBit_WEST), .A0N(n4871), .A1N(
        n6248), .Y(n4865) );
  OAI211XLTS U703 ( .A0(n3935), .A1(n344), .B0(n6191), .C0(n6190), .Y(n2871)
         );
  AOI22XLTS U704 ( .A0(n3409), .A1(n118), .B0(n3392), .B1(n4089), .Y(n6191) );
  OAI211XLTS U705 ( .A0(n3932), .A1(n344), .B0(n6193), .C0(n6192), .Y(n2872)
         );
  OAI211XLTS U706 ( .A0(n3929), .A1(n6205), .B0(n6195), .C0(n6194), .Y(n2873)
         );
  OAI211XLTS U707 ( .A0(n3926), .A1(n344), .B0(n6197), .C0(n6196), .Y(n2874)
         );
  OAI211XLTS U708 ( .A0(n3923), .A1(n6205), .B0(n6199), .C0(n6198), .Y(n2875)
         );
  OAI211XLTS U709 ( .A0(n3920), .A1(n344), .B0(n6204), .C0(n6203), .Y(n2876)
         );
  AOI22XLTS U710 ( .A0(n3408), .A1(n114), .B0(n3392), .B1(n4074), .Y(n6204) );
  OAI211XLTS U711 ( .A0(n3505), .A1(n23), .B0(n6211), .C0(n6210), .Y(n2879) );
  OAI211XLTS U712 ( .A0(n3504), .A1(n22), .B0(n6215), .C0(n6214), .Y(n2881) );
  OAI211XLTS U713 ( .A0(n3505), .A1(n19), .B0(n6207), .C0(n6206), .Y(n2877) );
  OAI211XLTS U714 ( .A0(n3504), .A1(n20), .B0(n6209), .C0(n6208), .Y(n2878) );
  OAI211XLTS U715 ( .A0(n3504), .A1(n21), .B0(n6213), .C0(n6212), .Y(n2880) );
  OAI211XLTS U716 ( .A0(n3505), .A1(n24), .B0(n6221), .C0(n6220), .Y(n2882) );
  OAI211XLTS U717 ( .A0(n3291), .A1(n6282), .B0(n6163), .C0(n6162), .Y(n2861)
         );
  OAI211XLTS U718 ( .A0(n3290), .A1(n6283), .B0(n6165), .C0(n6164), .Y(n2862)
         );
  OAI211XLTS U719 ( .A0(n3290), .A1(n6284), .B0(n6167), .C0(n6166), .Y(n2863)
         );
  OAI211XLTS U720 ( .A0(n3291), .A1(n6285), .B0(n6173), .C0(n6172), .Y(n2864)
         );
  OAI211XLTS U721 ( .A0(n3291), .A1(n6303), .B0(n6159), .C0(n6158), .Y(n2859)
         );
  OAI211XLTS U722 ( .A0(n3290), .A1(n6304), .B0(n6161), .C0(n6160), .Y(n2860)
         );
  OAI211XLTS U723 ( .A0(n3374), .A1(n6307), .B0(n6179), .C0(n6178), .Y(n2867)
         );
  OAI211XLTS U724 ( .A0(n3373), .A1(n6308), .B0(n6181), .C0(n6180), .Y(n2868)
         );
  OAI211XLTS U725 ( .A0(n3373), .A1(n6309), .B0(n6183), .C0(n6182), .Y(n2869)
         );
  OAI211XLTS U726 ( .A0(n3374), .A1(n6305), .B0(n6175), .C0(n6174), .Y(n2865)
         );
  OAI211XLTS U727 ( .A0(n3373), .A1(n6306), .B0(n6177), .C0(n6176), .Y(n2866)
         );
  OAI211XLTS U728 ( .A0(n3374), .A1(n6310), .B0(n6189), .C0(n6188), .Y(n2870)
         );
  OAI211XLTS U729 ( .A0(n771), .A1(n6289), .B0(n6118), .C0(n6117), .Y(n2843)
         );
  OAI211XLTS U730 ( .A0(n770), .A1(n6290), .B0(n6120), .C0(n6119), .Y(n2844)
         );
  OAI211XLTS U731 ( .A0(n770), .A1(n6291), .B0(n6122), .C0(n6121), .Y(n2845)
         );
  OAI211XLTS U732 ( .A0(n771), .A1(n6287), .B0(n6114), .C0(n6113), .Y(n2841)
         );
  OAI211XLTS U733 ( .A0(n770), .A1(n6288), .B0(n6116), .C0(n6115), .Y(n2842)
         );
  OAI211XLTS U734 ( .A0(n771), .A1(n6292), .B0(n6128), .C0(n6127), .Y(n2846)
         );
  OAI211XLTS U735 ( .A0(n4091), .A1(n3738), .B0(n6145), .C0(n6144), .Y(n2853)
         );
  OAI211XLTS U736 ( .A0(n4085), .A1(n3739), .B0(n6149), .C0(n6148), .Y(n2855)
         );
  OAI211XLTS U737 ( .A0(n4082), .A1(n3739), .B0(n6151), .C0(n6150), .Y(n2856)
         );
  OAI211XLTS U738 ( .A0(n4079), .A1(n3739), .B0(n6153), .C0(n6152), .Y(n2857)
         );
  OAI211XLTS U739 ( .A0(n4076), .A1(n3739), .B0(n6157), .C0(n6156), .Y(n2858)
         );
  OAI211XLTS U740 ( .A0(n4088), .A1(n3738), .B0(n6147), .C0(n6146), .Y(n2854)
         );
  OAI211XLTS U741 ( .A0(n4725), .A1(n3517), .B0(n5503), .C0(n5502), .Y(n2558)
         );
  INVXLTS U742 ( .A(n428), .Y(n3517) );
  OAI211XLTS U743 ( .A0(n4734), .A1(n576), .B0(n5479), .C0(n5478), .Y(n2545)
         );
  OAI211XLTS U744 ( .A0(n4745), .A1(n576), .B0(n5481), .C0(n5480), .Y(n2546)
         );
  OAI211XLTS U745 ( .A0(n4754), .A1(n575), .B0(n5483), .C0(n5482), .Y(n2547)
         );
  OAI211XLTS U746 ( .A0(n4763), .A1(n575), .B0(n5485), .C0(n5484), .Y(n2548)
         );
  OAI211XLTS U747 ( .A0(n4446), .A1(n574), .B0(n5655), .C0(n5654), .Y(n2613)
         );
  OAI211XLTS U748 ( .A0(n4496), .A1(n573), .B0(n5667), .C0(n5666), .Y(n2619)
         );
  OAI211XLTS U749 ( .A0(n4516), .A1(n572), .B0(n5671), .C0(n5670), .Y(n2621)
         );
  OAI211XLTS U750 ( .A0(n4523), .A1(n572), .B0(n5673), .C0(n5672), .Y(n2622)
         );
  OAI211XLTS U751 ( .A0(n4590), .A1(n570), .B0(n5687), .C0(n5686), .Y(n2629)
         );
  OAI211XLTS U752 ( .A0(n4601), .A1(n570), .B0(n5689), .C0(n5688), .Y(n2630)
         );
  OAI211XLTS U753 ( .A0(n4613), .A1(n569), .B0(n5693), .C0(n5692), .Y(n2632)
         );
  OAI211XLTS U754 ( .A0(n4649), .A1(n568), .B0(n5701), .C0(n5700), .Y(n2636)
         );
  OAI211XLTS U755 ( .A0(n4696), .A1(n567), .B0(n5711), .C0(n5710), .Y(n2641)
         );
  AOI22XLTS U756 ( .A0(n4137), .A1(n3422), .B0(n4294), .B1(n3698), .Y(n5711)
         );
  OAI211XLTS U757 ( .A0(n4427), .A1(n575), .B0(n5651), .C0(n5650), .Y(n2611)
         );
  OAI211XLTS U758 ( .A0(n4438), .A1(n575), .B0(n5653), .C0(n5652), .Y(n2612)
         );
  OAI211XLTS U759 ( .A0(n4454), .A1(n574), .B0(n5657), .C0(n5656), .Y(n2614)
         );
  OAI211XLTS U760 ( .A0(n4463), .A1(n574), .B0(n5659), .C0(n5658), .Y(n2615)
         );
  OAI211XLTS U761 ( .A0(n4474), .A1(n574), .B0(n5661), .C0(n5660), .Y(n2616)
         );
  OAI211XLTS U762 ( .A0(n4494), .A1(n573), .B0(n5665), .C0(n5664), .Y(n2618)
         );
  OAI211XLTS U763 ( .A0(n4512), .A1(n573), .B0(n5669), .C0(n5668), .Y(n2620)
         );
  OAI211XLTS U764 ( .A0(n4535), .A1(n572), .B0(n5675), .C0(n5674), .Y(n2623)
         );
  OAI211XLTS U765 ( .A0(n4557), .A1(n571), .B0(n5679), .C0(n5678), .Y(n2625)
         );
  OAI211XLTS U766 ( .A0(n4562), .A1(n571), .B0(n5681), .C0(n5680), .Y(n2626)
         );
  OAI211XLTS U767 ( .A0(n4575), .A1(n571), .B0(n5683), .C0(n5682), .Y(n2627)
         );
  OAI211XLTS U768 ( .A0(n4582), .A1(n570), .B0(n5685), .C0(n5684), .Y(n2628)
         );
  OAI211XLTS U769 ( .A0(n4611), .A1(n570), .B0(n5691), .C0(n5690), .Y(n2631)
         );
  OAI211XLTS U770 ( .A0(n4627), .A1(n569), .B0(n5695), .C0(n5694), .Y(n2633)
         );
  OAI211XLTS U771 ( .A0(n4638), .A1(n569), .B0(n5697), .C0(n5696), .Y(n2634)
         );
  OAI211XLTS U772 ( .A0(n4643), .A1(n569), .B0(n5699), .C0(n5698), .Y(n2635)
         );
  OAI211XLTS U773 ( .A0(n4661), .A1(n568), .B0(n5703), .C0(n5702), .Y(n2637)
         );
  OAI211XLTS U774 ( .A0(n4677), .A1(n568), .B0(n5707), .C0(n5706), .Y(n2639)
         );
  OAI211XLTS U775 ( .A0(n4692), .A1(n567), .B0(n5709), .C0(n5708), .Y(n2640)
         );
  OAI211XLTS U776 ( .A0(n4708), .A1(n572), .B0(n5713), .C0(n5712), .Y(n2642)
         );
  AOI22XLTS U777 ( .A0(n4134), .A1(n3422), .B0(n4291), .B1(n3698), .Y(n5713)
         );
  OAI211XLTS U778 ( .A0(n4484), .A1(n573), .B0(n5663), .C0(n5662), .Y(n2617)
         );
  OAI211XLTS U779 ( .A0(n4547), .A1(n571), .B0(n5677), .C0(n5676), .Y(n2624)
         );
  OAI211XLTS U780 ( .A0(n4673), .A1(n568), .B0(n5705), .C0(n5704), .Y(n2638)
         );
  OAI211XLTS U781 ( .A0(n4720), .A1(n567), .B0(n5475), .C0(n5474), .Y(n2543)
         );
  OAI211XLTS U782 ( .A0(n4731), .A1(n576), .B0(n5477), .C0(n5476), .Y(n2544)
         );
  OAI211XLTS U783 ( .A0(n4723), .A1(n3507), .B0(n5501), .C0(n5500), .Y(n2557)
         );
  OAI211XLTS U784 ( .A0(n4429), .A1(n3515), .B0(n5587), .C0(n5586), .Y(n2579)
         );
  OAI211XLTS U785 ( .A0(n4434), .A1(n3515), .B0(n5589), .C0(n5588), .Y(n2580)
         );
  OAI211XLTS U786 ( .A0(n4443), .A1(n3515), .B0(n5591), .C0(n5590), .Y(n2581)
         );
  OAI211XLTS U787 ( .A0(n4456), .A1(n3515), .B0(n5593), .C0(n5592), .Y(n2582)
         );
  OAI211XLTS U788 ( .A0(n4465), .A1(n3514), .B0(n5595), .C0(n5594), .Y(n2583)
         );
  OAI211XLTS U789 ( .A0(n4472), .A1(n3514), .B0(n5597), .C0(n5596), .Y(n2584)
         );
  OAI211XLTS U790 ( .A0(n4481), .A1(n3514), .B0(n5599), .C0(n5598), .Y(n2585)
         );
  OAI211XLTS U791 ( .A0(n4490), .A1(n3514), .B0(n5601), .C0(n5600), .Y(n2586)
         );
  OAI211XLTS U792 ( .A0(n4501), .A1(n3513), .B0(n5603), .C0(n5602), .Y(n2587)
         );
  OAI211XLTS U793 ( .A0(n4506), .A1(n3513), .B0(n5605), .C0(n5604), .Y(n2588)
         );
  OAI211XLTS U794 ( .A0(n4521), .A1(n3513), .B0(n5607), .C0(n5606), .Y(n2589)
         );
  OAI211XLTS U795 ( .A0(n4526), .A1(n3513), .B0(n5609), .C0(n5608), .Y(n2590)
         );
  OAI211XLTS U796 ( .A0(n4539), .A1(n3512), .B0(n5611), .C0(n5610), .Y(n2591)
         );
  OAI211XLTS U797 ( .A0(n4542), .A1(n3512), .B0(n5613), .C0(n5612), .Y(n2592)
         );
  OAI211XLTS U798 ( .A0(n4553), .A1(n3512), .B0(n5615), .C0(n5614), .Y(n2593)
         );
  OAI211XLTS U799 ( .A0(n4564), .A1(n3512), .B0(n5617), .C0(n5616), .Y(n2594)
         );
  OAI211XLTS U800 ( .A0(n4569), .A1(n3511), .B0(n5619), .C0(n5618), .Y(n2595)
         );
  OAI211XLTS U801 ( .A0(n4584), .A1(n3511), .B0(n5621), .C0(n5620), .Y(n2596)
         );
  OAI211XLTS U802 ( .A0(n4587), .A1(n3511), .B0(n5623), .C0(n5622), .Y(n2597)
         );
  OAI211XLTS U803 ( .A0(n4596), .A1(n3510), .B0(n5625), .C0(n5624), .Y(n2598)
         );
  OAI211XLTS U804 ( .A0(n4607), .A1(n3510), .B0(n5627), .C0(n5626), .Y(n2599)
         );
  OAI211XLTS U805 ( .A0(n4620), .A1(n3510), .B0(n5629), .C0(n5628), .Y(n2600)
         );
  OAI211XLTS U806 ( .A0(n4629), .A1(n3510), .B0(n5631), .C0(n5630), .Y(n2601)
         );
  OAI211XLTS U807 ( .A0(n4634), .A1(n3509), .B0(n5633), .C0(n5632), .Y(n2602)
         );
  OAI211XLTS U808 ( .A0(n4641), .A1(n3509), .B0(n5635), .C0(n5634), .Y(n2603)
         );
  OAI211XLTS U809 ( .A0(n4656), .A1(n3511), .B0(n5637), .C0(n5636), .Y(n2604)
         );
  OAI211XLTS U810 ( .A0(n4659), .A1(n3509), .B0(n5639), .C0(n5638), .Y(n2605)
         );
  OAI211XLTS U811 ( .A0(n4668), .A1(n3509), .B0(n5641), .C0(n5640), .Y(n2606)
         );
  OAI211XLTS U812 ( .A0(n4681), .A1(n3508), .B0(n5643), .C0(n5642), .Y(n2607)
         );
  OAI211XLTS U813 ( .A0(n4686), .A1(n3508), .B0(n5645), .C0(n5644), .Y(n2608)
         );
  OAI211XLTS U814 ( .A0(n4699), .A1(n3508), .B0(n5647), .C0(n5646), .Y(n2609)
         );
  OAI211XLTS U815 ( .A0(n4704), .A1(n3508), .B0(n5649), .C0(n5648), .Y(n2610)
         );
  OAI211XLTS U816 ( .A0(n4767), .A1(n3516), .B0(n5511), .C0(n5510), .Y(n2562)
         );
  OAI211XLTS U817 ( .A0(n4735), .A1(n3516), .B0(n5505), .C0(n5504), .Y(n2559)
         );
  OAI211XLTS U818 ( .A0(n4746), .A1(n3516), .B0(n5507), .C0(n5506), .Y(n2560)
         );
  OAI211XLTS U819 ( .A0(n4753), .A1(n3516), .B0(n5509), .C0(n5508), .Y(n2561)
         );
  OAI211XLTS U820 ( .A0(n4718), .A1(n3293), .B0(n5427), .C0(n5426), .Y(n2515)
         );
  OAI211XLTS U821 ( .A0(n4433), .A1(n3301), .B0(n5781), .C0(n5780), .Y(n2676)
         );
  OAI211XLTS U822 ( .A0(n4451), .A1(n3301), .B0(n5785), .C0(n5784), .Y(n2678)
         );
  OAI211XLTS U823 ( .A0(n4462), .A1(n3300), .B0(n5787), .C0(n5786), .Y(n2679)
         );
  OAI211XLTS U824 ( .A0(n4469), .A1(n3300), .B0(n5789), .C0(n5788), .Y(n2680)
         );
  OAI211XLTS U825 ( .A0(n4482), .A1(n3300), .B0(n5791), .C0(n5790), .Y(n2681)
         );
  OAI211XLTS U826 ( .A0(n4487), .A1(n3300), .B0(n5793), .C0(n5792), .Y(n2682)
         );
  OAI211XLTS U827 ( .A0(n4498), .A1(n3299), .B0(n5795), .C0(n5794), .Y(n2683)
         );
  OAI211XLTS U828 ( .A0(n4541), .A1(n3298), .B0(n5805), .C0(n5804), .Y(n2688)
         );
  OAI211XLTS U829 ( .A0(n4586), .A1(n3297), .B0(n5815), .C0(n5814), .Y(n2693)
         );
  OAI211XLTS U830 ( .A0(n4626), .A1(n3296), .B0(n5823), .C0(n5822), .Y(n2697)
         );
  OAI211XLTS U831 ( .A0(n4644), .A1(n3295), .B0(n5827), .C0(n5826), .Y(n2699)
         );
  OAI211XLTS U832 ( .A0(n4660), .A1(n3295), .B0(n5831), .C0(n5830), .Y(n2701)
         );
  OAI211XLTS U833 ( .A0(n4671), .A1(n3295), .B0(n5833), .C0(n5832), .Y(n2702)
         );
  OAI211XLTS U834 ( .A0(n4687), .A1(n3294), .B0(n5837), .C0(n5836), .Y(n2704)
         );
  OAI211XLTS U835 ( .A0(n4425), .A1(n3301), .B0(n5779), .C0(n5778), .Y(n2675)
         );
  OAI211XLTS U836 ( .A0(n4449), .A1(n3301), .B0(n5783), .C0(n5782), .Y(n2677)
         );
  OAI211XLTS U837 ( .A0(n4508), .A1(n3299), .B0(n5797), .C0(n5796), .Y(n2684)
         );
  OAI211XLTS U838 ( .A0(n4519), .A1(n3299), .B0(n5799), .C0(n5798), .Y(n2685)
         );
  OAI211XLTS U839 ( .A0(n4528), .A1(n3299), .B0(n5801), .C0(n5800), .Y(n2686)
         );
  OAI211XLTS U840 ( .A0(n4533), .A1(n3298), .B0(n5803), .C0(n5802), .Y(n2687)
         );
  OAI211XLTS U841 ( .A0(n4560), .A1(n3298), .B0(n5809), .C0(n5808), .Y(n2690)
         );
  OAI211XLTS U842 ( .A0(n4598), .A1(n3296), .B0(n5817), .C0(n5816), .Y(n2694)
         );
  OAI211XLTS U843 ( .A0(n4609), .A1(n3296), .B0(n5819), .C0(n5818), .Y(n2695)
         );
  OAI211XLTS U844 ( .A0(n4616), .A1(n3296), .B0(n5821), .C0(n5820), .Y(n2696)
         );
  OAI211XLTS U845 ( .A0(n4632), .A1(n3295), .B0(n5825), .C0(n5824), .Y(n2698)
         );
  OAI211XLTS U846 ( .A0(n4654), .A1(n3297), .B0(n5829), .C0(n5828), .Y(n2700)
         );
  OAI211XLTS U847 ( .A0(n4695), .A1(n3294), .B0(n5839), .C0(n5838), .Y(n2705)
         );
  OAI211XLTS U848 ( .A0(n4706), .A1(n3294), .B0(n5841), .C0(n5840), .Y(n2706)
         );
  OAI211XLTS U849 ( .A0(n4556), .A1(n3298), .B0(n5807), .C0(n5806), .Y(n2689)
         );
  OAI211XLTS U850 ( .A0(n4574), .A1(n3297), .B0(n5811), .C0(n5810), .Y(n2691)
         );
  OAI211XLTS U851 ( .A0(n4583), .A1(n3297), .B0(n5813), .C0(n5812), .Y(n2692)
         );
  OAI211XLTS U852 ( .A0(n4682), .A1(n3294), .B0(n5835), .C0(n5834), .Y(n2703)
         );
  OAI211XLTS U853 ( .A0(n4738), .A1(n3302), .B0(n5431), .C0(n5430), .Y(n2517)
         );
  OAI211XLTS U854 ( .A0(n4743), .A1(n3302), .B0(n5433), .C0(n5432), .Y(n2518)
         );
  OAI211XLTS U855 ( .A0(n4756), .A1(n3302), .B0(n5435), .C0(n5434), .Y(n2519)
         );
  OAI211XLTS U856 ( .A0(n4761), .A1(n3302), .B0(n5437), .C0(n5436), .Y(n2520)
         );
  OAI211XLTS U857 ( .A0(n4729), .A1(n3303), .B0(n5429), .C0(n5428), .Y(n2516)
         );
  INVXLTS U858 ( .A(n3305), .Y(n3303) );
  OAI211XLTS U859 ( .A0(n4721), .A1(n3376), .B0(n5451), .C0(n5450), .Y(n2529)
         );
  OAI211XLTS U860 ( .A0(n4428), .A1(n3384), .B0(n5715), .C0(n5714), .Y(n2643)
         );
  OAI211XLTS U861 ( .A0(n4563), .A1(n3381), .B0(n5745), .C0(n5744), .Y(n2658)
         );
  OAI211XLTS U862 ( .A0(n4568), .A1(n3380), .B0(n5747), .C0(n5746), .Y(n2659)
         );
  OAI211XLTS U863 ( .A0(n4606), .A1(n3379), .B0(n5755), .C0(n5754), .Y(n2663)
         );
  OAI211XLTS U864 ( .A0(n4698), .A1(n3377), .B0(n5775), .C0(n5774), .Y(n2673)
         );
  OAI211XLTS U865 ( .A0(n4436), .A1(n3384), .B0(n5717), .C0(n5716), .Y(n2644)
         );
  OAI211XLTS U866 ( .A0(n4447), .A1(n3384), .B0(n5719), .C0(n5718), .Y(n2645)
         );
  OAI211XLTS U867 ( .A0(n4458), .A1(n3384), .B0(n5721), .C0(n5720), .Y(n2646)
         );
  OAI211XLTS U868 ( .A0(n4461), .A1(n3383), .B0(n5723), .C0(n5722), .Y(n2647)
         );
  OAI211XLTS U869 ( .A0(n4470), .A1(n3383), .B0(n5725), .C0(n5724), .Y(n2648)
         );
  OAI211XLTS U870 ( .A0(n4485), .A1(n3383), .B0(n5727), .C0(n5726), .Y(n2649)
         );
  OAI211XLTS U871 ( .A0(n4492), .A1(n3383), .B0(n5729), .C0(n5728), .Y(n2650)
         );
  OAI211XLTS U872 ( .A0(n4499), .A1(n3382), .B0(n5731), .C0(n5730), .Y(n2651)
         );
  OAI211XLTS U873 ( .A0(n4510), .A1(n3382), .B0(n5733), .C0(n5732), .Y(n2652)
         );
  OAI211XLTS U874 ( .A0(n4517), .A1(n3382), .B0(n5735), .C0(n5734), .Y(n2653)
         );
  OAI211XLTS U875 ( .A0(n4524), .A1(n3382), .B0(n5737), .C0(n5736), .Y(n2654)
         );
  OAI211XLTS U876 ( .A0(n4537), .A1(n3381), .B0(n5739), .C0(n5738), .Y(n2655)
         );
  OAI211XLTS U877 ( .A0(n4544), .A1(n3381), .B0(n5741), .C0(n5740), .Y(n2656)
         );
  OAI211XLTS U878 ( .A0(n4555), .A1(n3381), .B0(n5743), .C0(n5742), .Y(n2657)
         );
  OAI211XLTS U879 ( .A0(n4578), .A1(n3380), .B0(n5749), .C0(n5748), .Y(n2660)
         );
  OAI211XLTS U880 ( .A0(n4591), .A1(n3380), .B0(n5751), .C0(n5750), .Y(n2661)
         );
  OAI211XLTS U881 ( .A0(n4600), .A1(n3379), .B0(n5753), .C0(n5752), .Y(n2662)
         );
  OAI211XLTS U882 ( .A0(n4614), .A1(n3379), .B0(n5757), .C0(n5756), .Y(n2664)
         );
  OAI211XLTS U883 ( .A0(n4625), .A1(n3379), .B0(n5759), .C0(n5758), .Y(n2665)
         );
  OAI211XLTS U884 ( .A0(n4636), .A1(n3378), .B0(n5761), .C0(n5760), .Y(n2666)
         );
  OAI211XLTS U885 ( .A0(n4645), .A1(n3378), .B0(n5763), .C0(n5762), .Y(n2667)
         );
  OAI211XLTS U886 ( .A0(n4652), .A1(n3380), .B0(n5765), .C0(n5764), .Y(n2668)
         );
  OAI211XLTS U887 ( .A0(n4665), .A1(n3378), .B0(n5767), .C0(n5766), .Y(n2669)
         );
  OAI211XLTS U888 ( .A0(n4672), .A1(n3378), .B0(n5769), .C0(n5768), .Y(n2670)
         );
  OAI211XLTS U889 ( .A0(n4683), .A1(n3377), .B0(n5771), .C0(n5770), .Y(n2671)
         );
  OAI211XLTS U890 ( .A0(n4688), .A1(n3377), .B0(n5773), .C0(n5772), .Y(n2672)
         );
  OAI211XLTS U891 ( .A0(n4710), .A1(n3377), .B0(n5777), .C0(n5776), .Y(n2674)
         );
  OAI211XLTS U892 ( .A0(n4717), .A1(n773), .B0(n5358), .C0(n5357), .Y(n2473)
         );
  OAI211XLTS U893 ( .A0(n4460), .A1(n781), .B0(n5979), .C0(n5978), .Y(n2775)
         );
  OAI211XLTS U894 ( .A0(n4509), .A1(n780), .B0(n5989), .C0(n5988), .Y(n2780)
         );
  OAI211XLTS U895 ( .A0(n4525), .A1(n780), .B0(n5993), .C0(n5992), .Y(n2782)
         );
  OAI211XLTS U896 ( .A0(n4536), .A1(n779), .B0(n5995), .C0(n5994), .Y(n2783)
         );
  OAI211XLTS U897 ( .A0(n4619), .A1(n776), .B0(n6013), .C0(n6012), .Y(n2792)
         );
  OAI211XLTS U898 ( .A0(n4633), .A1(n775), .B0(n6017), .C0(n6016), .Y(n2794)
         );
  OAI211XLTS U899 ( .A0(n4658), .A1(n775), .B0(n6023), .C0(n6022), .Y(n2797)
         );
  OAI211XLTS U900 ( .A0(n4685), .A1(n774), .B0(n6029), .C0(n6028), .Y(n2800)
         );
  OAI211XLTS U901 ( .A0(n4431), .A1(n782), .B0(n5971), .C0(n5970), .Y(n2771)
         );
  OAI211XLTS U902 ( .A0(n4440), .A1(n782), .B0(n5973), .C0(n5972), .Y(n2772)
         );
  OAI211XLTS U903 ( .A0(n4445), .A1(n782), .B0(n5975), .C0(n5974), .Y(n2773)
         );
  OAI211XLTS U904 ( .A0(n4452), .A1(n782), .B0(n5977), .C0(n5976), .Y(n2774)
         );
  OAI211XLTS U905 ( .A0(n4476), .A1(n781), .B0(n5981), .C0(n5980), .Y(n2776)
         );
  OAI211XLTS U906 ( .A0(n4483), .A1(n781), .B0(n5983), .C0(n5982), .Y(n2777)
         );
  OAI211XLTS U907 ( .A0(n4488), .A1(n781), .B0(n5985), .C0(n5984), .Y(n2778)
         );
  OAI211XLTS U908 ( .A0(n4497), .A1(n780), .B0(n5987), .C0(n5986), .Y(n2779)
         );
  OAI211XLTS U909 ( .A0(n4515), .A1(n780), .B0(n5991), .C0(n5990), .Y(n2781)
         );
  OAI211XLTS U910 ( .A0(n4548), .A1(n779), .B0(n5997), .C0(n5996), .Y(n2784)
         );
  OAI211XLTS U911 ( .A0(n4551), .A1(n779), .B0(n5999), .C0(n5998), .Y(n2785)
         );
  OAI211XLTS U912 ( .A0(n4566), .A1(n779), .B0(n6001), .C0(n6000), .Y(n2786)
         );
  OAI211XLTS U913 ( .A0(n4573), .A1(n777), .B0(n6003), .C0(n6002), .Y(n2787)
         );
  OAI211XLTS U914 ( .A0(n4580), .A1(n777), .B0(n6005), .C0(n6004), .Y(n2788)
         );
  OAI211XLTS U915 ( .A0(n4593), .A1(n777), .B0(n6007), .C0(n6006), .Y(n2789)
         );
  OAI211XLTS U916 ( .A0(n4602), .A1(n776), .B0(n6009), .C0(n6008), .Y(n2790)
         );
  OAI211XLTS U917 ( .A0(n4605), .A1(n776), .B0(n6011), .C0(n6010), .Y(n2791)
         );
  OAI211XLTS U918 ( .A0(n4623), .A1(n776), .B0(n6015), .C0(n6014), .Y(n2793)
         );
  OAI211XLTS U919 ( .A0(n4647), .A1(n775), .B0(n6019), .C0(n6018), .Y(n2795)
         );
  OAI211XLTS U920 ( .A0(n4650), .A1(n777), .B0(n6021), .C0(n6020), .Y(n2796)
         );
  OAI211XLTS U921 ( .A0(n4674), .A1(n775), .B0(n6025), .C0(n6024), .Y(n2798)
         );
  OAI211XLTS U922 ( .A0(n4679), .A1(n774), .B0(n6027), .C0(n6026), .Y(n2799)
         );
  OAI211XLTS U923 ( .A0(n4697), .A1(n774), .B0(n6031), .C0(n6030), .Y(n2801)
         );
  OAI211XLTS U924 ( .A0(n4709), .A1(n774), .B0(n6033), .C0(n6032), .Y(n2802)
         );
  OAI211XLTS U925 ( .A0(n4739), .A1(n3385), .B0(n5455), .C0(n5454), .Y(n2531)
         );
  OAI211XLTS U926 ( .A0(n4748), .A1(n3385), .B0(n5457), .C0(n5456), .Y(n2532)
         );
  OAI211XLTS U927 ( .A0(n4757), .A1(n3385), .B0(n5459), .C0(n5458), .Y(n2533)
         );
  OAI211XLTS U928 ( .A0(n4764), .A1(n3385), .B0(n5461), .C0(n5460), .Y(n2534)
         );
  OAI211XLTS U929 ( .A0(n4737), .A1(n783), .B0(n5362), .C0(n5361), .Y(n2475)
         );
  OAI211XLTS U930 ( .A0(n4750), .A1(n783), .B0(n5364), .C0(n5363), .Y(n2476)
         );
  OAI211XLTS U931 ( .A0(n4759), .A1(n783), .B0(n5366), .C0(n5365), .Y(n2477)
         );
  OAI211XLTS U932 ( .A0(n4768), .A1(n783), .B0(n5368), .C0(n5367), .Y(n2478)
         );
  OAI211XLTS U933 ( .A0(n4730), .A1(n3386), .B0(n5453), .C0(n5452), .Y(n2530)
         );
  INVXLTS U934 ( .A(n3387), .Y(n3386) );
  OAI211XLTS U935 ( .A0(n3731), .A1(n4106), .B0(n5407), .C0(n5406), .Y(n2502)
         );
  OAI211XLTS U936 ( .A0(n3731), .A1(n4103), .B0(n5409), .C0(n5408), .Y(n2503)
         );
  OAI211XLTS U937 ( .A0(n3731), .A1(n4100), .B0(n5411), .C0(n5410), .Y(n2504)
         );
  OAI211XLTS U938 ( .A0(n3731), .A1(n4109), .B0(n5405), .C0(n5404), .Y(n2501)
         );
  OAI211XLTS U939 ( .A0(n3738), .A1(n3983), .B0(n5903), .C0(n5902), .Y(n2737)
         );
  OAI211XLTS U940 ( .A0(n3738), .A1(n3980), .B0(n5905), .C0(n5904), .Y(n2738)
         );
  OAI211XLTS U941 ( .A0(n3741), .A1(n4097), .B0(n5413), .C0(n5412), .Y(n2505)
         );
  OAI211XLTS U942 ( .A0(n3742), .A1(n4094), .B0(n5415), .C0(n5414), .Y(n2506)
         );
  OAI211XLTS U943 ( .A0(n3742), .A1(n4073), .B0(n5843), .C0(n5842), .Y(n2707)
         );
  OAI211XLTS U944 ( .A0(n3744), .A1(n4070), .B0(n5845), .C0(n5844), .Y(n2708)
         );
  OAI211XLTS U945 ( .A0(n3743), .A1(n4067), .B0(n5847), .C0(n5846), .Y(n2709)
         );
  OAI211XLTS U946 ( .A0(n3743), .A1(n4064), .B0(n5849), .C0(n5848), .Y(n2710)
         );
  OAI211XLTS U947 ( .A0(n6343), .A1(n4061), .B0(n5851), .C0(n5850), .Y(n2711)
         );
  OAI211XLTS U948 ( .A0(n3743), .A1(n4058), .B0(n5853), .C0(n5852), .Y(n2712)
         );
  OAI211XLTS U949 ( .A0(n3732), .A1(n4052), .B0(n5857), .C0(n5856), .Y(n2714)
         );
  OAI211XLTS U950 ( .A0(n3732), .A1(n4046), .B0(n5861), .C0(n5860), .Y(n2716)
         );
  OAI211XLTS U951 ( .A0(n3733), .A1(n4043), .B0(n5863), .C0(n5862), .Y(n2717)
         );
  OAI211XLTS U952 ( .A0(n3733), .A1(n4037), .B0(n5867), .C0(n5866), .Y(n2719)
         );
  OAI211XLTS U953 ( .A0(n3734), .A1(n4031), .B0(n5871), .C0(n5870), .Y(n2721)
         );
  OAI211XLTS U954 ( .A0(n3734), .A1(n4028), .B0(n5873), .C0(n5872), .Y(n2722)
         );
  OAI211XLTS U955 ( .A0(n3734), .A1(n4022), .B0(n5877), .C0(n5876), .Y(n2724)
         );
  OAI211XLTS U956 ( .A0(n3735), .A1(n4016), .B0(n5881), .C0(n5880), .Y(n2726)
         );
  OAI211XLTS U957 ( .A0(n3735), .A1(n4013), .B0(n5883), .C0(n5882), .Y(n2727)
         );
  OAI211XLTS U958 ( .A0(n3735), .A1(n4010), .B0(n5885), .C0(n5884), .Y(n2728)
         );
  OAI211XLTS U959 ( .A0(n3736), .A1(n4007), .B0(n5887), .C0(n5886), .Y(n2729)
         );
  OAI211XLTS U960 ( .A0(n3736), .A1(n4004), .B0(n5889), .C0(n5888), .Y(n2730)
         );
  OAI211XLTS U961 ( .A0(n3736), .A1(n3998), .B0(n5893), .C0(n5892), .Y(n2732)
         );
  OAI211XLTS U962 ( .A0(n3737), .A1(n3989), .B0(n5899), .C0(n5898), .Y(n2735)
         );
  OAI211XLTS U963 ( .A0(n3732), .A1(n4055), .B0(n5855), .C0(n5854), .Y(n2713)
         );
  OAI211XLTS U964 ( .A0(n3732), .A1(n4049), .B0(n5859), .C0(n5858), .Y(n2715)
         );
  OAI211XLTS U965 ( .A0(n3733), .A1(n4040), .B0(n5865), .C0(n5864), .Y(n2718)
         );
  OAI211XLTS U966 ( .A0(n3733), .A1(n4034), .B0(n5869), .C0(n5868), .Y(n2720)
         );
  OAI211XLTS U967 ( .A0(n3734), .A1(n4025), .B0(n5875), .C0(n5874), .Y(n2723)
         );
  OAI211XLTS U968 ( .A0(n3735), .A1(n4019), .B0(n5879), .C0(n5878), .Y(n2725)
         );
  OAI211XLTS U969 ( .A0(n3737), .A1(n3995), .B0(n5895), .C0(n5894), .Y(n2733)
         );
  OAI211XLTS U970 ( .A0(n3737), .A1(n3992), .B0(n5897), .C0(n5896), .Y(n2734)
         );
  OAI211XLTS U971 ( .A0(n3737), .A1(n3986), .B0(n5901), .C0(n5900), .Y(n2736)
         );
  OAI211XLTS U972 ( .A0(n3736), .A1(n4001), .B0(n5891), .C0(n5890), .Y(n2731)
         );
  OAI2BB1XLTS U973 ( .A0N(n4843), .A1N(n4871), .B0(n4842), .Y(n4854) );
  AOI32XLTS U974 ( .A0(n336), .A1(n6236), .A2(n191), .B0(n340), .B1(n4841), 
        .Y(n4842) );
  XNOR2XLTS U975 ( .A(n6235), .B(n6248), .Y(n4841) );
  AOI32XLTS U976 ( .A0(n166), .A1(n5565), .A2(n5564), .B0(n3520), .B1(n104), 
        .Y(n2570) );
  AOI22XLTS U977 ( .A0(n3812), .A1(n5563), .B0(n3807), .B1(n5562), .Y(n5564)
         );
  AOI32XLTS U978 ( .A0(n112), .A1(n5544), .A2(n5543), .B0(n3304), .B1(n103), 
        .Y(n2567) );
  AOI32XLTS U979 ( .A0(n165), .A1(n5558), .A2(n5557), .B0(n579), .B1(n11), .Y(
        n2569) );
  NAND2XLTS U980 ( .A(n3806), .B(n5553), .Y(n5558) );
  INVXLTS U981 ( .A(selectBit_WEST), .Y(n6236) );
  AOI22XLTS U982 ( .A0(n5517), .A1(n5516), .B0(n184), .B1(n26), .Y(n2563) );
  AOI31XLTS U983 ( .A0(n5515), .A1(n169), .A2(readIn_SOUTH), .B0(n5514), .Y(
        n5516) );
  AOI21XLTS U984 ( .A0(n3819), .A1(n164), .B0(n6345), .Y(n5517) );
  OAI32XLTS U985 ( .A0(n3815), .A1(n6338), .A2(n5539), .B0(n5513), .B1(n3808), 
        .Y(n5514) );
  NAND2XLTS U986 ( .A(n172), .B(n120), .Y(n5439) );
  AOI32XLTS U987 ( .A0(n5536), .A1(n5535), .A2(n3812), .B0(n5534), .B1(n5533), 
        .Y(n5537) );
  AOI21XLTS U988 ( .A0(n3807), .A1(n6334), .B0(n173), .Y(n5538) );
  OAI22XLTS U989 ( .A0(n157), .A1(n193), .B0(n6323), .B1(n3821), .Y(n5533) );
  NAND3XLTS U990 ( .A(n4870), .B(n6250), .C(n341), .Y(n5305) );
  NAND3XLTS U991 ( .A(n422), .B(n4871), .C(n120), .Y(n5306) );
  NAND3XLTS U992 ( .A(n4870), .B(n189), .C(n119), .Y(n5304) );
  NAND4XLTS U993 ( .A(n340), .B(n422), .C(n6235), .D(n215), .Y(n5307) );
  NAND4XLTS U994 ( .A(n336), .B(n422), .C(n215), .D(n6236), .Y(n5303) );
  OAI31XLTS U995 ( .A0(n4835), .A1(n5314), .A2(n5313), .B0(n5312), .Y(n2450)
         );
  OAI31XLTS U996 ( .A0(n4833), .A1(n5314), .A2(n5313), .B0(n5297), .Y(n2449)
         );
  NOR3X1TS U997 ( .A(n195), .B(n3), .C(n276), .Y(n5287) );
  OAI2BB2XLTS U998 ( .B0(n6287), .B1(n3552), .A0N(
        \requesterAddressbuffer[2][5] ), .A1N(n180), .Y(n5130) );
  OAI2BB2XLTS U999 ( .B0(n6288), .B1(n3552), .A0N(
        \requesterAddressbuffer[2][4] ), .A1N(n180), .Y(n5138) );
  OAI2BB2XLTS U1000 ( .B0(n6290), .B1(n3551), .A0N(
        \requesterAddressbuffer[2][2] ), .A1N(n179), .Y(n5154) );
  OAI2BB2XLTS U1001 ( .B0(n6291), .B1(n3551), .A0N(
        \requesterAddressbuffer[2][1] ), .A1N(n179), .Y(n5162) );
  OAI2BB2XLTS U1002 ( .B0(n6289), .B1(n3551), .A0N(
        \requesterAddressbuffer[2][3] ), .A1N(n180), .Y(n5146) );
  OAI2BB2XLTS U1003 ( .B0(n6292), .B1(n3551), .A0N(
        \requesterAddressbuffer[2][0] ), .A1N(n180), .Y(n5170) );
  NAND2X1TS U1004 ( .A(n5), .B(n275), .Y(n6226) );
  AND2XLTS U1005 ( .A(n5512), .B(n5322), .Y(n421) );
  CLKBUFX2TS U1006 ( .A(n4872), .Y(n422) );
  CLKBUFX2TS U1007 ( .A(n3742), .Y(n3732) );
  CLKBUFX2TS U1008 ( .A(n3742), .Y(n3733) );
  CLKBUFX2TS U1009 ( .A(n3740), .Y(n3734) );
  CLKBUFX2TS U1010 ( .A(n3741), .Y(n3735) );
  CLKBUFX2TS U1011 ( .A(n3741), .Y(n3737) );
  CLKBUFX2TS U1012 ( .A(n3741), .Y(n3736) );
  CLKBUFX2TS U1013 ( .A(n3740), .Y(n3738) );
  CLKBUFX2TS U1014 ( .A(n3740), .Y(n3739) );
  CLKBUFX2TS U1015 ( .A(n3744), .Y(n3740) );
  CLKBUFX2TS U1016 ( .A(n6343), .Y(n3742) );
  CLKBUFX2TS U1017 ( .A(n3744), .Y(n3741) );
  CLKBUFX2TS U1018 ( .A(n3728), .Y(n3718) );
  CLKBUFX2TS U1019 ( .A(n3729), .Y(n3725) );
  CLKBUFX2TS U1020 ( .A(n3726), .Y(n3724) );
  CLKBUFX2TS U1021 ( .A(n3727), .Y(n3723) );
  CLKBUFX2TS U1022 ( .A(n3728), .Y(n3721) );
  CLKBUFX2TS U1023 ( .A(n3728), .Y(n3720) );
  CLKBUFX2TS U1024 ( .A(n3700), .Y(n3690) );
  CLKBUFX2TS U1025 ( .A(n3699), .Y(n3693) );
  CLKBUFX2TS U1026 ( .A(n3699), .Y(n3694) );
  CLKBUFX2TS U1027 ( .A(n3698), .Y(n3695) );
  CLKBUFX2TS U1028 ( .A(n3672), .Y(n3661) );
  CLKBUFX2TS U1029 ( .A(n3671), .Y(n3662) );
  CLKBUFX2TS U1030 ( .A(n3671), .Y(n3663) );
  CLKBUFX2TS U1031 ( .A(n3671), .Y(n3664) );
  CLKBUFX2TS U1032 ( .A(n3670), .Y(n3665) );
  CLKBUFX2TS U1033 ( .A(n3670), .Y(n3666) );
  CLKBUFX2TS U1034 ( .A(n3669), .Y(n3667) );
  CLKBUFX2TS U1035 ( .A(n3669), .Y(n3668) );
  CLKBUFX2TS U1036 ( .A(n3727), .Y(n3722) );
  CLKBUFX2TS U1037 ( .A(n3728), .Y(n3719) );
  CLKBUFX2TS U1038 ( .A(n3700), .Y(n3691) );
  CLKBUFX2TS U1039 ( .A(n3700), .Y(n3692) );
  CLKBUFX2TS U1040 ( .A(n3698), .Y(n3696) );
  CLKBUFX2TS U1041 ( .A(n3687), .Y(n3681) );
  CLKBUFX2TS U1042 ( .A(n3685), .Y(n3677) );
  CLKBUFX2TS U1043 ( .A(n3685), .Y(n3676) );
  CLKBUFX2TS U1044 ( .A(n3686), .Y(n3675) );
  CLKBUFX2TS U1045 ( .A(n3684), .Y(n3679) );
  CLKBUFX2TS U1046 ( .A(n3685), .Y(n3680) );
  CLKBUFX2TS U1047 ( .A(n3684), .Y(n3678) );
  CLKBUFX2TS U1048 ( .A(n3686), .Y(n3674) );
  CLKBUFX2TS U1049 ( .A(n6341), .Y(n3697) );
  CLKBUFX2TS U1050 ( .A(n228), .Y(n3791) );
  CLKBUFX2TS U1051 ( .A(n3800), .Y(n3792) );
  CLKBUFX2TS U1052 ( .A(n3798), .Y(n3797) );
  CLKBUFX2TS U1053 ( .A(n3798), .Y(n3796) );
  CLKBUFX2TS U1054 ( .A(n3799), .Y(n3795) );
  CLKBUFX2TS U1055 ( .A(n3799), .Y(n3794) );
  CLKBUFX2TS U1056 ( .A(n3800), .Y(n3793) );
  CLKBUFX2TS U1057 ( .A(n3688), .Y(n3682) );
  CLKBUFX2TS U1058 ( .A(n3786), .Y(n3782) );
  CLKBUFX2TS U1059 ( .A(n3786), .Y(n3783) );
  CLKBUFX2TS U1060 ( .A(n3788), .Y(n3778) );
  CLKBUFX2TS U1061 ( .A(n3788), .Y(n3779) );
  CLKBUFX2TS U1062 ( .A(n3787), .Y(n3780) );
  CLKBUFX2TS U1063 ( .A(n3787), .Y(n3781) );
  CLKBUFX2TS U1064 ( .A(n3785), .Y(n3784) );
  CLKBUFX2TS U1065 ( .A(n3743), .Y(n3731) );
  CLKBUFX2TS U1066 ( .A(n6343), .Y(n3743) );
  CLKBUFX2TS U1067 ( .A(n3688), .Y(n3683) );
  CLKBUFX2TS U1068 ( .A(n3802), .Y(n3798) );
  CLKBUFX2TS U1069 ( .A(n3802), .Y(n3799) );
  CLKBUFX2TS U1070 ( .A(n3802), .Y(n3800) );
  CLKBUFX2TS U1071 ( .A(n3730), .Y(n3726) );
  CLKBUFX2TS U1072 ( .A(n6341), .Y(n3699) );
  CLKBUFX2TS U1073 ( .A(n3687), .Y(n3685) );
  CLKBUFX2TS U1074 ( .A(n3673), .Y(n3671) );
  CLKBUFX2TS U1075 ( .A(n3673), .Y(n3670) );
  CLKBUFX2TS U1076 ( .A(n3673), .Y(n3669) );
  CLKBUFX2TS U1077 ( .A(n265), .Y(n3727) );
  CLKBUFX2TS U1078 ( .A(n3730), .Y(n3728) );
  CLKBUFX2TS U1079 ( .A(n3687), .Y(n3684) );
  CLKBUFX2TS U1080 ( .A(n3702), .Y(n3700) );
  CLKBUFX2TS U1081 ( .A(n3687), .Y(n3686) );
  CLKBUFX2TS U1082 ( .A(n6341), .Y(n3698) );
  CLKBUFX2TS U1083 ( .A(n6346), .Y(n3786) );
  CLKBUFX2TS U1084 ( .A(n6346), .Y(n3788) );
  CLKBUFX2TS U1085 ( .A(n6346), .Y(n3787) );
  CLKBUFX2TS U1086 ( .A(n6346), .Y(n3785) );
  CLKBUFX2TS U1087 ( .A(n6343), .Y(n3744) );
  CLKBUFX2TS U1088 ( .A(n3322), .Y(n3308) );
  CLKBUFX2TS U1089 ( .A(n3322), .Y(n3309) );
  CLKBUFX2TS U1090 ( .A(n3319), .Y(n3315) );
  CLKBUFX2TS U1091 ( .A(n3320), .Y(n3313) );
  CLKBUFX2TS U1092 ( .A(n3320), .Y(n3312) );
  CLKBUFX2TS U1093 ( .A(n3319), .Y(n3314) );
  CLKBUFX2TS U1094 ( .A(n3321), .Y(n3311) );
  CLKBUFX2TS U1095 ( .A(n3321), .Y(n3310) );
  CLKBUFX2TS U1096 ( .A(n3449), .Y(n3447) );
  CLKBUFX2TS U1097 ( .A(n3450), .Y(n3446) );
  CLKBUFX2TS U1098 ( .A(n3451), .Y(n3444) );
  CLKBUFX2TS U1099 ( .A(n3451), .Y(n3443) );
  CLKBUFX2TS U1100 ( .A(n3452), .Y(n3442) );
  CLKBUFX2TS U1101 ( .A(n3452), .Y(n3441) );
  CLKBUFX2TS U1102 ( .A(n3453), .Y(n3440) );
  CLKBUFX2TS U1103 ( .A(n3453), .Y(n3439) );
  CLKBUFX2TS U1104 ( .A(n3450), .Y(n3445) );
  CLKBUFX2TS U1105 ( .A(n803), .Y(n789) );
  CLKBUFX2TS U1106 ( .A(n3729), .Y(n3717) );
  CLKBUFX2TS U1107 ( .A(n3730), .Y(n3729) );
  CLKBUFX2TS U1108 ( .A(n3713), .Y(n3704) );
  CLKBUFX2TS U1109 ( .A(n3771), .Y(n3762) );
  CLKBUFX2TS U1110 ( .A(n803), .Y(n790) );
  CLKBUFX2TS U1111 ( .A(n801), .Y(n793) );
  CLKBUFX2TS U1112 ( .A(n3769), .Y(n3767) );
  CLKBUFX2TS U1113 ( .A(n3769), .Y(n3766) );
  CLKBUFX2TS U1114 ( .A(n3770), .Y(n3765) );
  CLKBUFX2TS U1115 ( .A(n3770), .Y(n3764) );
  CLKBUFX2TS U1116 ( .A(n3771), .Y(n3763) );
  CLKBUFX2TS U1117 ( .A(n798), .Y(n796) );
  CLKBUFX2TS U1118 ( .A(n3709), .Y(n3708) );
  CLKBUFX2TS U1119 ( .A(n3712), .Y(n3707) );
  CLKBUFX2TS U1120 ( .A(n3712), .Y(n3706) );
  CLKBUFX2TS U1121 ( .A(n3713), .Y(n3705) );
  CLKBUFX2TS U1122 ( .A(n800), .Y(n795) );
  CLKBUFX2TS U1123 ( .A(n801), .Y(n794) );
  CLKBUFX2TS U1124 ( .A(n802), .Y(n792) );
  CLKBUFX2TS U1125 ( .A(n802), .Y(n791) );
  CLKBUFX2TS U1126 ( .A(n3672), .Y(n3660) );
  CLKBUFX2TS U1127 ( .A(n6339), .Y(n3672) );
  CLKBUFX2TS U1128 ( .A(n3701), .Y(n3689) );
  CLKBUFX2TS U1129 ( .A(n3702), .Y(n3701) );
  CLKBUFX2TS U1130 ( .A(n767), .Y(n753) );
  CLKBUFX2TS U1131 ( .A(n3370), .Y(n3356) );
  CLKBUFX2TS U1132 ( .A(n3370), .Y(n3357) );
  CLKBUFX2TS U1133 ( .A(n767), .Y(n754) );
  CLKBUFX2TS U1134 ( .A(n3205), .Y(n1894) );
  CLKBUFX2TS U1135 ( .A(n3205), .Y(n3192) );
  CLKBUFX2TS U1136 ( .A(n3449), .Y(n3448) );
  CLKBUFX2TS U1137 ( .A(n3282), .Y(n3280) );
  CLKBUFX2TS U1138 ( .A(n769), .Y(n761) );
  CLKBUFX2TS U1139 ( .A(n764), .Y(n760) );
  CLKBUFX2TS U1140 ( .A(n765), .Y(n758) );
  CLKBUFX2TS U1141 ( .A(n765), .Y(n757) );
  CLKBUFX2TS U1142 ( .A(n764), .Y(n759) );
  CLKBUFX2TS U1143 ( .A(n766), .Y(n756) );
  CLKBUFX2TS U1144 ( .A(n766), .Y(n755) );
  CLKBUFX2TS U1145 ( .A(n3283), .Y(n3279) );
  CLKBUFX2TS U1146 ( .A(n3283), .Y(n3278) );
  CLKBUFX2TS U1147 ( .A(n3284), .Y(n3277) );
  CLKBUFX2TS U1148 ( .A(n3284), .Y(n3276) );
  CLKBUFX2TS U1149 ( .A(n3286), .Y(n3274) );
  CLKBUFX2TS U1150 ( .A(n3365), .Y(n3362) );
  CLKBUFX2TS U1151 ( .A(n3368), .Y(n3361) );
  CLKBUFX2TS U1152 ( .A(n3368), .Y(n3360) );
  CLKBUFX2TS U1153 ( .A(n3369), .Y(n3359) );
  CLKBUFX2TS U1154 ( .A(n3369), .Y(n3358) );
  CLKBUFX2TS U1155 ( .A(n685), .Y(n671) );
  CLKBUFX2TS U1156 ( .A(n685), .Y(n672) );
  CLKBUFX2TS U1157 ( .A(n837), .Y(n820) );
  CLKBUFX2TS U1158 ( .A(n837), .Y(n821) );
  CLKBUFX2TS U1159 ( .A(n3285), .Y(n3275) );
  CLKBUFX2TS U1160 ( .A(n3286), .Y(n3273) );
  CLKBUFX2TS U1161 ( .A(n836), .Y(n822) );
  CLKBUFX2TS U1162 ( .A(n3205), .Y(n3193) );
  CLKBUFX2TS U1163 ( .A(n835), .Y(n826) );
  CLKBUFX2TS U1164 ( .A(n835), .Y(n824) );
  CLKBUFX2TS U1165 ( .A(n832), .Y(n829) );
  CLKBUFX2TS U1166 ( .A(n834), .Y(n827) );
  CLKBUFX2TS U1167 ( .A(n834), .Y(n828) );
  CLKBUFX2TS U1168 ( .A(n836), .Y(n823) );
  CLKBUFX2TS U1169 ( .A(n3255), .Y(n3242) );
  CLKBUFX2TS U1170 ( .A(n683), .Y(n676) );
  CLKBUFX2TS U1171 ( .A(n3202), .Y(n3200) );
  CLKBUFX2TS U1172 ( .A(n3203), .Y(n3199) );
  CLKBUFX2TS U1173 ( .A(n3203), .Y(n3198) );
  CLKBUFX2TS U1174 ( .A(n3204), .Y(n3197) );
  CLKBUFX2TS U1175 ( .A(n3204), .Y(n3196) );
  CLKBUFX2TS U1176 ( .A(n3207), .Y(n3195) );
  CLKBUFX2TS U1177 ( .A(n3205), .Y(n3194) );
  CLKBUFX2TS U1178 ( .A(n682), .Y(n677) );
  CLKBUFX2TS U1179 ( .A(n683), .Y(n675) );
  CLKBUFX2TS U1180 ( .A(n684), .Y(n674) );
  CLKBUFX2TS U1181 ( .A(n832), .Y(n830) );
  CLKBUFX2TS U1182 ( .A(n3202), .Y(n3201) );
  CLKBUFX2TS U1183 ( .A(n3757), .Y(n3747) );
  CLKBUFX2TS U1184 ( .A(n3754), .Y(n3753) );
  CLKBUFX2TS U1185 ( .A(n3756), .Y(n3750) );
  CLKBUFX2TS U1186 ( .A(n3754), .Y(n3752) );
  CLKBUFX2TS U1187 ( .A(n3760), .Y(n3751) );
  CLKBUFX2TS U1188 ( .A(n3756), .Y(n3749) );
  CLKBUFX2TS U1189 ( .A(n3757), .Y(n3748) );
  CLKBUFX2TS U1190 ( .A(n3252), .Y(n3249) );
  CLKBUFX2TS U1191 ( .A(n3252), .Y(n3250) );
  CLKBUFX2TS U1192 ( .A(n3253), .Y(n3248) );
  CLKBUFX2TS U1193 ( .A(n3254), .Y(n3245) );
  CLKBUFX2TS U1194 ( .A(n3258), .Y(n3244) );
  CLKBUFX2TS U1195 ( .A(n3253), .Y(n3247) );
  CLKBUFX2TS U1196 ( .A(n3254), .Y(n3246) );
  CLKBUFX2TS U1197 ( .A(n3258), .Y(n3243) );
  CLKBUFX2TS U1198 ( .A(n3801), .Y(n3790) );
  CLKBUFX2TS U1199 ( .A(n3802), .Y(n3801) );
  CLKBUFX2TS U1200 ( .A(n3789), .Y(n3777) );
  CLKBUFX2TS U1201 ( .A(n3786), .Y(n3789) );
  INVX2TS U1202 ( .A(n1728), .Y(n1402) );
  INVX2TS U1203 ( .A(n1764), .Y(n986) );
  INVX2TS U1204 ( .A(n1654), .Y(n1602) );
  CLKBUFX2TS U1205 ( .A(n702), .Y(n688) );
  CLKBUFX2TS U1206 ( .A(n702), .Y(n689) );
  CLKBUFX2TS U1207 ( .A(n698), .Y(n697) );
  CLKBUFX2TS U1208 ( .A(n698), .Y(n696) );
  CLKBUFX2TS U1209 ( .A(n699), .Y(n695) );
  CLKBUFX2TS U1210 ( .A(n700), .Y(n693) );
  CLKBUFX2TS U1211 ( .A(n700), .Y(n692) );
  CLKBUFX2TS U1212 ( .A(n699), .Y(n694) );
  CLKBUFX2TS U1213 ( .A(n701), .Y(n691) );
  CLKBUFX2TS U1214 ( .A(n701), .Y(n690) );
  CLKBUFX2TS U1215 ( .A(n668), .Y(n661) );
  CLKBUFX2TS U1216 ( .A(n667), .Y(n662) );
  CLKBUFX2TS U1217 ( .A(n668), .Y(n627) );
  CLKBUFX2TS U1218 ( .A(n667), .Y(n659) );
  CLKBUFX2TS U1219 ( .A(n668), .Y(n660) );
  CLKBUFX2TS U1220 ( .A(n667), .Y(n663) );
  CLKBUFX2TS U1221 ( .A(n666), .Y(n664) );
  CLKBUFX2TS U1222 ( .A(n666), .Y(n665) );
  CLKBUFX2TS U1223 ( .A(n1822), .Y(n1654) );
  CLKBUFX2TS U1224 ( .A(n1822), .Y(n1728) );
  CLKBUFX2TS U1225 ( .A(n1822), .Y(n1764) );
  CLKBUFX2TS U1226 ( .A(n856), .Y(n851) );
  CLKBUFX2TS U1227 ( .A(n856), .Y(n853) );
  CLKBUFX2TS U1228 ( .A(n856), .Y(n852) );
  CLKBUFX2TS U1229 ( .A(n3288), .Y(n3287) );
  CLKBUFX2TS U1230 ( .A(n805), .Y(n799) );
  CLKBUFX2TS U1231 ( .A(n805), .Y(n800) );
  CLKBUFX2TS U1232 ( .A(n804), .Y(n801) );
  CLKBUFX2TS U1233 ( .A(n804), .Y(n802) );
  CLKBUFX2TS U1234 ( .A(n804), .Y(n803) );
  CLKBUFX2TS U1235 ( .A(n3288), .Y(n3285) );
  CLKBUFX2TS U1236 ( .A(n3288), .Y(n3286) );
  CLKBUFX2TS U1237 ( .A(n838), .Y(n835) );
  CLKBUFX2TS U1238 ( .A(n3760), .Y(n3754) );
  CLKBUFX2TS U1239 ( .A(n839), .Y(n832) );
  CLKBUFX2TS U1240 ( .A(n3760), .Y(n3755) );
  CLKBUFX2TS U1241 ( .A(n839), .Y(n833) );
  CLKBUFX2TS U1242 ( .A(n3759), .Y(n3756) );
  CLKBUFX2TS U1243 ( .A(n839), .Y(n834) );
  CLKBUFX2TS U1244 ( .A(n3759), .Y(n3757) );
  CLKBUFX2TS U1245 ( .A(n838), .Y(n836) );
  CLKBUFX2TS U1246 ( .A(n3256), .Y(n3255) );
  CLKBUFX2TS U1247 ( .A(n3372), .Y(n3365) );
  CLKBUFX2TS U1248 ( .A(n687), .Y(n680) );
  CLKBUFX2TS U1249 ( .A(n769), .Y(n763) );
  CLKBUFX2TS U1250 ( .A(n3774), .Y(n3768) );
  CLKBUFX2TS U1251 ( .A(n3774), .Y(n3769) );
  CLKBUFX2TS U1252 ( .A(n768), .Y(n765) );
  CLKBUFX2TS U1253 ( .A(n769), .Y(n764) );
  CLKBUFX2TS U1254 ( .A(n3773), .Y(n3770) );
  CLKBUFX2TS U1255 ( .A(n768), .Y(n766) );
  CLKBUFX2TS U1256 ( .A(n3206), .Y(n3202) );
  CLKBUFX2TS U1257 ( .A(n3206), .Y(n3203) );
  CLKBUFX2TS U1258 ( .A(n3206), .Y(n3204) );
  CLKBUFX2TS U1259 ( .A(n3257), .Y(n3252) );
  CLKBUFX2TS U1260 ( .A(n3324), .Y(n3317) );
  CLKBUFX2TS U1261 ( .A(n3716), .Y(n3709) );
  CLKBUFX2TS U1262 ( .A(n3372), .Y(n3366) );
  CLKBUFX2TS U1263 ( .A(n3324), .Y(n3318) );
  CLKBUFX2TS U1264 ( .A(n3716), .Y(n3710) );
  CLKBUFX2TS U1265 ( .A(n3716), .Y(n3711) );
  CLKBUFX2TS U1266 ( .A(n3371), .Y(n3368) );
  CLKBUFX2TS U1267 ( .A(n3323), .Y(n3320) );
  CLKBUFX2TS U1268 ( .A(n3372), .Y(n3367) );
  CLKBUFX2TS U1269 ( .A(n3324), .Y(n3319) );
  CLKBUFX2TS U1270 ( .A(n3715), .Y(n3712) );
  CLKBUFX2TS U1271 ( .A(n3371), .Y(n3369) );
  CLKBUFX2TS U1272 ( .A(n3323), .Y(n3321) );
  CLKBUFX2TS U1273 ( .A(n3715), .Y(n3713) );
  CLKBUFX2TS U1274 ( .A(n3371), .Y(n3370) );
  CLKBUFX2TS U1275 ( .A(n3323), .Y(n3322) );
  CLKBUFX2TS U1276 ( .A(n3454), .Y(n3451) );
  CLKBUFX2TS U1277 ( .A(n3454), .Y(n3452) );
  CLKBUFX2TS U1278 ( .A(n3454), .Y(n3453) );
  CLKBUFX2TS U1279 ( .A(n3455), .Y(n3450) );
  CLKBUFX2TS U1280 ( .A(n686), .Y(n685) );
  CLKBUFX2TS U1281 ( .A(n687), .Y(n681) );
  CLKBUFX2TS U1282 ( .A(n687), .Y(n682) );
  CLKBUFX2TS U1283 ( .A(n686), .Y(n683) );
  CLKBUFX2TS U1284 ( .A(n686), .Y(n684) );
  CLKBUFX2TS U1285 ( .A(n768), .Y(n767) );
  CLKBUFX2TS U1286 ( .A(n3773), .Y(n3771) );
  CLKBUFX2TS U1287 ( .A(n838), .Y(n837) );
  CLKBUFX2TS U1288 ( .A(n3257), .Y(n3253) );
  CLKBUFX2TS U1289 ( .A(n3257), .Y(n3254) );
  CLKBUFX2TS U1290 ( .A(n3289), .Y(n3283) );
  CLKBUFX2TS U1291 ( .A(n3289), .Y(n3284) );
  CLKBUFX2TS U1292 ( .A(n265), .Y(n3730) );
  CLKBUFX2TS U1293 ( .A(n421), .Y(n3802) );
  CLKBUFX2TS U1294 ( .A(n6341), .Y(n3702) );
  CLKBUFX2TS U1295 ( .A(n6340), .Y(n3687) );
  CLKBUFX2TS U1296 ( .A(n6339), .Y(n3673) );
  INVX2TS U1297 ( .A(n5576), .Y(n6343) );
  CLKBUFX2TS U1298 ( .A(n3240), .Y(n3225) );
  CLKBUFX2TS U1299 ( .A(n3240), .Y(n3226) );
  CLKBUFX2TS U1300 ( .A(n3236), .Y(n3234) );
  CLKBUFX2TS U1301 ( .A(n3236), .Y(n3233) );
  CLKBUFX2TS U1302 ( .A(n3237), .Y(n3232) );
  CLKBUFX2TS U1303 ( .A(n3237), .Y(n3231) );
  CLKBUFX2TS U1304 ( .A(n3239), .Y(n3228) );
  CLKBUFX2TS U1305 ( .A(n3433), .Y(n3429) );
  CLKBUFX2TS U1306 ( .A(n3434), .Y(n3427) );
  CLKBUFX2TS U1307 ( .A(n3435), .Y(n3425) );
  CLKBUFX2TS U1308 ( .A(n3435), .Y(n3424) );
  CLKBUFX2TS U1309 ( .A(n3436), .Y(n3422) );
  CLKBUFX2TS U1310 ( .A(n3238), .Y(n3230) );
  CLKBUFX2TS U1311 ( .A(n3238), .Y(n3229) );
  CLKBUFX2TS U1312 ( .A(n3239), .Y(n3227) );
  CLKBUFX2TS U1313 ( .A(n3433), .Y(n3428) );
  CLKBUFX2TS U1314 ( .A(n3434), .Y(n3426) );
  CLKBUFX2TS U1315 ( .A(n3436), .Y(n3423) );
  CLKBUFX2TS U1316 ( .A(n3406), .Y(n3391) );
  CLKBUFX2TS U1317 ( .A(n623), .Y(n584) );
  CLKBUFX2TS U1318 ( .A(n3714), .Y(n3703) );
  CLKBUFX2TS U1319 ( .A(n3715), .Y(n3714) );
  CLKBUFX2TS U1320 ( .A(n623), .Y(n585) );
  CLKBUFX2TS U1321 ( .A(n614), .Y(n607) );
  CLKBUFX2TS U1322 ( .A(n614), .Y(n594) );
  CLKBUFX2TS U1323 ( .A(n622), .Y(n587) );
  CLKBUFX2TS U1324 ( .A(n611), .Y(n609) );
  CLKBUFX2TS U1325 ( .A(n613), .Y(n608) );
  CLKBUFX2TS U1326 ( .A(n622), .Y(n586) );
  CLKBUFX2TS U1327 ( .A(n3323), .Y(n3316) );
  CLKBUFX2TS U1328 ( .A(n3498), .Y(n3495) );
  CLKBUFX2TS U1329 ( .A(n3499), .Y(n3494) );
  CLKBUFX2TS U1330 ( .A(n3499), .Y(n3493) );
  CLKBUFX2TS U1331 ( .A(n3501), .Y(n3492) );
  CLKBUFX2TS U1332 ( .A(n3501), .Y(n3491) );
  CLKBUFX2TS U1333 ( .A(n3502), .Y(n3490) );
  CLKBUFX2TS U1334 ( .A(n3502), .Y(n3489) );
  CLKBUFX2TS U1335 ( .A(n3503), .Y(n3488) );
  CLKBUFX2TS U1336 ( .A(n3503), .Y(n3487) );
  CLKBUFX2TS U1337 ( .A(n3471), .Y(n3456) );
  CLKBUFX2TS U1338 ( .A(n3471), .Y(n3457) );
  CLKBUFX2TS U1339 ( .A(n735), .Y(n705) );
  CLKBUFX2TS U1340 ( .A(n3339), .Y(n3325) );
  CLKBUFX2TS U1341 ( .A(n3339), .Y(n3326) );
  CLKBUFX2TS U1342 ( .A(n734), .Y(n706) );
  CLKBUFX2TS U1343 ( .A(n734), .Y(n707) );
  CLKBUFX2TS U1344 ( .A(n3470), .Y(n3458) );
  CLKBUFX2TS U1345 ( .A(n3402), .Y(n3400) );
  CLKBUFX2TS U1346 ( .A(n3403), .Y(n3398) );
  CLKBUFX2TS U1347 ( .A(n3404), .Y(n3396) );
  CLKBUFX2TS U1348 ( .A(n3404), .Y(n3395) );
  CLKBUFX2TS U1349 ( .A(n3405), .Y(n3393) );
  CLKBUFX2TS U1350 ( .A(n3467), .Y(n3464) );
  CLKBUFX2TS U1351 ( .A(n3468), .Y(n3462) );
  CLKBUFX2TS U1352 ( .A(n3469), .Y(n3461) );
  CLKBUFX2TS U1353 ( .A(n3469), .Y(n3460) );
  CLKBUFX2TS U1354 ( .A(n3470), .Y(n3459) );
  CLKBUFX2TS U1355 ( .A(n3468), .Y(n3463) );
  CLKBUFX2TS U1356 ( .A(n3402), .Y(n3399) );
  CLKBUFX2TS U1357 ( .A(n3403), .Y(n3397) );
  CLKBUFX2TS U1358 ( .A(n3405), .Y(n3394) );
  CLKBUFX2TS U1359 ( .A(n3498), .Y(n3496) );
  CLKBUFX2TS U1360 ( .A(n3258), .Y(n3251) );
  CLKBUFX2TS U1361 ( .A(n768), .Y(n762) );
  CLKBUFX2TS U1362 ( .A(n731), .Y(n716) );
  CLKBUFX2TS U1363 ( .A(n731), .Y(n715) );
  CLKBUFX2TS U1364 ( .A(n737), .Y(n714) );
  CLKBUFX2TS U1365 ( .A(n6124), .Y(n712) );
  CLKBUFX2TS U1366 ( .A(n733), .Y(n711) );
  CLKBUFX2TS U1367 ( .A(n3334), .Y(n3332) );
  CLKBUFX2TS U1368 ( .A(n3334), .Y(n3331) );
  CLKBUFX2TS U1369 ( .A(n3335), .Y(n3330) );
  CLKBUFX2TS U1370 ( .A(n3337), .Y(n3329) );
  CLKBUFX2TS U1371 ( .A(n3337), .Y(n3328) );
  CLKBUFX2TS U1372 ( .A(n733), .Y(n708) );
  CLKBUFX2TS U1373 ( .A(n3758), .Y(n3746) );
  CLKBUFX2TS U1374 ( .A(n3759), .Y(n3758) );
  INVX2TS U1375 ( .A(n1797), .Y(n871) );
  INVX2TS U1376 ( .A(n1817), .Y(n886) );
  INVX2TS U1377 ( .A(n1797), .Y(n970) );
  CLKBUFX2TS U1378 ( .A(n1822), .Y(n1797) );
  INVX2TS U1379 ( .A(n1817), .Y(n959) );
  CLKBUFX2TS U1380 ( .A(n424), .Y(n1817) );
  INVX2TS U1381 ( .A(n1817), .Y(n957) );
  INVX2TS U1382 ( .A(n1817), .Y(n955) );
  INVX2TS U1383 ( .A(n1797), .Y(n919) );
  INVX2TS U1384 ( .A(n1797), .Y(n936) );
  INVX2TS U1385 ( .A(n855), .Y(n844) );
  INVX2TS U1386 ( .A(n854), .Y(n840) );
  CLKBUFX2TS U1387 ( .A(n856), .Y(n854) );
  INVX2TS U1388 ( .A(n854), .Y(n842) );
  INVX2TS U1389 ( .A(n854), .Y(n846) );
  INVX2TS U1390 ( .A(n855), .Y(n841) );
  INVX2TS U1391 ( .A(n423), .Y(n843) );
  INVX2TS U1392 ( .A(n855), .Y(n845) );
  INVX2TS U1393 ( .A(n855), .Y(n847) );
  CLKBUFX2TS U1394 ( .A(n6123), .Y(n698) );
  CLKBUFX2TS U1395 ( .A(n703), .Y(n700) );
  CLKBUFX2TS U1396 ( .A(n6123), .Y(n699) );
  CLKBUFX2TS U1397 ( .A(n703), .Y(n701) );
  CLKBUFX2TS U1398 ( .A(n703), .Y(n702) );
  CLKBUFX2TS U1399 ( .A(n3772), .Y(n3761) );
  CLKBUFX2TS U1400 ( .A(n3773), .Y(n3772) );
  INVX2TS U1401 ( .A(n3223), .Y(n3209) );
  INVX2TS U1402 ( .A(n3224), .Y(n3208) );
  INVX2TS U1403 ( .A(n3219), .Y(n3210) );
  INVX2TS U1404 ( .A(n3219), .Y(n3211) );
  INVX2TS U1405 ( .A(n3220), .Y(n3212) );
  INVX2TS U1406 ( .A(n3221), .Y(n3213) );
  INVX2TS U1407 ( .A(n3221), .Y(n3214) );
  INVX2TS U1408 ( .A(n3222), .Y(n3216) );
  INVX2TS U1409 ( .A(n3222), .Y(n3215) );
  INVX2TS U1410 ( .A(n3220), .Y(n3218) );
  INVX2TS U1411 ( .A(n581), .Y(n575) );
  INVX2TS U1412 ( .A(n581), .Y(n574) );
  INVX2TS U1413 ( .A(n577), .Y(n570) );
  INVX2TS U1414 ( .A(n577), .Y(n569) );
  INVX2TS U1415 ( .A(n578), .Y(n572) );
  INVX2TS U1416 ( .A(n582), .Y(n573) );
  INVX2TS U1417 ( .A(n578), .Y(n571) );
  INVX2TS U1418 ( .A(n577), .Y(n568) );
  INVX2TS U1419 ( .A(n3304), .Y(n3300) );
  INVX2TS U1420 ( .A(n788), .Y(n781) );
  INVX2TS U1421 ( .A(n787), .Y(n780) );
  INVX2TS U1422 ( .A(n786), .Y(n779) );
  INVX2TS U1423 ( .A(n3304), .Y(n3299) );
  INVX2TS U1424 ( .A(n3388), .Y(n3383) );
  INVX2TS U1425 ( .A(n3389), .Y(n3382) );
  INVX2TS U1426 ( .A(n3390), .Y(n3381) );
  INVX2TS U1427 ( .A(n3521), .Y(n3514) );
  INVX2TS U1428 ( .A(n3520), .Y(n3513) );
  INVX2TS U1429 ( .A(n3519), .Y(n3512) );
  INVX2TS U1430 ( .A(n3304), .Y(n3298) );
  INVX2TS U1431 ( .A(n786), .Y(n772) );
  INVX2TS U1432 ( .A(n3388), .Y(n3375) );
  INVX2TS U1433 ( .A(n3519), .Y(n3506) );
  INVX2TS U1434 ( .A(n3307), .Y(n3292) );
  INVX2TS U1435 ( .A(n786), .Y(n773) );
  INVX2TS U1436 ( .A(n3388), .Y(n3376) );
  INVX2TS U1437 ( .A(n3519), .Y(n3507) );
  INVX2TS U1438 ( .A(n426), .Y(n3293) );
  INVX2TS U1439 ( .A(n785), .Y(n776) );
  INVX2TS U1440 ( .A(n785), .Y(n777) );
  INVX2TS U1441 ( .A(n785), .Y(n775) );
  INVX2TS U1442 ( .A(n3305), .Y(n3296) );
  INVX2TS U1443 ( .A(n3305), .Y(n3295) );
  INVX2TS U1444 ( .A(n3387), .Y(n3379) );
  INVX2TS U1445 ( .A(n3387), .Y(n3380) );
  INVX2TS U1446 ( .A(n3387), .Y(n3378) );
  INVX2TS U1447 ( .A(n3388), .Y(n3377) );
  INVX2TS U1448 ( .A(n3518), .Y(n3510) );
  INVX2TS U1449 ( .A(n3518), .Y(n3511) );
  INVX2TS U1450 ( .A(n3518), .Y(n3509) );
  INVX2TS U1451 ( .A(n3519), .Y(n3508) );
  INVX2TS U1452 ( .A(n786), .Y(n774) );
  INVX2TS U1453 ( .A(n3305), .Y(n3297) );
  INVX2TS U1454 ( .A(n426), .Y(n3294) );
  INVX2TS U1455 ( .A(n3223), .Y(n3217) );
  INVX2TS U1456 ( .A(n578), .Y(n576) );
  INVX2TS U1457 ( .A(n787), .Y(n770) );
  INVX2TS U1458 ( .A(n3389), .Y(n3373) );
  INVX2TS U1459 ( .A(n3306), .Y(n3290) );
  INVX2TS U1460 ( .A(n3520), .Y(n3504) );
  INVX2TS U1461 ( .A(n787), .Y(n771) );
  INVX2TS U1462 ( .A(n3306), .Y(n3291) );
  INVX2TS U1463 ( .A(n3389), .Y(n3374) );
  INVX2TS U1464 ( .A(n3520), .Y(n3505) );
  CLKBUFX2TS U1465 ( .A(n670), .Y(n668) );
  CLKBUFX2TS U1466 ( .A(n670), .Y(n667) );
  CLKBUFX2TS U1467 ( .A(n670), .Y(n666) );
  CLKBUFX2TS U1468 ( .A(n868), .Y(n857) );
  CLKBUFX2TS U1469 ( .A(n867), .Y(n859) );
  CLKBUFX2TS U1470 ( .A(n818), .Y(n806) );
  CLKBUFX2TS U1471 ( .A(n868), .Y(n858) );
  CLKBUFX2TS U1472 ( .A(n817), .Y(n807) );
  CLKBUFX2TS U1473 ( .A(n816), .Y(n809) );
  CLKBUFX2TS U1474 ( .A(n815), .Y(n811) );
  CLKBUFX2TS U1475 ( .A(n866), .Y(n862) );
  CLKBUFX2TS U1476 ( .A(n867), .Y(n860) );
  CLKBUFX2TS U1477 ( .A(n817), .Y(n808) );
  CLKBUFX2TS U1478 ( .A(n816), .Y(n810) );
  CLKBUFX2TS U1479 ( .A(n814), .Y(n812) );
  CLKBUFX2TS U1480 ( .A(n814), .Y(n813) );
  CLKBUFX2TS U1481 ( .A(n866), .Y(n861) );
  CLKBUFX2TS U1482 ( .A(n669), .Y(n626) );
  CLKBUFX2TS U1483 ( .A(n6109), .Y(n669) );
  CLKBUFX2TS U1484 ( .A(n3418), .Y(n3409) );
  CLKBUFX2TS U1485 ( .A(n749), .Y(n739) );
  CLKBUFX2TS U1486 ( .A(n748), .Y(n741) );
  CLKBUFX2TS U1487 ( .A(n749), .Y(n740) );
  CLKBUFX2TS U1488 ( .A(n747), .Y(n743) );
  CLKBUFX2TS U1489 ( .A(n3271), .Y(n3260) );
  CLKBUFX2TS U1490 ( .A(n3270), .Y(n3262) );
  CLKBUFX2TS U1491 ( .A(n3269), .Y(n3264) );
  CLKBUFX2TS U1492 ( .A(n3353), .Y(n3342) );
  CLKBUFX2TS U1493 ( .A(n3351), .Y(n3343) );
  CLKBUFX2TS U1494 ( .A(n3351), .Y(n3344) );
  CLKBUFX2TS U1495 ( .A(n3350), .Y(n3345) );
  CLKBUFX2TS U1496 ( .A(n3416), .Y(n3413) );
  CLKBUFX2TS U1497 ( .A(n3417), .Y(n3412) );
  CLKBUFX2TS U1498 ( .A(n3417), .Y(n3411) );
  CLKBUFX2TS U1499 ( .A(n3486), .Y(n3473) );
  CLKBUFX2TS U1500 ( .A(n3486), .Y(n3474) );
  CLKBUFX2TS U1501 ( .A(n3485), .Y(n3475) );
  CLKBUFX2TS U1502 ( .A(n3485), .Y(n3476) );
  CLKBUFX2TS U1503 ( .A(n3486), .Y(n3477) );
  CLKBUFX2TS U1504 ( .A(n3486), .Y(n3478) );
  CLKBUFX2TS U1505 ( .A(n3484), .Y(n3479) );
  CLKBUFX2TS U1506 ( .A(n3484), .Y(n3480) );
  CLKBUFX2TS U1507 ( .A(n3483), .Y(n3481) );
  CLKBUFX2TS U1508 ( .A(n3483), .Y(n3482) );
  CLKBUFX2TS U1509 ( .A(n748), .Y(n742) );
  CLKBUFX2TS U1510 ( .A(n3272), .Y(n3261) );
  CLKBUFX2TS U1511 ( .A(n3270), .Y(n3263) );
  CLKBUFX2TS U1512 ( .A(n3421), .Y(n3415) );
  CLKBUFX2TS U1513 ( .A(n3416), .Y(n3414) );
  CLKBUFX2TS U1514 ( .A(n3418), .Y(n3410) );
  CLKBUFX2TS U1515 ( .A(n3268), .Y(n3267) );
  CLKBUFX2TS U1516 ( .A(n3269), .Y(n3265) );
  CLKBUFX2TS U1517 ( .A(n3268), .Y(n3266) );
  CLKBUFX2TS U1518 ( .A(n3349), .Y(n3348) );
  CLKBUFX2TS U1519 ( .A(n3350), .Y(n3346) );
  CLKBUFX2TS U1520 ( .A(n3349), .Y(n3347) );
  CLKBUFX2TS U1521 ( .A(n3548), .Y(n3536) );
  CLKBUFX2TS U1522 ( .A(n3545), .Y(n3544) );
  CLKBUFX2TS U1523 ( .A(n3545), .Y(n3543) );
  CLKBUFX2TS U1524 ( .A(n3545), .Y(n3542) );
  CLKBUFX2TS U1525 ( .A(n3546), .Y(n3541) );
  CLKBUFX2TS U1526 ( .A(n3546), .Y(n3540) );
  CLKBUFX2TS U1527 ( .A(n3547), .Y(n3539) );
  CLKBUFX2TS U1528 ( .A(n3548), .Y(n3537) );
  CLKBUFX2TS U1529 ( .A(n3547), .Y(n3538) );
  CLKBUFX2TS U1530 ( .A(n3533), .Y(n3522) );
  CLKBUFX2TS U1531 ( .A(n3531), .Y(n3523) );
  CLKBUFX2TS U1532 ( .A(n3531), .Y(n3524) );
  CLKBUFX2TS U1533 ( .A(n3530), .Y(n3525) );
  CLKBUFX2TS U1534 ( .A(n3529), .Y(n3528) );
  CLKBUFX2TS U1535 ( .A(n3530), .Y(n3526) );
  CLKBUFX2TS U1536 ( .A(n3529), .Y(n3527) );
  CLKBUFX2TS U1537 ( .A(n3642), .Y(n3630) );
  CLKBUFX2TS U1538 ( .A(n3609), .Y(n3607) );
  CLKBUFX2TS U1539 ( .A(n3642), .Y(n3631) );
  CLKBUFX2TS U1540 ( .A(n3614), .Y(n3606) );
  CLKBUFX2TS U1541 ( .A(n3614), .Y(n3605) );
  CLKBUFX2TS U1542 ( .A(n3643), .Y(n3632) );
  CLKBUFX2TS U1543 ( .A(n3641), .Y(n3633) );
  CLKBUFX2TS U1544 ( .A(n3610), .Y(n3603) );
  CLKBUFX2TS U1545 ( .A(n3641), .Y(n3634) );
  CLKBUFX2TS U1546 ( .A(n3611), .Y(n3602) );
  CLKBUFX2TS U1547 ( .A(n3640), .Y(n3635) );
  CLKBUFX2TS U1548 ( .A(n3612), .Y(n3599) );
  CLKBUFX2TS U1549 ( .A(n3611), .Y(n3601) );
  CLKBUFX2TS U1550 ( .A(n3612), .Y(n3600) );
  CLKBUFX2TS U1551 ( .A(n3610), .Y(n3604) );
  CLKBUFX2TS U1552 ( .A(n3640), .Y(n3636) );
  CLKBUFX2TS U1553 ( .A(n3639), .Y(n3637) );
  CLKBUFX2TS U1554 ( .A(n3639), .Y(n3638) );
  CLKBUFX2TS U1555 ( .A(n419), .Y(n3223) );
  CLKBUFX2TS U1556 ( .A(n6139), .Y(n805) );
  CLKBUFX2TS U1557 ( .A(n6139), .Y(n804) );
  CLKBUFX2TS U1558 ( .A(n6171), .Y(n3288) );
  CLKBUFX2TS U1559 ( .A(n6200), .Y(n3405) );
  CLKBUFX2TS U1560 ( .A(n6200), .Y(n3406) );
  CLKBUFX2TS U1561 ( .A(n3407), .Y(n3404) );
  CLKBUFX2TS U1562 ( .A(n3472), .Y(n3471) );
  CLKBUFX2TS U1563 ( .A(n6217), .Y(n3466) );
  CLKBUFX2TS U1564 ( .A(n6217), .Y(n3467) );
  CLKBUFX2TS U1565 ( .A(n3472), .Y(n3469) );
  CLKBUFX2TS U1566 ( .A(n6217), .Y(n3468) );
  CLKBUFX2TS U1567 ( .A(n3407), .Y(n3402) );
  CLKBUFX2TS U1568 ( .A(n3407), .Y(n3403) );
  CLKBUFX2TS U1569 ( .A(n3472), .Y(n3470) );
  CLKBUFX2TS U1570 ( .A(n870), .Y(n863) );
  CLKBUFX2TS U1571 ( .A(n736), .Y(n735) );
  CLKBUFX2TS U1572 ( .A(n737), .Y(n731) );
  CLKBUFX2TS U1573 ( .A(n737), .Y(n732) );
  CLKBUFX2TS U1574 ( .A(n736), .Y(n734) );
  CLKBUFX2TS U1575 ( .A(n6168), .Y(n3237) );
  CLKBUFX2TS U1576 ( .A(n3241), .Y(n3240) );
  CLKBUFX2TS U1577 ( .A(n3340), .Y(n3339) );
  CLKBUFX2TS U1578 ( .A(n3341), .Y(n3334) );
  CLKBUFX2TS U1579 ( .A(n3341), .Y(n3335) );
  CLKBUFX2TS U1580 ( .A(n3341), .Y(n3336) );
  CLKBUFX2TS U1581 ( .A(n3340), .Y(n3337) );
  CLKBUFX2TS U1582 ( .A(n3340), .Y(n3338) );
  CLKBUFX2TS U1583 ( .A(n3437), .Y(n3435) );
  CLKBUFX2TS U1584 ( .A(n6219), .Y(n3499) );
  CLKBUFX2TS U1585 ( .A(n6219), .Y(n3501) );
  CLKBUFX2TS U1586 ( .A(n3499), .Y(n3502) );
  CLKBUFX2TS U1587 ( .A(n3498), .Y(n3503) );
  CLKBUFX2TS U1588 ( .A(n6219), .Y(n3500) );
  CLKBUFX2TS U1589 ( .A(n6168), .Y(n3236) );
  CLKBUFX2TS U1590 ( .A(n736), .Y(n733) );
  CLKBUFX2TS U1591 ( .A(n3241), .Y(n3238) );
  CLKBUFX2TS U1592 ( .A(n3241), .Y(n3239) );
  CLKBUFX2TS U1593 ( .A(n3438), .Y(n3433) );
  CLKBUFX2TS U1594 ( .A(n3437), .Y(n3434) );
  CLKBUFX2TS U1595 ( .A(n3437), .Y(n3436) );
  CLKBUFX2TS U1596 ( .A(n625), .Y(n611) );
  CLKBUFX2TS U1597 ( .A(n624), .Y(n614) );
  CLKBUFX2TS U1598 ( .A(n6155), .Y(n3207) );
  CLKBUFX2TS U1599 ( .A(n6169), .Y(n3258) );
  CLKBUFX2TS U1600 ( .A(n6123), .Y(n704) );
  CLKBUFX2TS U1601 ( .A(n625), .Y(n612) );
  CLKBUFX2TS U1602 ( .A(n625), .Y(n613) );
  CLKBUFX2TS U1603 ( .A(n624), .Y(n622) );
  CLKBUFX2TS U1604 ( .A(n624), .Y(n623) );
  CLKBUFX2TS U1605 ( .A(n6141), .Y(n839) );
  CLKBUFX2TS U1606 ( .A(n6141), .Y(n838) );
  CLKBUFX2TS U1607 ( .A(n6344), .Y(n3745) );
  CLKBUFX2TS U1608 ( .A(n158), .Y(n3775) );
  CLKBUFX2TS U1609 ( .A(n158), .Y(n3776) );
  CLKBUFX2TS U1610 ( .A(n6169), .Y(n3256) );
  CLKBUFX2TS U1611 ( .A(n6216), .Y(n3455) );
  CLKBUFX2TS U1612 ( .A(n6155), .Y(n3205) );
  CLKBUFX2TS U1613 ( .A(n6155), .Y(n3206) );
  CLKBUFX2TS U1614 ( .A(n6187), .Y(n3371) );
  CLKBUFX2TS U1615 ( .A(n6184), .Y(n3323) );
  CLKBUFX2TS U1616 ( .A(n6216), .Y(n3454) );
  CLKBUFX2TS U1617 ( .A(n6126), .Y(n768) );
  CLKBUFX2TS U1618 ( .A(n6169), .Y(n3257) );
  CLKBUFX2TS U1619 ( .A(n6110), .Y(n687) );
  CLKBUFX2TS U1620 ( .A(n6110), .Y(n686) );
  CLKBUFX2TS U1621 ( .A(n268), .Y(n3760) );
  CLKBUFX2TS U1622 ( .A(n268), .Y(n3759) );
  CLKBUFX2TS U1623 ( .A(n262), .Y(n3774) );
  CLKBUFX2TS U1624 ( .A(n6342), .Y(n3716) );
  CLKBUFX2TS U1625 ( .A(n6342), .Y(n3715) );
  CLKBUFX2TS U1626 ( .A(n262), .Y(n3773) );
  INVX2TS U1627 ( .A(n416), .Y(n6346) );
  CLKBUFX2TS U1628 ( .A(n6171), .Y(n3289) );
  INVX2TS U1629 ( .A(n5585), .Y(n6339) );
  INVX2TS U1630 ( .A(n5583), .Y(n6341) );
  CLKBUFX2TS U1631 ( .A(n423), .Y(n855) );
  CLKBUFX2TS U1632 ( .A(n423), .Y(n856) );
  CLKBUFX2TS U1633 ( .A(n424), .Y(n1822) );
  CLKBUFX2TS U1634 ( .A(n3438), .Y(n3431) );
  CLKBUFX2TS U1635 ( .A(n733), .Y(n729) );
  CLKBUFX2TS U1636 ( .A(n3337), .Y(n3333) );
  CLKBUFX2TS U1637 ( .A(n3224), .Y(n3222) );
  CLKBUFX2TS U1638 ( .A(n3224), .Y(n3219) );
  CLKBUFX2TS U1639 ( .A(n3224), .Y(n3220) );
  CLKBUFX2TS U1640 ( .A(n419), .Y(n3221) );
  CLKBUFX2TS U1641 ( .A(n788), .Y(n787) );
  CLKBUFX2TS U1642 ( .A(n3390), .Y(n3389) );
  CLKBUFX2TS U1643 ( .A(n3307), .Y(n3306) );
  CLKBUFX2TS U1644 ( .A(n3521), .Y(n3520) );
  CLKBUFX2TS U1645 ( .A(n6123), .Y(n703) );
  INVX2TS U1646 ( .A(n5462), .Y(n6328) );
  CLKBUFX2TS U1647 ( .A(n581), .Y(n579) );
  INVX2TS U1648 ( .A(n583), .Y(n565) );
  INVX2TS U1649 ( .A(n583), .Y(n566) );
  INVX2TS U1650 ( .A(n583), .Y(n567) );
  INVX2TS U1651 ( .A(n3306), .Y(n3302) );
  INVX2TS U1652 ( .A(n785), .Y(n783) );
  INVX2TS U1653 ( .A(n429), .Y(n782) );
  INVX2TS U1654 ( .A(n3306), .Y(n3301) );
  INVX2TS U1655 ( .A(n425), .Y(n3385) );
  INVX2TS U1656 ( .A(n425), .Y(n3384) );
  CLKBUFX2TS U1657 ( .A(n819), .Y(n815) );
  CLKBUFX2TS U1658 ( .A(n751), .Y(n749) );
  CLKBUFX2TS U1659 ( .A(n752), .Y(n747) );
  CLKBUFX2TS U1660 ( .A(n752), .Y(n746) );
  CLKBUFX2TS U1661 ( .A(n752), .Y(n745) );
  CLKBUFX2TS U1662 ( .A(n869), .Y(n868) );
  CLKBUFX2TS U1663 ( .A(n870), .Y(n864) );
  CLKBUFX2TS U1664 ( .A(n870), .Y(n865) );
  CLKBUFX2TS U1665 ( .A(n869), .Y(n867) );
  CLKBUFX2TS U1666 ( .A(n3272), .Y(n3269) );
  CLKBUFX2TS U1667 ( .A(n3272), .Y(n3268) );
  CLKBUFX2TS U1668 ( .A(n3354), .Y(n3353) );
  CLKBUFX2TS U1669 ( .A(n3355), .Y(n3351) );
  CLKBUFX2TS U1670 ( .A(n3354), .Y(n3352) );
  CLKBUFX2TS U1671 ( .A(n3355), .Y(n3350) );
  CLKBUFX2TS U1672 ( .A(n3355), .Y(n3349) );
  CLKBUFX2TS U1673 ( .A(n3420), .Y(n3417) );
  CLKBUFX2TS U1674 ( .A(n6218), .Y(n3486) );
  CLKBUFX2TS U1675 ( .A(n6218), .Y(n3485) );
  CLKBUFX2TS U1676 ( .A(n6218), .Y(n3484) );
  CLKBUFX2TS U1677 ( .A(n6218), .Y(n3483) );
  CLKBUFX2TS U1678 ( .A(n751), .Y(n748) );
  CLKBUFX2TS U1679 ( .A(n6140), .Y(n817) );
  CLKBUFX2TS U1680 ( .A(n819), .Y(n816) );
  CLKBUFX2TS U1681 ( .A(n819), .Y(n814) );
  CLKBUFX2TS U1682 ( .A(n869), .Y(n866) );
  CLKBUFX2TS U1683 ( .A(n3272), .Y(n3270) );
  CLKBUFX2TS U1684 ( .A(n3421), .Y(n3416) );
  CLKBUFX2TS U1685 ( .A(n3420), .Y(n3418) );
  CLKBUFX2TS U1686 ( .A(n6109), .Y(n670) );
  CLKBUFX2TS U1687 ( .A(n3419), .Y(n3408) );
  CLKBUFX2TS U1688 ( .A(n3420), .Y(n3419) );
  INVX2TS U1689 ( .A(n559), .Y(n541) );
  INVX2TS U1690 ( .A(n559), .Y(n543) );
  INVX2TS U1691 ( .A(n563), .Y(n557) );
  INVX2TS U1692 ( .A(n563), .Y(n556) );
  INVX2TS U1693 ( .A(n558), .Y(n555) );
  INVX2TS U1694 ( .A(n558), .Y(n554) );
  INVX2TS U1695 ( .A(n558), .Y(n551) );
  INVX2TS U1696 ( .A(n558), .Y(n546) );
  INVX2TS U1697 ( .A(n564), .Y(n545) );
  INVX2TS U1698 ( .A(n559), .Y(n548) );
  INVX2TS U1699 ( .A(n559), .Y(n544) );
  CLKBUFX2TS U1700 ( .A(n750), .Y(n738) );
  CLKBUFX2TS U1701 ( .A(n751), .Y(n750) );
  CLKBUFX2TS U1702 ( .A(n6140), .Y(n818) );
  CLKBUFX2TS U1703 ( .A(n3271), .Y(n3259) );
  CLKBUFX2TS U1704 ( .A(n6170), .Y(n3271) );
  CLKBUFX2TS U1705 ( .A(n492), .Y(n480) );
  CLKBUFX2TS U1706 ( .A(n490), .Y(n488) );
  CLKBUFX2TS U1707 ( .A(n489), .Y(n487) );
  CLKBUFX2TS U1708 ( .A(n489), .Y(n486) );
  CLKBUFX2TS U1709 ( .A(n490), .Y(n485) );
  CLKBUFX2TS U1710 ( .A(n490), .Y(n484) );
  CLKBUFX2TS U1711 ( .A(n492), .Y(n481) );
  CLKBUFX2TS U1712 ( .A(n491), .Y(n483) );
  CLKBUFX2TS U1713 ( .A(n491), .Y(n482) );
  INVX2TS U1714 ( .A(n458), .Y(n457) );
  INVX2TS U1715 ( .A(n459), .Y(n456) );
  INVX2TS U1716 ( .A(n460), .Y(n455) );
  CLKBUFX2TS U1717 ( .A(n3550), .Y(n3545) );
  CLKBUFX2TS U1718 ( .A(n3549), .Y(n3546) );
  CLKBUFX2TS U1719 ( .A(n3549), .Y(n3548) );
  CLKBUFX2TS U1720 ( .A(n3549), .Y(n3547) );
  CLKBUFX2TS U1721 ( .A(n3534), .Y(n3533) );
  CLKBUFX2TS U1722 ( .A(n3534), .Y(n3532) );
  CLKBUFX2TS U1723 ( .A(n3535), .Y(n3531) );
  CLKBUFX2TS U1724 ( .A(n3535), .Y(n3530) );
  CLKBUFX2TS U1725 ( .A(n3535), .Y(n3529) );
  CLKBUFX2TS U1726 ( .A(n444), .Y(n433) );
  CLKBUFX2TS U1727 ( .A(n442), .Y(n434) );
  CLKBUFX2TS U1728 ( .A(n442), .Y(n435) );
  CLKBUFX2TS U1729 ( .A(n441), .Y(n436) );
  CLKBUFX2TS U1730 ( .A(n440), .Y(n439) );
  CLKBUFX2TS U1731 ( .A(n441), .Y(n437) );
  CLKBUFX2TS U1732 ( .A(n440), .Y(n438) );
  CLKBUFX2TS U1733 ( .A(n477), .Y(n463) );
  CLKBUFX2TS U1734 ( .A(n475), .Y(n464) );
  CLKBUFX2TS U1735 ( .A(n475), .Y(n465) );
  CLKBUFX2TS U1736 ( .A(n474), .Y(n466) );
  CLKBUFX2TS U1737 ( .A(n474), .Y(n467) );
  CLKBUFX2TS U1738 ( .A(n473), .Y(n468) );
  CLKBUFX2TS U1739 ( .A(n472), .Y(n471) );
  CLKBUFX2TS U1740 ( .A(n473), .Y(n469) );
  CLKBUFX2TS U1741 ( .A(n472), .Y(n470) );
  INVX2TS U1742 ( .A(reset), .Y(n4422) );
  CLKBUFX2TS U1743 ( .A(n3580), .Y(n3568) );
  CLKBUFX2TS U1744 ( .A(n3624), .Y(n3621) );
  CLKBUFX2TS U1745 ( .A(n3580), .Y(n3569) );
  CLKBUFX2TS U1746 ( .A(n3658), .Y(n3645) );
  CLKBUFX2TS U1747 ( .A(n3657), .Y(n3646) );
  CLKBUFX2TS U1748 ( .A(n3625), .Y(n3620) );
  CLKBUFX2TS U1749 ( .A(n3625), .Y(n3619) );
  CLKBUFX2TS U1750 ( .A(n3657), .Y(n3647) );
  CLKBUFX2TS U1751 ( .A(n3581), .Y(n3570) );
  CLKBUFX2TS U1752 ( .A(n3626), .Y(n3618) );
  CLKBUFX2TS U1753 ( .A(n3656), .Y(n3648) );
  CLKBUFX2TS U1754 ( .A(n3579), .Y(n3571) );
  CLKBUFX2TS U1755 ( .A(n3626), .Y(n3617) );
  CLKBUFX2TS U1756 ( .A(n3656), .Y(n3649) );
  CLKBUFX2TS U1757 ( .A(n3579), .Y(n3572) );
  CLKBUFX2TS U1758 ( .A(n3627), .Y(n3616) );
  CLKBUFX2TS U1759 ( .A(n3655), .Y(n3650) );
  CLKBUFX2TS U1760 ( .A(n3578), .Y(n3573) );
  CLKBUFX2TS U1761 ( .A(n3627), .Y(n3615) );
  CLKBUFX2TS U1762 ( .A(n3566), .Y(n3551) );
  CLKBUFX2TS U1763 ( .A(n3566), .Y(n3552) );
  CLKBUFX2TS U1764 ( .A(n3594), .Y(n3584) );
  CLKBUFX2TS U1765 ( .A(n3562), .Y(n3558) );
  CLKBUFX2TS U1766 ( .A(n3563), .Y(n3557) );
  CLKBUFX2TS U1767 ( .A(n3592), .Y(n3588) );
  CLKBUFX2TS U1768 ( .A(n3564), .Y(n3556) );
  CLKBUFX2TS U1769 ( .A(n3592), .Y(n3587) );
  CLKBUFX2TS U1770 ( .A(n3564), .Y(n3555) );
  CLKBUFX2TS U1771 ( .A(n3593), .Y(n3586) );
  CLKBUFX2TS U1772 ( .A(n3565), .Y(n3554) );
  CLKBUFX2TS U1773 ( .A(n3593), .Y(n3585) );
  CLKBUFX2TS U1774 ( .A(n3565), .Y(n3553) );
  CLKBUFX2TS U1775 ( .A(n3578), .Y(n3574) );
  CLKBUFX2TS U1776 ( .A(n3655), .Y(n3651) );
  CLKBUFX2TS U1777 ( .A(n3577), .Y(n3576) );
  CLKBUFX2TS U1778 ( .A(n3614), .Y(n3609) );
  CLKBUFX2TS U1779 ( .A(n3643), .Y(n3642) );
  CLKBUFX2TS U1780 ( .A(n3644), .Y(n3641) );
  CLKBUFX2TS U1781 ( .A(n3644), .Y(n3640) );
  CLKBUFX2TS U1782 ( .A(n3613), .Y(n3611) );
  CLKBUFX2TS U1783 ( .A(n3613), .Y(n3612) );
  CLKBUFX2TS U1784 ( .A(n3613), .Y(n3610) );
  CLKBUFX2TS U1785 ( .A(n3644), .Y(n3639) );
  CLKBUFX2TS U1786 ( .A(n3562), .Y(n3559) );
  CLKBUFX2TS U1787 ( .A(n6316), .Y(n3608) );
  CLKBUFX2TS U1788 ( .A(n3577), .Y(n3575) );
  CLKBUFX2TS U1789 ( .A(n3624), .Y(n3622) );
  CLKBUFX2TS U1790 ( .A(n3654), .Y(n3652) );
  CLKBUFX2TS U1791 ( .A(n3626), .Y(n3623) );
  CLKBUFX2TS U1792 ( .A(n3654), .Y(n3653) );
  NAND2X1TS U1793 ( .A(n5542), .B(n5545), .Y(n5579) );
  NOR2X1TS U1794 ( .A(n5535), .B(n5531), .Y(n6155) );
  AND3X2TS U1795 ( .A(n172), .B(n5548), .C(n5552), .Y(n6187) );
  CLKBUFX2TS U1796 ( .A(n427), .Y(n583) );
  INVX2TS U1797 ( .A(n5574), .Y(n6344) );
  AND2X2TS U1798 ( .A(n5552), .B(n6333), .Y(n6184) );
  AND2X2TS U1799 ( .A(n5545), .B(n6337), .Y(n6169) );
  INVX2TS U1800 ( .A(n5535), .Y(n6334) );
  CLKBUFX2TS U1801 ( .A(n6168), .Y(n3241) );
  CLKBUFX2TS U1802 ( .A(n6124), .Y(n737) );
  CLKBUFX2TS U1803 ( .A(n6185), .Y(n3341) );
  CLKBUFX2TS U1804 ( .A(n6185), .Y(n3340) );
  CLKBUFX2TS U1805 ( .A(n6124), .Y(n736) );
  CLKBUFX2TS U1806 ( .A(n6200), .Y(n3407) );
  CLKBUFX2TS U1807 ( .A(n6217), .Y(n3472) );
  CLKBUFX2TS U1808 ( .A(n6202), .Y(n3438) );
  CLKBUFX2TS U1809 ( .A(n6202), .Y(n3437) );
  CLKBUFX2TS U1810 ( .A(n6154), .Y(n870) );
  INVX2TS U1811 ( .A(n5513), .Y(n6338) );
  INVX2TS U1812 ( .A(n5534), .Y(n6335) );
  CLKBUFX2TS U1813 ( .A(n6108), .Y(n624) );
  INVX2TS U1814 ( .A(n5536), .Y(n6329) );
  INVX2TS U1815 ( .A(n5581), .Y(n6342) );
  CLKBUFX2TS U1816 ( .A(n426), .Y(n3307) );
  CLKBUFX2TS U1817 ( .A(n427), .Y(n581) );
  CLKBUFX2TS U1818 ( .A(n427), .Y(n582) );
  CLKBUFX2TS U1819 ( .A(n425), .Y(n3390) );
  CLKBUFX2TS U1820 ( .A(n429), .Y(n788) );
  CLKBUFX2TS U1821 ( .A(n428), .Y(n3521) );
  CLKBUFX2TS U1822 ( .A(n419), .Y(n3224) );
  CLKBUFX2TS U1823 ( .A(n462), .Y(n458) );
  CLKBUFX2TS U1824 ( .A(n462), .Y(n459) );
  CLKBUFX2TS U1825 ( .A(n462), .Y(n460) );
  AND2X2TS U1826 ( .A(n5473), .B(n5356), .Y(n6109) );
  CLKBUFX2TS U1827 ( .A(n492), .Y(n489) );
  CLKBUFX2TS U1828 ( .A(n5282), .Y(n490) );
  CLKBUFX2TS U1829 ( .A(n494), .Y(n492) );
  CLKBUFX2TS U1830 ( .A(n494), .Y(n491) );
  CLKBUFX2TS U1831 ( .A(n6125), .Y(n752) );
  CLKBUFX2TS U1832 ( .A(n6186), .Y(n3354) );
  CLKBUFX2TS U1833 ( .A(n6186), .Y(n3355) );
  CLKBUFX2TS U1834 ( .A(n6125), .Y(n751) );
  CLKBUFX2TS U1835 ( .A(n6140), .Y(n819) );
  CLKBUFX2TS U1836 ( .A(n6154), .Y(n869) );
  CLKBUFX2TS U1837 ( .A(n6170), .Y(n3272) );
  CLKBUFX2TS U1838 ( .A(n6201), .Y(n3421) );
  CLKBUFX2TS U1839 ( .A(n6201), .Y(n3420) );
  CLKBUFX2TS U1840 ( .A(n563), .Y(n561) );
  CLKBUFX2TS U1841 ( .A(n563), .Y(n562) );
  CLKBUFX2TS U1842 ( .A(n493), .Y(n479) );
  CLKBUFX2TS U1843 ( .A(n494), .Y(n493) );
  INVX2TS U1844 ( .A(n461), .Y(n447) );
  CLKBUFX2TS U1845 ( .A(n462), .Y(n461) );
  INVX2TS U1846 ( .A(n430), .Y(n448) );
  INVX2TS U1847 ( .A(n461), .Y(n449) );
  INVX2TS U1848 ( .A(n430), .Y(n450) );
  INVX2TS U1849 ( .A(n430), .Y(n451) );
  INVX2TS U1850 ( .A(n461), .Y(n452) );
  INVX2TS U1851 ( .A(n461), .Y(n453) );
  INVX2TS U1852 ( .A(n460), .Y(n454) );
  CLKBUFX2TS U1853 ( .A(n445), .Y(n444) );
  CLKBUFX2TS U1854 ( .A(n477), .Y(n475) );
  CLKBUFX2TS U1855 ( .A(n445), .Y(n443) );
  CLKBUFX2TS U1856 ( .A(n478), .Y(n474) );
  CLKBUFX2TS U1857 ( .A(n446), .Y(n442) );
  CLKBUFX2TS U1858 ( .A(n478), .Y(n473) );
  CLKBUFX2TS U1859 ( .A(n446), .Y(n441) );
  CLKBUFX2TS U1860 ( .A(n478), .Y(n472) );
  CLKBUFX2TS U1861 ( .A(n446), .Y(n440) );
  CLKBUFX2TS U1862 ( .A(n6254), .Y(n3550) );
  CLKBUFX2TS U1863 ( .A(n6254), .Y(n3549) );
  CLKBUFX2TS U1864 ( .A(n5283), .Y(n3534) );
  CLKBUFX2TS U1865 ( .A(n5283), .Y(n3535) );
  CLKBUFX2TS U1866 ( .A(n477), .Y(n476) );
  CLKBUFX2TS U1867 ( .A(n4266), .Y(n4267) );
  CLKBUFX2TS U1868 ( .A(n4269), .Y(n4270) );
  CLKBUFX2TS U1869 ( .A(n4266), .Y(n4268) );
  CLKBUFX2TS U1870 ( .A(n4269), .Y(n4271) );
  INVX2TS U1871 ( .A(n3815), .Y(n3812) );
  CLKBUFX2TS U1872 ( .A(n3567), .Y(n3562) );
  CLKBUFX2TS U1873 ( .A(n3629), .Y(n3624) );
  CLKBUFX2TS U1874 ( .A(n3581), .Y(n3580) );
  CLKBUFX2TS U1875 ( .A(n6314), .Y(n3563) );
  CLKBUFX2TS U1876 ( .A(n3628), .Y(n3625) );
  CLKBUFX2TS U1877 ( .A(n3658), .Y(n3657) );
  CLKBUFX2TS U1878 ( .A(n3597), .Y(n3592) );
  CLKBUFX2TS U1879 ( .A(n3563), .Y(n3564) );
  CLKBUFX2TS U1880 ( .A(n3628), .Y(n3626) );
  CLKBUFX2TS U1881 ( .A(n3659), .Y(n3656) );
  CLKBUFX2TS U1882 ( .A(n3582), .Y(n3579) );
  CLKBUFX2TS U1883 ( .A(n3596), .Y(n3593) );
  CLKBUFX2TS U1884 ( .A(n3659), .Y(n3655) );
  CLKBUFX2TS U1885 ( .A(n3582), .Y(n3578) );
  CLKBUFX2TS U1886 ( .A(n6314), .Y(n3565) );
  CLKBUFX2TS U1887 ( .A(n3628), .Y(n3627) );
  CLKBUFX2TS U1888 ( .A(n3596), .Y(n3594) );
  CLKBUFX2TS U1889 ( .A(n3563), .Y(n3566) );
  CLKBUFX2TS U1890 ( .A(n3582), .Y(n3577) );
  CLKBUFX2TS U1891 ( .A(n516), .Y(n507) );
  CLKBUFX2TS U1892 ( .A(n514), .Y(n505) );
  CLKBUFX2TS U1893 ( .A(n514), .Y(n503) );
  CLKBUFX2TS U1894 ( .A(n516), .Y(n502) );
  CLKBUFX2TS U1895 ( .A(n517), .Y(n501) );
  CLKBUFX2TS U1896 ( .A(n517), .Y(n500) );
  CLKBUFX2TS U1897 ( .A(n526), .Y(n499) );
  CLKBUFX2TS U1898 ( .A(n526), .Y(n496) );
  CLKBUFX2TS U1899 ( .A(n3595), .Y(n3583) );
  CLKBUFX2TS U1900 ( .A(n3596), .Y(n3595) );
  INVX2TS U1901 ( .A(n5356), .Y(n6318) );
  CLKBUFX2TS U1902 ( .A(n3659), .Y(n3654) );
  CLKBUFX2TS U1903 ( .A(n6317), .Y(n3643) );
  CLKBUFX2TS U1904 ( .A(n6317), .Y(n3644) );
  CLKBUFX2TS U1905 ( .A(n6316), .Y(n3614) );
  CLKBUFX2TS U1906 ( .A(n6316), .Y(n3613) );
  CLKBUFX2TS U1907 ( .A(n3591), .Y(n3589) );
  CLKBUFX2TS U1908 ( .A(n3591), .Y(n3590) );
  CLKBUFX2TS U1909 ( .A(n3561), .Y(n3560) );
  AOI21X1TS U1910 ( .A0(n152), .A1(n6325), .B0(n6335), .Y(n5394) );
  OAI21X1TS U1911 ( .A0(n6326), .A1(n149), .B0(n5518), .Y(n5369) );
  NOR2X1TS U1912 ( .A(n5562), .B(n5563), .Y(n5560) );
  NOR2X1TS U1913 ( .A(n150), .B(n5390), .Y(n5536) );
  OAI2BB1X1TS U1914 ( .A0N(n159), .A1N(n5320), .B0(n5319), .Y(n5321) );
  AOI2BB1X1TS U1915 ( .A0N(n6323), .A1N(n5416), .B0(n5540), .Y(n5542) );
  NOR2X1TS U1916 ( .A(n5395), .B(n418), .Y(n6154) );
  OR2X2TS U1917 ( .A(n4862), .B(n4861), .Y(n4863) );
  INVX2TS U1918 ( .A(n170), .Y(n6327) );
  INVX2TS U1919 ( .A(n5561), .Y(n6324) );
  XNOR2X1TS U1920 ( .A(n6313), .B(n6234), .Y(n4860) );
  NAND2X1TS U1921 ( .A(n152), .B(n5489), .Y(n5395) );
  INVX2TS U1922 ( .A(n160), .Y(n6251) );
  NOR2BX1TS U1923 ( .AN(n5464), .B(n418), .Y(n5473) );
  AND2X2TS U1924 ( .A(n5473), .B(n152), .Y(n6140) );
  AND2X2TS U1925 ( .A(n5499), .B(n202), .Y(n6218) );
  AND2X2TS U1926 ( .A(n5499), .B(n200), .Y(n6125) );
  AND2X2TS U1927 ( .A(n5473), .B(n5498), .Y(n6201) );
  AND2X2TS U1928 ( .A(n5499), .B(n154), .Y(n6186) );
  AND2X2TS U1929 ( .A(n5473), .B(n5449), .Y(n6170) );
  CLKBUFX2TS U1930 ( .A(n564), .Y(n563) );
  CLKBUFX2TS U1931 ( .A(n5282), .Y(n494) );
  CLKBUFX2TS U1932 ( .A(n430), .Y(n462) );
  NAND2X1TS U1933 ( .A(n187), .B(n4422), .Y(n6232) );
  CLKBUFX2TS U1934 ( .A(destinationAddressIn_SOUTH[6]), .Y(n4266) );
  CLKBUFX2TS U1935 ( .A(destinationAddressIn_SOUTH[7]), .Y(n4269) );
  CLKBUFX2TS U1936 ( .A(n5281), .Y(n477) );
  CLKBUFX2TS U1937 ( .A(n5281), .Y(n478) );
  CLKBUFX2TS U1938 ( .A(n5218), .Y(n445) );
  CLKBUFX2TS U1939 ( .A(n5218), .Y(n446) );
  CLKBUFX2TS U1940 ( .A(n4293), .Y(n4294) );
  CLKBUFX2TS U1941 ( .A(n4404), .Y(n4405) );
  CLKBUFX2TS U1942 ( .A(n4377), .Y(n4378) );
  CLKBUFX2TS U1943 ( .A(n4359), .Y(n4360) );
  CLKBUFX2TS U1944 ( .A(n4353), .Y(n4354) );
  CLKBUFX2TS U1945 ( .A(n4350), .Y(n4351) );
  CLKBUFX2TS U1946 ( .A(n4329), .Y(n4330) );
  CLKBUFX2TS U1947 ( .A(n4326), .Y(n4327) );
  CLKBUFX2TS U1948 ( .A(n4320), .Y(n4321) );
  CLKBUFX2TS U1949 ( .A(n4308), .Y(n4309) );
  CLKBUFX2TS U1950 ( .A(n4383), .Y(n4384) );
  CLKBUFX2TS U1951 ( .A(n4380), .Y(n4381) );
  CLKBUFX2TS U1952 ( .A(n4374), .Y(n4375) );
  CLKBUFX2TS U1953 ( .A(n4371), .Y(n4372) );
  CLKBUFX2TS U1954 ( .A(n4368), .Y(n4369) );
  CLKBUFX2TS U1955 ( .A(n4362), .Y(n4363) );
  CLKBUFX2TS U1956 ( .A(n4356), .Y(n4357) );
  CLKBUFX2TS U1957 ( .A(n4347), .Y(n4348) );
  CLKBUFX2TS U1958 ( .A(n4338), .Y(n4339) );
  CLKBUFX2TS U1959 ( .A(n4323), .Y(n4324) );
  CLKBUFX2TS U1960 ( .A(n4317), .Y(n4318) );
  CLKBUFX2TS U1961 ( .A(n4314), .Y(n4315) );
  CLKBUFX2TS U1962 ( .A(n4311), .Y(n4312) );
  CLKBUFX2TS U1963 ( .A(n4305), .Y(n4306) );
  CLKBUFX2TS U1964 ( .A(n4296), .Y(n4297) );
  CLKBUFX2TS U1965 ( .A(n4419), .Y(n4420) );
  CLKBUFX2TS U1966 ( .A(n4413), .Y(n4414) );
  CLKBUFX2TS U1967 ( .A(n4410), .Y(n4411) );
  CLKBUFX2TS U1968 ( .A(n4407), .Y(n4408) );
  CLKBUFX2TS U1969 ( .A(n4290), .Y(n4291) );
  CLKBUFX2TS U1970 ( .A(n4341), .Y(n4342) );
  CLKBUFX2TS U1971 ( .A(n4335), .Y(n4336) );
  CLKBUFX2TS U1972 ( .A(n4332), .Y(n4333) );
  CLKBUFX2TS U1973 ( .A(n4299), .Y(n4300) );
  CLKBUFX2TS U1974 ( .A(n4416), .Y(n4417) );
  CLKBUFX2TS U1975 ( .A(n4365), .Y(n4366) );
  CLKBUFX2TS U1976 ( .A(n4344), .Y(n4345) );
  CLKBUFX2TS U1977 ( .A(n4302), .Y(n4303) );
  CLKBUFX2TS U1978 ( .A(n4401), .Y(n4402) );
  CLKBUFX2TS U1979 ( .A(n4398), .Y(n4399) );
  CLKBUFX2TS U1980 ( .A(n4392), .Y(n4393) );
  CLKBUFX2TS U1981 ( .A(n4395), .Y(n4396) );
  CLKBUFX2TS U1982 ( .A(n4389), .Y(n4390) );
  CLKBUFX2TS U1983 ( .A(n4386), .Y(n4387) );
  INVX2TS U1984 ( .A(n3917), .Y(n3915) );
  INVX2TS U1985 ( .A(n3914), .Y(n3912) );
  INVX2TS U1986 ( .A(n3911), .Y(n3909) );
  INVX2TS U1987 ( .A(n3908), .Y(n3906) );
  INVX2TS U1988 ( .A(n3905), .Y(n3903) );
  INVX2TS U1989 ( .A(n3902), .Y(n3900) );
  INVX2TS U1990 ( .A(n3899), .Y(n3897) );
  INVX2TS U1991 ( .A(n3896), .Y(n3894) );
  INVX2TS U1992 ( .A(n3893), .Y(n3891) );
  INVX2TS U1993 ( .A(n3890), .Y(n3888) );
  INVX2TS U1994 ( .A(n3887), .Y(n3885) );
  INVX2TS U1995 ( .A(n3884), .Y(n3882) );
  INVX2TS U1996 ( .A(n3881), .Y(n3879) );
  INVX2TS U1997 ( .A(n3878), .Y(n3876) );
  INVX2TS U1998 ( .A(n3875), .Y(n3873) );
  INVX2TS U1999 ( .A(n3872), .Y(n3870) );
  INVX2TS U2000 ( .A(n3869), .Y(n3867) );
  INVX2TS U2001 ( .A(n3866), .Y(n3864) );
  INVX2TS U2002 ( .A(n3863), .Y(n3861) );
  INVX2TS U2003 ( .A(n3860), .Y(n3858) );
  INVX2TS U2004 ( .A(n3857), .Y(n3855) );
  INVX2TS U2005 ( .A(n3854), .Y(n3852) );
  INVX2TS U2006 ( .A(n3851), .Y(n3849) );
  INVX2TS U2007 ( .A(n3848), .Y(n3846) );
  INVX2TS U2008 ( .A(n3845), .Y(n3843) );
  INVX2TS U2009 ( .A(n3842), .Y(n3840) );
  INVX2TS U2010 ( .A(n3839), .Y(n3837) );
  INVX2TS U2011 ( .A(n3836), .Y(n3834) );
  INVX2TS U2012 ( .A(n3833), .Y(n3831) );
  INVX2TS U2013 ( .A(n3830), .Y(n3828) );
  INVX2TS U2014 ( .A(n3827), .Y(n3825) );
  INVX2TS U2015 ( .A(n3824), .Y(n3822) );
  INVX2TS U2016 ( .A(n3938), .Y(n3936) );
  INVX2TS U2017 ( .A(n3953), .Y(n3951) );
  INVX2TS U2018 ( .A(n3947), .Y(n3945) );
  INVX2TS U2019 ( .A(n3944), .Y(n3942) );
  INVX2TS U2020 ( .A(n3941), .Y(n3939) );
  INVX2TS U2021 ( .A(n3950), .Y(n3948) );
  INVX2TS U2022 ( .A(n3935), .Y(n3933) );
  INVX2TS U2023 ( .A(n3932), .Y(n3930) );
  INVX2TS U2024 ( .A(n3926), .Y(n3924) );
  INVX2TS U2025 ( .A(n3929), .Y(n3927) );
  INVX2TS U2026 ( .A(n3923), .Y(n3921) );
  INVX2TS U2027 ( .A(n3920), .Y(n3918) );
  INVX2TS U2028 ( .A(n6222), .Y(n6254) );
  INVX2TS U2029 ( .A(n4088), .Y(n4086) );
  INVX2TS U2030 ( .A(n4091), .Y(n4089) );
  INVX2TS U2031 ( .A(n4082), .Y(n4080) );
  INVX2TS U2032 ( .A(n4085), .Y(n4083) );
  INVX2TS U2033 ( .A(n4079), .Y(n4077) );
  INVX2TS U2034 ( .A(n4076), .Y(n4074) );
  INVX2TS U2035 ( .A(n4241), .Y(n4239) );
  INVX2TS U2036 ( .A(n4238), .Y(n4236) );
  INVX2TS U2037 ( .A(n4235), .Y(n4233) );
  INVX2TS U2038 ( .A(n4232), .Y(n4230) );
  INVX2TS U2039 ( .A(n4247), .Y(n4245) );
  INVX2TS U2040 ( .A(n4244), .Y(n4242) );
  CLKBUFX2TS U2041 ( .A(n4419), .Y(n4421) );
  CLKBUFX2TS U2042 ( .A(n4416), .Y(n4418) );
  CLKBUFX2TS U2043 ( .A(n4413), .Y(n4415) );
  CLKBUFX2TS U2044 ( .A(n4407), .Y(n4409) );
  CLKBUFX2TS U2045 ( .A(n4404), .Y(n4406) );
  CLKBUFX2TS U2046 ( .A(n4410), .Y(n4412) );
  CLKBUFX2TS U2047 ( .A(n4380), .Y(n4382) );
  CLKBUFX2TS U2048 ( .A(n4377), .Y(n4379) );
  CLKBUFX2TS U2049 ( .A(n4368), .Y(n4370) );
  CLKBUFX2TS U2050 ( .A(n4365), .Y(n4367) );
  CLKBUFX2TS U2051 ( .A(n4353), .Y(n4355) );
  CLKBUFX2TS U2052 ( .A(n4347), .Y(n4349) );
  CLKBUFX2TS U2053 ( .A(n4344), .Y(n4346) );
  CLKBUFX2TS U2054 ( .A(n4341), .Y(n4343) );
  CLKBUFX2TS U2055 ( .A(n4335), .Y(n4337) );
  CLKBUFX2TS U2056 ( .A(n4332), .Y(n4334) );
  CLKBUFX2TS U2057 ( .A(n4329), .Y(n4331) );
  CLKBUFX2TS U2058 ( .A(n4326), .Y(n4328) );
  CLKBUFX2TS U2059 ( .A(n4323), .Y(n4325) );
  CLKBUFX2TS U2060 ( .A(n4320), .Y(n4322) );
  CLKBUFX2TS U2061 ( .A(n4314), .Y(n4316) );
  CLKBUFX2TS U2062 ( .A(n4302), .Y(n4304) );
  CLKBUFX2TS U2063 ( .A(n4299), .Y(n4301) );
  CLKBUFX2TS U2064 ( .A(n4374), .Y(n4376) );
  CLKBUFX2TS U2065 ( .A(n4371), .Y(n4373) );
  CLKBUFX2TS U2066 ( .A(n4359), .Y(n4361) );
  CLKBUFX2TS U2067 ( .A(n4350), .Y(n4352) );
  CLKBUFX2TS U2068 ( .A(n4317), .Y(n4319) );
  CLKBUFX2TS U2069 ( .A(n4305), .Y(n4307) );
  CLKBUFX2TS U2070 ( .A(n4293), .Y(n4295) );
  CLKBUFX2TS U2071 ( .A(n4383), .Y(n4385) );
  CLKBUFX2TS U2072 ( .A(n4362), .Y(n4364) );
  CLKBUFX2TS U2073 ( .A(n4356), .Y(n4358) );
  CLKBUFX2TS U2074 ( .A(n4338), .Y(n4340) );
  CLKBUFX2TS U2075 ( .A(n4308), .Y(n4310) );
  CLKBUFX2TS U2076 ( .A(n4296), .Y(n4298) );
  CLKBUFX2TS U2077 ( .A(n4290), .Y(n4292) );
  CLKBUFX2TS U2078 ( .A(n4311), .Y(n4313) );
  INVX2TS U2079 ( .A(n4013), .Y(n4011) );
  INVX2TS U2080 ( .A(n3983), .Y(n3981) );
  INVX2TS U2081 ( .A(n4070), .Y(n4068) );
  INVX2TS U2082 ( .A(n4067), .Y(n4065) );
  INVX2TS U2083 ( .A(n4064), .Y(n4062) );
  INVX2TS U2084 ( .A(n4061), .Y(n4059) );
  INVX2TS U2085 ( .A(n4058), .Y(n4056) );
  INVX2TS U2086 ( .A(n4055), .Y(n4053) );
  INVX2TS U2087 ( .A(n4049), .Y(n4047) );
  INVX2TS U2088 ( .A(n4043), .Y(n4041) );
  INVX2TS U2089 ( .A(n4040), .Y(n4038) );
  INVX2TS U2090 ( .A(n4037), .Y(n4035) );
  INVX2TS U2091 ( .A(n4034), .Y(n4032) );
  INVX2TS U2092 ( .A(n4019), .Y(n4017) );
  INVX2TS U2093 ( .A(n4016), .Y(n4014) );
  INVX2TS U2094 ( .A(n4010), .Y(n4008) );
  INVX2TS U2095 ( .A(n4007), .Y(n4005) );
  INVX2TS U2096 ( .A(n4004), .Y(n4002) );
  INVX2TS U2097 ( .A(n4001), .Y(n3999) );
  INVX2TS U2098 ( .A(n3995), .Y(n3993) );
  INVX2TS U2099 ( .A(n3992), .Y(n3990) );
  INVX2TS U2100 ( .A(n4073), .Y(n4071) );
  INVX2TS U2101 ( .A(n4052), .Y(n4050) );
  INVX2TS U2102 ( .A(n4046), .Y(n4044) );
  INVX2TS U2103 ( .A(n4028), .Y(n4026) );
  INVX2TS U2104 ( .A(n3998), .Y(n3996) );
  INVX2TS U2105 ( .A(n3986), .Y(n3984) );
  INVX2TS U2106 ( .A(n3980), .Y(n3978) );
  INVX2TS U2107 ( .A(n4031), .Y(n4029) );
  INVX2TS U2108 ( .A(n4025), .Y(n4023) );
  INVX2TS U2109 ( .A(n4022), .Y(n4020) );
  INVX2TS U2110 ( .A(n3989), .Y(n3987) );
  INVX2TS U2111 ( .A(n4109), .Y(n4107) );
  INVX2TS U2112 ( .A(n4106), .Y(n4104) );
  INVX2TS U2113 ( .A(n4103), .Y(n4101) );
  INVX2TS U2114 ( .A(n4100), .Y(n4098) );
  INVX2TS U2115 ( .A(n4097), .Y(n4095) );
  INVX2TS U2116 ( .A(n4094), .Y(n4092) );
  INVX2TS U2117 ( .A(n3821), .Y(n3819) );
  CLKBUFX2TS U2118 ( .A(n3972), .Y(n3973) );
  CLKBUFX2TS U2119 ( .A(n3960), .Y(n3961) );
  CLKBUFX2TS U2120 ( .A(n3954), .Y(n3955) );
  CLKBUFX2TS U2121 ( .A(n3969), .Y(n3970) );
  CLKBUFX2TS U2122 ( .A(n3963), .Y(n3964) );
  CLKBUFX2TS U2123 ( .A(n3975), .Y(n3976) );
  CLKBUFX2TS U2124 ( .A(n3966), .Y(n3967) );
  CLKBUFX2TS U2125 ( .A(n3957), .Y(n3958) );
  CLKBUFX2TS U2126 ( .A(n4284), .Y(n4285) );
  CLKBUFX2TS U2127 ( .A(n4278), .Y(n4279) );
  CLKBUFX2TS U2128 ( .A(n4275), .Y(n4276) );
  CLKBUFX2TS U2129 ( .A(n4287), .Y(n4288) );
  CLKBUFX2TS U2130 ( .A(n4281), .Y(n4282) );
  CLKBUFX2TS U2131 ( .A(n4272), .Y(n4273) );
  CLKBUFX2TS U2132 ( .A(n4131), .Y(n4132) );
  CLKBUFX2TS U2133 ( .A(n4128), .Y(n4129) );
  CLKBUFX2TS U2134 ( .A(n4122), .Y(n4123) );
  CLKBUFX2TS U2135 ( .A(n4116), .Y(n4117) );
  CLKBUFX2TS U2136 ( .A(n4110), .Y(n4111) );
  CLKBUFX2TS U2137 ( .A(n4125), .Y(n4126) );
  CLKBUFX2TS U2138 ( .A(n4119), .Y(n4120) );
  CLKBUFX2TS U2139 ( .A(n4113), .Y(n4114) );
  CLKBUFX2TS U2140 ( .A(n4128), .Y(n4130) );
  CLKBUFX2TS U2141 ( .A(n4110), .Y(n4112) );
  CLKBUFX2TS U2142 ( .A(n3972), .Y(n3974) );
  CLKBUFX2TS U2143 ( .A(n3966), .Y(n3968) );
  CLKBUFX2TS U2144 ( .A(n3954), .Y(n3956) );
  CLKBUFX2TS U2145 ( .A(n4122), .Y(n4124) );
  CLKBUFX2TS U2146 ( .A(n4119), .Y(n4121) );
  CLKBUFX2TS U2147 ( .A(n3963), .Y(n3965) );
  CLKBUFX2TS U2148 ( .A(n3975), .Y(n3977) );
  CLKBUFX2TS U2149 ( .A(n4131), .Y(n4133) );
  CLKBUFX2TS U2150 ( .A(n3969), .Y(n3971) );
  CLKBUFX2TS U2151 ( .A(n4125), .Y(n4127) );
  CLKBUFX2TS U2152 ( .A(n3960), .Y(n3962) );
  CLKBUFX2TS U2153 ( .A(n4116), .Y(n4118) );
  CLKBUFX2TS U2154 ( .A(n3957), .Y(n3959) );
  CLKBUFX2TS U2155 ( .A(n4113), .Y(n4115) );
  CLKBUFX2TS U2156 ( .A(n4284), .Y(n4286) );
  CLKBUFX2TS U2157 ( .A(n4272), .Y(n4274) );
  CLKBUFX2TS U2158 ( .A(n4281), .Y(n4283) );
  CLKBUFX2TS U2159 ( .A(n4275), .Y(n4277) );
  CLKBUFX2TS U2160 ( .A(n4287), .Y(n4289) );
  CLKBUFX2TS U2161 ( .A(n4278), .Y(n4280) );
  CLKBUFX2TS U2162 ( .A(n4398), .Y(n4400) );
  CLKBUFX2TS U2163 ( .A(n4389), .Y(n4391) );
  CLKBUFX2TS U2164 ( .A(n4386), .Y(n4388) );
  CLKBUFX2TS U2165 ( .A(n4401), .Y(n4403) );
  CLKBUFX2TS U2166 ( .A(n4395), .Y(n4397) );
  CLKBUFX2TS U2167 ( .A(n4392), .Y(n4394) );
  CLKBUFX2TS U2168 ( .A(n3815), .Y(n3814) );
  INVX2TS U2169 ( .A(n3805), .Y(n3803) );
  INVX2TS U2170 ( .A(n3818), .Y(n3816) );
  INVX2TS U2171 ( .A(n3811), .Y(n3809) );
  INVX2TS U2172 ( .A(n3863), .Y(n3862) );
  INVX2TS U2173 ( .A(n3911), .Y(n3910) );
  INVX2TS U2174 ( .A(n3887), .Y(n3886) );
  INVX2TS U2175 ( .A(n3860), .Y(n3859) );
  INVX2TS U2176 ( .A(n3854), .Y(n3853) );
  INVX2TS U2177 ( .A(n3842), .Y(n3841) );
  INVX2TS U2178 ( .A(n3917), .Y(n3916) );
  INVX2TS U2179 ( .A(n3914), .Y(n3913) );
  INVX2TS U2180 ( .A(n3902), .Y(n3901) );
  INVX2TS U2181 ( .A(n3896), .Y(n3895) );
  INVX2TS U2182 ( .A(n3890), .Y(n3889) );
  INVX2TS U2183 ( .A(n3881), .Y(n3880) );
  INVX2TS U2184 ( .A(n3872), .Y(n3871) );
  INVX2TS U2185 ( .A(n3857), .Y(n3856) );
  INVX2TS U2186 ( .A(n3848), .Y(n3847) );
  INVX2TS U2187 ( .A(n3908), .Y(n3907) );
  INVX2TS U2188 ( .A(n3905), .Y(n3904) );
  INVX2TS U2189 ( .A(n3893), .Y(n3892) );
  INVX2TS U2190 ( .A(n3884), .Y(n3883) );
  INVX2TS U2191 ( .A(n3851), .Y(n3850) );
  INVX2TS U2192 ( .A(n3839), .Y(n3838) );
  INVX2TS U2193 ( .A(n3830), .Y(n3829) );
  INVX2TS U2194 ( .A(n3827), .Y(n3826) );
  INVX2TS U2195 ( .A(n3824), .Y(n3823) );
  INVX2TS U2196 ( .A(n3845), .Y(n3844) );
  INVX2TS U2197 ( .A(n3875), .Y(n3874) );
  INVX2TS U2198 ( .A(n3869), .Y(n3868) );
  INVX2TS U2199 ( .A(n3866), .Y(n3865) );
  INVX2TS U2200 ( .A(n3833), .Y(n3832) );
  INVX2TS U2201 ( .A(n3899), .Y(n3898) );
  INVX2TS U2202 ( .A(n3878), .Y(n3877) );
  INVX2TS U2203 ( .A(n3836), .Y(n3835) );
  INVX2TS U2204 ( .A(n3953), .Y(n3952) );
  INVX2TS U2205 ( .A(n3950), .Y(n3949) );
  INVX2TS U2206 ( .A(n3947), .Y(n3946) );
  INVX2TS U2207 ( .A(n3941), .Y(n3940) );
  INVX2TS U2208 ( .A(n3938), .Y(n3937) );
  INVX2TS U2209 ( .A(n3944), .Y(n3943) );
  INVX2TS U2210 ( .A(n3805), .Y(n3804) );
  INVX2TS U2211 ( .A(n4262), .Y(n4261) );
  INVX2TS U2212 ( .A(n4250), .Y(n4249) );
  INVX2TS U2213 ( .A(n4265), .Y(n4264) );
  INVX2TS U2214 ( .A(n4259), .Y(n4258) );
  INVX2TS U2215 ( .A(n4256), .Y(n4255) );
  INVX2TS U2216 ( .A(n4253), .Y(n4252) );
  INVX2TS U2217 ( .A(n4226), .Y(n4225) );
  INVX2TS U2218 ( .A(n4223), .Y(n4222) );
  INVX2TS U2219 ( .A(n4220), .Y(n4219) );
  INVX2TS U2220 ( .A(n4217), .Y(n4216) );
  INVX2TS U2221 ( .A(n4214), .Y(n4213) );
  INVX2TS U2222 ( .A(n4211), .Y(n4210) );
  INVX2TS U2223 ( .A(n4205), .Y(n4204) );
  INVX2TS U2224 ( .A(n4199), .Y(n4198) );
  INVX2TS U2225 ( .A(n4196), .Y(n4195) );
  INVX2TS U2226 ( .A(n4193), .Y(n4192) );
  INVX2TS U2227 ( .A(n4190), .Y(n4189) );
  INVX2TS U2228 ( .A(n4187), .Y(n4186) );
  INVX2TS U2229 ( .A(n4181), .Y(n4180) );
  INVX2TS U2230 ( .A(n4178), .Y(n4177) );
  INVX2TS U2231 ( .A(n4175), .Y(n4174) );
  INVX2TS U2232 ( .A(n4172), .Y(n4171) );
  INVX2TS U2233 ( .A(n4169), .Y(n4168) );
  INVX2TS U2234 ( .A(n4166), .Y(n4165) );
  INVX2TS U2235 ( .A(n4163), .Y(n4162) );
  INVX2TS U2236 ( .A(n4160), .Y(n4159) );
  INVX2TS U2237 ( .A(n4157), .Y(n4156) );
  INVX2TS U2238 ( .A(n4151), .Y(n4150) );
  INVX2TS U2239 ( .A(n4148), .Y(n4147) );
  INVX2TS U2240 ( .A(n4145), .Y(n4144) );
  INVX2TS U2241 ( .A(n4139), .Y(n4138) );
  INVX2TS U2242 ( .A(n4229), .Y(n4228) );
  INVX2TS U2243 ( .A(n4208), .Y(n4207) );
  INVX2TS U2244 ( .A(n4202), .Y(n4201) );
  INVX2TS U2245 ( .A(n4184), .Y(n4183) );
  INVX2TS U2246 ( .A(n4154), .Y(n4153) );
  INVX2TS U2247 ( .A(n4142), .Y(n4141) );
  INVX2TS U2248 ( .A(n4136), .Y(n4135) );
  INVX2TS U2249 ( .A(n3818), .Y(n3817) );
  INVX2TS U2250 ( .A(n4247), .Y(n4246) );
  INVX2TS U2251 ( .A(n4244), .Y(n4243) );
  INVX2TS U2252 ( .A(n4238), .Y(n4237) );
  INVX2TS U2253 ( .A(n4241), .Y(n4240) );
  INVX2TS U2254 ( .A(n4235), .Y(n4234) );
  INVX2TS U2255 ( .A(n4232), .Y(n4231) );
  INVX2TS U2256 ( .A(n3811), .Y(n3810) );
  INVX2TS U2257 ( .A(n4073), .Y(n4072) );
  INVX2TS U2258 ( .A(n4070), .Y(n4069) );
  INVX2TS U2259 ( .A(n4067), .Y(n4066) );
  INVX2TS U2260 ( .A(n4064), .Y(n4063) );
  INVX2TS U2261 ( .A(n4061), .Y(n4060) );
  INVX2TS U2262 ( .A(n4058), .Y(n4057) );
  INVX2TS U2263 ( .A(n4052), .Y(n4051) );
  INVX2TS U2264 ( .A(n4049), .Y(n4048) );
  INVX2TS U2265 ( .A(n4046), .Y(n4045) );
  INVX2TS U2266 ( .A(n4043), .Y(n4042) );
  INVX2TS U2267 ( .A(n4040), .Y(n4039) );
  INVX2TS U2268 ( .A(n4037), .Y(n4036) );
  INVX2TS U2269 ( .A(n4031), .Y(n4030) );
  INVX2TS U2270 ( .A(n4028), .Y(n4027) );
  INVX2TS U2271 ( .A(n4025), .Y(n4024) );
  INVX2TS U2272 ( .A(n4022), .Y(n4021) );
  INVX2TS U2273 ( .A(n4019), .Y(n4018) );
  INVX2TS U2274 ( .A(n4016), .Y(n4015) );
  INVX2TS U2275 ( .A(n4013), .Y(n4012) );
  INVX2TS U2276 ( .A(n4010), .Y(n4009) );
  INVX2TS U2277 ( .A(n4007), .Y(n4006) );
  INVX2TS U2278 ( .A(n4004), .Y(n4003) );
  INVX2TS U2279 ( .A(n4001), .Y(n4000) );
  INVX2TS U2280 ( .A(n3998), .Y(n3997) );
  INVX2TS U2281 ( .A(n3995), .Y(n3994) );
  INVX2TS U2282 ( .A(n3989), .Y(n3988) );
  INVX2TS U2283 ( .A(n3986), .Y(n3985) );
  INVX2TS U2284 ( .A(n3983), .Y(n3982) );
  INVX2TS U2285 ( .A(n3980), .Y(n3979) );
  INVX2TS U2286 ( .A(n4055), .Y(n4054) );
  INVX2TS U2287 ( .A(n4034), .Y(n4033) );
  INVX2TS U2288 ( .A(n3992), .Y(n3991) );
  INVX2TS U2289 ( .A(n4094), .Y(n4093) );
  INVX2TS U2290 ( .A(n4109), .Y(n4108) );
  INVX2TS U2291 ( .A(n4103), .Y(n4102) );
  INVX2TS U2292 ( .A(n4100), .Y(n4099) );
  INVX2TS U2293 ( .A(n4097), .Y(n4096) );
  INVX2TS U2294 ( .A(n4106), .Y(n4105) );
  INVX2TS U2295 ( .A(n4091), .Y(n4090) );
  INVX2TS U2296 ( .A(n4088), .Y(n4087) );
  INVX2TS U2297 ( .A(n4085), .Y(n4084) );
  INVX2TS U2298 ( .A(n4082), .Y(n4081) );
  INVX2TS U2299 ( .A(n4079), .Y(n4078) );
  INVX2TS U2300 ( .A(n4076), .Y(n4075) );
  INVX2TS U2301 ( .A(n3929), .Y(n3928) );
  INVX2TS U2302 ( .A(n3926), .Y(n3925) );
  INVX2TS U2303 ( .A(n3923), .Y(n3922) );
  INVX2TS U2304 ( .A(n3920), .Y(n3919) );
  INVX2TS U2305 ( .A(n3935), .Y(n3934) );
  INVX2TS U2306 ( .A(n3932), .Y(n3931) );
  INVX2TS U2307 ( .A(n3821), .Y(n3820) );
  INVX2TS U2308 ( .A(n3808), .Y(n3806) );
  INVX2TS U2309 ( .A(n4265), .Y(n4263) );
  INVX2TS U2310 ( .A(n4259), .Y(n4257) );
  INVX2TS U2311 ( .A(n4253), .Y(n4251) );
  INVX2TS U2312 ( .A(n4250), .Y(n4248) );
  INVX2TS U2313 ( .A(n4256), .Y(n4254) );
  INVX2TS U2314 ( .A(n4175), .Y(n4173) );
  INVX2TS U2315 ( .A(n4223), .Y(n4221) );
  INVX2TS U2316 ( .A(n4199), .Y(n4197) );
  INVX2TS U2317 ( .A(n4172), .Y(n4170) );
  INVX2TS U2318 ( .A(n4166), .Y(n4164) );
  INVX2TS U2319 ( .A(n4154), .Y(n4152) );
  INVX2TS U2320 ( .A(n4229), .Y(n4227) );
  INVX2TS U2321 ( .A(n4226), .Y(n4224) );
  INVX2TS U2322 ( .A(n4214), .Y(n4212) );
  INVX2TS U2323 ( .A(n4208), .Y(n4206) );
  INVX2TS U2324 ( .A(n4202), .Y(n4200) );
  INVX2TS U2325 ( .A(n4193), .Y(n4191) );
  INVX2TS U2326 ( .A(n4184), .Y(n4182) );
  INVX2TS U2327 ( .A(n4169), .Y(n4167) );
  INVX2TS U2328 ( .A(n4160), .Y(n4158) );
  INVX2TS U2329 ( .A(n4220), .Y(n4218) );
  INVX2TS U2330 ( .A(n4217), .Y(n4215) );
  INVX2TS U2331 ( .A(n4205), .Y(n4203) );
  INVX2TS U2332 ( .A(n4196), .Y(n4194) );
  INVX2TS U2333 ( .A(n4163), .Y(n4161) );
  INVX2TS U2334 ( .A(n4151), .Y(n4149) );
  INVX2TS U2335 ( .A(n4142), .Y(n4140) );
  INVX2TS U2336 ( .A(n4139), .Y(n4137) );
  INVX2TS U2337 ( .A(n4136), .Y(n4134) );
  INVX2TS U2338 ( .A(n4157), .Y(n4155) );
  INVX2TS U2339 ( .A(n4187), .Y(n4185) );
  INVX2TS U2340 ( .A(n4181), .Y(n4179) );
  INVX2TS U2341 ( .A(n4178), .Y(n4176) );
  INVX2TS U2342 ( .A(n4145), .Y(n4143) );
  INVX2TS U2343 ( .A(n4262), .Y(n4260) );
  INVX2TS U2344 ( .A(n4211), .Y(n4209) );
  INVX2TS U2345 ( .A(n4190), .Y(n4188) );
  INVX2TS U2346 ( .A(n4148), .Y(n4146) );
  INVX2TS U2347 ( .A(n3808), .Y(n3807) );
  INVX2TS U2348 ( .A(n4848), .Y(n6320) );
  INVX2TS U2349 ( .A(n4845), .Y(n6319) );
  CLKBUFX2TS U2350 ( .A(n5301), .Y(n514) );
  CLKBUFX2TS U2351 ( .A(n536), .Y(n516) );
  CLKBUFX2TS U2352 ( .A(n536), .Y(n517) );
  CLKBUFX2TS U2353 ( .A(n536), .Y(n526) );
  CLKBUFX2TS U2354 ( .A(n9), .Y(n3658) );
  CLKBUFX2TS U2355 ( .A(n222), .Y(n3581) );
  CLKBUFX2TS U2356 ( .A(n9), .Y(n3659) );
  CLKBUFX2TS U2357 ( .A(n222), .Y(n3582) );
  CLKBUFX2TS U2358 ( .A(n6315), .Y(n3597) );
  CLKBUFX2TS U2359 ( .A(n1), .Y(n3629) );
  CLKBUFX2TS U2360 ( .A(n1), .Y(n3628) );
  CLKBUFX2TS U2361 ( .A(n6315), .Y(n3596) );
  INVX2TS U2362 ( .A(n5286), .Y(n6317) );
  CLKBUFX2TS U2363 ( .A(n3598), .Y(n3591) );
  CLKBUFX2TS U2364 ( .A(n6315), .Y(n3598) );
  CLKBUFX2TS U2365 ( .A(n3567), .Y(n3561) );
  CLKBUFX2TS U2366 ( .A(n6314), .Y(n3567) );
  INVX2TS U2367 ( .A(n5298), .Y(n6316) );
  CLKBUFX2TS U2368 ( .A(n511), .Y(n508) );
  CLKBUFX2TS U2369 ( .A(n511), .Y(n509) );
  AOI21X1TS U2370 ( .A0(n6250), .A1(n432), .B0(n5347), .Y(n5315) );
  XNOR2X1TS U2371 ( .A(n4858), .B(n4862), .Y(n6231) );
  XNOR2X1TS U2372 ( .A(n148), .B(n6231), .Y(n4859) );
  NOR2X1TS U2373 ( .A(n155), .B(n5316), .Y(n5317) );
  NOR3X1TS U2374 ( .A(n6321), .B(n5327), .C(n6249), .Y(n4861) );
  OAI211X1TS U2375 ( .A0(n4853), .A1(n4852), .B0(n4851), .C0(n4850), .Y(n4856)
         );
  NAND3BX1TS U2376 ( .AN(n6227), .B(n6225), .C(n4848), .Y(n4851) );
  OAI21X1TS U2377 ( .A0(n6251), .A1(n4865), .B0(n4849), .Y(n4850) );
  OAI32X1TS U2378 ( .A0(n4849), .A1(n6251), .A2(n4865), .B0(n6227), .B1(n4857), 
        .Y(n4852) );
  NOR2X1TS U2379 ( .A(n5346), .B(n6236), .Y(n5463) );
  INVX2TS U2380 ( .A(n5524), .Y(n6330) );
  AND2X2TS U2381 ( .A(n4871), .B(n331), .Y(n4870) );
  XOR2X1TS U2382 ( .A(n4867), .B(n4866), .Y(n6230) );
  XNOR2X1TS U2383 ( .A(n224), .B(n4864), .Y(n4867) );
  INVX2TS U2384 ( .A(n4843), .Y(n6248) );
  AND2X2TS U2385 ( .A(n422), .B(n4870), .Y(n5314) );
  INVX2TS U2386 ( .A(n5316), .Y(n6326) );
  INVX2TS U2387 ( .A(n4854), .Y(n6249) );
  OAI221XLTS U2388 ( .A0(n5581), .A1(n237), .B0(n3373), .B1(n18), .C0(n5580), 
        .Y(n2576) );
  AOI222XLTS U2389 ( .A0(n3803), .A1(n3317), .B0(n3817), .B1(n3327), .C0(n3809), .C1(n3363), .Y(n5580) );
  OAI221XLTS U2390 ( .A0(n5585), .A1(n237), .B0(n3504), .B1(n10), .C0(n5584), 
        .Y(n2578) );
  AOI222XLTS U2391 ( .A0(n3803), .A1(n3448), .B0(n3817), .B1(n3458), .C0(n3810), .C1(n3496), .Y(n5584) );
  NOR2X1TS U2392 ( .A(n6328), .B(n5326), .Y(n5555) );
  OAI33XLTS U2393 ( .A0(n6238), .A1(n6327), .A2(n5540), .B0(n3814), .B1(n6337), 
        .B2(n178), .Y(n5541) );
  XOR2X1TS U2394 ( .A(n4855), .B(n16), .Y(n6234) );
  NAND2X1TS U2395 ( .A(n3806), .B(n6336), .Y(n5522) );
  INVX2TS U2396 ( .A(n3814), .Y(n3813) );
  NAND2X1TS U2397 ( .A(n3806), .B(n6333), .Y(n5551) );
  NOR2X1TS U2398 ( .A(n5306), .B(n6252), .Y(n5282) );
  NOR2X1TS U2399 ( .A(n5307), .B(n6252), .Y(n5281) );
  OAI2BB2XLTS U2400 ( .B0(n217), .B1(n6238), .A0N(n217), .A1N(n3819), .Y(n5546) );
  INVX2TS U2401 ( .A(n5313), .Y(n564) );
  NAND4X1TS U2402 ( .A(n5307), .B(n5305), .C(n5303), .D(n4873), .Y(n5313) );
  AND3X2TS U2403 ( .A(n5295), .B(n5306), .C(n5304), .Y(n4873) );
  OAI222X1TS U2404 ( .A0(n3808), .A1(n5307), .B0(n3815), .B1(n5306), .C0(n193), 
        .C1(n5305), .Y(n5308) );
  OR2X2TS U2405 ( .A(n5304), .B(n6252), .Y(n430) );
  OAI211X1TS U2406 ( .A0(n3821), .A1(n5304), .B0(n5303), .C0(n6253), .Y(n5309)
         );
  INVX2TS U2407 ( .A(n5295), .Y(n6252) );
  NOR2X1TS U2408 ( .A(n6253), .B(reset), .Y(n6222) );
  NOR2X1TS U2409 ( .A(n5303), .B(n345), .Y(n5218) );
  INVX2TS U2410 ( .A(readIn_NORTH), .Y(n3821) );
  INVX2TS U2411 ( .A(writeIn_SOUTH), .Y(n3818) );
  INVX2TS U2412 ( .A(writeIn_WEST), .Y(n3805) );
  OAI221XLTS U2413 ( .A0(n236), .A1(n5304), .B0(n3811), .B1(n5306), .C0(n6253), 
        .Y(n5294) );
  INVX2TS U2414 ( .A(readIn_WEST), .Y(n3808) );
  INVX2TS U2415 ( .A(requesterAddressIn_WEST[4]), .Y(n3932) );
  INVX2TS U2416 ( .A(requesterAddressIn_WEST[1]), .Y(n3923) );
  INVX2TS U2417 ( .A(requesterAddressIn_WEST[0]), .Y(n3920) );
  INVX2TS U2418 ( .A(requesterAddressIn_WEST[5]), .Y(n3935) );
  INVX2TS U2419 ( .A(requesterAddressIn_WEST[3]), .Y(n3929) );
  INVX2TS U2420 ( .A(requesterAddressIn_WEST[2]), .Y(n3926) );
  INVX2TS U2421 ( .A(requesterAddressIn_EAST[5]), .Y(n4091) );
  INVX2TS U2422 ( .A(requesterAddressIn_EAST[3]), .Y(n4085) );
  INVX2TS U2423 ( .A(requesterAddressIn_EAST[4]), .Y(n4088) );
  INVX2TS U2424 ( .A(requesterAddressIn_EAST[2]), .Y(n4082) );
  INVX2TS U2425 ( .A(requesterAddressIn_EAST[1]), .Y(n4079) );
  INVX2TS U2426 ( .A(requesterAddressIn_EAST[0]), .Y(n4076) );
  INVX2TS U2427 ( .A(dataIn_EAST[31]), .Y(n4073) );
  INVX2TS U2428 ( .A(dataIn_EAST[30]), .Y(n4070) );
  INVX2TS U2429 ( .A(dataIn_EAST[29]), .Y(n4067) );
  INVX2TS U2430 ( .A(dataIn_EAST[26]), .Y(n4058) );
  INVX2TS U2431 ( .A(dataIn_EAST[24]), .Y(n4052) );
  INVX2TS U2432 ( .A(dataIn_EAST[22]), .Y(n4046) );
  INVX2TS U2433 ( .A(dataIn_EAST[21]), .Y(n4043) );
  INVX2TS U2434 ( .A(dataIn_EAST[19]), .Y(n4037) );
  INVX2TS U2435 ( .A(dataIn_EAST[17]), .Y(n4031) );
  INVX2TS U2436 ( .A(dataIn_EAST[16]), .Y(n4028) );
  INVX2TS U2437 ( .A(dataIn_EAST[14]), .Y(n4022) );
  INVX2TS U2438 ( .A(dataIn_EAST[12]), .Y(n4016) );
  INVX2TS U2439 ( .A(dataIn_EAST[11]), .Y(n4013) );
  INVX2TS U2440 ( .A(dataIn_EAST[10]), .Y(n4010) );
  INVX2TS U2441 ( .A(dataIn_EAST[8]), .Y(n4004) );
  INVX2TS U2442 ( .A(dataIn_EAST[6]), .Y(n3998) );
  INVX2TS U2443 ( .A(dataIn_EAST[3]), .Y(n3989) );
  INVX2TS U2444 ( .A(dataIn_EAST[25]), .Y(n4055) );
  INVX2TS U2445 ( .A(dataIn_EAST[18]), .Y(n4034) );
  INVX2TS U2446 ( .A(dataIn_EAST[15]), .Y(n4025) );
  INVX2TS U2447 ( .A(dataIn_EAST[13]), .Y(n4019) );
  INVX2TS U2448 ( .A(dataIn_EAST[4]), .Y(n3992) );
  INVX2TS U2449 ( .A(dataIn_EAST[28]), .Y(n4064) );
  INVX2TS U2450 ( .A(dataIn_EAST[27]), .Y(n4061) );
  INVX2TS U2451 ( .A(dataIn_EAST[23]), .Y(n4049) );
  INVX2TS U2452 ( .A(dataIn_EAST[20]), .Y(n4040) );
  INVX2TS U2453 ( .A(dataIn_EAST[9]), .Y(n4007) );
  INVX2TS U2454 ( .A(dataIn_EAST[5]), .Y(n3995) );
  INVX2TS U2455 ( .A(dataIn_EAST[2]), .Y(n3986) );
  INVX2TS U2456 ( .A(dataIn_EAST[1]), .Y(n3983) );
  INVX2TS U2457 ( .A(dataIn_EAST[0]), .Y(n3980) );
  INVX2TS U2458 ( .A(dataIn_EAST[7]), .Y(n4001) );
  INVX2TS U2459 ( .A(destinationAddressIn_EAST[5]), .Y(n4109) );
  INVX2TS U2460 ( .A(destinationAddressIn_EAST[3]), .Y(n4103) );
  INVX2TS U2461 ( .A(destinationAddressIn_EAST[1]), .Y(n4097) );
  INVX2TS U2462 ( .A(destinationAddressIn_EAST[4]), .Y(n4106) );
  INVX2TS U2463 ( .A(destinationAddressIn_EAST[0]), .Y(n4094) );
  INVX2TS U2464 ( .A(destinationAddressIn_EAST[2]), .Y(n4100) );
  INVX2TS U2465 ( .A(writeIn_EAST), .Y(n3811) );
  INVX2TS U2466 ( .A(destinationAddressIn_SOUTH[0]), .Y(n4250) );
  INVX2TS U2467 ( .A(requesterAddressIn_SOUTH[5]), .Y(n4247) );
  INVX2TS U2468 ( .A(requesterAddressIn_SOUTH[4]), .Y(n4244) );
  INVX2TS U2469 ( .A(requesterAddressIn_SOUTH[2]), .Y(n4238) );
  INVX2TS U2470 ( .A(destinationAddressIn_SOUTH[5]), .Y(n4265) );
  INVX2TS U2471 ( .A(destinationAddressIn_SOUTH[3]), .Y(n4259) );
  INVX2TS U2472 ( .A(destinationAddressIn_SOUTH[2]), .Y(n4256) );
  INVX2TS U2473 ( .A(destinationAddressIn_SOUTH[1]), .Y(n4253) );
  INVX2TS U2474 ( .A(dataIn_SOUTH[30]), .Y(n4226) );
  INVX2TS U2475 ( .A(dataIn_SOUTH[29]), .Y(n4223) );
  INVX2TS U2476 ( .A(dataIn_SOUTH[26]), .Y(n4214) );
  INVX2TS U2477 ( .A(dataIn_SOUTH[21]), .Y(n4199) );
  INVX2TS U2478 ( .A(dataIn_SOUTH[19]), .Y(n4193) );
  INVX2TS U2479 ( .A(dataIn_SOUTH[13]), .Y(n4175) );
  INVX2TS U2480 ( .A(dataIn_SOUTH[12]), .Y(n4172) );
  INVX2TS U2481 ( .A(dataIn_SOUTH[11]), .Y(n4169) );
  INVX2TS U2482 ( .A(dataIn_SOUTH[10]), .Y(n4166) );
  INVX2TS U2483 ( .A(dataIn_SOUTH[8]), .Y(n4160) );
  INVX2TS U2484 ( .A(requesterAddressIn_SOUTH[3]), .Y(n4241) );
  INVX2TS U2485 ( .A(requesterAddressIn_SOUTH[1]), .Y(n4235) );
  INVX2TS U2486 ( .A(requesterAddressIn_SOUTH[0]), .Y(n4232) );
  INVX2TS U2487 ( .A(dataIn_SOUTH[28]), .Y(n4220) );
  INVX2TS U2488 ( .A(dataIn_SOUTH[27]), .Y(n4217) );
  INVX2TS U2489 ( .A(dataIn_SOUTH[23]), .Y(n4205) );
  INVX2TS U2490 ( .A(dataIn_SOUTH[20]), .Y(n4196) );
  INVX2TS U2491 ( .A(dataIn_SOUTH[9]), .Y(n4163) );
  INVX2TS U2492 ( .A(dataIn_SOUTH[5]), .Y(n4151) );
  INVX2TS U2493 ( .A(dataIn_SOUTH[1]), .Y(n4139) );
  INVX2TS U2494 ( .A(dataIn_SOUTH[31]), .Y(n4229) );
  INVX2TS U2495 ( .A(dataIn_SOUTH[24]), .Y(n4208) );
  INVX2TS U2496 ( .A(dataIn_SOUTH[22]), .Y(n4202) );
  INVX2TS U2497 ( .A(dataIn_SOUTH[16]), .Y(n4184) );
  INVX2TS U2498 ( .A(dataIn_SOUTH[6]), .Y(n4154) );
  INVX2TS U2499 ( .A(dataIn_SOUTH[2]), .Y(n4142) );
  INVX2TS U2500 ( .A(dataIn_SOUTH[0]), .Y(n4136) );
  INVX2TS U2501 ( .A(dataIn_SOUTH[7]), .Y(n4157) );
  INVX2TS U2502 ( .A(dataIn_SOUTH[17]), .Y(n4187) );
  INVX2TS U2503 ( .A(dataIn_SOUTH[15]), .Y(n4181) );
  INVX2TS U2504 ( .A(dataIn_SOUTH[14]), .Y(n4178) );
  INVX2TS U2505 ( .A(dataIn_SOUTH[3]), .Y(n4145) );
  INVX2TS U2506 ( .A(destinationAddressIn_SOUTH[4]), .Y(n4262) );
  INVX2TS U2507 ( .A(dataIn_SOUTH[25]), .Y(n4211) );
  INVX2TS U2508 ( .A(dataIn_SOUTH[18]), .Y(n4190) );
  INVX2TS U2509 ( .A(dataIn_SOUTH[4]), .Y(n4148) );
  INVX2TS U2510 ( .A(dataIn_WEST[31]), .Y(n3917) );
  INVX2TS U2511 ( .A(dataIn_WEST[30]), .Y(n3914) );
  INVX2TS U2512 ( .A(dataIn_WEST[29]), .Y(n3911) );
  INVX2TS U2513 ( .A(dataIn_WEST[26]), .Y(n3902) );
  INVX2TS U2514 ( .A(dataIn_WEST[24]), .Y(n3896) );
  INVX2TS U2515 ( .A(dataIn_WEST[22]), .Y(n3890) );
  INVX2TS U2516 ( .A(dataIn_WEST[21]), .Y(n3887) );
  INVX2TS U2517 ( .A(dataIn_WEST[19]), .Y(n3881) );
  INVX2TS U2518 ( .A(dataIn_WEST[16]), .Y(n3872) );
  INVX2TS U2519 ( .A(dataIn_WEST[13]), .Y(n3863) );
  INVX2TS U2520 ( .A(dataIn_WEST[12]), .Y(n3860) );
  INVX2TS U2521 ( .A(dataIn_WEST[11]), .Y(n3857) );
  INVX2TS U2522 ( .A(dataIn_WEST[10]), .Y(n3854) );
  INVX2TS U2523 ( .A(dataIn_WEST[8]), .Y(n3848) );
  INVX2TS U2524 ( .A(dataIn_WEST[6]), .Y(n3842) );
  INVX2TS U2525 ( .A(dataIn_WEST[28]), .Y(n3908) );
  INVX2TS U2526 ( .A(dataIn_WEST[27]), .Y(n3905) );
  INVX2TS U2527 ( .A(dataIn_WEST[23]), .Y(n3893) );
  INVX2TS U2528 ( .A(dataIn_WEST[20]), .Y(n3884) );
  INVX2TS U2529 ( .A(dataIn_WEST[9]), .Y(n3851) );
  INVX2TS U2530 ( .A(dataIn_WEST[5]), .Y(n3839) );
  INVX2TS U2531 ( .A(dataIn_WEST[2]), .Y(n3830) );
  INVX2TS U2532 ( .A(dataIn_WEST[1]), .Y(n3827) );
  INVX2TS U2533 ( .A(dataIn_WEST[0]), .Y(n3824) );
  INVX2TS U2534 ( .A(dataIn_WEST[7]), .Y(n3845) );
  INVX2TS U2535 ( .A(dataIn_WEST[17]), .Y(n3875) );
  INVX2TS U2536 ( .A(dataIn_WEST[15]), .Y(n3869) );
  INVX2TS U2537 ( .A(dataIn_WEST[14]), .Y(n3866) );
  INVX2TS U2538 ( .A(dataIn_WEST[3]), .Y(n3833) );
  INVX2TS U2539 ( .A(dataIn_WEST[25]), .Y(n3899) );
  INVX2TS U2540 ( .A(dataIn_WEST[18]), .Y(n3878) );
  INVX2TS U2541 ( .A(dataIn_WEST[4]), .Y(n3836) );
  INVX2TS U2542 ( .A(destinationAddressIn_WEST[0]), .Y(n3938) );
  INVX2TS U2543 ( .A(destinationAddressIn_WEST[5]), .Y(n3953) );
  INVX2TS U2544 ( .A(destinationAddressIn_WEST[3]), .Y(n3947) );
  INVX2TS U2545 ( .A(destinationAddressIn_WEST[2]), .Y(n3944) );
  INVX2TS U2546 ( .A(destinationAddressIn_WEST[1]), .Y(n3941) );
  INVX2TS U2547 ( .A(destinationAddressIn_WEST[4]), .Y(n3950) );
  NOR2BX1TS U2548 ( .AN(n6233), .B(n6229), .Y(n2885) );
  AOI31X1TS U2549 ( .A0(n6228), .A1(n6320), .A2(n6227), .B0(n3549), .Y(n6229)
         );
  XNOR2X1TS U2550 ( .A(n6226), .B(n6225), .Y(n6228) );
  CLKBUFX2TS U2551 ( .A(destinationAddressIn_EAST[12]), .Y(n4128) );
  CLKBUFX2TS U2552 ( .A(destinationAddressIn_WEST[12]), .Y(n3972) );
  CLKBUFX2TS U2553 ( .A(destinationAddressIn_SOUTH[12]), .Y(n4284) );
  CLKBUFX2TS U2554 ( .A(destinationAddressIn_EAST[10]), .Y(n4122) );
  CLKBUFX2TS U2555 ( .A(destinationAddressIn_SOUTH[10]), .Y(n4278) );
  CLKBUFX2TS U2556 ( .A(destinationAddressIn_WEST[10]), .Y(n3966) );
  CLKBUFX2TS U2557 ( .A(destinationAddressIn_EAST[9]), .Y(n4119) );
  CLKBUFX2TS U2558 ( .A(destinationAddressIn_WEST[9]), .Y(n3963) );
  CLKBUFX2TS U2559 ( .A(destinationAddressIn_SOUTH[9]), .Y(n4275) );
  CLKBUFX2TS U2560 ( .A(destinationAddressIn_WEST[13]), .Y(n3975) );
  CLKBUFX2TS U2561 ( .A(destinationAddressIn_EAST[13]), .Y(n4131) );
  CLKBUFX2TS U2562 ( .A(destinationAddressIn_SOUTH[13]), .Y(n4287) );
  CLKBUFX2TS U2563 ( .A(destinationAddressIn_WEST[11]), .Y(n3969) );
  CLKBUFX2TS U2564 ( .A(destinationAddressIn_EAST[11]), .Y(n4125) );
  CLKBUFX2TS U2565 ( .A(destinationAddressIn_SOUTH[11]), .Y(n4281) );
  CLKBUFX2TS U2566 ( .A(destinationAddressIn_WEST[8]), .Y(n3960) );
  CLKBUFX2TS U2567 ( .A(destinationAddressIn_EAST[8]), .Y(n4116) );
  CLKBUFX2TS U2568 ( .A(destinationAddressIn_SOUTH[8]), .Y(n4272) );
  CLKBUFX2TS U2569 ( .A(destinationAddressIn_NORTH[0]), .Y(n4404) );
  CLKBUFX2TS U2570 ( .A(requesterAddressIn_NORTH[5]), .Y(n4401) );
  CLKBUFX2TS U2571 ( .A(requesterAddressIn_NORTH[4]), .Y(n4398) );
  CLKBUFX2TS U2572 ( .A(requesterAddressIn_NORTH[2]), .Y(n4392) );
  CLKBUFX2TS U2573 ( .A(destinationAddressIn_EAST[6]), .Y(n4110) );
  CLKBUFX2TS U2574 ( .A(destinationAddressIn_NORTH[5]), .Y(n4419) );
  CLKBUFX2TS U2575 ( .A(destinationAddressIn_NORTH[3]), .Y(n4413) );
  CLKBUFX2TS U2576 ( .A(destinationAddressIn_NORTH[2]), .Y(n4410) );
  CLKBUFX2TS U2577 ( .A(destinationAddressIn_NORTH[1]), .Y(n4407) );
  CLKBUFX2TS U2578 ( .A(dataIn_NORTH[30]), .Y(n4380) );
  CLKBUFX2TS U2579 ( .A(dataIn_NORTH[29]), .Y(n4377) );
  CLKBUFX2TS U2580 ( .A(dataIn_NORTH[26]), .Y(n4368) );
  CLKBUFX2TS U2581 ( .A(dataIn_NORTH[21]), .Y(n4353) );
  CLKBUFX2TS U2582 ( .A(dataIn_NORTH[19]), .Y(n4347) );
  CLKBUFX2TS U2583 ( .A(dataIn_NORTH[13]), .Y(n4329) );
  CLKBUFX2TS U2584 ( .A(dataIn_NORTH[12]), .Y(n4326) );
  CLKBUFX2TS U2585 ( .A(dataIn_NORTH[11]), .Y(n4323) );
  CLKBUFX2TS U2586 ( .A(dataIn_NORTH[10]), .Y(n4320) );
  CLKBUFX2TS U2587 ( .A(dataIn_NORTH[8]), .Y(n4314) );
  CLKBUFX2TS U2588 ( .A(requesterAddressIn_NORTH[3]), .Y(n4395) );
  CLKBUFX2TS U2589 ( .A(requesterAddressIn_NORTH[1]), .Y(n4389) );
  CLKBUFX2TS U2590 ( .A(requesterAddressIn_NORTH[0]), .Y(n4386) );
  CLKBUFX2TS U2591 ( .A(dataIn_NORTH[28]), .Y(n4374) );
  CLKBUFX2TS U2592 ( .A(dataIn_NORTH[27]), .Y(n4371) );
  CLKBUFX2TS U2593 ( .A(dataIn_NORTH[23]), .Y(n4359) );
  CLKBUFX2TS U2594 ( .A(dataIn_NORTH[20]), .Y(n4350) );
  CLKBUFX2TS U2595 ( .A(dataIn_NORTH[9]), .Y(n4317) );
  CLKBUFX2TS U2596 ( .A(dataIn_NORTH[5]), .Y(n4305) );
  CLKBUFX2TS U2597 ( .A(dataIn_NORTH[1]), .Y(n4293) );
  CLKBUFX2TS U2598 ( .A(destinationAddressIn_WEST[6]), .Y(n3954) );
  CLKBUFX2TS U2599 ( .A(dataIn_NORTH[31]), .Y(n4383) );
  CLKBUFX2TS U2600 ( .A(dataIn_NORTH[24]), .Y(n4362) );
  CLKBUFX2TS U2601 ( .A(dataIn_NORTH[22]), .Y(n4356) );
  CLKBUFX2TS U2602 ( .A(dataIn_NORTH[16]), .Y(n4338) );
  CLKBUFX2TS U2603 ( .A(dataIn_NORTH[6]), .Y(n4308) );
  CLKBUFX2TS U2604 ( .A(dataIn_NORTH[2]), .Y(n4296) );
  CLKBUFX2TS U2605 ( .A(dataIn_NORTH[0]), .Y(n4290) );
  CLKBUFX2TS U2606 ( .A(dataIn_NORTH[7]), .Y(n4311) );
  CLKBUFX2TS U2607 ( .A(dataIn_NORTH[17]), .Y(n4341) );
  CLKBUFX2TS U2608 ( .A(dataIn_NORTH[15]), .Y(n4335) );
  CLKBUFX2TS U2609 ( .A(dataIn_NORTH[14]), .Y(n4332) );
  CLKBUFX2TS U2610 ( .A(dataIn_NORTH[3]), .Y(n4299) );
  CLKBUFX2TS U2611 ( .A(destinationAddressIn_WEST[7]), .Y(n3957) );
  CLKBUFX2TS U2612 ( .A(destinationAddressIn_EAST[7]), .Y(n4113) );
  CLKBUFX2TS U2613 ( .A(destinationAddressIn_NORTH[4]), .Y(n4416) );
  CLKBUFX2TS U2614 ( .A(dataIn_NORTH[25]), .Y(n4365) );
  CLKBUFX2TS U2615 ( .A(dataIn_NORTH[18]), .Y(n4344) );
  CLKBUFX2TS U2616 ( .A(dataIn_NORTH[4]), .Y(n4302) );
  INVX2TS U2617 ( .A(readIn_EAST), .Y(n3815) );
  OAI21X1TS U2618 ( .A0(n6253), .A1(n6226), .B0(n4422), .Y(n6224) );
  OAI22X1TS U2619 ( .A0(n3536), .A1(n3619), .B0(n147), .B1(n6224), .Y(n2884)
         );
  XNOR2X1TS U2620 ( .A(n224), .B(n147), .Y(n6225) );
  AOI21X1TS U2621 ( .A0(n4), .A1(n121), .B0(n4845), .Y(n4848) );
  XNOR2X1TS U2622 ( .A(n6225), .B(n4847), .Y(n4849) );
  AOI21X1TS U2623 ( .A0(n5323), .A1(n6319), .B0(n4846), .Y(n4847) );
  AOI21X1TS U2624 ( .A0(n4845), .A1(n197), .B0(n148), .Y(n4846) );
  OAI22X1TS U2625 ( .A0(n6305), .A1(n501), .B0(n19), .B1(n3602), .Y(n5131) );
  OAI22X1TS U2626 ( .A0(n6306), .A1(n500), .B0(n20), .B1(n3601), .Y(n5139) );
  OAI22X1TS U2627 ( .A0(n6308), .A1(n500), .B0(n21), .B1(n3601), .Y(n5155) );
  OAI22X1TS U2628 ( .A0(n6309), .A1(n500), .B0(n22), .B1(n3601), .Y(n5163) );
  OAI22X1TS U2629 ( .A0(n6307), .A1(n500), .B0(n23), .B1(n3601), .Y(n5147) );
  OAI22X1TS U2630 ( .A0(n6310), .A1(n499), .B0(n24), .B1(n3600), .Y(n5171) );
  CLKBUFX2TS U2631 ( .A(n5301), .Y(n536) );
  INVX2TS U2632 ( .A(n5299), .Y(n6315) );
  INVX2TS U2633 ( .A(n5289), .Y(n6314) );
  NOR2X1TS U2634 ( .A(n6226), .B(n147), .Y(n5298) );
  INVX2TS U2635 ( .A(n275), .Y(n6313) );
  CLKBUFX2TS U2636 ( .A(n537), .Y(n511) );
  CLKBUFX2TS U2637 ( .A(n5301), .Y(n537) );
  AOI222XLTS U2638 ( .A0(n3961), .A1(n672), .B0(n4274), .B1(n610), .C0(n4117), 
        .C1(n415), .Y(n5331) );
  AOI222XLTS U2639 ( .A0(n3955), .A1(n672), .B0(n4268), .B1(n610), .C0(n4111), 
        .C1(n415), .Y(n5333) );
  AOI222XLTS U2640 ( .A0(n3803), .A1(n673), .B0(n3816), .B1(n610), .C0(n3809), 
        .C1(n415), .Y(n5568) );
  AOI222XLTS U2641 ( .A0(n3958), .A1(n672), .B0(n4271), .B1(n610), .C0(n4114), 
        .C1(n415), .Y(n5332) );
  AOI222XLTS U2642 ( .A0(n3973), .A1(n671), .B0(n4286), .B1(n612), .C0(n4129), 
        .C1(n416), .Y(n5325) );
  AOI222XLTS U2643 ( .A0(n4288), .A1(n820), .B0(destinationAddressIn_EAST[13]), 
        .B1(n804), .C0(n3977), .C1(n851), .Y(n5370) );
  AOI222XLTS U2644 ( .A0(n3976), .A1(n671), .B0(n4289), .B1(n624), .C0(n4132), 
        .C1(n417), .Y(n5324) );
  AOI222XLTS U2645 ( .A0(n3967), .A1(n671), .B0(n4280), .B1(n612), .C0(n4123), 
        .C1(n417), .Y(n5329) );
  AOI222XLTS U2646 ( .A0(n4282), .A1(n820), .B0(destinationAddressIn_EAST[11]), 
        .B1(n797), .C0(n3971), .C1(n851), .Y(n5372) );
  AOI222XLTS U2647 ( .A0(n4276), .A1(n821), .B0(destinationAddressIn_EAST[9]), 
        .B1(n797), .C0(n3965), .C1(n852), .Y(n5374) );
  AOI222XLTS U2648 ( .A0(n3816), .A1(n822), .B0(n3810), .B1(n798), .C0(n3804), 
        .C1(n853), .Y(n5573) );
  AOI222XLTS U2649 ( .A0(n3970), .A1(n671), .B0(n4283), .B1(n612), .C0(n4126), 
        .C1(n417), .Y(n5328) );
  AOI222XLTS U2650 ( .A0(n3964), .A1(n672), .B0(n4277), .B1(n611), .C0(n4120), 
        .C1(n417), .Y(n5330) );
  AOI222XLTS U2651 ( .A0(n4285), .A1(n820), .B0(destinationAddressIn_EAST[12]), 
        .B1(n797), .C0(n3974), .C1(n851), .Y(n5371) );
  AOI222XLTS U2652 ( .A0(n4279), .A1(n820), .B0(destinationAddressIn_EAST[10]), 
        .B1(n797), .C0(n3968), .C1(n852), .Y(n5373) );
  AOI222XLTS U2653 ( .A0(n4273), .A1(n821), .B0(destinationAddressIn_EAST[8]), 
        .B1(n798), .C0(n3962), .C1(n852), .Y(n5375) );
  AOI222XLTS U2654 ( .A0(n4267), .A1(n821), .B0(n4110), .B1(n798), .C0(n3956), 
        .C1(n853), .Y(n5377) );
  OAI221XLTS U2655 ( .A0(n269), .A1(n239), .B0(n4824), .B1(n329), .C0(n5376), 
        .Y(n2485) );
  AOI222XLTS U2656 ( .A0(n4270), .A1(n821), .B0(n4113), .B1(n800), .C0(n3959), 
        .C1(n853), .Y(n5376) );
  OAI2BB1X1TS U2657 ( .A0N(n4872), .A1N(selectBit_EAST), .B0(n4840), .Y(n4843)
         );
  INVX2TS U2658 ( .A(readReady), .Y(n6235) );
  NOR2X1TS U2659 ( .A(selectBit_WEST), .B(readReady), .Y(n4871) );
  NAND2X1TS U2660 ( .A(n4860), .B(n4859), .Y(n4869) );
  XNOR2X1TS U2661 ( .A(n194), .B(n6230), .Y(n4868) );
  OAI221XLTS U2662 ( .A0(n5583), .A1(n245), .B0(n4781), .B1(n565), .C0(n5466), 
        .Y(n2536) );
  AOI222XLTS U2663 ( .A0(n4285), .A1(n3430), .B0(n4130), .B1(n3392), .C0(n3974), .C1(n3683), .Y(n5466) );
  OAI221XLTS U2664 ( .A0(n328), .A1(n248), .B0(n4793), .B1(n566), .C0(n5468), 
        .Y(n2538) );
  AOI222XLTS U2665 ( .A0(n4279), .A1(n3430), .B0(n4124), .B1(n3392), .C0(n3968), .C1(n3682), .Y(n5468) );
  OAI221XLTS U2666 ( .A0(n327), .A1(n251), .B0(n4801), .B1(n566), .C0(n5469), 
        .Y(n2539) );
  AOI222XLTS U2667 ( .A0(n4276), .A1(n3438), .B0(n4121), .B1(n3402), .C0(n3965), .C1(n3682), .Y(n5469) );
  OAI221XLTS U2668 ( .A0(n328), .A1(n242), .B0(n4825), .B1(n567), .C0(n5472), 
        .Y(n2542) );
  AOI222XLTS U2669 ( .A0(n4267), .A1(n6202), .B0(n4112), .B1(n3406), .C0(n3956), .C1(n3683), .Y(n5472) );
  OAI221XLTS U2670 ( .A0(n327), .A1(n257), .B0(n4791), .B1(n565), .C0(n5467), 
        .Y(n2537) );
  AOI222XLTS U2671 ( .A0(n4282), .A1(n3430), .B0(n4127), .B1(n3404), .C0(n3971), .C1(n3683), .Y(n5467) );
  OAI221XLTS U2672 ( .A0(n328), .A1(n260), .B0(n4815), .B1(n566), .C0(n5470), 
        .Y(n2540) );
  AOI222XLTS U2673 ( .A0(n4273), .A1(n6202), .B0(n4118), .B1(n3405), .C0(n3962), .C1(n3682), .Y(n5470) );
  OAI221XLTS U2674 ( .A0(n327), .A1(n239), .B0(n4821), .B1(n566), .C0(n5471), 
        .Y(n2541) );
  AOI222XLTS U2675 ( .A0(n4270), .A1(n3432), .B0(n4115), .B1(n3403), .C0(n3959), .C1(n3682), .Y(n5471) );
  OAI221XLTS U2676 ( .A0(n263), .A1(n255), .B0(n4770), .B1(n772), .C0(n5348), 
        .Y(n2465) );
  AOI222XLTS U2677 ( .A0(n4132), .A1(n703), .B0(destinationAddressIn_SOUTH[13]), .B1(n735), .C0(n3977), .C1(n764), .Y(n5348) );
  OAI221XLTS U2678 ( .A0(n264), .A1(n246), .B0(n4778), .B1(n771), .C0(n5349), 
        .Y(n2466) );
  AOI222XLTS U2679 ( .A0(n4129), .A1(n704), .B0(destinationAddressIn_SOUTH[12]), .B1(n733), .C0(n3974), .C1(n762), .Y(n5349) );
  OAI221XLTS U2680 ( .A0(n5572), .A1(n258), .B0(n4788), .B1(n772), .C0(n5350), 
        .Y(n2467) );
  AOI222XLTS U2681 ( .A0(n4126), .A1(n704), .B0(destinationAddressIn_SOUTH[11]), .B1(n731), .C0(n3971), .C1(n762), .Y(n5350) );
  OAI221XLTS U2682 ( .A0(n264), .A1(n249), .B0(n4794), .B1(n772), .C0(n5351), 
        .Y(n2468) );
  AOI222XLTS U2683 ( .A0(n4123), .A1(n704), .B0(destinationAddressIn_SOUTH[10]), .B1(n734), .C0(n3968), .C1(n762), .Y(n5351) );
  OAI221XLTS U2684 ( .A0(n5572), .A1(n252), .B0(n4806), .B1(n773), .C0(n5352), 
        .Y(n2469) );
  AOI222XLTS U2685 ( .A0(n4120), .A1(n704), .B0(destinationAddressIn_SOUTH[9]), 
        .B1(n705), .C0(n3965), .C1(n762), .Y(n5352) );
  OAI221XLTS U2686 ( .A0(n264), .A1(n260), .B0(n4810), .B1(n773), .C0(n5353), 
        .Y(n2470) );
  AOI222XLTS U2687 ( .A0(n4117), .A1(n701), .B0(destinationAddressIn_SOUTH[8]), 
        .B1(n705), .C0(n3962), .C1(n766), .Y(n5353) );
  OAI221XLTS U2688 ( .A0(n5572), .A1(n6241), .B0(n4818), .B1(n773), .C0(n5354), 
        .Y(n2471) );
  AOI222XLTS U2689 ( .A0(n4114), .A1(n702), .B0(n4269), .B1(n705), .C0(n3959), 
        .C1(n764), .Y(n5354) );
  OAI221XLTS U2690 ( .A0(n264), .A1(n242), .B0(n4830), .B1(n772), .C0(n5355), 
        .Y(n2472) );
  AOI222XLTS U2691 ( .A0(n4111), .A1(n702), .B0(n4266), .B1(n705), .C0(n3956), 
        .C1(n763), .Y(n5355) );
  OAI221XLTS U2692 ( .A0(n263), .A1(n237), .B0(n770), .B1(n6286), .C0(n5571), 
        .Y(n2572) );
  AOI222XLTS U2693 ( .A0(n3809), .A1(n700), .B0(n3817), .B1(n706), .C0(n3804), 
        .C1(n767), .Y(n5571) );
  OAI221XLTS U2694 ( .A0(n328), .A1(n254), .B0(n4771), .B1(n565), .C0(n5465), 
        .Y(n2535) );
  AOI222XLTS U2695 ( .A0(n4288), .A1(n3433), .B0(n4133), .B1(n3404), .C0(n3977), .C1(n3683), .Y(n5465) );
  OAI221XLTS U2696 ( .A0(n327), .A1(n6239), .B0(n565), .B1(n106), .C0(n5582), 
        .Y(n2577) );
  AOI222XLTS U2697 ( .A0(n3816), .A1(n3436), .B0(n3810), .B1(n3406), .C0(n3804), .C1(n3688), .Y(n5582) );
  OAI221XLTS U2698 ( .A0(n1764), .A1(n236), .B0(n3223), .B1(n108), .C0(n5577), 
        .Y(n2574) );
  AOI222XLTS U2699 ( .A0(n3803), .A1(n3193), .B0(n3817), .B1(n232), .C0(n3810), 
        .C1(n413), .Y(n5577) );
  OAI221XLTS U2700 ( .A0(n266), .A1(n236), .B0(n3290), .B1(n107), .C0(n5578), 
        .Y(n2575) );
  OAI221XLTS U2701 ( .A0(n1654), .A1(n6245), .B0(n4787), .B1(n3222), .C0(n5398), .Y(n2495) );
  AOI222XLTS U2702 ( .A0(n3970), .A1(n1894), .B0(n4283), .B1(n285), .C0(n4127), 
        .C1(n5576), .Y(n5398) );
  OAI221XLTS U2703 ( .A0(n1764), .A1(n6240), .B0(n4827), .B1(n3222), .C0(n5403), .Y(n2500) );
  AOI222XLTS U2704 ( .A0(n3955), .A1(n3192), .B0(n4268), .B1(n233), .C0(n4112), 
        .C1(n413), .Y(n5403) );
  OAI221XLTS U2705 ( .A0(n267), .A1(n245), .B0(n4779), .B1(n3291), .C0(n5419), 
        .Y(n2508) );
  AOI222XLTS U2706 ( .A0(n4285), .A1(n3240), .B0(n3974), .B1(n3242), .C0(n4130), .C1(n3288), .Y(n5419) );
  OAI221XLTS U2707 ( .A0(n5579), .A1(n258), .B0(n4785), .B1(n3292), .C0(n5420), 
        .Y(n2509) );
  AOI222XLTS U2708 ( .A0(n4282), .A1(n3237), .B0(n3971), .B1(n3242), .C0(n4127), .C1(n6171), .Y(n5420) );
  OAI221XLTS U2709 ( .A0(n266), .A1(n248), .B0(n4795), .B1(n3292), .C0(n5421), 
        .Y(n2510) );
  AOI222XLTS U2710 ( .A0(n4279), .A1(n3239), .B0(n3968), .B1(n3242), .C0(n4124), .C1(n6171), .Y(n5421) );
  OAI221XLTS U2711 ( .A0(n267), .A1(n260), .B0(n4813), .B1(n3293), .C0(n5423), 
        .Y(n2512) );
  AOI222XLTS U2712 ( .A0(n4273), .A1(n3235), .B0(n3962), .B1(n3255), .C0(n4118), .C1(n3281), .Y(n5423) );
  OAI221XLTS U2713 ( .A0(n267), .A1(n239), .B0(n4817), .B1(n3293), .C0(n5424), 
        .Y(n2513) );
  AOI222XLTS U2714 ( .A0(n4270), .A1(n3235), .B0(n3959), .B1(n3253), .C0(n4115), .C1(n3281), .Y(n5424) );
  OAI221XLTS U2715 ( .A0(n266), .A1(n243), .B0(n4829), .B1(n3292), .C0(n5425), 
        .Y(n2514) );
  AOI222XLTS U2716 ( .A0(n4267), .A1(n3235), .B0(n3956), .B1(n3252), .C0(n4112), .C1(n3281), .Y(n5425) );
  OAI221XLTS U2717 ( .A0(n324), .A1(n251), .B0(n4805), .B1(n3507), .C0(n5494), 
        .Y(n2553) );
  AOI222XLTS U2718 ( .A0(n3964), .A1(n3455), .B0(n4277), .B1(n3457), .C0(n4121), .C1(n3497), .Y(n5494) );
  OAI221XLTS U2719 ( .A0(n1654), .A1(n246), .B0(n4780), .B1(n3219), .C0(n5397), 
        .Y(n2494) );
  OAI221XLTS U2720 ( .A0(n1728), .A1(n252), .B0(n4802), .B1(n3220), .C0(n5400), 
        .Y(n2497) );
  AOI222XLTS U2721 ( .A0(n3964), .A1(n3192), .B0(n4277), .B1(n233), .C0(n4121), 
        .C1(n414), .Y(n5400) );
  OAI221XLTS U2722 ( .A0(n1728), .A1(n261), .B0(n4816), .B1(n3221), .C0(n5401), 
        .Y(n2498) );
  AOI222XLTS U2723 ( .A0(n3961), .A1(n3192), .B0(n4274), .B1(n232), .C0(n4118), 
        .C1(n413), .Y(n5401) );
  OAI221XLTS U2724 ( .A0(n326), .A1(n6247), .B0(n4774), .B1(n3375), .C0(n5441), 
        .Y(n2521) );
  OAI221XLTS U2725 ( .A0(n325), .A1(n245), .B0(n4784), .B1(n3374), .C0(n5442), 
        .Y(n2522) );
  AOI222XLTS U2726 ( .A0(n3973), .A1(n3316), .B0(n4286), .B1(n3325), .C0(n4129), .C1(n3364), .Y(n5442) );
  OAI221XLTS U2727 ( .A0(n326), .A1(n257), .B0(n4790), .B1(n3375), .C0(n5443), 
        .Y(n2523) );
  AOI222XLTS U2728 ( .A0(n3970), .A1(n3316), .B0(n4283), .B1(n3325), .C0(n4126), .C1(n3364), .Y(n5443) );
  OAI221XLTS U2729 ( .A0(n325), .A1(n249), .B0(n4800), .B1(n3375), .C0(n5444), 
        .Y(n2524) );
  AOI222XLTS U2730 ( .A0(n3967), .A1(n3316), .B0(n4280), .B1(n3325), .C0(n4123), .C1(n3364), .Y(n5444) );
  OAI221XLTS U2731 ( .A0(n326), .A1(n251), .B0(n4804), .B1(n3376), .C0(n5445), 
        .Y(n2525) );
  AOI222XLTS U2732 ( .A0(n3964), .A1(n3316), .B0(n4277), .B1(n3326), .C0(n4120), .C1(n3364), .Y(n5445) );
  OAI221XLTS U2733 ( .A0(n325), .A1(n260), .B0(n4814), .B1(n3376), .C0(n5446), 
        .Y(n2526) );
  AOI222XLTS U2734 ( .A0(n3961), .A1(n3317), .B0(n4274), .B1(n3326), .C0(n4117), .C1(n3363), .Y(n5446) );
  OAI221XLTS U2735 ( .A0(n326), .A1(n240), .B0(n4820), .B1(n3376), .C0(n5447), 
        .Y(n2527) );
  AOI222XLTS U2736 ( .A0(n3958), .A1(n3324), .B0(n4271), .B1(n3326), .C0(n4114), .C1(n3363), .Y(n5447) );
  OAI221XLTS U2737 ( .A0(n325), .A1(n242), .B0(n4826), .B1(n3375), .C0(n5448), 
        .Y(n2528) );
  AOI222XLTS U2738 ( .A0(n3955), .A1(n3319), .B0(n4268), .B1(n3326), .C0(n4111), .C1(n3363), .Y(n5448) );
  OAI221XLTS U2739 ( .A0(n323), .A1(n255), .B0(n4772), .B1(n3506), .C0(n5490), 
        .Y(n2549) );
  AOI222XLTS U2740 ( .A0(n3976), .A1(n3454), .B0(n4289), .B1(n3456), .C0(n4133), .C1(n3501), .Y(n5490) );
  OAI221XLTS U2741 ( .A0(n324), .A1(n6246), .B0(n4782), .B1(n3505), .C0(n5491), 
        .Y(n2550) );
  AOI222XLTS U2742 ( .A0(n3973), .A1(n3450), .B0(n4286), .B1(n3456), .C0(n4130), .C1(n3497), .Y(n5491) );
  OAI221XLTS U2743 ( .A0(n323), .A1(n257), .B0(n4786), .B1(n3506), .C0(n5492), 
        .Y(n2551) );
  AOI222XLTS U2744 ( .A0(n3970), .A1(n6216), .B0(n4283), .B1(n3456), .C0(n4127), .C1(n3497), .Y(n5492) );
  OAI221XLTS U2745 ( .A0(n324), .A1(n248), .B0(n4796), .B1(n3506), .C0(n5493), 
        .Y(n2552) );
  AOI222XLTS U2746 ( .A0(n3967), .A1(n3450), .B0(n4280), .B1(n3456), .C0(n4124), .C1(n3497), .Y(n5493) );
  OAI221XLTS U2747 ( .A0(n323), .A1(n6242), .B0(n4812), .B1(n3507), .C0(n5495), 
        .Y(n2554) );
  AOI222XLTS U2748 ( .A0(n3961), .A1(n3448), .B0(n4274), .B1(n3457), .C0(n4118), .C1(n3496), .Y(n5495) );
  OAI221XLTS U2749 ( .A0(n324), .A1(n239), .B0(n4822), .B1(n3507), .C0(n5496), 
        .Y(n2555) );
  AOI222XLTS U2750 ( .A0(n3958), .A1(n3448), .B0(n4271), .B1(n3457), .C0(n4115), .C1(n3496), .Y(n5496) );
  OAI221XLTS U2751 ( .A0(n323), .A1(n242), .B0(n4828), .B1(n3506), .C0(n5497), 
        .Y(n2556) );
  AOI222XLTS U2752 ( .A0(n3955), .A1(n3448), .B0(n4268), .B1(n3457), .C0(n4112), .C1(n3496), .Y(n5497) );
  OAI221XLTS U2753 ( .A0(n1654), .A1(n254), .B0(n4773), .B1(n3219), .C0(n5396), 
        .Y(n2493) );
  AOI222XLTS U2754 ( .A0(n3976), .A1(n1894), .B0(n4289), .B1(n232), .C0(n4133), 
        .C1(n414), .Y(n5396) );
  OAI221XLTS U2755 ( .A0(n1728), .A1(n6244), .B0(n4799), .B1(n3220), .C0(n5399), .Y(n2496) );
  AOI222XLTS U2756 ( .A0(n3967), .A1(n1894), .B0(n4280), .B1(n232), .C0(n4124), 
        .C1(n414), .Y(n5399) );
  OAI221XLTS U2757 ( .A0(n1764), .A1(n6241), .B0(n4823), .B1(n3221), .C0(n5402), .Y(n2499) );
  AOI222XLTS U2758 ( .A0(n3958), .A1(n3192), .B0(n4271), .B1(n233), .C0(n4115), 
        .C1(n413), .Y(n5402) );
  OAI221XLTS U2759 ( .A0(n267), .A1(n254), .B0(n4775), .B1(n3292), .C0(n5418), 
        .Y(n2507) );
  AOI222XLTS U2760 ( .A0(n4288), .A1(n3241), .B0(n3977), .B1(n3242), .C0(n4133), .C1(n3285), .Y(n5418) );
  OAI221XLTS U2761 ( .A0(n5579), .A1(n6243), .B0(n4807), .B1(n3293), .C0(n5422), .Y(n2511) );
  AOI222XLTS U2762 ( .A0(n4276), .A1(n3237), .B0(n3965), .B1(n3254), .C0(n4121), .C1(n3282), .Y(n5422) );
  AOI22X1TS U2763 ( .A0(n3225), .A1(n4239), .B0(n3717), .B1(n4396), .Y(n6163)
         );
  AOI222XLTS U2764 ( .A0(n3287), .A1(n4084), .B0(n3265), .B1(n117), .C0(n6169), 
        .C1(n3928), .Y(n6162) );
  AOI22X1TS U2765 ( .A0(n3225), .A1(n4236), .B0(n3717), .B1(n4393), .Y(n6165)
         );
  AOI222XLTS U2766 ( .A0(n3287), .A1(n4081), .B0(n3265), .B1(n116), .C0(n3256), 
        .C1(n3925), .Y(n6164) );
  AOI22X1TS U2767 ( .A0(n3225), .A1(n4233), .B0(n3717), .B1(n4390), .Y(n6167)
         );
  AOI222XLTS U2768 ( .A0(n3286), .A1(n4078), .B0(n3265), .B1(n115), .C0(n3252), 
        .C1(n3922), .Y(n6166) );
  AOI22X1TS U2769 ( .A0(n3226), .A1(n4230), .B0(n3717), .B1(n4387), .Y(n6173)
         );
  AOI222XLTS U2770 ( .A0(n3286), .A1(n4075), .B0(n3266), .B1(n114), .C0(n3254), 
        .C1(n3919), .Y(n6172) );
  AOI22X1TS U2771 ( .A0(n3226), .A1(n4245), .B0(n3718), .B1(n4402), .Y(n6159)
         );
  AOI222XLTS U2772 ( .A0(n3285), .A1(n4090), .B0(n3266), .B1(n118), .C0(n3256), 
        .C1(n3934), .Y(n6158) );
  AOI22X1TS U2773 ( .A0(n3225), .A1(n4242), .B0(n3718), .B1(n4399), .Y(n6161)
         );
  AOI222XLTS U2774 ( .A0(n3285), .A1(n4087), .B0(n3266), .B1(n141), .C0(n3257), 
        .C1(n3931), .Y(n6160) );
  AOI22X1TS U2775 ( .A0(n3309), .A1(n3933), .B0(n3704), .B1(n4402), .Y(n6175)
         );
  AOI222XLTS U2776 ( .A0(n3357), .A1(n4090), .B0(n3347), .B1(n146), .C0(n3338), 
        .C1(n4246), .Y(n6174) );
  AOI22X1TS U2777 ( .A0(n3308), .A1(n3930), .B0(n3704), .B1(n4399), .Y(n6177)
         );
  AOI222XLTS U2778 ( .A0(n3356), .A1(n4087), .B0(n3347), .B1(n142), .C0(n3340), 
        .C1(n4243), .Y(n6176) );
  AOI22X1TS U2779 ( .A0(n3308), .A1(n3927), .B0(n3703), .B1(n4396), .Y(n6179)
         );
  AOI222XLTS U2780 ( .A0(n3356), .A1(n4084), .B0(n3346), .B1(n137), .C0(n3327), 
        .C1(n4240), .Y(n6178) );
  AOI22X1TS U2781 ( .A0(n3308), .A1(n3924), .B0(n3703), .B1(n4393), .Y(n6181)
         );
  AOI222XLTS U2782 ( .A0(n3356), .A1(n4081), .B0(n3346), .B1(n133), .C0(n3327), 
        .C1(n4237), .Y(n6180) );
  AOI22X1TS U2783 ( .A0(n3308), .A1(n3921), .B0(n3703), .B1(n4390), .Y(n6183)
         );
  AOI222XLTS U2784 ( .A0(n3356), .A1(n4078), .B0(n3346), .B1(n129), .C0(n3327), 
        .C1(n4234), .Y(n6182) );
  AOI22X1TS U2785 ( .A0(n3309), .A1(n3918), .B0(n3703), .B1(n4387), .Y(n6189)
         );
  AOI222XLTS U2786 ( .A0(n3357), .A1(n4075), .B0(n3347), .B1(n125), .C0(n3339), 
        .C1(n4231), .Y(n6188) );
  AOI22X1TS U2787 ( .A0(n859), .A1(n145), .B0(n214), .B1(n4245), .Y(n6145) );
  AOI222XLTS U2788 ( .A0(\requesterAddressbuffer[3][5] ), .A1(n3217), .B0(
        n3201), .B1(n3934), .C0(n886), .C1(n4403), .Y(n6144) );
  AOI22X1TS U2789 ( .A0(n859), .A1(n140), .B0(n211), .B1(n4242), .Y(n6147) );
  AOI222XLTS U2790 ( .A0(\requesterAddressbuffer[3][4] ), .A1(n3217), .B0(
        n3207), .B1(n3931), .C0(n886), .C1(n4400), .Y(n6146) );
  AOI22X1TS U2791 ( .A0(n859), .A1(n136), .B0(n209), .B1(n4239), .Y(n6149) );
  AOI222XLTS U2792 ( .A0(\requesterAddressbuffer[3][3] ), .A1(n3218), .B0(
        n3207), .B1(n3928), .C0(n871), .C1(n4397), .Y(n6148) );
  AOI22X1TS U2793 ( .A0(n858), .A1(n132), .B0(n218), .B1(n4236), .Y(n6151) );
  AOI222XLTS U2794 ( .A0(\requesterAddressbuffer[3][2] ), .A1(n3218), .B0(
        n3203), .B1(n3925), .C0(n871), .C1(n4394), .Y(n6150) );
  AOI22X1TS U2795 ( .A0(n857), .A1(n128), .B0(n213), .B1(n4233), .Y(n6153) );
  AOI222XLTS U2796 ( .A0(\requesterAddressbuffer[3][1] ), .A1(n3218), .B0(
        n3204), .B1(n3922), .C0(n871), .C1(n4391), .Y(n6152) );
  AOI22X1TS U2797 ( .A0(n859), .A1(n124), .B0(n219), .B1(n4230), .Y(n6157) );
  AOI222XLTS U2798 ( .A0(\requesterAddressbuffer[3][0] ), .A1(n3218), .B0(
        n6155), .B1(n3919), .C0(n871), .C1(n4388), .Y(n6156) );
  AOI22X1TS U2799 ( .A0(n689), .A1(n4089), .B0(n3762), .B1(n4402), .Y(n6114)
         );
  AOI222XLTS U2800 ( .A0(n754), .A1(n3933), .B0(n745), .B1(n144), .C0(n707), 
        .C1(n4246), .Y(n6113) );
  AOI22X1TS U2801 ( .A0(n688), .A1(n4086), .B0(n3762), .B1(n4399), .Y(n6116)
         );
  AOI222XLTS U2802 ( .A0(n753), .A1(n3930), .B0(n752), .B1(n139), .C0(n707), 
        .C1(n4243), .Y(n6115) );
  AOI22X1TS U2803 ( .A0(n688), .A1(n4083), .B0(n3761), .B1(n4396), .Y(n6118)
         );
  AOI222XLTS U2804 ( .A0(n753), .A1(n3927), .B0(n746), .B1(n135), .C0(n706), 
        .C1(n4240), .Y(n6117) );
  AOI22X1TS U2805 ( .A0(n688), .A1(n4080), .B0(n3761), .B1(n4393), .Y(n6120)
         );
  AOI222XLTS U2806 ( .A0(n753), .A1(n3924), .B0(n748), .B1(n131), .C0(n706), 
        .C1(n4237), .Y(n6119) );
  AOI22X1TS U2807 ( .A0(n688), .A1(n4077), .B0(n3761), .B1(n4390), .Y(n6122)
         );
  AOI222XLTS U2808 ( .A0(n753), .A1(n3921), .B0(n746), .B1(n127), .C0(n706), 
        .C1(n4234), .Y(n6121) );
  AOI22X1TS U2809 ( .A0(n689), .A1(n4074), .B0(n3761), .B1(n4387), .Y(n6128)
         );
  AOI222XLTS U2810 ( .A0(n754), .A1(n3918), .B0(n750), .B1(n123), .C0(n707), 
        .C1(n4231), .Y(n6127) );
  AOI222XLTS U2811 ( .A0(\requesterAddressbuffer[6][5] ), .A1(n578), .B0(n3430), .B1(n4245), .C0(n3702), .C1(n4403), .Y(n6190) );
  AOI22X1TS U2812 ( .A0(n3409), .A1(n141), .B0(n3391), .B1(n4086), .Y(n6193)
         );
  AOI222XLTS U2813 ( .A0(\requesterAddressbuffer[6][4] ), .A1(n577), .B0(n3431), .B1(n4242), .C0(n3699), .C1(n4400), .Y(n6192) );
  AOI22X1TS U2814 ( .A0(n3408), .A1(n133), .B0(n3391), .B1(n4080), .Y(n6197)
         );
  AOI222XLTS U2815 ( .A0(\requesterAddressbuffer[6][2] ), .A1(n581), .B0(n3431), .B1(n4236), .C0(n3697), .C1(n4394), .Y(n6196) );
  AOI22X1TS U2816 ( .A0(n4263), .A1(n3428), .B0(n4420), .B1(n3689), .Y(n5475)
         );
  AOI222XLTS U2817 ( .A0(n3951), .A1(n3688), .B0(n3416), .B1(n144), .C0(n4108), 
        .C1(n6200), .Y(n5474) );
  AOI22X1TS U2818 ( .A0(n4257), .A1(n3435), .B0(n4414), .B1(n3689), .Y(n5479)
         );
  AOI222XLTS U2819 ( .A0(n3945), .A1(n3686), .B0(n3416), .B1(n135), .C0(n4102), 
        .C1(n3401), .Y(n5478) );
  AOI22X1TS U2820 ( .A0(n4254), .A1(n3434), .B0(n4411), .B1(n3689), .Y(n5481)
         );
  AOI222XLTS U2821 ( .A0(n3942), .A1(n3685), .B0(n3418), .B1(n131), .C0(n4099), 
        .C1(n3401), .Y(n5480) );
  AOI22X1TS U2822 ( .A0(n4251), .A1(n3433), .B0(n4408), .B1(n3700), .Y(n5483)
         );
  AOI222XLTS U2823 ( .A0(n3939), .A1(n3684), .B0(n6201), .B1(n127), .C0(n4096), 
        .C1(n3401), .Y(n5482) );
  AOI22X1TS U2824 ( .A0(n4248), .A1(n3435), .B0(n4405), .B1(n3699), .Y(n5485)
         );
  AOI222XLTS U2825 ( .A0(n3936), .A1(n3686), .B0(n3417), .B1(n123), .C0(n4093), 
        .C1(n3401), .Y(n5484) );
  AOI22X1TS U2826 ( .A0(n4221), .A1(n3429), .B0(n4378), .B1(n3690), .Y(n5655)
         );
  AOI22X1TS U2827 ( .A0(n4203), .A1(n3427), .B0(n4360), .B1(n3691), .Y(n5667)
         );
  AOI22X1TS U2828 ( .A0(n4197), .A1(n3427), .B0(n4354), .B1(n3692), .Y(n5671)
         );
  AOI22X1TS U2829 ( .A0(n4194), .A1(n3427), .B0(n4351), .B1(n3692), .Y(n5673)
         );
  AOI22X1TS U2830 ( .A0(n4173), .A1(n3425), .B0(n4330), .B1(n3694), .Y(n5687)
         );
  AOI22X1TS U2831 ( .A0(n4170), .A1(n3425), .B0(n4327), .B1(n3694), .Y(n5689)
         );
  AOI22X1TS U2832 ( .A0(n4164), .A1(n3424), .B0(n4321), .B1(n3694), .Y(n5693)
         );
  AOI22X1TS U2833 ( .A0(n4152), .A1(n3423), .B0(n4309), .B1(n3695), .Y(n5701)
         );
  AOI22X1TS U2834 ( .A0(n3948), .A1(n3447), .B0(n4417), .B1(n3660), .Y(n5503)
         );
  AOI222XLTS U2835 ( .A0(n4105), .A1(n3495), .B0(n142), .B1(n3483), .C0(n4261), 
        .C1(n3467), .Y(n5502) );
  AOI22X1TS U2836 ( .A0(n3936), .A1(n3451), .B0(n4405), .B1(n3661), .Y(n5511)
         );
  AOI222XLTS U2837 ( .A0(n4093), .A1(n3494), .B0(n125), .B1(n3473), .C0(n4249), 
        .C1(n3465), .Y(n5510) );
  AOI22X1TS U2838 ( .A0(n4227), .A1(n3434), .B0(n4384), .B1(n3702), .Y(n5651)
         );
  AOI22X1TS U2839 ( .A0(n4224), .A1(n3429), .B0(n4381), .B1(n3701), .Y(n5653)
         );
  AOI22X1TS U2840 ( .A0(n4218), .A1(n3429), .B0(n4375), .B1(n3690), .Y(n5657)
         );
  AOI22X1TS U2841 ( .A0(n4215), .A1(n3429), .B0(n4372), .B1(n3690), .Y(n5659)
         );
  AOI22X1TS U2842 ( .A0(n4212), .A1(n3428), .B0(n4369), .B1(n3690), .Y(n5661)
         );
  AOI22X1TS U2843 ( .A0(n4206), .A1(n3428), .B0(n4363), .B1(n3691), .Y(n5665)
         );
  AOI22X1TS U2844 ( .A0(n4200), .A1(n3427), .B0(n4357), .B1(n3691), .Y(n5669)
         );
  AOI22X1TS U2845 ( .A0(n4191), .A1(n3426), .B0(n4348), .B1(n3692), .Y(n5675)
         );
  AOI22X1TS U2846 ( .A0(n4185), .A1(n3426), .B0(n4342), .B1(n3693), .Y(n5679)
         );
  AOI22X1TS U2847 ( .A0(n4182), .A1(n3426), .B0(n4339), .B1(n3693), .Y(n5681)
         );
  AOI22X1TS U2848 ( .A0(n4179), .A1(n3425), .B0(n4336), .B1(n3693), .Y(n5683)
         );
  AOI22X1TS U2849 ( .A0(n4176), .A1(n3425), .B0(n4333), .B1(n3693), .Y(n5685)
         );
  AOI22X1TS U2850 ( .A0(n4167), .A1(n3424), .B0(n4324), .B1(n3694), .Y(n5691)
         );
  AOI22X1TS U2851 ( .A0(n4161), .A1(n3424), .B0(n4318), .B1(n3695), .Y(n5695)
         );
  AOI22X1TS U2852 ( .A0(n4158), .A1(n3424), .B0(n4315), .B1(n3695), .Y(n5697)
         );
  AOI22X1TS U2853 ( .A0(n4155), .A1(n3423), .B0(n4312), .B1(n3695), .Y(n5699)
         );
  AOI22X1TS U2854 ( .A0(n4149), .A1(n3423), .B0(n4306), .B1(n3696), .Y(n5703)
         );
  AOI22X1TS U2855 ( .A0(n4143), .A1(n3422), .B0(n4300), .B1(n3696), .Y(n5707)
         );
  AOI22X1TS U2856 ( .A0(n4140), .A1(n3422), .B0(n4297), .B1(n3696), .Y(n5709)
         );
  AOI22X1TS U2857 ( .A0(n3951), .A1(n3447), .B0(n4420), .B1(n3660), .Y(n5501)
         );
  AOI222XLTS U2858 ( .A0(n4108), .A1(n3495), .B0(n145), .B1(n3485), .C0(n4264), 
        .C1(n3458), .Y(n5500) );
  AOI22X1TS U2859 ( .A0(n3945), .A1(n3447), .B0(n4414), .B1(n3660), .Y(n5505)
         );
  AOI222XLTS U2860 ( .A0(n4102), .A1(n3495), .B0(n137), .B1(n3483), .C0(n4258), 
        .C1(n3465), .Y(n5504) );
  AOI22X1TS U2861 ( .A0(n3942), .A1(n3447), .B0(n4411), .B1(n3660), .Y(n5507)
         );
  AOI222XLTS U2862 ( .A0(n4099), .A1(n3495), .B0(n133), .B1(n3485), .C0(n4255), 
        .C1(n3465), .Y(n5506) );
  AOI22X1TS U2863 ( .A0(n3939), .A1(n3453), .B0(n4408), .B1(n3661), .Y(n5509)
         );
  AOI222XLTS U2864 ( .A0(n4096), .A1(n3494), .B0(n129), .B1(n3473), .C0(n4252), 
        .C1(n3465), .Y(n5508) );
  AOI22X1TS U2865 ( .A0(n3915), .A1(n6216), .B0(n4385), .B1(n3661), .Y(n5587)
         );
  AOI22X1TS U2866 ( .A0(n3912), .A1(n3455), .B0(n4382), .B1(n3661), .Y(n5589)
         );
  AOI22X1TS U2867 ( .A0(n3909), .A1(n3452), .B0(n4379), .B1(n3662), .Y(n5591)
         );
  AOI22X1TS U2868 ( .A0(n3906), .A1(n3451), .B0(n4376), .B1(n3662), .Y(n5593)
         );
  AOI22X1TS U2869 ( .A0(n3903), .A1(n3453), .B0(n4373), .B1(n3662), .Y(n5595)
         );
  AOI22X1TS U2870 ( .A0(n3900), .A1(n3452), .B0(n4370), .B1(n3662), .Y(n5597)
         );
  AOI22X1TS U2871 ( .A0(n3897), .A1(n3446), .B0(n4367), .B1(n3672), .Y(n5599)
         );
  AOI22X1TS U2872 ( .A0(n3894), .A1(n3446), .B0(n4364), .B1(n3669), .Y(n5601)
         );
  AOI22X1TS U2873 ( .A0(n3891), .A1(n3446), .B0(n4361), .B1(n6339), .Y(n5603)
         );
  AOI22X1TS U2874 ( .A0(n3888), .A1(n3446), .B0(n4358), .B1(n3670), .Y(n5605)
         );
  AOI22X1TS U2875 ( .A0(n3885), .A1(n3445), .B0(n4355), .B1(n3663), .Y(n5607)
         );
  AOI22X1TS U2876 ( .A0(n3882), .A1(n3445), .B0(n4352), .B1(n3663), .Y(n5609)
         );
  AOI22X1TS U2877 ( .A0(n3879), .A1(n3445), .B0(n4349), .B1(n3663), .Y(n5611)
         );
  AOI22X1TS U2878 ( .A0(n3876), .A1(n3444), .B0(n4346), .B1(n3663), .Y(n5613)
         );
  AOI22X1TS U2879 ( .A0(n3873), .A1(n3444), .B0(n4343), .B1(n3664), .Y(n5615)
         );
  AOI22X1TS U2880 ( .A0(n3870), .A1(n3444), .B0(n4340), .B1(n3664), .Y(n5617)
         );
  AOI22X1TS U2881 ( .A0(n3867), .A1(n3444), .B0(n4337), .B1(n3664), .Y(n5619)
         );
  AOI22X1TS U2882 ( .A0(n3864), .A1(n3443), .B0(n4334), .B1(n3664), .Y(n5621)
         );
  AOI22X1TS U2883 ( .A0(n3861), .A1(n3443), .B0(n4331), .B1(n3670), .Y(n5623)
         );
  AOI22X1TS U2884 ( .A0(n3858), .A1(n3443), .B0(n4328), .B1(n3672), .Y(n5625)
         );
  AOI22X1TS U2885 ( .A0(n3855), .A1(n3443), .B0(n4325), .B1(n3671), .Y(n5627)
         );
  AOI22X1TS U2886 ( .A0(n3852), .A1(n3442), .B0(n4322), .B1(n3669), .Y(n5629)
         );
  AOI22X1TS U2887 ( .A0(n3849), .A1(n3442), .B0(n4319), .B1(n3665), .Y(n5631)
         );
  AOI22X1TS U2888 ( .A0(n3846), .A1(n3442), .B0(n4316), .B1(n3665), .Y(n5633)
         );
  AOI22X1TS U2889 ( .A0(n3843), .A1(n3442), .B0(n4313), .B1(n3665), .Y(n5635)
         );
  AOI22X1TS U2890 ( .A0(n3840), .A1(n3441), .B0(n4310), .B1(n3665), .Y(n5637)
         );
  AOI22X1TS U2891 ( .A0(n3837), .A1(n3441), .B0(n4307), .B1(n3666), .Y(n5639)
         );
  AOI22X1TS U2892 ( .A0(n3834), .A1(n3441), .B0(n4304), .B1(n3666), .Y(n5641)
         );
  AOI22X1TS U2893 ( .A0(n3831), .A1(n3441), .B0(n4301), .B1(n3666), .Y(n5643)
         );
  AOI22X1TS U2894 ( .A0(n3828), .A1(n3440), .B0(n4298), .B1(n3666), .Y(n5645)
         );
  AOI22X1TS U2895 ( .A0(n3825), .A1(n3440), .B0(n4295), .B1(n3667), .Y(n5647)
         );
  AOI22X1TS U2896 ( .A0(n3822), .A1(n3440), .B0(n4292), .B1(n3667), .Y(n5649)
         );
  AOI22X1TS U2897 ( .A0(n4260), .A1(n3436), .B0(n4417), .B1(n3689), .Y(n5477)
         );
  AOI222XLTS U2898 ( .A0(n3948), .A1(n6340), .B0(n6201), .B1(
        readRequesterAddress[4]), .C0(n4105), .C1(n3403), .Y(n5476) );
  AOI22X1TS U2899 ( .A0(n4209), .A1(n3428), .B0(n4366), .B1(n3691), .Y(n5663)
         );
  AOI22X1TS U2900 ( .A0(n4188), .A1(n3426), .B0(n4345), .B1(n3692), .Y(n5677)
         );
  AOI22X1TS U2901 ( .A0(n4146), .A1(n3423), .B0(n4303), .B1(n3696), .Y(n5705)
         );
  AOI22X1TS U2902 ( .A0(n4059), .A1(n696), .B0(n4372), .B1(n3768), .Y(n5979)
         );
  AOI22X1TS U2903 ( .A0(n4044), .A1(n695), .B0(n4357), .B1(n3772), .Y(n5989)
         );
  AOI22X1TS U2904 ( .A0(n4038), .A1(n694), .B0(n4351), .B1(n3767), .Y(n5993)
         );
  AOI22X1TS U2905 ( .A0(n4035), .A1(n694), .B0(n4348), .B1(n3767), .Y(n5995)
         );
  AOI22X1TS U2906 ( .A0(n4008), .A1(n691), .B0(n4321), .B1(n3765), .Y(n6013)
         );
  AOI22X1TS U2907 ( .A0(n4002), .A1(n691), .B0(n4315), .B1(n3764), .Y(n6017)
         );
  AOI22X1TS U2908 ( .A0(n3993), .A1(n690), .B0(n4306), .B1(n3763), .Y(n6023)
         );
  AOI22X1TS U2909 ( .A0(n3984), .A1(n690), .B0(n4297), .B1(n3763), .Y(n6029)
         );
  AOI22X1TS U2910 ( .A0(n4263), .A1(n3234), .B0(n4421), .B1(n3725), .Y(n5427)
         );
  AOI222XLTS U2911 ( .A0(n4107), .A1(n3280), .B0(n3265), .B1(n145), .C0(n3952), 
        .C1(n3253), .Y(n5426) );
  AOI22X1TS U2912 ( .A0(n4260), .A1(n3234), .B0(n4418), .B1(n3725), .Y(n5429)
         );
  AOI222XLTS U2913 ( .A0(n4104), .A1(n3280), .B0(n3267), .B1(n139), .C0(n3949), 
        .C1(n3258), .Y(n5428) );
  AOI22X1TS U2914 ( .A0(n4257), .A1(n3234), .B0(n4415), .B1(n3725), .Y(n5431)
         );
  AOI222XLTS U2915 ( .A0(n4101), .A1(n3280), .B0(n3267), .B1(n136), .C0(n3946), 
        .C1(n3251), .Y(n5430) );
  AOI22X1TS U2916 ( .A0(n4254), .A1(n3234), .B0(n4412), .B1(n3725), .Y(n5433)
         );
  AOI222XLTS U2917 ( .A0(n4098), .A1(n3280), .B0(n3267), .B1(n132), .C0(n3943), 
        .C1(n3251), .Y(n5432) );
  AOI22X1TS U2918 ( .A0(n4251), .A1(n3240), .B0(n4409), .B1(n3729), .Y(n5435)
         );
  AOI222XLTS U2919 ( .A0(n4095), .A1(n3279), .B0(n3267), .B1(n128), .C0(n3940), 
        .C1(n3251), .Y(n5434) );
  AOI22X1TS U2920 ( .A0(n4248), .A1(n3238), .B0(n4406), .B1(n3726), .Y(n5437)
         );
  AOI222XLTS U2921 ( .A0(n4092), .A1(n3279), .B0(n3266), .B1(n124), .C0(n3937), 
        .C1(n3251), .Y(n5436) );
  AOI22X1TS U2922 ( .A0(n4224), .A1(n3238), .B0(n4381), .B1(n3727), .Y(n5781)
         );
  AOI222XLTS U2923 ( .A0(n4068), .A1(n3279), .B0(cacheDataOut[30]), .B1(n3259), 
        .C0(n3913), .C1(n3250), .Y(n5780) );
  AOI22X1TS U2924 ( .A0(n4218), .A1(n3233), .B0(n4375), .B1(n3724), .Y(n5785)
         );
  AOI222XLTS U2925 ( .A0(n4062), .A1(n3278), .B0(cacheDataOut[28]), .B1(n3259), 
        .C0(n3907), .C1(n3250), .Y(n5784) );
  AOI22X1TS U2926 ( .A0(n4215), .A1(n3233), .B0(n4372), .B1(n3724), .Y(n5787)
         );
  AOI222XLTS U2927 ( .A0(n4059), .A1(n3278), .B0(cacheDataOut[27]), .B1(n3259), 
        .C0(n3904), .C1(n3249), .Y(n5786) );
  AOI22X1TS U2928 ( .A0(n4212), .A1(n3233), .B0(n4369), .B1(n3724), .Y(n5789)
         );
  AOI222XLTS U2929 ( .A0(n4056), .A1(n3278), .B0(cacheDataOut[26]), .B1(n3261), 
        .C0(n3901), .C1(n3249), .Y(n5788) );
  AOI22X1TS U2930 ( .A0(n4209), .A1(n3232), .B0(n4366), .B1(n3726), .Y(n5791)
         );
  AOI222XLTS U2931 ( .A0(n4053), .A1(n3277), .B0(cacheDataOut[25]), .B1(n3261), 
        .C0(n3898), .C1(n3249), .Y(n5790) );
  AOI22X1TS U2932 ( .A0(n4206), .A1(n3232), .B0(n4363), .B1(n3726), .Y(n5793)
         );
  AOI222XLTS U2933 ( .A0(n4050), .A1(n3277), .B0(cacheDataOut[24]), .B1(n3260), 
        .C0(n3895), .C1(n3249), .Y(n5792) );
  AOI22X1TS U2934 ( .A0(n4203), .A1(n3232), .B0(n4360), .B1(n3729), .Y(n5795)
         );
  AOI222XLTS U2935 ( .A0(n4047), .A1(n3277), .B0(cacheDataOut[23]), .B1(n3268), 
        .C0(n3892), .C1(n3248), .Y(n5794) );
  AOI22X1TS U2936 ( .A0(n4188), .A1(n3230), .B0(n4345), .B1(n3723), .Y(n5805)
         );
  AOI222XLTS U2937 ( .A0(n4032), .A1(n3283), .B0(cacheDataOut[18]), .B1(n3261), 
        .C0(n3877), .C1(n3247), .Y(n5804) );
  AOI22X1TS U2938 ( .A0(n4173), .A1(n3229), .B0(n4330), .B1(n3721), .Y(n5815)
         );
  AOI222XLTS U2939 ( .A0(n4017), .A1(n3275), .B0(cacheDataOut[13]), .B1(n3262), 
        .C0(n3862), .C1(n3246), .Y(n5814) );
  AOI22X1TS U2940 ( .A0(n4161), .A1(n3231), .B0(n4318), .B1(n3720), .Y(n5823)
         );
  AOI222XLTS U2941 ( .A0(n4005), .A1(n3276), .B0(cacheDataOut[9]), .B1(n3262), 
        .C0(n3850), .C1(n3245), .Y(n5822) );
  AOI22X1TS U2942 ( .A0(n4155), .A1(n3228), .B0(n4312), .B1(n3720), .Y(n5827)
         );
  AOI222XLTS U2943 ( .A0(n3999), .A1(n3274), .B0(cacheDataOut[7]), .B1(n3262), 
        .C0(n3844), .C1(n3244), .Y(n5826) );
  AOI22X1TS U2944 ( .A0(n4149), .A1(n3227), .B0(n4306), .B1(n3719), .Y(n5831)
         );
  AOI222XLTS U2945 ( .A0(n3993), .A1(n3273), .B0(cacheDataOut[5]), .B1(n3264), 
        .C0(n3838), .C1(n3244), .Y(n5830) );
  AOI22X1TS U2946 ( .A0(n4146), .A1(n3227), .B0(n4303), .B1(n3719), .Y(n5833)
         );
  AOI222XLTS U2947 ( .A0(n3990), .A1(n3273), .B0(cacheDataOut[4]), .B1(n3264), 
        .C0(n3835), .C1(n3244), .Y(n5832) );
  AOI22X1TS U2948 ( .A0(n4140), .A1(n3227), .B0(n4297), .B1(n3719), .Y(n5837)
         );
  AOI222XLTS U2949 ( .A0(n3984), .A1(n3273), .B0(cacheDataOut[2]), .B1(n3264), 
        .C0(n3829), .C1(n3243), .Y(n5836) );
  AOI22X1TS U2950 ( .A0(n3915), .A1(n3318), .B0(n4384), .B1(n3714), .Y(n5715)
         );
  AOI22X1TS U2951 ( .A0(n3870), .A1(n3313), .B0(n4339), .B1(n3714), .Y(n5745)
         );
  AOI22X1TS U2952 ( .A0(n3867), .A1(n3313), .B0(n4336), .B1(n3711), .Y(n5747)
         );
  AOI22X1TS U2953 ( .A0(n3855), .A1(n3312), .B0(n4324), .B1(n3707), .Y(n5755)
         );
  AOI22X1TS U2954 ( .A0(n3825), .A1(n3309), .B0(n4294), .B1(n3704), .Y(n5775)
         );
  AOI22X1TS U2955 ( .A0(n4107), .A1(n699), .B0(n4420), .B1(n3768), .Y(n5358)
         );
  AOI222XLTS U2956 ( .A0(n3952), .A1(n763), .B0(n748), .B1(n118), .C0(n4264), 
        .C1(n707), .Y(n5357) );
  OAI211X1TS U2957 ( .A0(n4726), .A1(n784), .B0(n5360), .C0(n5359), .Y(n2474)
         );
  INVX2TS U2958 ( .A(n429), .Y(n784) );
  AOI22X1TS U2959 ( .A0(n4104), .A1(n698), .B0(n4417), .B1(n3768), .Y(n5360)
         );
  AOI222XLTS U2960 ( .A0(n3949), .A1(n763), .B0(n745), .B1(
        readRequesterAddress[4]), .C0(n4261), .C1(n737), .Y(n5359) );
  AOI22X1TS U2961 ( .A0(n4101), .A1(n698), .B0(n4414), .B1(n3771), .Y(n5362)
         );
  AOI222XLTS U2962 ( .A0(n3946), .A1(n763), .B0(n745), .B1(n117), .C0(n4258), 
        .C1(n729), .Y(n5361) );
  AOI22X1TS U2963 ( .A0(n4098), .A1(n699), .B0(n4411), .B1(n3774), .Y(n5364)
         );
  AOI222XLTS U2964 ( .A0(n3943), .A1(n766), .B0(n745), .B1(n116), .C0(n4255), 
        .C1(n729), .Y(n5363) );
  AOI22X1TS U2965 ( .A0(n4095), .A1(n697), .B0(n4408), .B1(n3773), .Y(n5366)
         );
  AOI222XLTS U2966 ( .A0(n3940), .A1(n765), .B0(n749), .B1(n115), .C0(n4252), 
        .C1(n729), .Y(n5365) );
  AOI22X1TS U2967 ( .A0(n4092), .A1(n697), .B0(n4405), .B1(n3768), .Y(n5368)
         );
  AOI222XLTS U2968 ( .A0(n3937), .A1(n767), .B0(n750), .B1(n114), .C0(n4249), 
        .C1(n729), .Y(n5367) );
  AOI22X1TS U2969 ( .A0(n4071), .A1(n697), .B0(n4384), .B1(n3770), .Y(n5971)
         );
  AOI22X1TS U2970 ( .A0(n4068), .A1(n697), .B0(n4381), .B1(n3772), .Y(n5973)
         );
  AOI22X1TS U2971 ( .A0(n4065), .A1(n696), .B0(n4378), .B1(n3771), .Y(n5975)
         );
  AOI22X1TS U2972 ( .A0(n4062), .A1(n696), .B0(n4375), .B1(n3769), .Y(n5977)
         );
  AOI22X1TS U2973 ( .A0(n4056), .A1(n696), .B0(n4369), .B1(n3770), .Y(n5981)
         );
  AOI22X1TS U2974 ( .A0(n4053), .A1(n695), .B0(n4366), .B1(n3769), .Y(n5983)
         );
  AOI22X1TS U2975 ( .A0(n4050), .A1(n695), .B0(n4363), .B1(n3772), .Y(n5985)
         );
  AOI22X1TS U2976 ( .A0(n4047), .A1(n695), .B0(n4360), .B1(n3774), .Y(n5987)
         );
  AOI22X1TS U2977 ( .A0(n4041), .A1(n694), .B0(n4354), .B1(n3767), .Y(n5991)
         );
  AOI22X1TS U2978 ( .A0(n4032), .A1(n693), .B0(n4345), .B1(n3767), .Y(n5997)
         );
  AOI22X1TS U2979 ( .A0(n4029), .A1(n693), .B0(n4342), .B1(n3766), .Y(n5999)
         );
  AOI22X1TS U2980 ( .A0(n4026), .A1(n693), .B0(n4339), .B1(n3766), .Y(n6001)
         );
  AOI22X1TS U2981 ( .A0(n4023), .A1(n693), .B0(n4336), .B1(n3766), .Y(n6003)
         );
  AOI22X1TS U2982 ( .A0(n4020), .A1(n692), .B0(n4333), .B1(n3766), .Y(n6005)
         );
  AOI22X1TS U2983 ( .A0(n4017), .A1(n692), .B0(n4330), .B1(n3765), .Y(n6007)
         );
  AOI22X1TS U2984 ( .A0(n4014), .A1(n692), .B0(n4327), .B1(n3765), .Y(n6009)
         );
  AOI22X1TS U2985 ( .A0(n4011), .A1(n692), .B0(n4324), .B1(n3765), .Y(n6011)
         );
  AOI22X1TS U2986 ( .A0(n4005), .A1(n694), .B0(n4318), .B1(n3764), .Y(n6015)
         );
  AOI22X1TS U2987 ( .A0(n3999), .A1(n691), .B0(n4312), .B1(n3764), .Y(n6019)
         );
  AOI22X1TS U2988 ( .A0(n3996), .A1(n691), .B0(n4309), .B1(n3764), .Y(n6021)
         );
  AOI22X1TS U2989 ( .A0(n3990), .A1(n690), .B0(n4303), .B1(n3763), .Y(n6025)
         );
  AOI22X1TS U2990 ( .A0(n3987), .A1(n690), .B0(n4300), .B1(n3763), .Y(n6027)
         );
  AOI22X1TS U2991 ( .A0(n3981), .A1(n689), .B0(n4294), .B1(n3762), .Y(n6031)
         );
  AOI22X1TS U2992 ( .A0(n4227), .A1(n3239), .B0(n4384), .B1(n3727), .Y(n5779)
         );
  AOI222XLTS U2993 ( .A0(n4071), .A1(n3279), .B0(cacheDataOut[31]), .B1(n3260), 
        .C0(n3916), .C1(n3250), .Y(n5778) );
  AOI22X1TS U2994 ( .A0(n4221), .A1(n3233), .B0(n4378), .B1(n3724), .Y(n5783)
         );
  AOI222XLTS U2995 ( .A0(n4065), .A1(n3278), .B0(cacheDataOut[29]), .B1(n3260), 
        .C0(n3910), .C1(n3250), .Y(n5782) );
  AOI22X1TS U2996 ( .A0(n4200), .A1(n3232), .B0(n4357), .B1(n3730), .Y(n5797)
         );
  AOI222XLTS U2997 ( .A0(n4044), .A1(n3277), .B0(cacheDataOut[22]), .B1(n6170), 
        .C0(n3889), .C1(n3248), .Y(n5796) );
  AOI22X1TS U2998 ( .A0(n4197), .A1(n3231), .B0(n4354), .B1(n3723), .Y(n5799)
         );
  AOI222XLTS U2999 ( .A0(n4041), .A1(n3276), .B0(cacheDataOut[21]), .B1(n3260), 
        .C0(n3886), .C1(n3248), .Y(n5798) );
  AOI22X1TS U3000 ( .A0(n4194), .A1(n3231), .B0(n4351), .B1(n3723), .Y(n5801)
         );
  AOI222XLTS U3001 ( .A0(n4038), .A1(n3276), .B0(cacheDataOut[20]), .B1(n3271), 
        .C0(n3883), .C1(n3248), .Y(n5800) );
  AOI22X1TS U3002 ( .A0(n4191), .A1(n3231), .B0(n4348), .B1(n3723), .Y(n5803)
         );
  AOI222XLTS U3003 ( .A0(n4035), .A1(n3276), .B0(cacheDataOut[19]), .B1(n3271), 
        .C0(n3880), .C1(n3247), .Y(n5802) );
  AOI22X1TS U3004 ( .A0(n4182), .A1(n3230), .B0(n4339), .B1(n3722), .Y(n5809)
         );
  AOI222XLTS U3005 ( .A0(n4026), .A1(n3284), .B0(cacheDataOut[16]), .B1(n3259), 
        .C0(n3871), .C1(n3247), .Y(n5808) );
  AOI22X1TS U3006 ( .A0(n4170), .A1(n3229), .B0(n4327), .B1(n3721), .Y(n5817)
         );
  AOI222XLTS U3007 ( .A0(n4014), .A1(n3275), .B0(cacheDataOut[12]), .B1(n3269), 
        .C0(n3859), .C1(n3245), .Y(n5816) );
  AOI22X1TS U3008 ( .A0(n4167), .A1(n3229), .B0(n4324), .B1(n3721), .Y(n5819)
         );
  AOI222XLTS U3009 ( .A0(n4011), .A1(n3275), .B0(cacheDataOut[11]), .B1(n3263), 
        .C0(n3856), .C1(n3245), .Y(n5818) );
  AOI22X1TS U3010 ( .A0(n4164), .A1(n3228), .B0(n4321), .B1(n3721), .Y(n5821)
         );
  AOI222XLTS U3011 ( .A0(n4008), .A1(n3274), .B0(cacheDataOut[10]), .B1(n3263), 
        .C0(n3853), .C1(n3245), .Y(n5820) );
  AOI22X1TS U3012 ( .A0(n4158), .A1(n3228), .B0(n4315), .B1(n3720), .Y(n5825)
         );
  AOI222XLTS U3013 ( .A0(n4002), .A1(n3274), .B0(cacheDataOut[8]), .B1(n3263), 
        .C0(n3847), .C1(n3244), .Y(n5824) );
  AOI22X1TS U3014 ( .A0(n4152), .A1(n3228), .B0(n4309), .B1(n3720), .Y(n5829)
         );
  AOI222XLTS U3015 ( .A0(n3996), .A1(n3274), .B0(cacheDataOut[6]), .B1(n3262), 
        .C0(n3841), .C1(n3246), .Y(n5828) );
  AOI22X1TS U3016 ( .A0(n4137), .A1(n3226), .B0(n4294), .B1(n3718), .Y(n5839)
         );
  AOI222XLTS U3017 ( .A0(n3981), .A1(n3287), .B0(cacheDataOut[1]), .B1(n3264), 
        .C0(n3826), .C1(n3243), .Y(n5838) );
  AOI22X1TS U3018 ( .A0(n4134), .A1(n3226), .B0(n4291), .B1(n3718), .Y(n5841)
         );
  AOI222XLTS U3019 ( .A0(n3978), .A1(n3287), .B0(cacheDataOut[0]), .B1(n3270), 
        .C0(n3823), .C1(n3243), .Y(n5840) );
  AOI22X1TS U3020 ( .A0(n3951), .A1(n3320), .B0(n4420), .B1(n3708), .Y(n5451)
         );
  AOI222XLTS U3021 ( .A0(n4107), .A1(n3362), .B0(n3346), .B1(n146), .C0(n4264), 
        .C1(n3338), .Y(n5450) );
  AOI22X1TS U3022 ( .A0(n3948), .A1(n3321), .B0(n4417), .B1(n3708), .Y(n5453)
         );
  AOI222XLTS U3023 ( .A0(n4104), .A1(n3362), .B0(n3348), .B1(n140), .C0(n4261), 
        .C1(n3341), .Y(n5452) );
  AOI22X1TS U3024 ( .A0(n3945), .A1(n3317), .B0(n4414), .B1(n3708), .Y(n5455)
         );
  AOI222XLTS U3025 ( .A0(n4101), .A1(n3362), .B0(n3348), .B1(n136), .C0(n4258), 
        .C1(n3333), .Y(n5454) );
  AOI22X1TS U3026 ( .A0(n3942), .A1(n3317), .B0(n4411), .B1(n3708), .Y(n5457)
         );
  AOI222XLTS U3027 ( .A0(n4098), .A1(n3362), .B0(n3348), .B1(n132), .C0(n4255), 
        .C1(n3333), .Y(n5456) );
  AOI22X1TS U3028 ( .A0(n3939), .A1(n3322), .B0(n4408), .B1(n3709), .Y(n5459)
         );
  AOI222XLTS U3029 ( .A0(n4095), .A1(n6187), .B0(n3348), .B1(n128), .C0(n4252), 
        .C1(n3333), .Y(n5458) );
  AOI22X1TS U3030 ( .A0(n3936), .A1(n3322), .B0(n4405), .B1(n6342), .Y(n5461)
         );
  AOI222XLTS U3031 ( .A0(n4092), .A1(n6187), .B0(n3347), .B1(n125), .C0(n4249), 
        .C1(n3333), .Y(n5460) );
  AOI22X1TS U3032 ( .A0(n3912), .A1(n3318), .B0(n4381), .B1(n3709), .Y(n5717)
         );
  AOI22X1TS U3033 ( .A0(n3909), .A1(n3318), .B0(n4378), .B1(n3710), .Y(n5719)
         );
  AOI22X1TS U3034 ( .A0(n3906), .A1(n3318), .B0(n4375), .B1(n3710), .Y(n5721)
         );
  AOI22X1TS U3035 ( .A0(n3903), .A1(n3320), .B0(n4372), .B1(n3712), .Y(n5723)
         );
  AOI22X1TS U3036 ( .A0(n3900), .A1(n3321), .B0(n4369), .B1(n3709), .Y(n5725)
         );
  AOI22X1TS U3037 ( .A0(n3897), .A1(n3315), .B0(n4366), .B1(n3713), .Y(n5727)
         );
  AOI22X1TS U3038 ( .A0(n3894), .A1(n3315), .B0(n4363), .B1(n3710), .Y(n5729)
         );
  AOI22X1TS U3039 ( .A0(n3891), .A1(n3315), .B0(n4360), .B1(n3713), .Y(n5731)
         );
  AOI22X1TS U3040 ( .A0(n3888), .A1(n3315), .B0(n4357), .B1(n3710), .Y(n5733)
         );
  AOI22X1TS U3041 ( .A0(n3885), .A1(n3314), .B0(n4354), .B1(n3711), .Y(n5735)
         );
  AOI22X1TS U3042 ( .A0(n3882), .A1(n3314), .B0(n4351), .B1(n3711), .Y(n5737)
         );
  AOI22X1TS U3043 ( .A0(n3879), .A1(n3314), .B0(n4348), .B1(n3716), .Y(n5739)
         );
  AOI22X1TS U3044 ( .A0(n3876), .A1(n3313), .B0(n4345), .B1(n3712), .Y(n5741)
         );
  AOI22X1TS U3045 ( .A0(n3873), .A1(n3313), .B0(n4342), .B1(n3714), .Y(n5743)
         );
  AOI22X1TS U3046 ( .A0(n3864), .A1(n3312), .B0(n4333), .B1(n3711), .Y(n5749)
         );
  AOI22X1TS U3047 ( .A0(n3861), .A1(n3312), .B0(n4330), .B1(n3707), .Y(n5751)
         );
  AOI22X1TS U3048 ( .A0(n3858), .A1(n3312), .B0(n4327), .B1(n3707), .Y(n5753)
         );
  AOI22X1TS U3049 ( .A0(n3852), .A1(n3311), .B0(n4321), .B1(n3707), .Y(n5757)
         );
  AOI22X1TS U3050 ( .A0(n3849), .A1(n3314), .B0(n4318), .B1(n3706), .Y(n5759)
         );
  AOI22X1TS U3051 ( .A0(n3846), .A1(n3311), .B0(n4315), .B1(n3706), .Y(n5761)
         );
  AOI22X1TS U3052 ( .A0(n3843), .A1(n3311), .B0(n4312), .B1(n3706), .Y(n5763)
         );
  AOI22X1TS U3053 ( .A0(n3840), .A1(n3311), .B0(n4309), .B1(n3706), .Y(n5765)
         );
  AOI22X1TS U3054 ( .A0(n3837), .A1(n3310), .B0(n4306), .B1(n3705), .Y(n5767)
         );
  AOI22X1TS U3055 ( .A0(n3834), .A1(n3310), .B0(n4303), .B1(n3705), .Y(n5769)
         );
  AOI22X1TS U3056 ( .A0(n3831), .A1(n3310), .B0(n4300), .B1(n3705), .Y(n5771)
         );
  AOI22X1TS U3057 ( .A0(n3828), .A1(n3310), .B0(n4297), .B1(n3705), .Y(n5773)
         );
  AOI22X1TS U3058 ( .A0(n3822), .A1(n3309), .B0(n4291), .B1(n3704), .Y(n5777)
         );
  AOI22X1TS U3059 ( .A0(n3978), .A1(n689), .B0(n4291), .B1(n3762), .Y(n6033)
         );
  AOI22X1TS U3060 ( .A0(n4185), .A1(n3230), .B0(n4342), .B1(n3722), .Y(n5807)
         );
  AOI222XLTS U3061 ( .A0(n4029), .A1(n3283), .B0(cacheDataOut[17]), .B1(n6170), 
        .C0(n3874), .C1(n3247), .Y(n5806) );
  AOI22X1TS U3062 ( .A0(n4179), .A1(n3230), .B0(n4336), .B1(n3722), .Y(n5811)
         );
  AOI222XLTS U3063 ( .A0(n4023), .A1(n3284), .B0(cacheDataOut[15]), .B1(n3268), 
        .C0(n3868), .C1(n3246), .Y(n5810) );
  AOI22X1TS U3064 ( .A0(n4176), .A1(n3229), .B0(n4333), .B1(n3722), .Y(n5813)
         );
  AOI222XLTS U3065 ( .A0(n4020), .A1(n3275), .B0(cacheDataOut[14]), .B1(n3261), 
        .C0(n3865), .C1(n3246), .Y(n5812) );
  AOI22X1TS U3066 ( .A0(n4143), .A1(n3227), .B0(n4300), .B1(n3719), .Y(n5835)
         );
  AOI222XLTS U3067 ( .A0(n3987), .A1(n3273), .B0(cacheDataOut[3]), .B1(n3263), 
        .C0(n3832), .C1(n3243), .Y(n5834) );
  AOI22X1TS U3068 ( .A0(n817), .A1(n129), .B0(n789), .B1(n4077), .Y(n6138) );
  AOI222XLTS U3069 ( .A0(\requesterAddressbuffer[2][1] ), .A1(n289), .B0(n831), 
        .B1(n4234), .C0(n3746), .C1(n4391), .Y(n6137) );
  AOI22X1TS U3070 ( .A0(n6140), .A1(n114), .B0(n790), .B1(n4074), .Y(n6143) );
  AOI222XLTS U3071 ( .A0(\requesterAddressbuffer[2][0] ), .A1(n272), .B0(n831), 
        .B1(n4231), .C0(n3746), .C1(n4388), .Y(n6142) );
  AOI22X1TS U3072 ( .A0(n817), .A1(n137), .B0(n789), .B1(n4083), .Y(n6134) );
  AOI222XLTS U3073 ( .A0(\requesterAddressbuffer[2][3] ), .A1(n273), .B0(n831), 
        .B1(n4240), .C0(n3746), .C1(n4397), .Y(n6133) );
  AOI22X1TS U3074 ( .A0(n818), .A1(n131), .B0(n789), .B1(n4080), .Y(n6136) );
  AOI222XLTS U3075 ( .A0(\requesterAddressbuffer[2][2] ), .A1(n234), .B0(n831), 
        .B1(n4237), .C0(n3746), .C1(n4394), .Y(n6135) );
  AOI22X1TS U3076 ( .A0(n814), .A1(n142), .B0(n789), .B1(n4086), .Y(n6132) );
  AOI222XLTS U3077 ( .A0(\requesterAddressbuffer[2][4] ), .A1(n186), .B0(n837), 
        .B1(n4243), .C0(n3747), .C1(n4400), .Y(n6131) );
  AOI22X1TS U3078 ( .A0(n819), .A1(n118), .B0(n790), .B1(n4089), .Y(n6130) );
  AOI222XLTS U3079 ( .A0(\requesterAddressbuffer[2][5] ), .A1(n290), .B0(n830), 
        .B1(n4246), .C0(n3747), .C1(n4403), .Y(n6129) );
  AOI22X1TS U3080 ( .A0(n3408), .A1(n135), .B0(n3391), .B1(n4083), .Y(n6195)
         );
  AOI222XLTS U3081 ( .A0(\requesterAddressbuffer[6][3] ), .A1(n579), .B0(n3431), .B1(n4239), .C0(n3697), .C1(n4397), .Y(n6194) );
  AOI22X1TS U3082 ( .A0(n3408), .A1(n127), .B0(n3391), .B1(n4077), .Y(n6199)
         );
  AOI222XLTS U3083 ( .A0(\requesterAddressbuffer[6][1] ), .A1(n579), .B0(n3431), .B1(n4233), .C0(n3697), .C1(n4391), .Y(n6198) );
  AOI222XLTS U3084 ( .A0(\requesterAddressbuffer[6][0] ), .A1(n579), .B0(n3437), .B1(n4230), .C0(n3697), .C1(n4388), .Y(n6203) );
  AOI22X1TS U3085 ( .A0(n669), .A1(n144), .B0(n585), .B1(n4245), .Y(n6099) );
  AOI222XLTS U3086 ( .A0(\requesterAddressbuffer[0][5] ), .A1(n207), .B0(n678), 
        .B1(n3934), .C0(n3791), .C1(n4403), .Y(n6098) );
  AOI22X1TS U3087 ( .A0(n626), .A1(n135), .B0(n584), .B1(n4239), .Y(n6103) );
  AOI222XLTS U3088 ( .A0(\requesterAddressbuffer[0][3] ), .A1(n3776), .B0(n679), .B1(n3928), .C0(n3790), .C1(n4397), .Y(n6102) );
  AOI22X1TS U3089 ( .A0(n669), .A1(n140), .B0(n584), .B1(n4242), .Y(n6101) );
  AOI222XLTS U3090 ( .A0(\requesterAddressbuffer[0][4] ), .A1(n278), .B0(n685), 
        .B1(n3931), .C0(n3791), .C1(n4400), .Y(n6100) );
  AOI22X1TS U3091 ( .A0(n626), .A1(n131), .B0(n584), .B1(n4236), .Y(n6105) );
  AOI222XLTS U3092 ( .A0(\requesterAddressbuffer[0][2] ), .A1(n278), .B0(n679), 
        .B1(n3925), .C0(n3790), .C1(n4394), .Y(n6104) );
  AOI22X1TS U3093 ( .A0(n626), .A1(n127), .B0(n584), .B1(n4233), .Y(n6107) );
  AOI222XLTS U3094 ( .A0(\requesterAddressbuffer[0][1] ), .A1(n207), .B0(n679), 
        .B1(n3922), .C0(n3790), .C1(n4391), .Y(n6106) );
  AOI22X1TS U3095 ( .A0(n666), .A1(n123), .B0(n585), .B1(n4230), .Y(n6112) );
  AOI222XLTS U3096 ( .A0(\requesterAddressbuffer[0][0] ), .A1(n282), .B0(n679), 
        .B1(n3919), .C0(n3790), .C1(n4388), .Y(n6111) );
  AOI22X1TS U3097 ( .A0(n626), .A1(readRequesterAddress[5]), .B0(n4263), .B1(
        n609), .Y(n5335) );
  AOI222XLTS U3098 ( .A0(n280), .A1(n27), .B0(n3952), .B1(n673), .C0(n4421), 
        .C1(n3797), .Y(n5334) );
  AOI22X1TS U3099 ( .A0(n6109), .A1(n117), .B0(n4257), .B1(n609), .Y(n5339) );
  AOI222XLTS U3100 ( .A0(n278), .A1(n28), .B0(n3946), .B1(n678), .C0(n4415), 
        .C1(n3797), .Y(n5338) );
  AOI22X1TS U3101 ( .A0(n669), .A1(n116), .B0(n4254), .B1(n609), .Y(n5341) );
  AOI222XLTS U3102 ( .A0(n3776), .A1(n29), .B0(n3943), .B1(n678), .C0(n4412), 
        .C1(n3797), .Y(n5340) );
  AOI22X1TS U3103 ( .A0(n668), .A1(n115), .B0(n4251), .B1(n614), .Y(n5343) );
  AOI222XLTS U3104 ( .A0(n184), .A1(n30), .B0(n3940), .B1(n680), .C0(n4409), 
        .C1(n3796), .Y(n5342) );
  AOI22X1TS U3105 ( .A0(n347), .A1(n665), .B0(n4227), .B1(n612), .Y(n6035) );
  AOI222XLTS U3106 ( .A0(n207), .A1(n31), .B0(n3916), .B1(n680), .C0(n4385), 
        .C1(n3796), .Y(n6034) );
  AOI22X1TS U3107 ( .A0(n349), .A1(n627), .B0(n4224), .B1(n625), .Y(n6037) );
  AOI222XLTS U3108 ( .A0(n279), .A1(n32), .B0(n3913), .B1(n687), .C0(n4382), 
        .C1(n3796), .Y(n6036) );
  AOI22X1TS U3109 ( .A0(n351), .A1(n627), .B0(n4221), .B1(n622), .Y(n6039) );
  AOI222XLTS U3110 ( .A0(n206), .A1(n33), .B0(n3910), .B1(n681), .C0(n4379), 
        .C1(n3795), .Y(n6038) );
  AOI22X1TS U3111 ( .A0(n357), .A1(n662), .B0(n4212), .B1(n623), .Y(n6045) );
  AOI222XLTS U3112 ( .A0(n280), .A1(n34), .B0(n3901), .B1(n680), .C0(n4370), 
        .C1(n3795), .Y(n6044) );
  AOI22X1TS U3113 ( .A0(n359), .A1(n627), .B0(n4209), .B1(n613), .Y(n6047) );
  AOI222XLTS U3114 ( .A0(n208), .A1(n35), .B0(n3898), .B1(n681), .C0(n4367), 
        .C1(n3794), .Y(n6046) );
  AOI22X1TS U3115 ( .A0(n361), .A1(n659), .B0(n4206), .B1(n613), .Y(n6049) );
  AOI222XLTS U3116 ( .A0(n184), .A1(n36), .B0(n3895), .B1(n684), .C0(n4364), 
        .C1(n3794), .Y(n6048) );
  AOI22X1TS U3117 ( .A0(n365), .A1(n659), .B0(n4200), .B1(n613), .Y(n6053) );
  AOI222XLTS U3118 ( .A0(n280), .A1(n37), .B0(n3889), .B1(n681), .C0(n4358), 
        .C1(n3794), .Y(n6052) );
  AOI22X1TS U3119 ( .A0(n367), .A1(n660), .B0(n4197), .B1(n608), .Y(n6055) );
  AOI222XLTS U3120 ( .A0(n185), .A1(n38), .B0(n3886), .B1(n677), .C0(n4355), 
        .C1(n3793), .Y(n6054) );
  AOI22X1TS U3121 ( .A0(n371), .A1(n660), .B0(n4191), .B1(n608), .Y(n6059) );
  AOI222XLTS U3122 ( .A0(n207), .A1(n39), .B0(n3880), .B1(n677), .C0(n4349), 
        .C1(n3793), .Y(n6058) );
  AOI22X1TS U3123 ( .A0(n373), .A1(n661), .B0(n4188), .B1(n607), .Y(n6061) );
  AOI222XLTS U3124 ( .A0(n279), .A1(n40), .B0(n3877), .B1(n682), .C0(n4346), 
        .C1(n3793), .Y(n6060) );
  AOI22X1TS U3125 ( .A0(n375), .A1(n660), .B0(n4185), .B1(n607), .Y(n6063) );
  AOI222XLTS U3126 ( .A0(n158), .A1(n41), .B0(n3874), .B1(n682), .C0(n4343), 
        .C1(n3792), .Y(n6062) );
  AOI22X1TS U3127 ( .A0(n377), .A1(n661), .B0(n4182), .B1(n607), .Y(n6065) );
  AOI222XLTS U3128 ( .A0(n206), .A1(n42), .B0(n3871), .B1(n681), .C0(n4340), 
        .C1(n3792), .Y(n6064) );
  AOI22X1TS U3129 ( .A0(n379), .A1(n662), .B0(n4179), .B1(n607), .Y(n6067) );
  AOI222XLTS U3130 ( .A0(n283), .A1(n43), .B0(n3868), .B1(n683), .C0(n4337), 
        .C1(n3792), .Y(n6066) );
  AOI22X1TS U3131 ( .A0(n381), .A1(n661), .B0(n4176), .B1(n594), .Y(n6069) );
  AOI222XLTS U3132 ( .A0(n279), .A1(n44), .B0(n3865), .B1(n676), .C0(n4334), 
        .C1(n3792), .Y(n6068) );
  AOI22X1TS U3133 ( .A0(n383), .A1(n661), .B0(n4173), .B1(n594), .Y(n6071) );
  AOI222XLTS U3134 ( .A0(n185), .A1(n45), .B0(n3862), .B1(n676), .C0(n4331), 
        .C1(n3798), .Y(n6070) );
  AOI22X1TS U3135 ( .A0(n385), .A1(n662), .B0(n4170), .B1(n594), .Y(n6073) );
  AOI222XLTS U3136 ( .A0(n279), .A1(n46), .B0(n3859), .B1(n676), .C0(n4328), 
        .C1(n421), .Y(n6072) );
  AOI22X1TS U3137 ( .A0(n387), .A1(n662), .B0(n4167), .B1(n594), .Y(n6075) );
  AOI222XLTS U3138 ( .A0(n208), .A1(n47), .B0(n3856), .B1(n676), .C0(n4325), 
        .C1(n3799), .Y(n6074) );
  AOI22X1TS U3139 ( .A0(n389), .A1(n665), .B0(n4164), .B1(n587), .Y(n6077) );
  AOI222XLTS U3140 ( .A0(n208), .A1(n48), .B0(n3853), .B1(n675), .C0(n4322), 
        .C1(n3800), .Y(n6076) );
  AOI22X1TS U3141 ( .A0(n393), .A1(n663), .B0(n4158), .B1(n587), .Y(n6081) );
  AOI222XLTS U3142 ( .A0(n206), .A1(n49), .B0(n3847), .B1(n675), .C0(n4316), 
        .C1(n3801), .Y(n6080) );
  AOI22X1TS U3143 ( .A0(n395), .A1(n663), .B0(n4155), .B1(n587), .Y(n6083) );
  AOI222XLTS U3144 ( .A0(n3775), .A1(n50), .B0(n3844), .B1(n675), .C0(n4313), 
        .C1(n3801), .Y(n6082) );
  AOI22X1TS U3145 ( .A0(n397), .A1(n664), .B0(n4152), .B1(n587), .Y(n6085) );
  AOI222XLTS U3146 ( .A0(n208), .A1(n51), .B0(n3841), .B1(n677), .C0(n4310), 
        .C1(n3801), .Y(n6084) );
  AOI22X1TS U3147 ( .A0(n401), .A1(n664), .B0(n4146), .B1(n586), .Y(n6089) );
  AOI222XLTS U3148 ( .A0(n184), .A1(n52), .B0(n3835), .B1(n674), .C0(n4304), 
        .C1(n228), .Y(n6088) );
  AOI22X1TS U3149 ( .A0(n403), .A1(n665), .B0(n4143), .B1(n586), .Y(n6091) );
  AOI222XLTS U3150 ( .A0(n185), .A1(n53), .B0(n3832), .B1(n674), .C0(n4301), 
        .C1(n3799), .Y(n6090) );
  AOI22X1TS U3151 ( .A0(n6109), .A1(n142), .B0(n4260), .B1(n609), .Y(n5337) );
  AOI22X1TS U3152 ( .A0(n670), .A1(readRequesterAddress[0]), .B0(n4248), .B1(
        n6108), .Y(n5345) );
  AOI222XLTS U3153 ( .A0(n282), .A1(n55), .B0(n3937), .B1(n686), .C0(n4406), 
        .C1(n3796), .Y(n5344) );
  AOI22X1TS U3154 ( .A0(n353), .A1(n627), .B0(n4218), .B1(n622), .Y(n6041) );
  AOI222XLTS U3155 ( .A0(n282), .A1(n56), .B0(n3907), .B1(n683), .C0(n4376), 
        .C1(n3795), .Y(n6040) );
  AOI22X1TS U3156 ( .A0(n355), .A1(n659), .B0(n4215), .B1(n623), .Y(n6043) );
  AOI222XLTS U3157 ( .A0(n3776), .A1(n57), .B0(n3904), .B1(n682), .C0(n4373), 
        .C1(n3795), .Y(n6042) );
  AOI22X1TS U3158 ( .A0(n363), .A1(n659), .B0(n4203), .B1(n614), .Y(n6051) );
  AOI222XLTS U3159 ( .A0(n280), .A1(n58), .B0(n3892), .B1(n684), .C0(n4361), 
        .C1(n3794), .Y(n6050) );
  AOI22X1TS U3160 ( .A0(n369), .A1(n660), .B0(n4194), .B1(n608), .Y(n6057) );
  AOI222XLTS U3161 ( .A0(n283), .A1(n59), .B0(n3883), .B1(n677), .C0(n4352), 
        .C1(n3793), .Y(n6056) );
  AOI22X1TS U3162 ( .A0(n391), .A1(n663), .B0(n4161), .B1(n608), .Y(n6079) );
  AOI222XLTS U3163 ( .A0(n283), .A1(n60), .B0(n3850), .B1(n675), .C0(n4319), 
        .C1(n421), .Y(n6078) );
  AOI22X1TS U3164 ( .A0(n399), .A1(n663), .B0(n4149), .B1(n586), .Y(n6087) );
  AOI222XLTS U3165 ( .A0(n282), .A1(n61), .B0(n3838), .B1(n674), .C0(n4307), 
        .C1(n3800), .Y(n6086) );
  AOI22X1TS U3166 ( .A0(n405), .A1(n664), .B0(n4140), .B1(n586), .Y(n6093) );
  AOI222XLTS U3167 ( .A0(n3775), .A1(n62), .B0(n3829), .B1(n674), .C0(n4298), 
        .C1(n3798), .Y(n6092) );
  AOI22X1TS U3168 ( .A0(n407), .A1(n664), .B0(n4137), .B1(n585), .Y(n6095) );
  AOI222XLTS U3169 ( .A0(n185), .A1(n63), .B0(n3826), .B1(n673), .C0(n4295), 
        .C1(n3791), .Y(n6094) );
  AOI22X1TS U3170 ( .A0(n409), .A1(n665), .B0(n4134), .B1(n585), .Y(n6097) );
  AOI222XLTS U3171 ( .A0(n283), .A1(n64), .B0(n3823), .B1(n673), .C0(n4292), 
        .C1(n3791), .Y(n6096) );
  AOI22X1TS U3172 ( .A0(n857), .A1(readRequesterAddress[5]), .B0(n4263), .B1(
        n288), .Y(n5405) );
  AOI222XLTS U3173 ( .A0(n3208), .A1(n6255), .B0(n3952), .B1(n3193), .C0(n4421), .C1(n1602), .Y(n5404) );
  AOI22X1TS U3174 ( .A0(n857), .A1(n139), .B0(n4260), .B1(n221), .Y(n5407) );
  AOI222XLTS U3175 ( .A0(n3208), .A1(n6256), .B0(n3949), .B1(n3201), .C0(n4418), .C1(n1602), .Y(n5406) );
  AOI22X1TS U3176 ( .A0(n857), .A1(readRequesterAddress[3]), .B0(n4257), .B1(
        n288), .Y(n5409) );
  AOI222XLTS U3177 ( .A0(n3208), .A1(n6257), .B0(n3946), .B1(n3201), .C0(n4415), .C1(n1602), .Y(n5408) );
  AOI22X1TS U3178 ( .A0(n858), .A1(readRequesterAddress[1]), .B0(n4251), .B1(
        n287), .Y(n5413) );
  AOI222XLTS U3179 ( .A0(n3209), .A1(n6258), .B0(n3940), .B1(n3200), .C0(n4409), .C1(n1402), .Y(n5412) );
  AOI22X1TS U3180 ( .A0(n858), .A1(readRequesterAddress[0]), .B0(n4248), .B1(
        n287), .Y(n5415) );
  AOI222XLTS U3181 ( .A0(n3209), .A1(n6259), .B0(n3937), .B1(n3200), .C0(n4406), .C1(n1402), .Y(n5414) );
  AOI22X1TS U3182 ( .A0(n347), .A1(n863), .B0(n4227), .B1(n213), .Y(n5843) );
  AOI222XLTS U3183 ( .A0(n3209), .A1(n6260), .B0(n3916), .B1(n3200), .C0(n4385), .C1(n1402), .Y(n5842) );
  AOI22X1TS U3184 ( .A0(n349), .A1(n870), .B0(n4224), .B1(n209), .Y(n5845) );
  AOI222XLTS U3185 ( .A0(n3209), .A1(n6261), .B0(n3913), .B1(n3200), .C0(n4382), .C1(n1402), .Y(n5844) );
  AOI22X1TS U3186 ( .A0(n351), .A1(n6154), .B0(n4221), .B1(n214), .Y(n5847) );
  AOI222XLTS U3187 ( .A0(n3210), .A1(n6262), .B0(n3910), .B1(n3199), .C0(n4379), .C1(n986), .Y(n5846) );
  AOI22X1TS U3188 ( .A0(n353), .A1(n864), .B0(n4218), .B1(n211), .Y(n5849) );
  AOI222XLTS U3189 ( .A0(n3210), .A1(n6263), .B0(n3907), .B1(n3199), .C0(n4376), .C1(n986), .Y(n5848) );
  AOI22X1TS U3190 ( .A0(n355), .A1(n6154), .B0(n4215), .B1(n219), .Y(n5851) );
  AOI222XLTS U3191 ( .A0(n3210), .A1(n6264), .B0(n3904), .B1(n3199), .C0(n4373), .C1(n986), .Y(n5850) );
  AOI22X1TS U3192 ( .A0(n357), .A1(n863), .B0(n4212), .B1(n218), .Y(n5853) );
  AOI222XLTS U3193 ( .A0(n3210), .A1(n6265), .B0(n3901), .B1(n3199), .C0(n4370), .C1(n986), .Y(n5852) );
  AOI22X1TS U3194 ( .A0(n361), .A1(n864), .B0(n4206), .B1(n209), .Y(n5857) );
  AOI222XLTS U3195 ( .A0(n3211), .A1(n6266), .B0(n3895), .B1(n3198), .C0(n4364), .C1(n970), .Y(n5856) );
  AOI22X1TS U3196 ( .A0(n365), .A1(n868), .B0(n4200), .B1(n221), .Y(n5861) );
  AOI222XLTS U3197 ( .A0(n3211), .A1(n6267), .B0(n3889), .B1(n3198), .C0(n4358), .C1(n970), .Y(n5860) );
  AOI22X1TS U3198 ( .A0(n367), .A1(n867), .B0(n4197), .B1(n286), .Y(n5863) );
  AOI222XLTS U3199 ( .A0(n3212), .A1(n6268), .B0(n3886), .B1(n3197), .C0(n4355), .C1(n959), .Y(n5862) );
  AOI22X1TS U3200 ( .A0(n371), .A1(n864), .B0(n4191), .B1(n288), .Y(n5867) );
  AOI222XLTS U3201 ( .A0(n3212), .A1(n6269), .B0(n3880), .B1(n3197), .C0(n4349), .C1(n959), .Y(n5866) );
  AOI22X1TS U3202 ( .A0(n375), .A1(n865), .B0(n4185), .B1(n286), .Y(n5871) );
  AOI222XLTS U3203 ( .A0(n3213), .A1(n6270), .B0(n3874), .B1(n3196), .C0(n4343), .C1(n957), .Y(n5870) );
  AOI22X1TS U3204 ( .A0(n377), .A1(n865), .B0(n4182), .B1(n287), .Y(n5873) );
  AOI222XLTS U3205 ( .A0(n3213), .A1(n6271), .B0(n3871), .B1(n3196), .C0(n4340), .C1(n957), .Y(n5872) );
  AOI22X1TS U3206 ( .A0(n381), .A1(n865), .B0(n4176), .B1(n220), .Y(n5877) );
  AOI222XLTS U3207 ( .A0(n3213), .A1(n6272), .B0(n3865), .B1(n3195), .C0(n4334), .C1(n957), .Y(n5876) );
  AOI22X1TS U3208 ( .A0(n385), .A1(n868), .B0(n4170), .B1(n288), .Y(n5881) );
  AOI222XLTS U3209 ( .A0(n3214), .A1(n6273), .B0(n3859), .B1(n3195), .C0(n4328), .C1(n955), .Y(n5880) );
  AOI22X1TS U3210 ( .A0(n387), .A1(n862), .B0(n4167), .B1(n221), .Y(n5883) );
  AOI222XLTS U3211 ( .A0(n3214), .A1(n6274), .B0(n3856), .B1(n3195), .C0(n4325), .C1(n955), .Y(n5882) );
  AOI22X1TS U3212 ( .A0(n389), .A1(n862), .B0(n4164), .B1(n218), .Y(n5885) );
  AOI222XLTS U3213 ( .A0(n3214), .A1(n6275), .B0(n3853), .B1(n3207), .C0(n4322), .C1(n955), .Y(n5884) );
  AOI22X1TS U3214 ( .A0(n391), .A1(n862), .B0(n4161), .B1(n220), .Y(n5887) );
  AOI222XLTS U3215 ( .A0(n3215), .A1(n6276), .B0(n3850), .B1(n3202), .C0(n4319), .C1(n936), .Y(n5886) );
  AOI22X1TS U3216 ( .A0(n393), .A1(n862), .B0(n4158), .B1(n213), .Y(n5889) );
  AOI222XLTS U3217 ( .A0(n3215), .A1(n6277), .B0(n3847), .B1(n3202), .C0(n4316), .C1(n936), .Y(n5888) );
  AOI22X1TS U3218 ( .A0(n397), .A1(n861), .B0(n4152), .B1(n211), .Y(n5893) );
  AOI222XLTS U3219 ( .A0(n3215), .A1(n6278), .B0(n3841), .B1(n3197), .C0(n4310), .C1(n936), .Y(n5892) );
  AOI22X1TS U3220 ( .A0(n403), .A1(n860), .B0(n4143), .B1(n214), .Y(n5899) );
  AOI222XLTS U3221 ( .A0(n3216), .A1(n6279), .B0(n3832), .B1(n3194), .C0(n4301), .C1(n919), .Y(n5898) );
  AOI22X1TS U3222 ( .A0(n407), .A1(n860), .B0(n4137), .B1(n285), .Y(n5903) );
  AOI222XLTS U3223 ( .A0(n3217), .A1(n6280), .B0(n3826), .B1(n3193), .C0(n4295), .C1(n886), .Y(n5902) );
  AOI22X1TS U3224 ( .A0(n409), .A1(n860), .B0(n4134), .B1(n213), .Y(n5905) );
  AOI222XLTS U3225 ( .A0(n3217), .A1(n6281), .B0(n3823), .B1(n3193), .C0(n4292), .C1(n886), .Y(n5904) );
  AOI22X1TS U3226 ( .A0(n858), .A1(readRequesterAddress[2]), .B0(n4254), .B1(
        n220), .Y(n5411) );
  AOI222XLTS U3227 ( .A0(n3208), .A1(n6293), .B0(n3943), .B1(n3201), .C0(n4412), .C1(n1602), .Y(n5410) );
  AOI22X1TS U3228 ( .A0(n359), .A1(n867), .B0(n4209), .B1(n286), .Y(n5855) );
  AOI222XLTS U3229 ( .A0(n3211), .A1(n6294), .B0(n3898), .B1(n3198), .C0(n4367), .C1(n970), .Y(n5854) );
  AOI22X1TS U3230 ( .A0(n363), .A1(n866), .B0(n4203), .B1(n219), .Y(n5859) );
  AOI222XLTS U3231 ( .A0(n3211), .A1(n6295), .B0(n3892), .B1(n3198), .C0(n4361), .C1(n970), .Y(n5858) );
  AOI22X1TS U3232 ( .A0(n369), .A1(n866), .B0(n4194), .B1(n219), .Y(n5865) );
  AOI222XLTS U3233 ( .A0(n3212), .A1(n6296), .B0(n3883), .B1(n3197), .C0(n4352), .C1(n959), .Y(n5864) );
  AOI22X1TS U3234 ( .A0(n373), .A1(n865), .B0(n4188), .B1(n287), .Y(n5869) );
  AOI222XLTS U3235 ( .A0(n3212), .A1(n6297), .B0(n3877), .B1(n3196), .C0(n4346), .C1(n959), .Y(n5868) );
  AOI22X1TS U3236 ( .A0(n379), .A1(n864), .B0(n4179), .B1(n220), .Y(n5875) );
  AOI222XLTS U3237 ( .A0(n3213), .A1(n6298), .B0(n3868), .B1(n3196), .C0(n4337), .C1(n957), .Y(n5874) );
  AOI22X1TS U3238 ( .A0(n383), .A1(n869), .B0(n4173), .B1(n286), .Y(n5879) );
  AOI222XLTS U3239 ( .A0(n3214), .A1(n6299), .B0(n3862), .B1(n3195), .C0(n4331), .C1(n955), .Y(n5878) );
  AOI22X1TS U3240 ( .A0(n399), .A1(n861), .B0(n4149), .B1(n211), .Y(n5895) );
  AOI222XLTS U3241 ( .A0(n3216), .A1(n6300), .B0(n3838), .B1(n3194), .C0(n4307), .C1(n919), .Y(n5894) );
  AOI22X1TS U3242 ( .A0(n401), .A1(n861), .B0(n4146), .B1(n214), .Y(n5897) );
  AOI222XLTS U3243 ( .A0(n3216), .A1(n6301), .B0(n3835), .B1(n3194), .C0(n4304), .C1(n919), .Y(n5896) );
  AOI22X1TS U3244 ( .A0(n405), .A1(n860), .B0(n4140), .B1(n218), .Y(n5901) );
  AOI222XLTS U3245 ( .A0(n3216), .A1(n6302), .B0(n3829), .B1(n3194), .C0(n4298), .C1(n919), .Y(n5900) );
  AOI22X1TS U3246 ( .A0(n395), .A1(n861), .B0(n4155), .B1(n209), .Y(n5891) );
  AOI222XLTS U3247 ( .A0(n3215), .A1(n6312), .B0(n3844), .B1(n3206), .C0(n4313), .C1(n936), .Y(n5890) );
  AOI22X1TS U3248 ( .A0(n806), .A1(readRequesterAddress[2]), .B0(n4098), .B1(
        n796), .Y(n5385) );
  AOI222XLTS U3249 ( .A0(n226), .A1(n65), .B0(n4255), .B1(n830), .C0(n4412), 
        .C1(n3753), .Y(n5384) );
  AOI22X1TS U3250 ( .A0(n350), .A1(n807), .B0(n4068), .B1(n801), .Y(n5909) );
  AOI222XLTS U3251 ( .A0(n186), .A1(n66), .B0(n4225), .B1(n829), .C0(n4382), 
        .C1(n3752), .Y(n5908) );
  AOI22X1TS U3252 ( .A0(n352), .A1(n807), .B0(n4065), .B1(n799), .Y(n5911) );
  AOI222XLTS U3253 ( .A0(n289), .A1(n67), .B0(n4222), .B1(n833), .C0(n4379), 
        .C1(n3755), .Y(n5910) );
  AOI22X1TS U3254 ( .A0(n354), .A1(n807), .B0(n4062), .B1(n799), .Y(n5913) );
  AOI222XLTS U3255 ( .A0(n272), .A1(n68), .B0(n4219), .B1(n833), .C0(n4376), 
        .C1(n3755), .Y(n5912) );
  AOI22X1TS U3256 ( .A0(n358), .A1(n815), .B0(n4056), .B1(n802), .Y(n5917) );
  AOI222XLTS U3257 ( .A0(n227), .A1(n69), .B0(n4213), .B1(n836), .C0(n4370), 
        .C1(n3755), .Y(n5916) );
  AOI22X1TS U3258 ( .A0(n360), .A1(n807), .B0(n4053), .B1(n795), .Y(n5919) );
  AOI222XLTS U3259 ( .A0(n234), .A1(n70), .B0(n4210), .B1(n833), .C0(n4367), 
        .C1(n3756), .Y(n5918) );
  AOI22X1TS U3260 ( .A0(n364), .A1(n808), .B0(n4047), .B1(n795), .Y(n5923) );
  AOI222XLTS U3261 ( .A0(n273), .A1(n71), .B0(n4204), .B1(n833), .C0(n4361), 
        .C1(n3755), .Y(n5922) );
  AOI22X1TS U3262 ( .A0(n368), .A1(n809), .B0(n4041), .B1(n800), .Y(n5927) );
  AOI222XLTS U3263 ( .A0(n234), .A1(n72), .B0(n4198), .B1(n828), .C0(n4355), 
        .C1(n3758), .Y(n5926) );
  AOI22X1TS U3264 ( .A0(n370), .A1(n809), .B0(n4038), .B1(n800), .Y(n5929) );
  AOI222XLTS U3265 ( .A0(n272), .A1(n73), .B0(n4195), .B1(n828), .C0(n4352), 
        .C1(n3758), .Y(n5928) );
  AOI22X1TS U3266 ( .A0(n372), .A1(n809), .B0(n4035), .B1(n799), .Y(n5931) );
  AOI222XLTS U3267 ( .A0(n226), .A1(n74), .B0(n4192), .B1(n828), .C0(n4349), 
        .C1(n3758), .Y(n5930) );
  AOI22X1TS U3268 ( .A0(n374), .A1(n810), .B0(n4032), .B1(n794), .Y(n5933) );
  AOI222XLTS U3269 ( .A0(n198), .A1(n75), .B0(n4189), .B1(n827), .C0(n4346), 
        .C1(n3760), .Y(n5932) );
  AOI22X1TS U3270 ( .A0(n376), .A1(n809), .B0(n4029), .B1(n794), .Y(n5935) );
  AOI222XLTS U3271 ( .A0(n186), .A1(n76), .B0(n4186), .B1(n827), .C0(n4343), 
        .C1(n3751), .Y(n5934) );
  AOI22X1TS U3272 ( .A0(n380), .A1(n816), .B0(n4023), .B1(n794), .Y(n5939) );
  AOI222XLTS U3273 ( .A0(n227), .A1(n77), .B0(n4180), .B1(n827), .C0(n4337), 
        .C1(n3751), .Y(n5938) );
  AOI22X1TS U3274 ( .A0(n382), .A1(n810), .B0(n4020), .B1(n793), .Y(n5941) );
  AOI222XLTS U3275 ( .A0(n3745), .A1(n78), .B0(n4177), .B1(n826), .C0(n4334), 
        .C1(n3751), .Y(n5940) );
  AOI22X1TS U3276 ( .A0(n384), .A1(n810), .B0(n4017), .B1(n793), .Y(n5943) );
  AOI222XLTS U3277 ( .A0(n226), .A1(n79), .B0(n4174), .B1(n826), .C0(n4331), 
        .C1(n3750), .Y(n5942) );
  AOI22X1TS U3278 ( .A0(n386), .A1(n815), .B0(n4014), .B1(n793), .Y(n5945) );
  AOI222XLTS U3279 ( .A0(n272), .A1(n80), .B0(n4171), .B1(n826), .C0(n4328), 
        .C1(n3750), .Y(n5944) );
  AOI22X1TS U3280 ( .A0(n388), .A1(n816), .B0(n4011), .B1(n793), .Y(n5947) );
  AOI222XLTS U3281 ( .A0(n6344), .A1(n81), .B0(n4168), .B1(n826), .C0(n4325), 
        .C1(n3750), .Y(n5946) );
  AOI22X1TS U3282 ( .A0(n392), .A1(n811), .B0(n4005), .B1(n802), .Y(n5951) );
  AOI222XLTS U3283 ( .A0(n3745), .A1(n82), .B0(n4162), .B1(n824), .C0(n4319), 
        .C1(n3749), .Y(n5950) );
  AOI22X1TS U3284 ( .A0(n394), .A1(n811), .B0(n4002), .B1(n792), .Y(n5953) );
  AOI222XLTS U3285 ( .A0(n183), .A1(n83), .B0(n4159), .B1(n824), .C0(n4316), 
        .C1(n3749), .Y(n5952) );
  AOI22X1TS U3286 ( .A0(n396), .A1(n811), .B0(n3999), .B1(n792), .Y(n5955) );
  AOI222XLTS U3287 ( .A0(n273), .A1(n84), .B0(n4156), .B1(n824), .C0(n4313), 
        .C1(n3749), .Y(n5954) );
  AOI22X1TS U3288 ( .A0(n400), .A1(n811), .B0(n3993), .B1(n791), .Y(n5959) );
  AOI222XLTS U3289 ( .A0(n274), .A1(n85), .B0(n4150), .B1(n823), .C0(n4307), 
        .C1(n3748), .Y(n5958) );
  AOI22X1TS U3290 ( .A0(n402), .A1(n812), .B0(n3990), .B1(n791), .Y(n5961) );
  AOI222XLTS U3291 ( .A0(n290), .A1(n86), .B0(n4147), .B1(n823), .C0(n4304), 
        .C1(n3748), .Y(n5960) );
  AOI22X1TS U3292 ( .A0(n404), .A1(n813), .B0(n3987), .B1(n791), .Y(n5963) );
  AOI222XLTS U3293 ( .A0(n3745), .A1(n87), .B0(n4144), .B1(n823), .C0(n4301), 
        .C1(n3748), .Y(n5962) );
  AOI22X1TS U3294 ( .A0(n3933), .A1(n3440), .B0(n4402), .B1(n3667), .Y(n6207)
         );
  AOI222XLTS U3295 ( .A0(n4089), .A1(n3488), .B0(n146), .B1(n3481), .C0(n4246), 
        .C1(n3459), .Y(n6206) );
  AOI22X1TS U3296 ( .A0(n3930), .A1(n3439), .B0(n4399), .B1(n3667), .Y(n6209)
         );
  AOI222XLTS U3297 ( .A0(n4086), .A1(n3487), .B0(n141), .B1(n3481), .C0(n4243), 
        .C1(n3459), .Y(n6208) );
  AOI22X1TS U3298 ( .A0(n3924), .A1(n3439), .B0(n4393), .B1(n3668), .Y(n6213)
         );
  AOI222XLTS U3299 ( .A0(n4080), .A1(n3487), .B0(n133), .B1(n3482), .C0(n4237), 
        .C1(n3459), .Y(n6212) );
  AOI22X1TS U3300 ( .A0(n818), .A1(n144), .B0(n4107), .B1(n796), .Y(n5379) );
  AOI222XLTS U3301 ( .A0(n227), .A1(n88), .B0(n4264), .B1(n822), .C0(n4421), 
        .C1(n3753), .Y(n5378) );
  AOI22X1TS U3302 ( .A0(n806), .A1(n139), .B0(n4104), .B1(n796), .Y(n5381) );
  AOI222XLTS U3303 ( .A0(n183), .A1(n89), .B0(n4261), .B1(n830), .C0(n4418), 
        .C1(n3753), .Y(n5380) );
  AOI22X1TS U3304 ( .A0(n806), .A1(readRequesterAddress[3]), .B0(n4101), .B1(
        n796), .Y(n5383) );
  AOI222XLTS U3305 ( .A0(n289), .A1(n90), .B0(n4258), .B1(n830), .C0(n4415), 
        .C1(n3753), .Y(n5382) );
  AOI22X1TS U3306 ( .A0(n818), .A1(readRequesterAddress[1]), .B0(n4095), .B1(
        n803), .Y(n5387) );
  AOI222XLTS U3307 ( .A0(n290), .A1(n91), .B0(n4252), .B1(n829), .C0(n4409), 
        .C1(n3752), .Y(n5386) );
  AOI22X1TS U3308 ( .A0(n806), .A1(n123), .B0(n4092), .B1(n799), .Y(n5389) );
  AOI222XLTS U3309 ( .A0(n226), .A1(n92), .B0(n4249), .B1(n829), .C0(n4406), 
        .C1(n3752), .Y(n5388) );
  AOI22X1TS U3310 ( .A0(n356), .A1(n808), .B0(n4059), .B1(n803), .Y(n5915) );
  AOI222XLTS U3311 ( .A0(n183), .A1(n93), .B0(n4216), .B1(n832), .C0(n4373), 
        .C1(n3754), .Y(n5914) );
  AOI22X1TS U3312 ( .A0(n390), .A1(n813), .B0(n4008), .B1(n792), .Y(n5949) );
  AOI222XLTS U3313 ( .A0(n273), .A1(n94), .B0(n4165), .B1(n824), .C0(n4322), 
        .C1(n3750), .Y(n5948) );
  AOI22X1TS U3314 ( .A0(n408), .A1(n812), .B0(n3981), .B1(n790), .Y(n5967) );
  AOI222XLTS U3315 ( .A0(n274), .A1(n95), .B0(n4138), .B1(n822), .C0(n4295), 
        .C1(n3747), .Y(n5966) );
  AOI22X1TS U3316 ( .A0(n3927), .A1(n3439), .B0(n4396), .B1(n3668), .Y(n6211)
         );
  AOI222XLTS U3317 ( .A0(n4083), .A1(n3487), .B0(n137), .B1(n3482), .C0(n4240), 
        .C1(n3458), .Y(n6210) );
  AOI22X1TS U3318 ( .A0(n3921), .A1(n3439), .B0(n4390), .B1(n3668), .Y(n6215)
         );
  AOI222XLTS U3319 ( .A0(n4077), .A1(n3487), .B0(n129), .B1(n3482), .C0(n4234), 
        .C1(n3458), .Y(n6214) );
  AOI22X1TS U3320 ( .A0(n3918), .A1(n3445), .B0(n4387), .B1(n3668), .Y(n6221)
         );
  AOI222XLTS U3321 ( .A0(n4074), .A1(n3499), .B0(n124), .B1(n3482), .C0(n4231), 
        .C1(n3463), .Y(n6220) );
  AOI22X1TS U3322 ( .A0(n348), .A1(n813), .B0(n4071), .B1(n801), .Y(n5907) );
  AOI222XLTS U3323 ( .A0(n234), .A1(n96), .B0(n4228), .B1(n829), .C0(n4385), 
        .C1(n3752), .Y(n5906) );
  AOI22X1TS U3324 ( .A0(n362), .A1(n808), .B0(n4050), .B1(n795), .Y(n5921) );
  AOI222XLTS U3325 ( .A0(n289), .A1(n97), .B0(n4207), .B1(n834), .C0(n4364), 
        .C1(n3757), .Y(n5920) );
  AOI22X1TS U3326 ( .A0(n366), .A1(n808), .B0(n4044), .B1(n795), .Y(n5925) );
  AOI222XLTS U3327 ( .A0(n290), .A1(n98), .B0(n4201), .B1(n835), .C0(n4358), 
        .C1(n3759), .Y(n5924) );
  AOI22X1TS U3328 ( .A0(n378), .A1(n810), .B0(n4026), .B1(n794), .Y(n5937) );
  AOI222XLTS U3329 ( .A0(n186), .A1(n99), .B0(n4183), .B1(n827), .C0(n4340), 
        .C1(n3751), .Y(n5936) );
  AOI22X1TS U3330 ( .A0(n398), .A1(n812), .B0(n3996), .B1(n792), .Y(n5957) );
  AOI222XLTS U3331 ( .A0(n274), .A1(n100), .B0(n4153), .B1(n828), .C0(n4310), 
        .C1(n3749), .Y(n5956) );
  AOI22X1TS U3332 ( .A0(n406), .A1(n812), .B0(n3984), .B1(n791), .Y(n5965) );
  AOI222XLTS U3333 ( .A0(n274), .A1(n101), .B0(n4141), .B1(n823), .C0(n4298), 
        .C1(n3748), .Y(n5964) );
  AOI22X1TS U3334 ( .A0(n410), .A1(n813), .B0(n3978), .B1(n790), .Y(n5969) );
  AOI222XLTS U3335 ( .A0(n227), .A1(n102), .B0(n4135), .B1(n822), .C0(n4292), 
        .C1(n3747), .Y(n5968) );
  OAI22X1TS U3336 ( .A0(n332), .A1(n6231), .B0(n155), .B1(n6232), .Y(n2887) );
  OAI22X1TS U3337 ( .A0(n6234), .A1(n6233), .B0(n432), .B1(n6232), .Y(n2888)
         );
  CLKBUFX2TS U3338 ( .A(n5327), .Y(n432) );
  AOI2BB2X1TS U3339 ( .B0(n5538), .B1(n5537), .A0N(n419), .A1N(
        readOutbuffer[3]), .Y(n2566) );
  OAI221XLTS U3340 ( .A0(readIn_SOUTH), .A1(n6324), .B0(n3820), .B1(n5561), 
        .C0(n5560), .Y(n5565) );
  NAND2X1TS U3341 ( .A(n3806), .B(n6337), .Y(n5544) );
  AOI222XLTS U3342 ( .A0(n3812), .A1(n5556), .B0(readIn_SOUTH), .B1(n5555), 
        .C0(n3820), .C1(n5554), .Y(n5557) );
  OAI22X1TS U3343 ( .A0(n543), .A1(n4711), .B0(n5134), .B1(n3539), .Y(n5135)
         );
  NOR4XLTS U3344 ( .A(n5133), .B(n5132), .C(n5131), .D(n5130), .Y(n5134) );
  AO22X1TS U3345 ( .A0(n231), .A1(\requesterAddressbuffer[3][5] ), .B0(
        \requesterAddressbuffer[6][5] ), .B1(n5286), .Y(n5132) );
  OAI2BB2XLTS U3346 ( .B0(n6303), .B1(n3584), .A0N(
        \requesterAddressbuffer[0][5] ), .A1N(n223), .Y(n5133) );
  OAI22X1TS U3347 ( .A0(n543), .A1(n4712), .B0(n5142), .B1(n3539), .Y(n5143)
         );
  NOR4XLTS U3348 ( .A(n5141), .B(n5140), .C(n5139), .D(n5138), .Y(n5142) );
  AO22X1TS U3349 ( .A0(n181), .A1(\requesterAddressbuffer[3][4] ), .B0(
        \requesterAddressbuffer[6][4] ), .B1(n5286), .Y(n5140) );
  OAI2BB2XLTS U3350 ( .B0(n6304), .B1(n3584), .A0N(
        \requesterAddressbuffer[0][4] ), .A1N(n5287), .Y(n5141) );
  OAI22X1TS U3351 ( .A0(n541), .A1(n4713), .B0(n5158), .B1(n3538), .Y(n5159)
         );
  NOR4XLTS U3352 ( .A(n5157), .B(n5156), .C(n5155), .D(n5154), .Y(n5158) );
  AO22X1TS U3353 ( .A0(n231), .A1(\requesterAddressbuffer[3][2] ), .B0(
        \requesterAddressbuffer[6][2] ), .B1(n5286), .Y(n5156) );
  OAI2BB2XLTS U3354 ( .B0(n6283), .B1(n3583), .A0N(
        \requesterAddressbuffer[0][2] ), .A1N(n223), .Y(n5157) );
  OAI22X1TS U3355 ( .A0(n541), .A1(n4714), .B0(n5166), .B1(n3538), .Y(n5167)
         );
  NOR4XLTS U3356 ( .A(n5165), .B(n5164), .C(n5163), .D(n5162), .Y(n5166) );
  AO22X1TS U3357 ( .A0(n181), .A1(\requesterAddressbuffer[3][1] ), .B0(
        \requesterAddressbuffer[6][1] ), .B1(n346), .Y(n5164) );
  OAI2BB2XLTS U3358 ( .B0(n6284), .B1(n3583), .A0N(
        \requesterAddressbuffer[0][1] ), .A1N(n5287), .Y(n5165) );
  OAI22X1TS U3359 ( .A0(n541), .A1(n4838), .B0(n5150), .B1(n3538), .Y(n5151)
         );
  NOR4XLTS U3360 ( .A(n5149), .B(n5148), .C(n5147), .D(n5146), .Y(n5150) );
  AO22X1TS U3361 ( .A0(n231), .A1(\requesterAddressbuffer[3][3] ), .B0(
        \requesterAddressbuffer[6][3] ), .B1(n346), .Y(n5148) );
  OAI2BB2XLTS U3362 ( .B0(n6282), .B1(n3583), .A0N(
        \requesterAddressbuffer[0][3] ), .A1N(n223), .Y(n5149) );
  OAI22X1TS U3363 ( .A0(n541), .A1(n4837), .B0(n5174), .B1(n3538), .Y(n5175)
         );
  NOR4XLTS U3364 ( .A(n5173), .B(n5172), .C(n5171), .D(n5170), .Y(n5174) );
  AO22X1TS U3365 ( .A0(n181), .A1(\requesterAddressbuffer[3][0] ), .B0(
        \requesterAddressbuffer[6][0] ), .B1(n346), .Y(n5172) );
  OAI2BB2XLTS U3366 ( .B0(n6285), .B1(n3583), .A0N(
        \requesterAddressbuffer[0][0] ), .A1N(n5287), .Y(n5173) );
  OAI22X1TS U3367 ( .A0(n4423), .A1(n543), .B0(n4878), .B1(n3536), .Y(n4879)
         );
  NOR4XLTS U3368 ( .A(n4877), .B(n4876), .C(n4875), .D(n4874), .Y(n4878) );
  OAI22X1TS U3369 ( .A0(n4424), .A1(n3568), .B0(n4425), .B1(n3587), .Y(n4877)
         );
  OAI22X1TS U3370 ( .A0(n4426), .A1(n3615), .B0(n4427), .B1(n3630), .Y(n4876)
         );
  OAI22X1TS U3371 ( .A0(n4432), .A1(n557), .B0(n4886), .B1(n3550), .Y(n4887)
         );
  NOR4XLTS U3372 ( .A(n4885), .B(n4884), .C(n4883), .D(n4882), .Y(n4886) );
  OAI22X1TS U3373 ( .A0(n4437), .A1(n3568), .B0(n4433), .B1(n3597), .Y(n4885)
         );
  OAI22X1TS U3374 ( .A0(n4439), .A1(n3624), .B0(n4438), .B1(n3630), .Y(n4884)
         );
  OAI22X1TS U3375 ( .A0(n4441), .A1(n557), .B0(n4894), .B1(n3550), .Y(n4895)
         );
  NOR4XLTS U3376 ( .A(n4893), .B(n4892), .C(n4891), .D(n4890), .Y(n4894) );
  OAI22X1TS U3377 ( .A0(n4448), .A1(n3568), .B0(n4449), .B1(n6315), .Y(n4893)
         );
  OAI22X1TS U3378 ( .A0(n4444), .A1(n3629), .B0(n4446), .B1(n3630), .Y(n4892)
         );
  OAI22X1TS U3379 ( .A0(n4450), .A1(n557), .B0(n4902), .B1(n3548), .Y(n4903)
         );
  NOR4XLTS U3380 ( .A(n4901), .B(n4900), .C(n4899), .D(n4898), .Y(n4902) );
  OAI22X1TS U3381 ( .A0(n4457), .A1(n3568), .B0(n4451), .B1(n3594), .Y(n4901)
         );
  OAI22X1TS U3382 ( .A0(n4455), .A1(n3629), .B0(n4454), .B1(n3630), .Y(n4900)
         );
  OAI22X1TS U3383 ( .A0(n4459), .A1(n557), .B0(n4910), .B1(n3546), .Y(n4911)
         );
  NOR4XLTS U3384 ( .A(n4909), .B(n4908), .C(n4907), .D(n4906), .Y(n4910) );
  OAI22X1TS U3385 ( .A0(n4466), .A1(n3569), .B0(n4462), .B1(n3593), .Y(n4909)
         );
  OAI22X1TS U3386 ( .A0(n4464), .A1(n3621), .B0(n4463), .B1(n3631), .Y(n4908)
         );
  OAI22X1TS U3387 ( .A0(n4468), .A1(n556), .B0(n4918), .B1(n3547), .Y(n4919)
         );
  NOR4XLTS U3388 ( .A(n4917), .B(n4916), .C(n4915), .D(n4914), .Y(n4918) );
  OAI22X1TS U3389 ( .A0(n4473), .A1(n3569), .B0(n4469), .B1(n3596), .Y(n4917)
         );
  OAI22X1TS U3390 ( .A0(n4475), .A1(n3621), .B0(n4474), .B1(n3631), .Y(n4916)
         );
  OAI22X1TS U3391 ( .A0(n4477), .A1(n556), .B0(n4926), .B1(n3550), .Y(n4927)
         );
  NOR4XLTS U3392 ( .A(n4925), .B(n4924), .C(n4923), .D(n4922), .Y(n4926) );
  OAI22X1TS U3393 ( .A0(n4480), .A1(n3569), .B0(n4482), .B1(n3592), .Y(n4925)
         );
  OAI22X1TS U3394 ( .A0(n4479), .A1(n3621), .B0(n4484), .B1(n3631), .Y(n4924)
         );
  OAI22X1TS U3395 ( .A0(n4486), .A1(n556), .B0(n4934), .B1(n3547), .Y(n4935)
         );
  NOR4XLTS U3396 ( .A(n4933), .B(n4932), .C(n4931), .D(n4930), .Y(n4934) );
  OAI22X1TS U3397 ( .A0(n4489), .A1(n3569), .B0(n4487), .B1(n3597), .Y(n4933)
         );
  OAI22X1TS U3398 ( .A0(n4491), .A1(n3621), .B0(n4494), .B1(n3631), .Y(n4932)
         );
  OAI22X1TS U3399 ( .A0(n4495), .A1(n556), .B0(n4942), .B1(n3548), .Y(n4943)
         );
  NOR4XLTS U3400 ( .A(n4941), .B(n4940), .C(n4939), .D(n4938), .Y(n4942) );
  OAI22X1TS U3401 ( .A0(n4502), .A1(n3581), .B0(n4498), .B1(n3597), .Y(n4941)
         );
  OAI22X1TS U3402 ( .A0(n4503), .A1(n3626), .B0(n4496), .B1(n3643), .Y(n4940)
         );
  OAI22X1TS U3403 ( .A0(n4504), .A1(n555), .B0(n4950), .B1(n3545), .Y(n4951)
         );
  NOR4XLTS U3404 ( .A(n4949), .B(n4948), .C(n4947), .D(n4946), .Y(n4950) );
  OAI22X1TS U3405 ( .A0(n4505), .A1(n3578), .B0(n4508), .B1(n3591), .Y(n4949)
         );
  OAI22X1TS U3406 ( .A0(n4507), .A1(n3627), .B0(n4512), .B1(n3640), .Y(n4948)
         );
  OAI22X1TS U3407 ( .A0(n4513), .A1(n555), .B0(n4958), .B1(n3546), .Y(n4959)
         );
  NOR4XLTS U3408 ( .A(n4957), .B(n4956), .C(n4955), .D(n4954), .Y(n4958) );
  OAI22X1TS U3409 ( .A0(n4520), .A1(n3579), .B0(n4519), .B1(n3595), .Y(n4957)
         );
  OAI22X1TS U3410 ( .A0(n4518), .A1(n3627), .B0(n4516), .B1(n3642), .Y(n4956)
         );
  OAI22X1TS U3411 ( .A0(n4522), .A1(n555), .B0(n4966), .B1(n3544), .Y(n4967)
         );
  NOR4XLTS U3412 ( .A(n4965), .B(n4964), .C(n4963), .D(n4962), .Y(n4966) );
  OAI22X1TS U3413 ( .A0(n4529), .A1(n3576), .B0(n4528), .B1(n3595), .Y(n4965)
         );
  OAI22X1TS U3414 ( .A0(n4530), .A1(n3625), .B0(n4523), .B1(n3638), .Y(n4964)
         );
  OAI22X1TS U3415 ( .A0(n4531), .A1(n555), .B0(n4974), .B1(n3544), .Y(n4975)
         );
  NOR4XLTS U3416 ( .A(n4973), .B(n4972), .C(n4971), .D(n4970), .Y(n4974) );
  OAI22X1TS U3417 ( .A0(n4534), .A1(n3580), .B0(n4533), .B1(n3595), .Y(n4973)
         );
  OAI22X1TS U3418 ( .A0(n4538), .A1(n3623), .B0(n4535), .B1(n3641), .Y(n4972)
         );
  OAI22X1TS U3419 ( .A0(n4540), .A1(n554), .B0(n4982), .B1(n3544), .Y(n4983)
         );
  NOR4XLTS U3420 ( .A(n4981), .B(n4980), .C(n4979), .D(n4978), .Y(n4982) );
  OAI22X1TS U3421 ( .A0(n4543), .A1(n3578), .B0(n4541), .B1(n3598), .Y(n4981)
         );
  OAI22X1TS U3422 ( .A0(n4546), .A1(n3625), .B0(n4547), .B1(n6317), .Y(n4980)
         );
  OAI22X1TS U3423 ( .A0(n4549), .A1(n554), .B0(n4990), .B1(n3544), .Y(n4991)
         );
  NOR4XLTS U3424 ( .A(n4989), .B(n4988), .C(n4987), .D(n4986), .Y(n4990) );
  OAI22X1TS U3425 ( .A0(n4552), .A1(n3580), .B0(n4556), .B1(n3598), .Y(n4989)
         );
  OAI22X1TS U3426 ( .A0(n4550), .A1(n3628), .B0(n4557), .B1(n3640), .Y(n4988)
         );
  OAI22X1TS U3427 ( .A0(n4558), .A1(n554), .B0(n4998), .B1(n3543), .Y(n4999)
         );
  NOR4XLTS U3428 ( .A(n4997), .B(n4996), .C(n4995), .D(n4994), .Y(n4998) );
  OAI22X1TS U3429 ( .A0(n4561), .A1(n3579), .B0(n4560), .B1(n3598), .Y(n4997)
         );
  OAI22X1TS U3430 ( .A0(n4559), .A1(n3624), .B0(n4562), .B1(n3641), .Y(n4996)
         );
  OAI22X1TS U3431 ( .A0(n4567), .A1(n554), .B0(n5006), .B1(n3543), .Y(n5007)
         );
  NOR4XLTS U3432 ( .A(n5005), .B(n5004), .C(n5003), .D(n5002), .Y(n5006) );
  OAI22X1TS U3433 ( .A0(n4572), .A1(n3577), .B0(n4574), .B1(n3591), .Y(n5005)
         );
  OAI22X1TS U3434 ( .A0(n4571), .A1(n3620), .B0(n4575), .B1(n3639), .Y(n5004)
         );
  OAI22X1TS U3435 ( .A0(n4576), .A1(n551), .B0(n5014), .B1(n3543), .Y(n5015)
         );
  NOR4XLTS U3436 ( .A(n5013), .B(n5012), .C(n5011), .D(n5010), .Y(n5014) );
  OAI22X1TS U3437 ( .A0(n4579), .A1(n3577), .B0(n4583), .B1(n3588), .Y(n5013)
         );
  OAI22X1TS U3438 ( .A0(n4581), .A1(n3620), .B0(n4582), .B1(n3639), .Y(n5012)
         );
  OAI22X1TS U3439 ( .A0(n4585), .A1(n551), .B0(n5022), .B1(n3543), .Y(n5023)
         );
  NOR4XLTS U3440 ( .A(n5021), .B(n5020), .C(n5019), .D(n5018), .Y(n5022) );
  OAI22X1TS U3441 ( .A0(n4592), .A1(n3581), .B0(n4586), .B1(n3588), .Y(n5021)
         );
  OAI22X1TS U3442 ( .A0(n4589), .A1(n3620), .B0(n4590), .B1(n3642), .Y(n5020)
         );
  OAI22X1TS U3443 ( .A0(n4594), .A1(n551), .B0(n5030), .B1(n3542), .Y(n5031)
         );
  NOR4XLTS U3444 ( .A(n5029), .B(n5028), .C(n5027), .D(n5026), .Y(n5030) );
  OAI22X1TS U3445 ( .A0(n4599), .A1(n3582), .B0(n4598), .B1(n3588), .Y(n5029)
         );
  OAI22X1TS U3446 ( .A0(n4597), .A1(n3620), .B0(n4601), .B1(n3643), .Y(n5028)
         );
  OAI22X1TS U3447 ( .A0(n4603), .A1(n551), .B0(n5038), .B1(n3542), .Y(n5039)
         );
  NOR4XLTS U3448 ( .A(n5037), .B(n5036), .C(n5035), .D(n5034), .Y(n5038) );
  OAI22X1TS U3449 ( .A0(n4604), .A1(n3570), .B0(n4609), .B1(n3588), .Y(n5037)
         );
  OAI22X1TS U3450 ( .A0(n4608), .A1(n3619), .B0(n4611), .B1(n3632), .Y(n5036)
         );
  OAI22X1TS U3451 ( .A0(n4612), .A1(n548), .B0(n5046), .B1(n3542), .Y(n5047)
         );
  NOR4XLTS U3452 ( .A(n5045), .B(n5044), .C(n5043), .D(n5042), .Y(n5046) );
  OAI22X1TS U3453 ( .A0(n4617), .A1(n3570), .B0(n4616), .B1(n3587), .Y(n5045)
         );
  OAI22X1TS U3454 ( .A0(n4615), .A1(n3619), .B0(n4613), .B1(n3632), .Y(n5044)
         );
  OAI22X1TS U3455 ( .A0(n4621), .A1(n548), .B0(n5054), .B1(n3542), .Y(n5055)
         );
  NOR4XLTS U3456 ( .A(n5053), .B(n5052), .C(n5051), .D(n5050), .Y(n5054) );
  OAI22X1TS U3457 ( .A0(n4628), .A1(n3570), .B0(n4626), .B1(n3587), .Y(n5053)
         );
  OAI22X1TS U3458 ( .A0(n4624), .A1(n3619), .B0(n4627), .B1(n3632), .Y(n5052)
         );
  OAI22X1TS U3459 ( .A0(n4630), .A1(n548), .B0(n5062), .B1(n3541), .Y(n5063)
         );
  NOR4XLTS U3460 ( .A(n5061), .B(n5060), .C(n5059), .D(n5058), .Y(n5062) );
  OAI22X1TS U3461 ( .A0(n4637), .A1(n3570), .B0(n4632), .B1(n3587), .Y(n5061)
         );
  OAI22X1TS U3462 ( .A0(n4631), .A1(n3618), .B0(n4638), .B1(n3632), .Y(n5060)
         );
  OAI22X1TS U3463 ( .A0(n4639), .A1(n546), .B0(n5070), .B1(n3541), .Y(n5071)
         );
  NOR4XLTS U3464 ( .A(n5069), .B(n5068), .C(n5067), .D(n5066), .Y(n5070) );
  OAI22X1TS U3465 ( .A0(n4642), .A1(n3571), .B0(n4644), .B1(n3586), .Y(n5069)
         );
  OAI22X1TS U3466 ( .A0(n4646), .A1(n3618), .B0(n4643), .B1(n3633), .Y(n5068)
         );
  OAI22X1TS U3467 ( .A0(n4648), .A1(n546), .B0(n5078), .B1(n3541), .Y(n5079)
         );
  NOR4XLTS U3468 ( .A(n5077), .B(n5076), .C(n5075), .D(n5074), .Y(n5078) );
  OAI22X1TS U3469 ( .A0(n4651), .A1(n3571), .B0(n4654), .B1(n3586), .Y(n5077)
         );
  OAI22X1TS U3470 ( .A0(n4653), .A1(n3618), .B0(n4649), .B1(n3633), .Y(n5076)
         );
  OAI22X1TS U3471 ( .A0(n4657), .A1(n546), .B0(n5086), .B1(n3540), .Y(n5087)
         );
  NOR4XLTS U3472 ( .A(n5085), .B(n5084), .C(n5083), .D(n5082), .Y(n5086) );
  OAI22X1TS U3473 ( .A0(n4664), .A1(n3571), .B0(n4660), .B1(n3586), .Y(n5085)
         );
  OAI22X1TS U3474 ( .A0(n4663), .A1(n3618), .B0(n4661), .B1(n3633), .Y(n5084)
         );
  OAI22X1TS U3475 ( .A0(n4666), .A1(n546), .B0(n5094), .B1(n3540), .Y(n5095)
         );
  NOR4XLTS U3476 ( .A(n5093), .B(n5092), .C(n5091), .D(n5090), .Y(n5094) );
  OAI22X1TS U3477 ( .A0(n4667), .A1(n3571), .B0(n4671), .B1(n3586), .Y(n5093)
         );
  OAI22X1TS U3478 ( .A0(n4670), .A1(n3617), .B0(n4673), .B1(n3633), .Y(n5092)
         );
  OAI22X1TS U3479 ( .A0(n4675), .A1(n545), .B0(n5102), .B1(n3540), .Y(n5103)
         );
  NOR4XLTS U3480 ( .A(n5101), .B(n5100), .C(n5099), .D(n5098), .Y(n5102) );
  OAI22X1TS U3481 ( .A0(n4678), .A1(n3572), .B0(n4682), .B1(n3585), .Y(n5101)
         );
  OAI22X1TS U3482 ( .A0(n4680), .A1(n3617), .B0(n4677), .B1(n3634), .Y(n5100)
         );
  OAI22X1TS U3483 ( .A0(n4684), .A1(n545), .B0(n5110), .B1(n3540), .Y(n5111)
         );
  NOR4XLTS U3484 ( .A(n5109), .B(n5108), .C(n5107), .D(n5106), .Y(n5110) );
  OAI22X1TS U3485 ( .A0(n4691), .A1(n3572), .B0(n4687), .B1(n3585), .Y(n5109)
         );
  OAI22X1TS U3486 ( .A0(n4690), .A1(n3617), .B0(n4692), .B1(n3634), .Y(n5108)
         );
  OAI22X1TS U3487 ( .A0(n4693), .A1(n545), .B0(n5118), .B1(n3539), .Y(n5119)
         );
  NOR4XLTS U3488 ( .A(n5117), .B(n5116), .C(n5115), .D(n5114), .Y(n5118) );
  OAI22X1TS U3489 ( .A0(n4700), .A1(n3572), .B0(n4695), .B1(n3585), .Y(n5117)
         );
  OAI22X1TS U3490 ( .A0(n4694), .A1(n3617), .B0(n4696), .B1(n3634), .Y(n5116)
         );
  OAI22X1TS U3491 ( .A0(n4702), .A1(n545), .B0(n5126), .B1(n3539), .Y(n5127)
         );
  NOR4XLTS U3492 ( .A(n5125), .B(n5124), .C(n5123), .D(n5122), .Y(n5126) );
  OAI22X1TS U3493 ( .A0(n4707), .A1(n3572), .B0(n4706), .B1(n3585), .Y(n5125)
         );
  OAI22X1TS U3494 ( .A0(n4703), .A1(n3616), .B0(n4708), .B1(n3634), .Y(n5124)
         );
  OAI22X1TS U3495 ( .A0(n4715), .A1(n544), .B0(n5182), .B1(n3537), .Y(n5183)
         );
  NOR4XLTS U3496 ( .A(n5181), .B(n5180), .C(n5179), .D(n5178), .Y(n5182) );
  OAI22X1TS U3497 ( .A0(n4716), .A1(n3573), .B0(n4718), .B1(n3594), .Y(n5181)
         );
  OAI22X1TS U3498 ( .A0(n4722), .A1(n3616), .B0(n4720), .B1(n3635), .Y(n5180)
         );
  OAI22X1TS U3499 ( .A0(n4724), .A1(n544), .B0(n5190), .B1(n3537), .Y(n5191)
         );
  NOR4XLTS U3500 ( .A(n5189), .B(n5188), .C(n5187), .D(n5186), .Y(n5190) );
  OAI22X1TS U3501 ( .A0(n4728), .A1(n3573), .B0(n4729), .B1(n3594), .Y(n5189)
         );
  OAI22X1TS U3502 ( .A0(n4727), .A1(n3616), .B0(n4731), .B1(n3635), .Y(n5188)
         );
  OAI22X1TS U3503 ( .A0(n4733), .A1(n548), .B0(n5198), .B1(n3537), .Y(n5199)
         );
  NOR4XLTS U3504 ( .A(n5197), .B(n5196), .C(n5195), .D(n5194), .Y(n5198) );
  OAI22X1TS U3505 ( .A0(n4736), .A1(n3573), .B0(n4738), .B1(n3593), .Y(n5197)
         );
  OAI22X1TS U3506 ( .A0(n4740), .A1(n3616), .B0(n4734), .B1(n3635), .Y(n5196)
         );
  OAI22X1TS U3507 ( .A0(n4742), .A1(n544), .B0(n5206), .B1(n3537), .Y(n5207)
         );
  NOR4XLTS U3508 ( .A(n5205), .B(n5204), .C(n5203), .D(n5202), .Y(n5206) );
  OAI22X1TS U3509 ( .A0(n4747), .A1(n3573), .B0(n4743), .B1(n3584), .Y(n5205)
         );
  OAI22X1TS U3510 ( .A0(n4744), .A1(n3615), .B0(n4745), .B1(n3635), .Y(n5204)
         );
  OAI22X1TS U3511 ( .A0(n4751), .A1(n543), .B0(n5214), .B1(n3536), .Y(n5215)
         );
  NOR4XLTS U3512 ( .A(n5213), .B(n5212), .C(n5211), .D(n5210), .Y(n5214) );
  OAI22X1TS U3513 ( .A0(n4752), .A1(n3574), .B0(n4756), .B1(n3592), .Y(n5213)
         );
  OAI22X1TS U3514 ( .A0(n4758), .A1(n3615), .B0(n4754), .B1(n3636), .Y(n5212)
         );
  OAI22X1TS U3515 ( .A0(n4760), .A1(n544), .B0(n5223), .B1(n3536), .Y(n5224)
         );
  NOR4XLTS U3516 ( .A(n5222), .B(n5221), .C(n5220), .D(n5219), .Y(n5223) );
  OAI22X1TS U3517 ( .A0(n4766), .A1(n3574), .B0(n4761), .B1(n3584), .Y(n5222)
         );
  OAI22X1TS U3518 ( .A0(n4765), .A1(n3615), .B0(n4763), .B1(n3636), .Y(n5221)
         );
  OAI221XLTS U3519 ( .A0(n5311), .A1(n5310), .B0(n5309), .B1(n5308), .C0(n4422), .Y(n5312) );
  OAI211X1TS U3520 ( .A0(n3567), .A1(n17), .B0(n4834), .C0(n5302), .Y(n5310)
         );
  OAI221XLTS U3521 ( .A0(n3576), .A1(n26), .B0(n3638), .B1(n11), .C0(n5300), 
        .Y(n5311) );
  OAI211X1TS U3522 ( .A0(n255), .A1(n458), .B0(n5233), .C0(n5232), .Y(n2441)
         );
  AOI22X1TS U3523 ( .A0(n411), .A1(n5231), .B0(n561), .B1(
        destinationAddressOut[13]), .Y(n5233) );
  AOI222XLTS U3524 ( .A0(n339), .A1(n4288), .B0(n480), .B1(n4132), .C0(n472), 
        .C1(destinationAddressIn_WEST[13]), .Y(n5232) );
  NAND4X1TS U3525 ( .A(n5230), .B(n5229), .C(n5228), .D(n5227), .Y(n5231) );
  OAI211X1TS U3526 ( .A0(n246), .A1(n458), .B0(n5240), .C0(n5239), .Y(n2442)
         );
  AOI22X1TS U3527 ( .A0(n412), .A1(n5238), .B0(n561), .B1(
        destinationAddressOut[12]), .Y(n5240) );
  AOI222XLTS U3528 ( .A0(n338), .A1(n4285), .B0(n480), .B1(n4129), .C0(n475), 
        .C1(destinationAddressIn_WEST[12]), .Y(n5239) );
  NAND4X1TS U3529 ( .A(n5237), .B(n5236), .C(n5235), .D(n5234), .Y(n5238) );
  OAI211X1TS U3530 ( .A0(n258), .A1(n458), .B0(n5247), .C0(n5246), .Y(n2443)
         );
  AOI22X1TS U3531 ( .A0(n412), .A1(n5245), .B0(n561), .B1(
        destinationAddressOut[11]), .Y(n5247) );
  AOI222XLTS U3532 ( .A0(n339), .A1(n4282), .B0(n480), .B1(n4126), .C0(n475), 
        .C1(destinationAddressIn_WEST[11]), .Y(n5246) );
  NAND4X1TS U3533 ( .A(n5244), .B(n5243), .C(n5242), .D(n5241), .Y(n5245) );
  OAI211X1TS U3534 ( .A0(n249), .A1(n459), .B0(n5254), .C0(n5253), .Y(n2444)
         );
  AOI22X1TS U3535 ( .A0(n411), .A1(n5252), .B0(n561), .B1(
        destinationAddressOut[10]), .Y(n5254) );
  AOI222XLTS U3536 ( .A0(n338), .A1(n4279), .B0(n480), .B1(n4123), .C0(n474), 
        .C1(destinationAddressIn_WEST[10]), .Y(n5253) );
  NAND4X1TS U3537 ( .A(n5251), .B(n5250), .C(n5249), .D(n5248), .Y(n5252) );
  OAI211X1TS U3538 ( .A0(n252), .A1(n459), .B0(n5261), .C0(n5260), .Y(n2445)
         );
  AOI22X1TS U3539 ( .A0(n412), .A1(n5259), .B0(n562), .B1(
        destinationAddressOut[9]), .Y(n5261) );
  AOI222XLTS U3540 ( .A0(n339), .A1(n4276), .B0(n479), .B1(n4120), .C0(n478), 
        .C1(destinationAddressIn_WEST[9]), .Y(n5260) );
  NAND4X1TS U3541 ( .A(n5258), .B(n5257), .C(n5256), .D(n5255), .Y(n5259) );
  OAI211X1TS U3542 ( .A0(n261), .A1(n459), .B0(n5268), .C0(n5267), .Y(n2446)
         );
  AOI22X1TS U3543 ( .A0(n411), .A1(n5266), .B0(n562), .B1(
        destinationAddressOut[8]), .Y(n5268) );
  AOI222XLTS U3544 ( .A0(n338), .A1(n4273), .B0(n479), .B1(n4117), .C0(n477), 
        .C1(destinationAddressIn_WEST[8]), .Y(n5267) );
  NAND4X1TS U3545 ( .A(n5265), .B(n5264), .C(n5263), .D(n5262), .Y(n5266) );
  OAI211X1TS U3546 ( .A0(n240), .A1(n460), .B0(n5275), .C0(n5274), .Y(n2447)
         );
  AOI22X1TS U3547 ( .A0(n411), .A1(n5273), .B0(n562), .B1(
        destinationAddressOut[7]), .Y(n5275) );
  AOI222XLTS U3548 ( .A0(n339), .A1(n4270), .B0(n479), .B1(n4114), .C0(n476), 
        .C1(n3957), .Y(n5274) );
  NAND4X1TS U3549 ( .A(n5272), .B(n5271), .C(n5270), .D(n5269), .Y(n5273) );
  OAI211X1TS U3550 ( .A0(n243), .A1(n460), .B0(n5285), .C0(n5284), .Y(n2448)
         );
  AOI22X1TS U3551 ( .A0(n412), .A1(n5280), .B0(n562), .B1(
        destinationAddressOut[6]), .Y(n5285) );
  AOI222XLTS U3552 ( .A0(n338), .A1(n4267), .B0(n479), .B1(n4111), .C0(n473), 
        .C1(n3954), .Y(n5284) );
  NAND4X1TS U3553 ( .A(n5279), .B(n5278), .C(n5277), .D(n5276), .Y(n5280) );
  OAI211X1TS U3554 ( .A0(n4229), .A1(n3533), .B0(n4881), .C0(n4880), .Y(n2397)
         );
  AOI22X1TS U3555 ( .A0(n444), .A1(n348), .B0(n476), .B1(n3915), .Y(n4881) );
  AOI221X1TS U3556 ( .A0(n447), .A1(n4383), .B0(n493), .B1(n4072), .C0(n4879), 
        .Y(n4880) );
  OAI211X1TS U3557 ( .A0(n4226), .A1(n3532), .B0(n4889), .C0(n4888), .Y(n2398)
         );
  AOI22X1TS U3558 ( .A0(n443), .A1(n350), .B0(n472), .B1(n3912), .Y(n4889) );
  AOI221X1TS U3559 ( .A0(n447), .A1(n4380), .B0(n491), .B1(n4069), .C0(n4887), 
        .Y(n4888) );
  OAI211X1TS U3560 ( .A0(n4223), .A1(n3534), .B0(n4897), .C0(n4896), .Y(n2399)
         );
  AOI22X1TS U3561 ( .A0(n445), .A1(n352), .B0(n474), .B1(n3909), .Y(n4897) );
  AOI221X1TS U3562 ( .A0(n447), .A1(n4377), .B0(n491), .B1(n4066), .C0(n4895), 
        .Y(n4896) );
  OAI211X1TS U3563 ( .A0(n4220), .A1(n3535), .B0(n4905), .C0(n4904), .Y(n2400)
         );
  AOI22X1TS U3564 ( .A0(n5218), .A1(n354), .B0(n476), .B1(n3906), .Y(n4905) );
  AOI221X1TS U3565 ( .A0(n447), .A1(n4374), .B0(n5282), .B1(n4063), .C0(n4903), 
        .Y(n4904) );
  OAI211X1TS U3566 ( .A0(n4217), .A1(n3522), .B0(n4913), .C0(n4912), .Y(n2401)
         );
  AOI22X1TS U3567 ( .A0(n433), .A1(n356), .B0(n476), .B1(n3903), .Y(n4913) );
  AOI221X1TS U3568 ( .A0(n448), .A1(n4371), .B0(n5282), .B1(n4060), .C0(n4911), 
        .Y(n4912) );
  OAI211X1TS U3569 ( .A0(n4214), .A1(n3522), .B0(n4921), .C0(n4920), .Y(n2402)
         );
  AOI22X1TS U3570 ( .A0(n433), .A1(n358), .B0(n473), .B1(n3900), .Y(n4921) );
  AOI221X1TS U3571 ( .A0(n448), .A1(n4368), .B0(n492), .B1(n4057), .C0(n4919), 
        .Y(n4920) );
  OAI211X1TS U3572 ( .A0(n4211), .A1(n3522), .B0(n4929), .C0(n4928), .Y(n2403)
         );
  AOI22X1TS U3573 ( .A0(n433), .A1(n360), .B0(n5281), .B1(n3897), .Y(n4929) );
  AOI221X1TS U3574 ( .A0(n448), .A1(n4365), .B0(n493), .B1(n4054), .C0(n4927), 
        .Y(n4928) );
  OAI211X1TS U3575 ( .A0(n4208), .A1(n3522), .B0(n4937), .C0(n4936), .Y(n2404)
         );
  AOI22X1TS U3576 ( .A0(n433), .A1(n362), .B0(n5281), .B1(n3894), .Y(n4937) );
  AOI221X1TS U3577 ( .A0(n448), .A1(n4362), .B0(n494), .B1(n4051), .C0(n4935), 
        .Y(n4936) );
  OAI211X1TS U3578 ( .A0(n4205), .A1(n3531), .B0(n4945), .C0(n4944), .Y(n2405)
         );
  AOI22X1TS U3579 ( .A0(n444), .A1(n364), .B0(n463), .B1(n3891), .Y(n4945) );
  AOI221X1TS U3580 ( .A0(n449), .A1(n4359), .B0(n489), .B1(n4048), .C0(n4943), 
        .Y(n4944) );
  OAI211X1TS U3581 ( .A0(n4202), .A1(n3530), .B0(n4953), .C0(n4952), .Y(n2406)
         );
  AOI22X1TS U3582 ( .A0(n5218), .A1(n366), .B0(n463), .B1(n3888), .Y(n4953) );
  AOI221X1TS U3583 ( .A0(n449), .A1(n4356), .B0(n490), .B1(n4045), .C0(n4951), 
        .Y(n4952) );
  OAI211X1TS U3584 ( .A0(n4199), .A1(n3529), .B0(n4961), .C0(n4960), .Y(n2407)
         );
  AOI22X1TS U3585 ( .A0(n441), .A1(n368), .B0(n463), .B1(n3885), .Y(n4961) );
  AOI221X1TS U3586 ( .A0(n449), .A1(n4353), .B0(n493), .B1(n4042), .C0(n4959), 
        .Y(n4960) );
  OAI211X1TS U3587 ( .A0(n4196), .A1(n3533), .B0(n4969), .C0(n4968), .Y(n2408)
         );
  AOI22X1TS U3588 ( .A0(n440), .A1(n370), .B0(n463), .B1(n3882), .Y(n4969) );
  AOI221X1TS U3589 ( .A0(n449), .A1(n4350), .B0(n489), .B1(n4039), .C0(n4967), 
        .Y(n4968) );
  OAI211X1TS U3590 ( .A0(n4193), .A1(n3532), .B0(n4977), .C0(n4976), .Y(n2409)
         );
  AOI22X1TS U3591 ( .A0(n443), .A1(n372), .B0(n464), .B1(n3879), .Y(n4977) );
  AOI221X1TS U3592 ( .A0(n450), .A1(n4347), .B0(n488), .B1(n4036), .C0(n4975), 
        .Y(n4976) );
  OAI211X1TS U3593 ( .A0(n4190), .A1(n3532), .B0(n4985), .C0(n4984), .Y(n2410)
         );
  AOI22X1TS U3594 ( .A0(n443), .A1(n374), .B0(n464), .B1(n3876), .Y(n4985) );
  AOI221X1TS U3595 ( .A0(n450), .A1(n4344), .B0(n488), .B1(n4033), .C0(n4983), 
        .Y(n4984) );
  OAI211X1TS U3596 ( .A0(n4187), .A1(n3533), .B0(n4993), .C0(n4992), .Y(n2411)
         );
  AOI22X1TS U3597 ( .A0(n442), .A1(n376), .B0(n464), .B1(n3873), .Y(n4993) );
  AOI221X1TS U3598 ( .A0(n450), .A1(n4341), .B0(n488), .B1(n4030), .C0(n4991), 
        .Y(n4992) );
  OAI211X1TS U3599 ( .A0(n4184), .A1(n3534), .B0(n5001), .C0(n5000), .Y(n2412)
         );
  AOI22X1TS U3600 ( .A0(n445), .A1(n378), .B0(n464), .B1(n3870), .Y(n5001) );
  AOI221X1TS U3601 ( .A0(n450), .A1(n4338), .B0(n488), .B1(n4027), .C0(n4999), 
        .Y(n5000) );
  OAI211X1TS U3602 ( .A0(n4181), .A1(n3532), .B0(n5009), .C0(n5008), .Y(n2413)
         );
  AOI22X1TS U3603 ( .A0(n446), .A1(n380), .B0(n465), .B1(n3867), .Y(n5009) );
  AOI221X1TS U3604 ( .A0(n451), .A1(n4335), .B0(n487), .B1(n4024), .C0(n5007), 
        .Y(n5008) );
  OAI211X1TS U3605 ( .A0(n4178), .A1(n3531), .B0(n5017), .C0(n5016), .Y(n2414)
         );
  AOI22X1TS U3606 ( .A0(n443), .A1(n382), .B0(n465), .B1(n3864), .Y(n5017) );
  AOI221X1TS U3607 ( .A0(n451), .A1(n4332), .B0(n487), .B1(n4021), .C0(n5015), 
        .Y(n5016) );
  OAI211X1TS U3608 ( .A0(n4175), .A1(n3530), .B0(n5025), .C0(n5024), .Y(n2415)
         );
  AOI22X1TS U3609 ( .A0(n441), .A1(n384), .B0(n465), .B1(n3861), .Y(n5025) );
  AOI221X1TS U3610 ( .A0(n451), .A1(n4329), .B0(n487), .B1(n4018), .C0(n5023), 
        .Y(n5024) );
  OAI211X1TS U3611 ( .A0(n4172), .A1(n3529), .B0(n5033), .C0(n5032), .Y(n2416)
         );
  AOI22X1TS U3612 ( .A0(n440), .A1(n386), .B0(n465), .B1(n3858), .Y(n5033) );
  AOI221X1TS U3613 ( .A0(n451), .A1(n4326), .B0(n487), .B1(n4015), .C0(n5031), 
        .Y(n5032) );
  OAI211X1TS U3614 ( .A0(n4169), .A1(n3523), .B0(n5041), .C0(n5040), .Y(n2417)
         );
  AOI22X1TS U3615 ( .A0(n434), .A1(n388), .B0(n466), .B1(n3855), .Y(n5041) );
  AOI221X1TS U3616 ( .A0(n452), .A1(n4323), .B0(n486), .B1(n4012), .C0(n5039), 
        .Y(n5040) );
  OAI211X1TS U3617 ( .A0(n4166), .A1(n3523), .B0(n5049), .C0(n5048), .Y(n2418)
         );
  AOI22X1TS U3618 ( .A0(n434), .A1(n390), .B0(n466), .B1(n3852), .Y(n5049) );
  AOI221X1TS U3619 ( .A0(n452), .A1(n4320), .B0(n486), .B1(n4009), .C0(n5047), 
        .Y(n5048) );
  OAI211X1TS U3620 ( .A0(n4163), .A1(n3523), .B0(n5057), .C0(n5056), .Y(n2419)
         );
  AOI22X1TS U3621 ( .A0(n434), .A1(n392), .B0(n466), .B1(n3849), .Y(n5057) );
  AOI221X1TS U3622 ( .A0(n452), .A1(n4317), .B0(n486), .B1(n4006), .C0(n5055), 
        .Y(n5056) );
  OAI211X1TS U3623 ( .A0(n4160), .A1(n3523), .B0(n5065), .C0(n5064), .Y(n2420)
         );
  AOI22X1TS U3624 ( .A0(n434), .A1(n394), .B0(n466), .B1(n3846), .Y(n5065) );
  AOI221X1TS U3625 ( .A0(n452), .A1(n4314), .B0(n486), .B1(n4003), .C0(n5063), 
        .Y(n5064) );
  OAI211X1TS U3626 ( .A0(n4157), .A1(n3524), .B0(n5073), .C0(n5072), .Y(n2421)
         );
  AOI22X1TS U3627 ( .A0(n435), .A1(n396), .B0(n467), .B1(n3843), .Y(n5073) );
  AOI221X1TS U3628 ( .A0(n453), .A1(n4311), .B0(n485), .B1(n4000), .C0(n5071), 
        .Y(n5072) );
  OAI211X1TS U3629 ( .A0(n4154), .A1(n3524), .B0(n5081), .C0(n5080), .Y(n2422)
         );
  AOI22X1TS U3630 ( .A0(n435), .A1(n398), .B0(n467), .B1(n3840), .Y(n5081) );
  AOI221X1TS U3631 ( .A0(n453), .A1(n4308), .B0(n485), .B1(n3997), .C0(n5079), 
        .Y(n5080) );
  OAI211X1TS U3632 ( .A0(n4151), .A1(n3524), .B0(n5089), .C0(n5088), .Y(n2423)
         );
  AOI22X1TS U3633 ( .A0(n435), .A1(n400), .B0(n467), .B1(n3837), .Y(n5089) );
  AOI221X1TS U3634 ( .A0(n453), .A1(n4305), .B0(n485), .B1(n3994), .C0(n5087), 
        .Y(n5088) );
  OAI211X1TS U3635 ( .A0(n4148), .A1(n3524), .B0(n5097), .C0(n5096), .Y(n2424)
         );
  AOI22X1TS U3636 ( .A0(n435), .A1(n402), .B0(n467), .B1(n3834), .Y(n5097) );
  AOI221X1TS U3637 ( .A0(n453), .A1(n4302), .B0(n485), .B1(n3991), .C0(n5095), 
        .Y(n5096) );
  OAI211X1TS U3638 ( .A0(n4145), .A1(n3525), .B0(n5105), .C0(n5104), .Y(n2425)
         );
  AOI22X1TS U3639 ( .A0(n436), .A1(n404), .B0(n468), .B1(n3831), .Y(n5105) );
  AOI221X1TS U3640 ( .A0(n454), .A1(n4299), .B0(n484), .B1(n3988), .C0(n5103), 
        .Y(n5104) );
  OAI211X1TS U3641 ( .A0(n4142), .A1(n3525), .B0(n5113), .C0(n5112), .Y(n2426)
         );
  AOI22X1TS U3642 ( .A0(n436), .A1(n406), .B0(n468), .B1(n3828), .Y(n5113) );
  AOI221X1TS U3643 ( .A0(n454), .A1(n4296), .B0(n484), .B1(n3985), .C0(n5111), 
        .Y(n5112) );
  OAI211X1TS U3644 ( .A0(n4139), .A1(n3525), .B0(n5121), .C0(n5120), .Y(n2427)
         );
  AOI22X1TS U3645 ( .A0(n436), .A1(n408), .B0(n468), .B1(n3825), .Y(n5121) );
  AOI221X1TS U3646 ( .A0(n454), .A1(n4293), .B0(n484), .B1(n3982), .C0(n5119), 
        .Y(n5120) );
  OAI211X1TS U3647 ( .A0(n4136), .A1(n3525), .B0(n5129), .C0(n5128), .Y(n2428)
         );
  AOI22X1TS U3648 ( .A0(n436), .A1(n410), .B0(n468), .B1(n3822), .Y(n5129) );
  AOI221X1TS U3649 ( .A0(n454), .A1(n4290), .B0(n484), .B1(n3979), .C0(n5127), 
        .Y(n5128) );
  OAI211X1TS U3650 ( .A0(n4247), .A1(n3526), .B0(n5137), .C0(n5136), .Y(n2429)
         );
  AOI22X1TS U3651 ( .A0(n437), .A1(n145), .B0(n469), .B1(n3933), .Y(n5137) );
  AOI221X1TS U3652 ( .A0(n455), .A1(n4401), .B0(n483), .B1(n4090), .C0(n5135), 
        .Y(n5136) );
  OAI211X1TS U3653 ( .A0(n4244), .A1(n3526), .B0(n5145), .C0(n5144), .Y(n2430)
         );
  AOI22X1TS U3654 ( .A0(n437), .A1(n140), .B0(n469), .B1(n3930), .Y(n5145) );
  AOI221X1TS U3655 ( .A0(n455), .A1(n4398), .B0(n483), .B1(n4087), .C0(n5143), 
        .Y(n5144) );
  OAI211X1TS U3656 ( .A0(n4238), .A1(n3526), .B0(n5161), .C0(n5160), .Y(n2432)
         );
  AOI22X1TS U3657 ( .A0(n437), .A1(n116), .B0(n469), .B1(n3924), .Y(n5161) );
  AOI221X1TS U3658 ( .A0(n455), .A1(n4392), .B0(n483), .B1(n4081), .C0(n5159), 
        .Y(n5160) );
  OAI211X1TS U3659 ( .A0(n4235), .A1(n3527), .B0(n5169), .C0(n5168), .Y(n2433)
         );
  AOI22X1TS U3660 ( .A0(n438), .A1(n115), .B0(n470), .B1(n3921), .Y(n5169) );
  AOI221X1TS U3661 ( .A0(n456), .A1(n4389), .B0(n482), .B1(n4078), .C0(n5167), 
        .Y(n5168) );
  OAI211X1TS U3662 ( .A0(n4265), .A1(n3527), .B0(n5185), .C0(n5184), .Y(n2435)
         );
  AOI22X1TS U3663 ( .A0(n438), .A1(n146), .B0(n470), .B1(n3951), .Y(n5185) );
  AOI221X1TS U3664 ( .A0(n456), .A1(n4419), .B0(n482), .B1(n4108), .C0(n5183), 
        .Y(n5184) );
  OAI211X1TS U3665 ( .A0(n4262), .A1(n3527), .B0(n5193), .C0(n5192), .Y(n2436)
         );
  AOI22X1TS U3666 ( .A0(n438), .A1(n141), .B0(n470), .B1(n3948), .Y(n5193) );
  AOI221X1TS U3667 ( .A0(n456), .A1(n4416), .B0(n482), .B1(n4105), .C0(n5191), 
        .Y(n5192) );
  OAI211X1TS U3668 ( .A0(n4259), .A1(n3528), .B0(n5201), .C0(n5200), .Y(n2437)
         );
  AOI22X1TS U3669 ( .A0(n439), .A1(n117), .B0(n471), .B1(n3945), .Y(n5201) );
  AOI221X1TS U3670 ( .A0(n457), .A1(n4413), .B0(n481), .B1(n4102), .C0(n5199), 
        .Y(n5200) );
  OAI211X1TS U3671 ( .A0(n4256), .A1(n3528), .B0(n5209), .C0(n5208), .Y(n2438)
         );
  AOI22X1TS U3672 ( .A0(n439), .A1(n132), .B0(n471), .B1(n3942), .Y(n5209) );
  AOI221X1TS U3673 ( .A0(n457), .A1(n4410), .B0(n481), .B1(n4099), .C0(n5207), 
        .Y(n5208) );
  OAI211X1TS U3674 ( .A0(n4253), .A1(n3528), .B0(n5217), .C0(n5216), .Y(n2439)
         );
  AOI22X1TS U3675 ( .A0(n439), .A1(n128), .B0(n471), .B1(n3939), .Y(n5217) );
  AOI221X1TS U3676 ( .A0(n457), .A1(n4407), .B0(n481), .B1(n4096), .C0(n5215), 
        .Y(n5216) );
  OAI211X1TS U3677 ( .A0(n4250), .A1(n3528), .B0(n5226), .C0(n5225), .Y(n2440)
         );
  AOI22X1TS U3678 ( .A0(n439), .A1(n124), .B0(n471), .B1(n3936), .Y(n5226) );
  AOI221X1TS U3679 ( .A0(n457), .A1(n4404), .B0(n481), .B1(n4093), .C0(n5224), 
        .Y(n5225) );
  OAI211X1TS U3680 ( .A0(n4241), .A1(n3526), .B0(n5153), .C0(n5152), .Y(n2431)
         );
  AOI22X1TS U3681 ( .A0(n437), .A1(n136), .B0(n469), .B1(n3927), .Y(n5153) );
  AOI221X1TS U3682 ( .A0(n455), .A1(n4395), .B0(n483), .B1(n4084), .C0(n5151), 
        .Y(n5152) );
  OAI211X1TS U3683 ( .A0(n4232), .A1(n3527), .B0(n5177), .C0(n5176), .Y(n2434)
         );
  AOI22X1TS U3684 ( .A0(n438), .A1(n125), .B0(n470), .B1(n3918), .Y(n5177) );
  AOI221X1TS U3685 ( .A0(n456), .A1(n4386), .B0(n482), .B1(n4075), .C0(n5175), 
        .Y(n5176) );
  NOR2X1TS U3686 ( .A(reset), .B(n4834), .Y(n5295) );
  INVX2TS U3687 ( .A(readIn_SOUTH), .Y(n6238) );
  INVX2TS U3688 ( .A(writeIn_NORTH), .Y(n6239) );
  OAI22X1TS U3689 ( .A0(n5296), .A1(n5295), .B0(n5294), .B1(n5293), .Y(n5297)
         );
  AOI31X1TS U3690 ( .A0(n5292), .A1(n5291), .A2(n5290), .B0(reset), .Y(n5296)
         );
  OAI22X1TS U3691 ( .A0(n3818), .A1(n5305), .B0(n3805), .B1(n5307), .Y(n5293)
         );
  OAI22X1TS U3692 ( .A0(n345), .A1(n6313), .B0(n4), .B1(n3541), .Y(n2889) );
  INVX2TS U3693 ( .A(destinationAddressIn_NORTH[7]), .Y(n6241) );
  INVX2TS U3694 ( .A(destinationAddressIn_NORTH[6]), .Y(n6240) );
  INVX2TS U3695 ( .A(destinationAddressIn_NORTH[12]), .Y(n6246) );
  INVX2TS U3696 ( .A(destinationAddressIn_NORTH[10]), .Y(n6244) );
  INVX2TS U3697 ( .A(destinationAddressIn_NORTH[9]), .Y(n6243) );
  INVX2TS U3698 ( .A(destinationAddressIn_NORTH[13]), .Y(n6247) );
  INVX2TS U3699 ( .A(destinationAddressIn_NORTH[11]), .Y(n6245) );
  INVX2TS U3700 ( .A(destinationAddressIn_NORTH[8]), .Y(n6242) );
  NOR2X1TS U3701 ( .A(n6223), .B(n6224), .Y(n2883) );
  AOI21X1TS U3702 ( .A0(n275), .A1(n6222), .B0(n5), .Y(n6223) );
  XNOR2X1TS U3703 ( .A(n4844), .B(n6319), .Y(n6227) );
  XNOR2X1TS U3704 ( .A(n195), .B(n5323), .Y(n4844) );
  OAI22X1TS U3705 ( .A0(n4430), .A1(n3658), .B0(n4431), .B1(n3556), .Y(n4874)
         );
  OAI22X1TS U3706 ( .A0(n4435), .A1(n3653), .B0(n4440), .B1(n3558), .Y(n4882)
         );
  OAI22X1TS U3707 ( .A0(n4442), .A1(n3657), .B0(n4445), .B1(n3558), .Y(n4890)
         );
  OAI22X1TS U3708 ( .A0(n4453), .A1(n3655), .B0(n4452), .B1(n3558), .Y(n4898)
         );
  OAI22X1TS U3709 ( .A0(n4467), .A1(n3655), .B0(n4460), .B1(n3558), .Y(n4906)
         );
  OAI22X1TS U3710 ( .A0(n4471), .A1(n3657), .B0(n4476), .B1(n3557), .Y(n4914)
         );
  OAI22X1TS U3711 ( .A0(n4478), .A1(n3656), .B0(n4483), .B1(n3557), .Y(n4922)
         );
  OAI22X1TS U3712 ( .A0(n4493), .A1(n3653), .B0(n4488), .B1(n3557), .Y(n4930)
         );
  OAI22X1TS U3713 ( .A0(n4500), .A1(n3654), .B0(n4497), .B1(n3557), .Y(n4938)
         );
  OAI22X1TS U3714 ( .A0(n4511), .A1(n3654), .B0(n4509), .B1(n3565), .Y(n4946)
         );
  OAI22X1TS U3715 ( .A0(n4514), .A1(n3656), .B0(n4515), .B1(n3565), .Y(n4954)
         );
  OAI22X1TS U3716 ( .A0(n4527), .A1(n3659), .B0(n4525), .B1(n3564), .Y(n4962)
         );
  OAI22X1TS U3717 ( .A0(n4532), .A1(n3645), .B0(n4536), .B1(n3563), .Y(n4970)
         );
  OAI22X1TS U3718 ( .A0(n4545), .A1(n3645), .B0(n4548), .B1(n3564), .Y(n4978)
         );
  OAI22X1TS U3719 ( .A0(n4554), .A1(n3645), .B0(n4551), .B1(n3566), .Y(n4986)
         );
  OAI22X1TS U3720 ( .A0(n4565), .A1(n3645), .B0(n4566), .B1(n3566), .Y(n4994)
         );
  OAI22X1TS U3721 ( .A0(n4570), .A1(n3646), .B0(n4573), .B1(n3567), .Y(n5002)
         );
  OAI22X1TS U3722 ( .A0(n4577), .A1(n3646), .B0(n4580), .B1(n3561), .Y(n5010)
         );
  OAI22X1TS U3723 ( .A0(n4588), .A1(n3646), .B0(n4593), .B1(n3561), .Y(n5018)
         );
  OAI22X1TS U3724 ( .A0(n4595), .A1(n3646), .B0(n4602), .B1(n3561), .Y(n5026)
         );
  OAI22X1TS U3725 ( .A0(n4610), .A1(n3647), .B0(n4605), .B1(n6314), .Y(n5034)
         );
  OAI22X1TS U3726 ( .A0(n4618), .A1(n3647), .B0(n4619), .B1(n3556), .Y(n5042)
         );
  OAI22X1TS U3727 ( .A0(n4622), .A1(n3647), .B0(n4623), .B1(n3556), .Y(n5050)
         );
  OAI22X1TS U3728 ( .A0(n4635), .A1(n3647), .B0(n4633), .B1(n3556), .Y(n5058)
         );
  OAI22X1TS U3729 ( .A0(n4640), .A1(n3648), .B0(n4647), .B1(n3555), .Y(n5066)
         );
  OAI22X1TS U3730 ( .A0(n4655), .A1(n3648), .B0(n4650), .B1(n3555), .Y(n5074)
         );
  OAI22X1TS U3731 ( .A0(n4662), .A1(n3648), .B0(n4658), .B1(n3555), .Y(n5082)
         );
  OAI22X1TS U3732 ( .A0(n4669), .A1(n3648), .B0(n4674), .B1(n3555), .Y(n5090)
         );
  OAI22X1TS U3733 ( .A0(n4676), .A1(n3649), .B0(n4679), .B1(n3554), .Y(n5098)
         );
  OAI22X1TS U3734 ( .A0(n4689), .A1(n3649), .B0(n4685), .B1(n3554), .Y(n5106)
         );
  OAI22X1TS U3735 ( .A0(n4701), .A1(n3649), .B0(n4697), .B1(n3554), .Y(n5114)
         );
  OAI22X1TS U3736 ( .A0(n4705), .A1(n3649), .B0(n4709), .B1(n3554), .Y(n5122)
         );
  OAI22X1TS U3737 ( .A0(n4719), .A1(n3650), .B0(n4717), .B1(n3553), .Y(n5178)
         );
  OAI22X1TS U3738 ( .A0(n4732), .A1(n3650), .B0(n4726), .B1(n3553), .Y(n5186)
         );
  OAI22X1TS U3739 ( .A0(n4741), .A1(n3650), .B0(n4737), .B1(n3553), .Y(n5194)
         );
  OAI22X1TS U3740 ( .A0(n4749), .A1(n3650), .B0(n4750), .B1(n3552), .Y(n5202)
         );
  OAI22X1TS U3741 ( .A0(n4755), .A1(n3651), .B0(n4759), .B1(n3553), .Y(n5210)
         );
  OAI22X1TS U3742 ( .A0(n4762), .A1(n3651), .B0(n4768), .B1(n3552), .Y(n5219)
         );
  OAI22X1TS U3743 ( .A0(n4428), .A1(n502), .B0(n4429), .B1(n3599), .Y(n4875)
         );
  OAI22X1TS U3744 ( .A0(n4436), .A1(n511), .B0(n4434), .B1(n3609), .Y(n4883)
         );
  OAI22X1TS U3745 ( .A0(n4447), .A1(n536), .B0(n4443), .B1(n3607), .Y(n4891)
         );
  OAI22X1TS U3746 ( .A0(n4458), .A1(n517), .B0(n4456), .B1(n3607), .Y(n4899)
         );
  OAI22X1TS U3747 ( .A0(n4461), .A1(n526), .B0(n4465), .B1(n3607), .Y(n4907)
         );
  OAI22X1TS U3748 ( .A0(n4470), .A1(n517), .B0(n4472), .B1(n3607), .Y(n4915)
         );
  OAI22X1TS U3749 ( .A0(n4485), .A1(n537), .B0(n4481), .B1(n3614), .Y(n4923)
         );
  OAI22X1TS U3750 ( .A0(n4492), .A1(n537), .B0(n4490), .B1(n3611), .Y(n4931)
         );
  OAI22X1TS U3751 ( .A0(n4499), .A1(n537), .B0(n4501), .B1(n3609), .Y(n4939)
         );
  OAI22X1TS U3752 ( .A0(n4510), .A1(n511), .B0(n4506), .B1(n3610), .Y(n4947)
         );
  OAI22X1TS U3753 ( .A0(n4517), .A1(n507), .B0(n4521), .B1(n3613), .Y(n4955)
         );
  OAI22X1TS U3754 ( .A0(n4524), .A1(n507), .B0(n4526), .B1(n3612), .Y(n4963)
         );
  OAI22X1TS U3755 ( .A0(n4537), .A1(n507), .B0(n4539), .B1(n6316), .Y(n4971)
         );
  OAI22X1TS U3756 ( .A0(n4544), .A1(n507), .B0(n4542), .B1(n3611), .Y(n4979)
         );
  OAI22X1TS U3757 ( .A0(n4555), .A1(n505), .B0(n4553), .B1(n3606), .Y(n4987)
         );
  OAI22X1TS U3758 ( .A0(n4563), .A1(n505), .B0(n4564), .B1(n3606), .Y(n4995)
         );
  OAI22X1TS U3759 ( .A0(n4568), .A1(n505), .B0(n4569), .B1(n3606), .Y(n5003)
         );
  OAI22X1TS U3760 ( .A0(n4578), .A1(n505), .B0(n4584), .B1(n3606), .Y(n5011)
         );
  OAI22X1TS U3761 ( .A0(n4591), .A1(n503), .B0(n4587), .B1(n3605), .Y(n5019)
         );
  OAI22X1TS U3762 ( .A0(n4600), .A1(n503), .B0(n4596), .B1(n3605), .Y(n5027)
         );
  OAI22X1TS U3763 ( .A0(n4606), .A1(n503), .B0(n4607), .B1(n3605), .Y(n5035)
         );
  OAI22X1TS U3764 ( .A0(n4614), .A1(n503), .B0(n4620), .B1(n3605), .Y(n5043)
         );
  OAI22X1TS U3765 ( .A0(n4625), .A1(n502), .B0(n4629), .B1(n3604), .Y(n5051)
         );
  OAI22X1TS U3766 ( .A0(n4636), .A1(n502), .B0(n4634), .B1(n3604), .Y(n5059)
         );
  OAI22X1TS U3767 ( .A0(n4645), .A1(n502), .B0(n4641), .B1(n3604), .Y(n5067)
         );
  OAI22X1TS U3768 ( .A0(n4652), .A1(n514), .B0(n4656), .B1(n3603), .Y(n5075)
         );
  OAI22X1TS U3769 ( .A0(n4665), .A1(n514), .B0(n4659), .B1(n3603), .Y(n5083)
         );
  OAI22X1TS U3770 ( .A0(n4672), .A1(n516), .B0(n4668), .B1(n3603), .Y(n5091)
         );
  OAI22X1TS U3771 ( .A0(n4683), .A1(n516), .B0(n4681), .B1(n3603), .Y(n5099)
         );
  OAI22X1TS U3772 ( .A0(n4688), .A1(n501), .B0(n4686), .B1(n3602), .Y(n5107)
         );
  OAI22X1TS U3773 ( .A0(n4698), .A1(n501), .B0(n4699), .B1(n3602), .Y(n5115)
         );
  OAI22X1TS U3774 ( .A0(n4710), .A1(n501), .B0(n4704), .B1(n3602), .Y(n5123)
         );
  OAI22X1TS U3775 ( .A0(n4721), .A1(n499), .B0(n4723), .B1(n3600), .Y(n5179)
         );
  OAI22X1TS U3776 ( .A0(n4730), .A1(n499), .B0(n4725), .B1(n3600), .Y(n5187)
         );
  OAI22X1TS U3777 ( .A0(n4739), .A1(n499), .B0(n4735), .B1(n3600), .Y(n5195)
         );
  OAI22X1TS U3778 ( .A0(n4748), .A1(n496), .B0(n4746), .B1(n3599), .Y(n5203)
         );
  OAI22X1TS U3779 ( .A0(n4757), .A1(n496), .B0(n4753), .B1(n3599), .Y(n5211)
         );
  OAI22X1TS U3780 ( .A0(n4764), .A1(n496), .B0(n4767), .B1(n3599), .Y(n5220)
         );
  NOR3X1TS U3781 ( .A(n4), .B(n195), .C(n147), .Y(n5299) );
  NOR3X1TS U3782 ( .A(n5), .B(n194), .C(n6313), .Y(n5289) );
  NAND3X1TS U3783 ( .A(n276), .B(n335), .C(n3), .Y(n5301) );
  AOI2BB2X1TS U3784 ( .B0(readOutbuffer[3]), .B1(n231), .A0N(n25), .A1N(n509), 
        .Y(n5302) );
  AOI222XLTS U3785 ( .A0(readOutbuffer[4]), .A1(n5299), .B0(readOutbuffer[7]), 
        .B1(n5298), .C0(readOutbuffer[2]), .C1(n179), .Y(n5300) );
  AOI221X1TS U3786 ( .A0(n5289), .A1(writeOutbuffer[1]), .B0(n179), .B1(
        writeOutbuffer[2]), .C0(n5288), .Y(n5290) );
  OAI22X1TS U3787 ( .A0(n18), .A1(n496), .B0(n10), .B1(n3604), .Y(n5288) );
  OA22X1TS U3788 ( .A0(n3559), .A1(n4770), .B0(n3651), .B1(n4769), .Y(n5230)
         );
  OA22X1TS U3789 ( .A0(n3559), .A1(n4778), .B0(n3651), .B1(n4783), .Y(n5237)
         );
  OA22X1TS U3790 ( .A0(n3559), .A1(n4788), .B0(n3652), .B1(n4792), .Y(n5244)
         );
  OA22X1TS U3791 ( .A0(n3559), .A1(n4794), .B0(n3652), .B1(n4797), .Y(n5251)
         );
  OA22X1TS U3792 ( .A0(n3560), .A1(n4806), .B0(n3652), .B1(n4808), .Y(n5258)
         );
  OA22X1TS U3793 ( .A0(n3560), .A1(n4810), .B0(n3652), .B1(n4811), .Y(n5265)
         );
  OA22X1TS U3794 ( .A0(n3560), .A1(n4818), .B0(n3653), .B1(n4824), .Y(n5272)
         );
  OA22X1TS U3795 ( .A0(n3560), .A1(n4830), .B0(n3653), .B1(n4831), .Y(n5279)
         );
  OA22X1TS U3796 ( .A0(n3589), .A1(n4775), .B0(n3574), .B1(n4776), .Y(n5227)
         );
  OA22X1TS U3797 ( .A0(n3589), .A1(n4779), .B0(n3574), .B1(n4777), .Y(n5234)
         );
  OA22X1TS U3798 ( .A0(n3589), .A1(n4785), .B0(n3575), .B1(n4789), .Y(n5241)
         );
  OA22X1TS U3799 ( .A0(n3589), .A1(n4795), .B0(n3575), .B1(n4798), .Y(n5248)
         );
  OA22X1TS U3800 ( .A0(n3590), .A1(n4807), .B0(n3575), .B1(n4803), .Y(n5255)
         );
  OA22X1TS U3801 ( .A0(n3590), .A1(n4813), .B0(n3575), .B1(n4809), .Y(n5262)
         );
  OA22X1TS U3802 ( .A0(n3590), .A1(n4817), .B0(n3576), .B1(n4819), .Y(n5269)
         );
  OA22X1TS U3803 ( .A0(n3590), .A1(n4829), .B0(n3576), .B1(n4832), .Y(n5276)
         );
  OA22X1TS U3804 ( .A0(n3609), .A1(n4772), .B0(n509), .B1(n4774), .Y(n5229) );
  OA22X1TS U3805 ( .A0(n3610), .A1(n4782), .B0(n508), .B1(n4784), .Y(n5236) );
  OA22X1TS U3806 ( .A0(n3612), .A1(n4786), .B0(n5301), .B1(n4790), .Y(n5243)
         );
  AOI2BB2X1TS U3807 ( .B0(n5298), .B1(n431), .A0N(n509), .A1N(n4800), .Y(n5250) );
  OA22X1TS U3808 ( .A0(n3608), .A1(n4805), .B0(n508), .B1(n4804), .Y(n5257) );
  OA22X1TS U3809 ( .A0(n3608), .A1(n4812), .B0(n508), .B1(n4814), .Y(n5264) );
  OA22X1TS U3810 ( .A0(n3608), .A1(n4822), .B0(n508), .B1(n4820), .Y(n5271) );
  OA22X1TS U3811 ( .A0(n3608), .A1(n4828), .B0(n509), .B1(n4826), .Y(n5278) );
  OA22X1TS U3812 ( .A0(n3636), .A1(n4771), .B0(n1), .B1(n4773), .Y(n5228) );
  OA22X1TS U3813 ( .A0(n3636), .A1(n4781), .B0(n3622), .B1(n4780), .Y(n5235)
         );
  OA22X1TS U3814 ( .A0(n3637), .A1(n4791), .B0(n3622), .B1(n4787), .Y(n5242)
         );
  OA22X1TS U3815 ( .A0(n3637), .A1(n4793), .B0(n3623), .B1(n4799), .Y(n5249)
         );
  OA22X1TS U3816 ( .A0(n3637), .A1(n4801), .B0(n3622), .B1(n4802), .Y(n5256)
         );
  OA22X1TS U3817 ( .A0(n3637), .A1(n4815), .B0(n3622), .B1(n4816), .Y(n5263)
         );
  OA22X1TS U3818 ( .A0(n3638), .A1(n4821), .B0(n3623), .B1(n4823), .Y(n5270)
         );
  OA22X1TS U3819 ( .A0(n3638), .A1(n4825), .B0(n3623), .B1(n4827), .Y(n5277)
         );
  AOI22X1TS U3820 ( .A0(n346), .A1(writeOutbuffer[6]), .B0(writeOutbuffer[3]), 
        .B1(n181), .Y(n5292) );
  AOI22X1TS U3821 ( .A0(n5299), .A1(writeOutbuffer[4]), .B0(n223), .B1(
        writeOutbuffer[0]), .Y(n5291) );
  AOI32X1TS U3822 ( .A0(n331), .A1(n189), .A2(n119), .B0(n4839), .B1(
        selectBit_SOUTH), .Y(n4840) );
  AOI21XLTS U3823 ( .A0(n3819), .A1(n5542), .B0(n5541), .Y(n5543) );
  OAI221XLTS U3824 ( .A0(n229), .A1(n237), .B0(n330), .B1(n109), .C0(n5568), 
        .Y(n2571) );
  OAI221XLTS U3825 ( .A0(n5570), .A1(n243), .B0(n4832), .B1(n281), .C0(n5333), 
        .Y(n2458) );
  OAI221XLTS U3826 ( .A0(n230), .A1(n240), .B0(n4819), .B1(n5569), .C0(n5332), 
        .Y(n2457) );
  OAI221XLTS U3827 ( .A0(n229), .A1(n261), .B0(n4809), .B1(n330), .C0(n5331), 
        .Y(n2456) );
  OAI221XLTS U3828 ( .A0(n230), .A1(n251), .B0(n4803), .B1(n5569), .C0(n5330), 
        .Y(n2455) );
  OAI221XLTS U3829 ( .A0(n229), .A1(n248), .B0(n4798), .B1(n330), .C0(n5329), 
        .Y(n2454) );
  OAI221XLTS U3830 ( .A0(n5570), .A1(n257), .B0(n4789), .B1(n5569), .C0(n5328), 
        .Y(n2453) );
  OAI221XLTS U3831 ( .A0(n230), .A1(n245), .B0(n4777), .B1(n330), .C0(n5325), 
        .Y(n2452) );
  OAI221XLTS U3832 ( .A0(n5570), .A1(n254), .B0(n4776), .B1(n205), .C0(n5324), 
        .Y(n2451) );
  NOR2X1TS U3833 ( .A(n5524), .B(n5487), .Y(n5556) );
  NOR2X1TS U3834 ( .A(n6329), .B(n5487), .Y(n5563) );
  AOI32XLTS U3835 ( .A0(n162), .A1(n5529), .A2(n5528), .B0(n198), .B1(n105), 
        .Y(n2565) );
  OAI221XLTS U3836 ( .A0(n270), .A1(n6239), .B0(n199), .B1(n6311), .C0(n5573), 
        .Y(n2573) );
  OAI221XLTS U3837 ( .A0(n5575), .A1(n6240), .B0(n4831), .B1(n5574), .C0(n5377), .Y(n2486) );
  OAI221XLTS U3838 ( .A0(n270), .A1(n6242), .B0(n4811), .B1(n199), .C0(n5375), 
        .Y(n2484) );
  OAI221XLTS U3839 ( .A0(n5575), .A1(n6243), .B0(n4808), .B1(n5574), .C0(n5374), .Y(n2483) );
  OAI221XLTS U3840 ( .A0(n270), .A1(n6244), .B0(n4797), .B1(n329), .C0(n5373), 
        .Y(n2482) );
  OAI221XLTS U3841 ( .A0(n5575), .A1(n6245), .B0(n4792), .B1(n5574), .C0(n5372), .Y(n2481) );
  OAI221XLTS U3842 ( .A0(n270), .A1(n6246), .B0(n4783), .B1(n199), .C0(n5371), 
        .Y(n2480) );
  OAI221XLTS U3843 ( .A0(n269), .A1(n6247), .B0(n4769), .B1(n329), .C0(n5370), 
        .Y(n2479) );
endmodule


module router ( clk, reset, localRouterAddress, destinationAddressIn_NORTH, 
        requesterAddressIn_NORTH, readIn_NORTH, writeIn_NORTH, dataIn_NORTH, 
        destinationAddressOut_NORTH, requesterAddressOut_NORTH, readOut_NORTH, 
        writeOut_NORTH, dataOut_NORTH, destinationAddressIn_SOUTH, 
        requesterAddressIn_SOUTH, readIn_SOUTH, writeIn_SOUTH, dataIn_SOUTH, 
        destinationAddressOut_SOUTH, requesterAddressOut_SOUTH, readOut_SOUTH, 
        writeOut_SOUTH, dataOut_SOUTH, destinationAddressIn_EAST, 
        requesterAddressIn_EAST, readIn_EAST, writeIn_EAST, dataIn_EAST, 
        destinationAddressOut_EAST, requesterAddressOut_EAST, readOut_EAST, 
        writeOut_EAST, dataOut_EAST, destinationAddressIn_WEST, 
        requesterAddressIn_WEST, readIn_WEST, writeIn_WEST, dataIn_WEST, 
        destinationAddressOut_WEST, requesterAddressOut_WEST, readOut_WEST, 
        writeOut_WEST, dataOut_WEST, cacheDataIn_A, cacheAddressIn_A, 
        cacheDataOut_A, memWrite_A, portA_writtenTo, cacheDataIn_B, 
        cacheAddressIn_B, cacheDataOut_B, memWrite_B, portB_writtenTo );
  input [5:0] localRouterAddress;
  input [13:0] destinationAddressIn_NORTH;
  input [5:0] requesterAddressIn_NORTH;
  input [31:0] dataIn_NORTH;
  output [13:0] destinationAddressOut_NORTH;
  output [5:0] requesterAddressOut_NORTH;
  output [31:0] dataOut_NORTH;
  input [13:0] destinationAddressIn_SOUTH;
  input [5:0] requesterAddressIn_SOUTH;
  input [31:0] dataIn_SOUTH;
  output [13:0] destinationAddressOut_SOUTH;
  output [5:0] requesterAddressOut_SOUTH;
  output [31:0] dataOut_SOUTH;
  input [13:0] destinationAddressIn_EAST;
  input [5:0] requesterAddressIn_EAST;
  input [31:0] dataIn_EAST;
  output [13:0] destinationAddressOut_EAST;
  output [5:0] requesterAddressOut_EAST;
  output [31:0] dataOut_EAST;
  input [13:0] destinationAddressIn_WEST;
  input [5:0] requesterAddressIn_WEST;
  input [31:0] dataIn_WEST;
  output [13:0] destinationAddressOut_WEST;
  output [5:0] requesterAddressOut_WEST;
  output [31:0] dataOut_WEST;
  output [31:0] cacheDataIn_A;
  output [7:0] cacheAddressIn_A;
  input [31:0] cacheDataOut_A;
  output [31:0] cacheDataIn_B;
  output [7:0] cacheAddressIn_B;
  input [31:0] cacheDataOut_B;
  input clk, reset, readIn_NORTH, writeIn_NORTH, readIn_SOUTH, writeIn_SOUTH,
         readIn_EAST, writeIn_EAST, readIn_WEST, writeIn_WEST, portA_writtenTo,
         portB_writtenTo;
  output readOut_NORTH, writeOut_NORTH, readOut_SOUTH, writeOut_SOUTH,
         readOut_EAST, writeOut_EAST, readOut_WEST, writeOut_WEST, memWrite_A,
         memWrite_B;
  wire   memRead_NORTH, memWrite_NORTH, memRead_SOUTH, memWrite_SOUTH,
         memRead_EAST, memWrite_EAST, memRead_WEST, memWrite_WEST,
         readReady_NORTH, readReady_SOUTH, readReady_EAST, readReady_WEST,
         readInBuffer_NORTH, writeInBuffer_NORTH, writeInBuffer_SOUTH,
         readInBuffer_EAST, writeInBuffer_EAST, readInBuffer_WEST,
         writeInBuffer_WEST, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366;
  wire   [3:0] outputPortSelect_NORTH;
  wire   [3:0] outputPortSelect_SOUTH;
  wire   [3:0] outputPortSelect_EAST;
  wire   [3:0] outputPortSelect_WEST;
  wire   [13:0] destinationAddressInBuffer_NORTH;
  wire   [5:0] requesterAddressInBuffer_NORTH;
  wire   [31:0] dataInBuffer_NORTH;
  wire   [5:0] cacheRequesterAddress_NORTH;
  wire   [31:0] cacheDataOut_NORTH;
  wire   [13:0] destinationAddressInBuffer_SOUTH;
  wire   [5:0] requesterAddressInBuffer_SOUTH;
  wire   [31:0] dataInBuffer_SOUTH;
  wire   [5:0] cacheRequesterAddress_SOUTH;
  wire   [31:0] cacheDataOut_SOUTH;
  wire   [13:0] destinationAddressInBuffer_EAST;
  wire   [5:0] requesterAddressInBuffer_EAST;
  wire   [31:0] dataInBuffer_EAST;
  wire   [5:0] cacheRequesterAddress_EAST;
  wire   [31:0] cacheDataOut_EAST;
  wire   [13:0] destinationAddressInBuffer_WEST;
  wire   [5:0] requesterAddressInBuffer_WEST;
  wire   [31:0] dataInBuffer_WEST;
  wire   [5:0] cacheRequesterAddress_WEST;
  wire   [31:0] cacheDataOut_WEST;

  incomingPortHandler_0 inNorth ( .clk(clk), .reset(n364), 
        .localRouterAddress({n112, n125, n123, n118, n115, n85}), 
        .destinationAddressIn({destinationAddressIn_NORTH[13:12], n109, 
        destinationAddressIn_NORTH[10:9], n83, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .requesterAddressIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .readIn(n93), .writeIn(n101), .outputPortSelect(
        outputPortSelect_NORTH), .memRead(memRead_NORTH), .memWrite(
        memWrite_NORTH) );
  incomingPortHandler_3 inSouth ( .clk(clk), .reset(n366), 
        .localRouterAddress({n111, n126, n120, n117, n114, n85}), 
        .destinationAddressIn({destinationAddressIn_SOUTH[13:12], n107, 
        destinationAddressIn_SOUTH[10:9], n81, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .requesterAddressIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .readIn(n91), .writeIn(n99), .outputPortSelect(
        outputPortSelect_SOUTH), .memRead(memRead_SOUTH), .memWrite(
        memWrite_SOUTH) );
  incomingPortHandler_2 inEast ( .clk(clk), .reset(n364), .localRouterAddress(
        {n112, n127, n121, n118, n115, n85}), .destinationAddressIn({
        destinationAddressIn_EAST[13:12], n105, 
        destinationAddressIn_EAST[10:9], n79, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .requesterAddressIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .readIn(n89), .writeIn(n97), .outputPortSelect(
        outputPortSelect_EAST), .memRead(memRead_EAST), .memWrite(
        memWrite_EAST) );
  incomingPortHandler_1 inWest ( .clk(clk), .reset(n366), .localRouterAddress(
        {n111, n128, n122, n117, n114, n85}), .destinationAddressIn({
        destinationAddressIn_WEST[13:12], n103, 
        destinationAddressIn_WEST[10:9], n77, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .requesterAddressIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .readIn(n87), .writeIn(n95), .outputPortSelect(
        outputPortSelect_WEST), .memRead(memRead_WEST), .memWrite(
        memWrite_WEST) );
  cacheAccessArbiter cacheController ( .clk(clk), .reset(n75), 
        .cacheAddressIn_NORTH({n6, n7, n360, n359, n358, n357, n356, n355}), 
        .requesterAddressIn_NORTH({n354, n353, n352, n351, n350, n349}), 
        .memRead_NORTH(memRead_NORTH), .memWrite_NORTH(memWrite_NORTH), 
        .dataIn_NORTH({n348, n347, n346, n345, n344, n343, n342, n341, n340, 
        n339, n338, n337, n336, n335, n334, n333, n332, n331, n330, n329, n328, 
        n327, n326, n325, n324, n323, n322, n321, n320, n319, n318, n317}), 
        .readReady_NORTH(readReady_NORTH), .requesterAddressOut_NORTH(
        cacheRequesterAddress_NORTH), .cacheDataOut_NORTH(cacheDataOut_NORTH), 
        .cacheAddressIn_SOUTH({n304, n303, 
        destinationAddressInBuffer_SOUTH[5:0]}), .requesterAddressIn_SOUTH(
        requesterAddressInBuffer_SOUTH), .memRead_SOUTH(memRead_SOUTH), 
        .memWrite_SOUTH(memWrite_SOUTH), .dataIn_SOUTH(dataInBuffer_SOUTH), 
        .readReady_SOUTH(readReady_SOUTH), .requesterAddressOut_SOUTH(
        cacheRequesterAddress_SOUTH), .cacheDataOut_SOUTH(cacheDataOut_SOUTH), 
        .cacheAddressIn_EAST({n245, n243, n242, n241, n240, n239, n238, n237}), 
        .requesterAddressIn_EAST({n236, n235, n234, n233, n232, n231}), 
        .memRead_EAST(memRead_EAST), .memWrite_EAST(memWrite_EAST), 
        .dataIn_EAST(dataInBuffer_EAST), .readReady_EAST(readReady_EAST), 
        .requesterAddressOut_EAST(cacheRequesterAddress_EAST), 
        .cacheDataOut_EAST(cacheDataOut_EAST), .cacheAddressIn_WEST({n185, 
        n183, n182, n181, n180, n179, n178, n177}), .requesterAddressIn_WEST({
        n176, n175, n174, n173, n172, n171}), .memRead_WEST(memRead_WEST), 
        .memWrite_WEST(memWrite_WEST), .dataIn_WEST(dataInBuffer_WEST), 
        .readReady_WEST(readReady_WEST), .requesterAddressOut_WEST(
        cacheRequesterAddress_WEST), .cacheDataOut_WEST(cacheDataOut_WEST), 
        .cacheDataIn_A(cacheDataIn_A), .cacheAddressIn_A(cacheAddressIn_A), 
        .cacheDataOut_A(cacheDataOut_A), .memWrite_A(memWrite_A), 
        .cacheDataIn_B(cacheDataIn_B), .cacheAddressIn_B(cacheAddressIn_B), 
        .cacheDataOut_B(cacheDataOut_B), .memWrite_B(memWrite_B) );
  outputPortArbiter_0 outNorth ( .clk(clk), .reset(n365), .selectBit_NORTH(
        outputPortSelect_NORTH[0]), .destinationAddressIn_NORTH({
        destinationAddressInBuffer_NORTH[13:8], n2, n7, 
        destinationAddressInBuffer_NORTH[5], n359, 
        destinationAddressInBuffer_NORTH[3], n357, n356, n355}), 
        .requesterAddressIn_NORTH({requesterAddressInBuffer_NORTH[5], n353, 
        n352, requesterAddressInBuffer_NORTH[2], n350, n349}), .readIn_NORTH(
        readInBuffer_NORTH), .writeIn_NORTH(writeInBuffer_NORTH), 
        .dataIn_NORTH({n348, n347, dataInBuffer_NORTH[29], n345, n344, 
        dataInBuffer_NORTH[26], n342, n341, n340, n339, n338, 
        dataInBuffer_NORTH[20], n336, n335, n334, n333, n332, 
        dataInBuffer_NORTH[14], n330, n329, n328, n327, n326, n325, n324, n323, 
        dataInBuffer_NORTH[5], n321, dataInBuffer_NORTH[3], n319, n318, 
        dataInBuffer_NORTH[0]}), .selectBit_SOUTH(outputPortSelect_SOUTH[0]), 
        .destinationAddressIn_SOUTH({n315, n313, n311, n309, n307, n305, 
        destinationAddressInBuffer_SOUTH[7:6], n302, n301, n300, n299, n298, 
        n297}), .requesterAddressIn_SOUTH({n296, n295, n294, n293, n292, n291}), .readIn_SOUTH(n5), .writeIn_SOUTH(writeInBuffer_SOUTH), .dataIn_SOUTH({n290, 
        n289, n288, n287, n286, n285, n284, n283, n282, n281, n280, n279, n278, 
        n277, n276, n275, n274, n273, n272, n271, n270, n269, n268, n267, n266, 
        n265, n264, n263, n262, n261, n260, n259}), .selectBit_EAST(
        outputPortSelect_EAST[0]), .destinationAddressIn_EAST({n257, n255, 
        n253, n251, n249, n247, n245, n243, n242, n241, n240, n239, n238, n237}), .requesterAddressIn_EAST({requesterAddressInBuffer_EAST[5], n235, n234, 
        requesterAddressInBuffer_EAST[2:0]}), .readIn_EAST(readInBuffer_EAST), 
        .writeIn_EAST(writeInBuffer_EAST), .dataIn_EAST({n230, n229, n228, 
        n227, n226, n225, n224, n223, n222, n221, n220, n219, n218, n217, n216, 
        n215, n214, n213, n212, n211, n210, n209, n208, n207, n206, n205, n204, 
        n203, n202, n201, n200, n199}), .selectBit_WEST(
        outputPortSelect_WEST[0]), .destinationAddressIn_WEST({n197, n195, 
        n193, n191, n189, n187, n185, n183, n182, n181, n180, n179, n178, n177}), .requesterAddressIn_WEST({n176, n175, n174, n173, n172, n171}), 
        .readIn_WEST(readInBuffer_WEST), .writeIn_WEST(writeInBuffer_WEST), 
        .dataIn_WEST({n170, n169, n168, n167, n166, n165, n164, n163, n162, 
        n161, n160, n159, n158, n157, n156, n155, n154, n153, n152, n151, n150, 
        n149, n148, n147, n146, n145, n144, n143, n142, n141, n140, n139}), 
        .readReady(readReady_NORTH), .readRequesterAddress(
        cacheRequesterAddress_NORTH), .cacheDataOut(cacheDataOut_NORTH), 
        .destinationAddressOut(destinationAddressOut_NORTH), 
        .requesterAddressOut(requesterAddressOut_NORTH), .readOut(
        readOut_NORTH), .writeOut(writeOut_NORTH), .dataOut(dataOut_NORTH) );
  outputPortArbiter_3 outSouth ( .clk(clk), .reset(n361), .selectBit_NORTH(
        outputPortSelect_NORTH[1]), .destinationAddressIn_NORTH({
        destinationAddressInBuffer_NORTH[13:8], n6, n7, n360, 
        destinationAddressInBuffer_NORTH[4], n358, 
        destinationAddressInBuffer_NORTH[2:0]}), .requesterAddressIn_NORTH({
        n354, requesterAddressInBuffer_NORTH[4:3], n351, 
        requesterAddressInBuffer_NORTH[1:0]}), .readIn_NORTH(
        readInBuffer_NORTH), .writeIn_NORTH(writeInBuffer_NORTH), 
        .dataIn_NORTH({dataInBuffer_NORTH[31:30], n346, 
        dataInBuffer_NORTH[28:27], n343, dataInBuffer_NORTH[25:21], n337, 
        dataInBuffer_NORTH[19:15], n331, dataInBuffer_NORTH[13:6], n322, 
        dataInBuffer_NORTH[4], n320, dataInBuffer_NORTH[2:1], n317}), 
        .selectBit_SOUTH(outputPortSelect_SOUTH[1]), 
        .destinationAddressIn_SOUTH({n316, n314, n312, n310, n308, n306, 
        destinationAddressInBuffer_SOUTH[7:6], n302, n301, n300, n299, n298, 
        n297}), .requesterAddressIn_SOUTH({n296, n295, n294, n293, n292, n291}), .readIn_SOUTH(n136), .writeIn_SOUTH(writeInBuffer_SOUTH), .dataIn_SOUTH({
        n290, n289, n288, n287, n286, n285, n284, n283, n282, n281, n280, n279, 
        n278, n277, n276, n275, n274, n273, n272, n271, n270, n269, n268, n267, 
        n266, n265, n264, n263, n262, n261, n260, n259}), .selectBit_EAST(
        outputPortSelect_EAST[1]), .destinationAddressIn_EAST({n258, n256, 
        n254, n252, n250, n248, destinationAddressInBuffer_EAST[7:0]}), 
        .requesterAddressIn_EAST({n236, requesterAddressInBuffer_EAST[4:3], 
        n233, n232, n231}), .readIn_EAST(readInBuffer_EAST), .writeIn_EAST(
        writeInBuffer_EAST), .dataIn_EAST({n230, n229, n228, n227, n226, n225, 
        n224, n223, n222, n221, n220, n219, n218, n217, n216, n215, n214, n213, 
        n212, n211, n210, n209, n208, n207, n206, n205, n204, n203, n202, n201, 
        n200, n199}), .selectBit_WEST(outputPortSelect_WEST[1]), 
        .destinationAddressIn_WEST({n198, n196, n194, n192, n190, n188, 
        destinationAddressInBuffer_WEST[7:0]}), .requesterAddressIn_WEST(
        requesterAddressInBuffer_WEST), .readIn_WEST(readInBuffer_WEST), 
        .writeIn_WEST(writeInBuffer_WEST), .dataIn_WEST({n170, n169, n168, 
        n167, n166, n165, n164, n163, n162, n161, n160, n159, n158, n157, n156, 
        n155, n154, n153, n152, n151, n150, n149, n148, n147, n146, n145, n144, 
        n143, n142, n141, n140, n139}), .readReady(readReady_SOUTH), 
        .readRequesterAddress(cacheRequesterAddress_SOUTH), .cacheDataOut(
        cacheDataOut_SOUTH), .destinationAddressOut(
        destinationAddressOut_SOUTH), .requesterAddressOut(
        requesterAddressOut_SOUTH), .readOut(readOut_SOUTH), .writeOut(
        writeOut_SOUTH), .dataOut(dataOut_SOUTH) );
  outputPortArbiter_2 outEast ( .clk(clk), .reset(n362), .selectBit_NORTH(
        outputPortSelect_NORTH[2]), .destinationAddressIn_NORTH({
        destinationAddressInBuffer_NORTH[13:8], n2, n1, n360, 
        destinationAddressInBuffer_NORTH[4], n358, 
        destinationAddressInBuffer_NORTH[2:0]}), .requesterAddressIn_NORTH({
        n354, requesterAddressInBuffer_NORTH[4:3], n351, 
        requesterAddressInBuffer_NORTH[1:0]}), .readIn_NORTH(
        readInBuffer_NORTH), .writeIn_NORTH(writeInBuffer_NORTH), 
        .dataIn_NORTH({dataInBuffer_NORTH[31:30], n346, 
        dataInBuffer_NORTH[28:27], n343, dataInBuffer_NORTH[25:21], n337, 
        dataInBuffer_NORTH[19:15], n331, dataInBuffer_NORTH[13:6], n322, 
        dataInBuffer_NORTH[4], n320, dataInBuffer_NORTH[2:1], n317}), 
        .selectBit_SOUTH(outputPortSelect_SOUTH[2]), 
        .destinationAddressIn_SOUTH({n316, n314, n312, n310, n308, n306, n304, 
        n303, n302, n301, n300, n299, n298, n297}), .requesterAddressIn_SOUTH(
        {n296, n295, n294, n293, n292, n291}), .readIn_SOUTH(n137), 
        .writeIn_SOUTH(writeInBuffer_SOUTH), .dataIn_SOUTH({n290, n289, n288, 
        n287, n286, n285, n284, n283, n282, n281, n280, n279, n278, n277, n276, 
        n275, n274, n273, n272, n271, n270, n269, n268, n267, n266, n265, n264, 
        n263, n262, n261, n260, n259}), .selectBit_EAST(
        outputPortSelect_EAST[2]), .destinationAddressIn_EAST({n258, n256, 
        n254, n252, n250, n248, n246, n244, 
        destinationAddressInBuffer_EAST[5:0]}), .requesterAddressIn_EAST({n236, 
        requesterAddressInBuffer_EAST[4:3], n233, n232, n231}), .readIn_EAST(
        readInBuffer_EAST), .writeIn_EAST(writeInBuffer_EAST), .dataIn_EAST({
        n230, n229, n228, n227, n226, n225, n224, n223, n222, n221, n220, n219, 
        n218, n217, n216, n215, n214, n213, n212, n211, n210, n209, n208, n207, 
        n206, n205, n204, n203, n202, n201, n200, n199}), .selectBit_WEST(
        outputPortSelect_WEST[2]), .destinationAddressIn_WEST({n198, n196, 
        n194, n192, n190, n188, n186, n184, 
        destinationAddressInBuffer_WEST[5:0]}), .requesterAddressIn_WEST(
        requesterAddressInBuffer_WEST), .readIn_WEST(readInBuffer_WEST), 
        .writeIn_WEST(writeInBuffer_WEST), .dataIn_WEST({n170, n169, n168, 
        n167, n166, n165, n164, n163, n162, n161, n160, n159, n158, n157, n156, 
        n155, n154, n153, n152, n151, n150, n149, n148, n147, n146, n145, n144, 
        n143, n142, n141, n140, n139}), .readReady(readReady_EAST), 
        .readRequesterAddress(cacheRequesterAddress_EAST), .cacheDataOut(
        cacheDataOut_EAST), .destinationAddressOut(destinationAddressOut_EAST), 
        .requesterAddressOut(requesterAddressOut_EAST), .readOut(readOut_EAST), 
        .writeOut(writeOut_EAST), .dataOut(dataOut_EAST) );
  outputPortArbiter_1 outWest ( .clk(clk), .reset(n363), .selectBit_NORTH(
        outputPortSelect_NORTH[3]), .destinationAddressIn_NORTH({
        destinationAddressInBuffer_NORTH[13:8], n6, n1, n360, 
        destinationAddressInBuffer_NORTH[4], n358, 
        destinationAddressInBuffer_NORTH[2:0]}), .requesterAddressIn_NORTH({
        n354, requesterAddressInBuffer_NORTH[4:3], n351, 
        requesterAddressInBuffer_NORTH[1:0]}), .readIn_NORTH(
        readInBuffer_NORTH), .writeIn_NORTH(writeInBuffer_NORTH), 
        .dataIn_NORTH({dataInBuffer_NORTH[31:30], n346, 
        dataInBuffer_NORTH[28:27], n343, dataInBuffer_NORTH[25:21], n337, 
        dataInBuffer_NORTH[19:15], n331, dataInBuffer_NORTH[13:6], n322, 
        dataInBuffer_NORTH[4], n320, dataInBuffer_NORTH[2:1], n317}), 
        .selectBit_SOUTH(outputPortSelect_SOUTH[3]), 
        .destinationAddressIn_SOUTH({n315, n313, n311, n309, n307, n305, n304, 
        n303, n302, n301, n300, n299, n298, n297}), .requesterAddressIn_SOUTH(
        {n296, n295, n294, n293, n292, n291}), .readIn_SOUTH(n135), 
        .writeIn_SOUTH(writeInBuffer_SOUTH), .dataIn_SOUTH({n290, n289, n288, 
        n287, n286, n285, n284, n283, n282, n281, n280, n279, n278, n277, n276, 
        n275, n274, n273, n272, n271, n270, n269, n268, n267, n266, n265, n264, 
        n263, n262, n261, n260, n259}), .selectBit_EAST(
        outputPortSelect_EAST[3]), .destinationAddressIn_EAST({n257, n255, 
        n253, n251, n249, n247, n246, n244, 
        destinationAddressInBuffer_EAST[5:0]}), .requesterAddressIn_EAST({
        requesterAddressInBuffer_EAST[5], n235, n234, 
        requesterAddressInBuffer_EAST[2:0]}), .readIn_EAST(readInBuffer_EAST), 
        .writeIn_EAST(writeInBuffer_EAST), .dataIn_EAST({n230, n229, n228, 
        n227, n226, n225, n224, n223, n222, n221, n220, n219, n218, n217, n216, 
        n215, n214, n213, n212, n211, n210, n209, n208, n207, n206, n205, n204, 
        n203, n202, n201, n200, n199}), .selectBit_WEST(
        outputPortSelect_WEST[3]), .destinationAddressIn_WEST({n197, n195, 
        n193, n191, n189, n187, n186, n184, 
        destinationAddressInBuffer_WEST[5:0]}), .requesterAddressIn_WEST(
        requesterAddressInBuffer_WEST), .readIn_WEST(readInBuffer_WEST), 
        .writeIn_WEST(writeInBuffer_WEST), .dataIn_WEST({n170, n169, n168, 
        n167, n166, n165, n164, n163, n162, n161, n160, n159, n158, n157, n156, 
        n155, n154, n153, n152, n151, n150, n149, n148, n147, n146, n145, n144, 
        n143, n142, n141, n140, n139}), .readReady(readReady_WEST), 
        .readRequesterAddress(cacheRequesterAddress_WEST), .cacheDataOut(
        cacheDataOut_WEST), .destinationAddressOut(destinationAddressOut_WEST), 
        .requesterAddressOut(requesterAddressOut_WEST), .readOut(readOut_WEST), 
        .writeOut(writeOut_WEST), .dataOut(dataOut_WEST) );
  DFFTRX2TS \dataInBuffer_WEST_reg[9]  ( .D(dataIn_WEST[9]), .RN(n40), .CK(clk), .Q(dataInBuffer_WEST[9]) );
  DFFTRX2TS \requesterAddressInBuffer_NORTH_reg[3]  ( .D(
        requesterAddressIn_NORTH[3]), .RN(n62), .CK(clk), .Q(
        requesterAddressInBuffer_NORTH[3]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[22]  ( .D(dataIn_WEST[22]), .RN(n55), .CK(
        clk), .Q(dataInBuffer_WEST[22]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[21]  ( .D(dataIn_WEST[21]), .RN(n47), .CK(
        clk), .Q(dataInBuffer_WEST[21]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[20]  ( .D(dataIn_WEST[20]), .RN(n35), .CK(
        clk), .Q(dataInBuffer_WEST[20]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[19]  ( .D(dataIn_WEST[19]), .RN(n26), .CK(
        clk), .Q(dataInBuffer_WEST[19]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[18]  ( .D(dataIn_WEST[18]), .RN(n51), .CK(
        clk), .Q(dataInBuffer_WEST[18]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[17]  ( .D(dataIn_WEST[17]), .RN(n44), .CK(
        clk), .Q(dataInBuffer_WEST[17]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[16]  ( .D(dataIn_WEST[16]), .RN(n30), .CK(
        clk), .Q(dataInBuffer_WEST[16]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[15]  ( .D(dataIn_WEST[15]), .RN(n41), .CK(
        clk), .Q(dataInBuffer_WEST[15]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[14]  ( .D(dataIn_WEST[14]), .RN(n32), .CK(
        clk), .Q(dataInBuffer_WEST[14]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[13]  ( .D(dataIn_WEST[13]), .RN(n30), .CK(
        clk), .Q(dataInBuffer_WEST[13]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[12]  ( .D(dataIn_WEST[12]), .RN(n18), .CK(
        clk), .Q(dataInBuffer_WEST[12]) );
  DFFTRX2TS writeInBuffer_WEST_reg ( .D(n95), .RN(n29), .CK(clk), .Q(
        writeInBuffer_WEST) );
  DFFTRX2TS \requesterAddressInBuffer_WEST_reg[5]  ( .D(
        requesterAddressIn_WEST[5]), .RN(n28), .CK(clk), .Q(
        requesterAddressInBuffer_WEST[5]) );
  DFFTRX2TS \requesterAddressInBuffer_WEST_reg[4]  ( .D(
        requesterAddressIn_WEST[4]), .RN(n24), .CK(clk), .Q(
        requesterAddressInBuffer_WEST[4]) );
  DFFTRX2TS \requesterAddressInBuffer_WEST_reg[3]  ( .D(
        requesterAddressIn_WEST[3]), .RN(n39), .CK(clk), .Q(
        requesterAddressInBuffer_WEST[3]) );
  DFFTRX2TS \requesterAddressInBuffer_WEST_reg[2]  ( .D(
        requesterAddressIn_WEST[2]), .RN(n61), .CK(clk), .Q(
        requesterAddressInBuffer_WEST[2]) );
  DFFTRX2TS \requesterAddressInBuffer_WEST_reg[1]  ( .D(
        requesterAddressIn_WEST[1]), .RN(n54), .CK(clk), .Q(
        requesterAddressInBuffer_WEST[1]) );
  DFFTRX2TS \requesterAddressInBuffer_WEST_reg[0]  ( .D(
        requesterAddressIn_WEST[0]), .RN(n72), .CK(clk), .Q(
        requesterAddressInBuffer_WEST[0]) );
  DFFTRX2TS \requesterAddressInBuffer_NORTH_reg[0]  ( .D(
        requesterAddressIn_NORTH[0]), .RN(n34), .CK(clk), .Q(
        requesterAddressInBuffer_NORTH[0]) );
  DFFTRX2TS readInBuffer_WEST_reg ( .D(n87), .RN(n28), .CK(clk), .Q(
        readInBuffer_WEST) );
  DFFTRX2TS \destinationAddressInBuffer_WEST_reg[13]  ( .D(
        destinationAddressIn_WEST[13]), .RN(n50), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[13]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[1]  ( .D(dataIn_WEST[1]), .RN(n43), .CK(clk), .Q(dataInBuffer_WEST[1]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[0]  ( .D(dataIn_WEST[0]), .RN(n18), .CK(clk), .Q(dataInBuffer_WEST[0]) );
  DFFTRX2TS \requesterAddressInBuffer_NORTH_reg[2]  ( .D(
        requesterAddressIn_NORTH[2]), .RN(n29), .CK(clk), .Q(
        requesterAddressInBuffer_NORTH[2]) );
  DFFTRX2TS \destinationAddressInBuffer_NORTH_reg[6]  ( .D(
        destinationAddressIn_NORTH[6]), .RN(n26), .CK(clk), .Q(n1), .QN(n3) );
  DFFTRX2TS \dataInBuffer_WEST_reg[11]  ( .D(dataIn_WEST[11]), .RN(n24), .CK(
        clk), .Q(dataInBuffer_WEST[11]) );
  DFFTRX2TS writeInBuffer_SOUTH_reg ( .D(n99), .RN(n9), .CK(clk), .Q(
        writeInBuffer_SOUTH) );
  DFFTRX2TS writeInBuffer_NORTH_reg ( .D(n101), .RN(n13), .CK(clk), .Q(
        writeInBuffer_NORTH) );
  DFFTRX2TS writeInBuffer_EAST_reg ( .D(n97), .RN(n31), .CK(clk), .Q(
        writeInBuffer_EAST) );
  DFFTRX2TS \requesterAddressInBuffer_SOUTH_reg[5]  ( .D(
        requesterAddressIn_SOUTH[5]), .RN(n27), .CK(clk), .Q(
        requesterAddressInBuffer_SOUTH[5]) );
  DFFTRX2TS \requesterAddressInBuffer_SOUTH_reg[4]  ( .D(
        requesterAddressIn_SOUTH[4]), .RN(n42), .CK(clk), .Q(
        requesterAddressInBuffer_SOUTH[4]) );
  DFFTRX2TS \requesterAddressInBuffer_SOUTH_reg[3]  ( .D(
        requesterAddressIn_SOUTH[3]), .RN(n64), .CK(clk), .Q(
        requesterAddressInBuffer_SOUTH[3]) );
  DFFTRX2TS \requesterAddressInBuffer_SOUTH_reg[2]  ( .D(
        requesterAddressIn_SOUTH[2]), .RN(n57), .CK(clk), .Q(
        requesterAddressInBuffer_SOUTH[2]) );
  DFFTRX2TS \requesterAddressInBuffer_SOUTH_reg[1]  ( .D(
        requesterAddressIn_SOUTH[1]), .RN(n49), .CK(clk), .Q(
        requesterAddressInBuffer_SOUTH[1]) );
  DFFTRX2TS \requesterAddressInBuffer_SOUTH_reg[0]  ( .D(
        requesterAddressIn_SOUTH[0]), .RN(n37), .CK(clk), .Q(
        requesterAddressInBuffer_SOUTH[0]) );
  DFFTRX2TS \requesterAddressInBuffer_NORTH_reg[5]  ( .D(
        requesterAddressIn_NORTH[5]), .RN(n60), .CK(clk), .Q(
        requesterAddressInBuffer_NORTH[5]) );
  DFFTRX2TS \requesterAddressInBuffer_NORTH_reg[4]  ( .D(
        requesterAddressIn_NORTH[4]), .RN(n53), .CK(clk), .Q(
        requesterAddressInBuffer_NORTH[4]) );
  DFFTRX2TS \requesterAddressInBuffer_EAST_reg[5]  ( .D(
        requesterAddressIn_EAST[5]), .RN(n46), .CK(clk), .Q(
        requesterAddressInBuffer_EAST[5]) );
  DFFTRX2TS \requesterAddressInBuffer_EAST_reg[4]  ( .D(
        requesterAddressIn_EAST[4]), .RN(n18), .CK(clk), .Q(
        requesterAddressInBuffer_EAST[4]) );
  DFFTRX2TS \requesterAddressInBuffer_EAST_reg[3]  ( .D(
        requesterAddressIn_EAST[3]), .RN(n36), .CK(clk), .Q(
        requesterAddressInBuffer_EAST[3]) );
  DFFTRX2TS \requesterAddressInBuffer_EAST_reg[2]  ( .D(
        requesterAddressIn_EAST[2]), .RN(n10), .CK(clk), .Q(
        requesterAddressInBuffer_EAST[2]) );
  DFFTRX2TS \requesterAddressInBuffer_EAST_reg[1]  ( .D(
        requesterAddressIn_EAST[1]), .RN(n14), .CK(clk), .Q(
        requesterAddressInBuffer_EAST[1]) );
  DFFTRX2TS \requesterAddressInBuffer_EAST_reg[0]  ( .D(
        requesterAddressIn_EAST[0]), .RN(n9), .CK(clk), .Q(
        requesterAddressInBuffer_EAST[0]) );
  DFFTRX2TS readInBuffer_SOUTH_reg ( .D(n91), .RN(n46), .CK(clk), .Q(n5), .QN(
        n134) );
  DFFTRX2TS readInBuffer_NORTH_reg ( .D(n93), .RN(n11), .CK(clk), .Q(
        readInBuffer_NORTH) );
  DFFTRX2TS readInBuffer_EAST_reg ( .D(n89), .RN(n10), .CK(clk), .Q(
        readInBuffer_EAST) );
  DFFTRX2TS \destinationAddressInBuffer_WEST_reg[12]  ( .D(
        destinationAddressIn_WEST[12]), .RN(n41), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[12]) );
  DFFTRX2TS \destinationAddressInBuffer_WEST_reg[11]  ( .D(n103), .RN(n63), 
        .CK(clk), .Q(destinationAddressInBuffer_WEST[11]) );
  DFFTRX2TS \destinationAddressInBuffer_WEST_reg[10]  ( .D(
        destinationAddressIn_WEST[10]), .RN(n56), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[10]) );
  DFFTRX2TS \destinationAddressInBuffer_WEST_reg[9]  ( .D(
        destinationAddressIn_WEST[9]), .RN(n48), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[9]) );
  DFFTRX2TS \destinationAddressInBuffer_WEST_reg[8]  ( .D(n77), .RN(n36), .CK(
        clk), .Q(destinationAddressInBuffer_WEST[8]) );
  DFFTRX2TS \destinationAddressInBuffer_WEST_reg[7]  ( .D(
        destinationAddressIn_WEST[7]), .RN(n59), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[7]) );
  DFFTRX2TS \destinationAddressInBuffer_WEST_reg[6]  ( .D(
        destinationAddressIn_WEST[6]), .RN(n52), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[6]) );
  DFFTRX2TS \destinationAddressInBuffer_WEST_reg[5]  ( .D(
        destinationAddressIn_WEST[5]), .RN(n45), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[5]) );
  DFFTRX2TS \destinationAddressInBuffer_WEST_reg[4]  ( .D(
        destinationAddressIn_WEST[4]), .RN(n19), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[4]) );
  DFFTRX2TS \destinationAddressInBuffer_WEST_reg[3]  ( .D(
        destinationAddressIn_WEST[3]), .RN(n14), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[3]) );
  DFFTRX2TS \destinationAddressInBuffer_WEST_reg[2]  ( .D(
        destinationAddressIn_WEST[2]), .RN(n27), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[2]) );
  DFFTRX2TS \destinationAddressInBuffer_WEST_reg[1]  ( .D(
        destinationAddressIn_WEST[1]), .RN(n25), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[1]) );
  DFFTRX2TS \destinationAddressInBuffer_WEST_reg[0]  ( .D(
        destinationAddressIn_WEST[0]), .RN(n67), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[0]) );
  DFFTRX2TS \destinationAddressInBuffer_SOUTH_reg[13]  ( .D(
        destinationAddressIn_SOUTH[13]), .RN(n28), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[13]) );
  DFFTRX2TS \destinationAddressInBuffer_SOUTH_reg[12]  ( .D(
        destinationAddressIn_SOUTH[12]), .RN(n72), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[12]) );
  DFFTRX2TS \destinationAddressInBuffer_SOUTH_reg[11]  ( .D(n107), .RN(n70), 
        .CK(clk), .Q(destinationAddressInBuffer_SOUTH[11]) );
  DFFTRX2TS \destinationAddressInBuffer_SOUTH_reg[10]  ( .D(
        destinationAddressIn_SOUTH[10]), .RN(n40), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[10]) );
  DFFTRX2TS \destinationAddressInBuffer_SOUTH_reg[9]  ( .D(
        destinationAddressIn_SOUTH[9]), .RN(n62), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[9]) );
  DFFTRX2TS \destinationAddressInBuffer_SOUTH_reg[8]  ( .D(n81), .RN(n55), 
        .CK(clk), .Q(destinationAddressInBuffer_SOUTH[8]) );
  DFFTRX2TS \destinationAddressInBuffer_SOUTH_reg[7]  ( .D(
        destinationAddressIn_SOUTH[7]), .RN(n47), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[7]) );
  DFFTRX2TS \destinationAddressInBuffer_SOUTH_reg[6]  ( .D(
        destinationAddressIn_SOUTH[6]), .RN(n35), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[6]) );
  DFFTRX2TS \destinationAddressInBuffer_SOUTH_reg[5]  ( .D(
        destinationAddressIn_SOUTH[5]), .RN(n133), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[5]) );
  DFFTRX2TS \destinationAddressInBuffer_SOUTH_reg[4]  ( .D(
        destinationAddressIn_SOUTH[4]), .RN(n51), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[4]) );
  DFFTRX2TS \destinationAddressInBuffer_SOUTH_reg[3]  ( .D(
        destinationAddressIn_SOUTH[3]), .RN(n44), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[3]) );
  DFFTRX2TS \destinationAddressInBuffer_SOUTH_reg[2]  ( .D(
        destinationAddressIn_SOUTH[2]), .RN(n66), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[2]) );
  DFFTRX2TS \destinationAddressInBuffer_SOUTH_reg[1]  ( .D(
        destinationAddressIn_SOUTH[1]), .RN(n13), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[1]) );
  DFFTRX2TS \destinationAddressInBuffer_SOUTH_reg[0]  ( .D(
        destinationAddressIn_SOUTH[0]), .RN(n71), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[0]) );
  DFFTRX2TS \destinationAddressInBuffer_NORTH_reg[13]  ( .D(
        destinationAddressIn_NORTH[13]), .RN(n69), .CK(clk), .Q(
        destinationAddressInBuffer_NORTH[13]) );
  DFFTRX2TS \destinationAddressInBuffer_NORTH_reg[12]  ( .D(
        destinationAddressIn_NORTH[12]), .RN(n67), .CK(clk), .Q(
        destinationAddressInBuffer_NORTH[12]) );
  DFFTRX2TS \destinationAddressInBuffer_NORTH_reg[11]  ( .D(n109), .RN(n132), 
        .CK(clk), .Q(destinationAddressInBuffer_NORTH[11]) );
  DFFTRX2TS \destinationAddressInBuffer_NORTH_reg[10]  ( .D(
        destinationAddressIn_NORTH[10]), .RN(n72), .CK(clk), .Q(
        destinationAddressInBuffer_NORTH[10]) );
  DFFTRX2TS \destinationAddressInBuffer_NORTH_reg[9]  ( .D(
        destinationAddressIn_NORTH[9]), .RN(n70), .CK(clk), .Q(
        destinationAddressInBuffer_NORTH[9]) );
  DFFTRX2TS \destinationAddressInBuffer_NORTH_reg[8]  ( .D(n83), .RN(n39), 
        .CK(clk), .Q(destinationAddressInBuffer_NORTH[8]) );
  DFFTRX2TS \destinationAddressInBuffer_NORTH_reg[7]  ( .D(
        destinationAddressIn_NORTH[7]), .RN(n61), .CK(clk), .Q(n2), .QN(n4) );
  DFFTRX2TS \destinationAddressInBuffer_NORTH_reg[5]  ( .D(
        destinationAddressIn_NORTH[5]), .RN(n54), .CK(clk), .Q(
        destinationAddressInBuffer_NORTH[5]) );
  DFFTRX2TS \destinationAddressInBuffer_NORTH_reg[4]  ( .D(
        destinationAddressIn_NORTH[4]), .RN(n31), .CK(clk), .Q(
        destinationAddressInBuffer_NORTH[4]) );
  DFFTRX2TS \destinationAddressInBuffer_NORTH_reg[3]  ( .D(
        destinationAddressIn_NORTH[3]), .RN(n34), .CK(clk), .Q(
        destinationAddressInBuffer_NORTH[3]) );
  DFFTRX2TS \destinationAddressInBuffer_NORTH_reg[2]  ( .D(
        destinationAddressIn_NORTH[2]), .RN(n28), .CK(clk), .Q(
        destinationAddressInBuffer_NORTH[2]) );
  DFFTRX2TS \destinationAddressInBuffer_NORTH_reg[1]  ( .D(
        destinationAddressIn_NORTH[1]), .RN(n50), .CK(clk), .Q(
        destinationAddressInBuffer_NORTH[1]) );
  DFFTRX2TS \destinationAddressInBuffer_NORTH_reg[0]  ( .D(
        destinationAddressIn_NORTH[0]), .RN(n43), .CK(clk), .Q(
        destinationAddressInBuffer_NORTH[0]) );
  DFFTRX2TS \destinationAddressInBuffer_EAST_reg[13]  ( .D(
        destinationAddressIn_EAST[13]), .RN(n131), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[13]) );
  DFFTRX2TS \destinationAddressInBuffer_EAST_reg[12]  ( .D(
        destinationAddressIn_EAST[12]), .RN(n60), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[12]) );
  DFFTRX2TS \destinationAddressInBuffer_EAST_reg[11]  ( .D(n105), .RN(n63), 
        .CK(clk), .Q(destinationAddressInBuffer_EAST[11]) );
  DFFTRX2TS \destinationAddressInBuffer_EAST_reg[10]  ( .D(
        destinationAddressIn_EAST[10]), .RN(n138), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[10]) );
  DFFTRX2TS \destinationAddressInBuffer_EAST_reg[9]  ( .D(
        destinationAddressIn_EAST[9]), .RN(n20), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[9]) );
  DFFTRX2TS \destinationAddressInBuffer_EAST_reg[8]  ( .D(n79), .RN(n74), .CK(
        clk), .Q(destinationAddressInBuffer_EAST[8]) );
  DFFTRX2TS \destinationAddressInBuffer_EAST_reg[7]  ( .D(
        destinationAddressIn_EAST[7]), .RN(n11), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[7]) );
  DFFTRX2TS \destinationAddressInBuffer_EAST_reg[6]  ( .D(
        destinationAddressIn_EAST[6]), .RN(n29), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[6]) );
  DFFTRX2TS \destinationAddressInBuffer_EAST_reg[5]  ( .D(
        destinationAddressIn_EAST[5]), .RN(n42), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[5]) );
  DFFTRX2TS \destinationAddressInBuffer_EAST_reg[4]  ( .D(
        destinationAddressIn_EAST[4]), .RN(n64), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[4]) );
  DFFTRX2TS \destinationAddressInBuffer_EAST_reg[3]  ( .D(
        destinationAddressIn_EAST[3]), .RN(n57), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[3]) );
  DFFTRX2TS \destinationAddressInBuffer_EAST_reg[2]  ( .D(
        destinationAddressIn_EAST[2]), .RN(n49), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[2]) );
  DFFTRX2TS \destinationAddressInBuffer_EAST_reg[1]  ( .D(
        destinationAddressIn_EAST[1]), .RN(n37), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[1]) );
  DFFTRX2TS \destinationAddressInBuffer_EAST_reg[0]  ( .D(
        destinationAddressIn_EAST[0]), .RN(n60), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[0]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[31]  ( .D(dataIn_WEST[31]), .RN(n53), .CK(
        clk), .Q(dataInBuffer_WEST[31]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[30]  ( .D(dataIn_WEST[30]), .RN(n46), .CK(
        clk), .Q(dataInBuffer_WEST[30]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[29]  ( .D(dataIn_WEST[29]), .RN(n66), .CK(
        clk), .Q(dataInBuffer_WEST[29]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[28]  ( .D(dataIn_WEST[28]), .RN(n73), .CK(
        clk), .Q(dataInBuffer_WEST[28]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[27]  ( .D(dataIn_WEST[27]), .RN(n71), .CK(
        clk), .Q(dataInBuffer_WEST[27]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[26]  ( .D(dataIn_WEST[26]), .RN(n69), .CK(
        clk), .Q(dataInBuffer_WEST[26]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[25]  ( .D(dataIn_WEST[25]), .RN(n19), .CK(
        clk), .Q(dataInBuffer_WEST[25]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[24]  ( .D(dataIn_WEST[24]), .RN(n20), .CK(
        clk), .Q(dataInBuffer_WEST[24]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[23]  ( .D(dataIn_WEST[23]), .RN(n27), .CK(
        clk), .Q(dataInBuffer_WEST[23]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[10]  ( .D(dataIn_WEST[10]), .RN(n25), .CK(
        clk), .Q(dataInBuffer_WEST[10]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[31]  ( .D(dataIn_SOUTH[31]), .RN(n41), 
        .CK(clk), .Q(dataInBuffer_SOUTH[31]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[30]  ( .D(dataIn_SOUTH[30]), .RN(n63), 
        .CK(clk), .Q(dataInBuffer_SOUTH[30]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[29]  ( .D(dataIn_SOUTH[29]), .RN(n56), 
        .CK(clk), .Q(dataInBuffer_SOUTH[29]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[28]  ( .D(dataIn_SOUTH[28]), .RN(n48), 
        .CK(clk), .Q(dataInBuffer_SOUTH[28]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[27]  ( .D(dataIn_SOUTH[27]), .RN(n36), 
        .CK(clk), .Q(dataInBuffer_SOUTH[27]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[26]  ( .D(dataIn_SOUTH[26]), .RN(n59), 
        .CK(clk), .Q(dataInBuffer_SOUTH[26]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[25]  ( .D(dataIn_SOUTH[25]), .RN(n52), 
        .CK(clk), .Q(dataInBuffer_SOUTH[25]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[24]  ( .D(dataIn_SOUTH[24]), .RN(n45), 
        .CK(clk), .Q(dataInBuffer_SOUTH[24]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[23]  ( .D(dataIn_SOUTH[23]), .RN(n9), .CK(
        clk), .Q(dataInBuffer_SOUTH[23]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[22]  ( .D(dataIn_SOUTH[22]), .RN(n73), 
        .CK(clk), .Q(dataInBuffer_SOUTH[22]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[21]  ( .D(dataIn_SOUTH[21]), .RN(n11), 
        .CK(clk), .Q(dataInBuffer_SOUTH[21]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[20]  ( .D(dataIn_SOUTH[20]), .RN(n10), 
        .CK(clk), .Q(dataInBuffer_SOUTH[20]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[19]  ( .D(dataIn_SOUTH[19]), .RN(n32), 
        .CK(clk), .Q(dataInBuffer_SOUTH[19]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[18]  ( .D(dataIn_SOUTH[18]), .RN(n132), 
        .CK(clk), .Q(dataInBuffer_SOUTH[18]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[17]  ( .D(dataIn_SOUTH[17]), .RN(n30), 
        .CK(clk), .Q(dataInBuffer_SOUTH[17]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[16]  ( .D(dataIn_SOUTH[16]), .RN(n57), 
        .CK(clk), .Q(dataInBuffer_SOUTH[16]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[15]  ( .D(dataIn_SOUTH[15]), .RN(n40), 
        .CK(clk), .Q(dataInBuffer_SOUTH[15]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[14]  ( .D(dataIn_SOUTH[14]), .RN(n62), 
        .CK(clk), .Q(dataInBuffer_SOUTH[14]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[13]  ( .D(dataIn_SOUTH[13]), .RN(n55), 
        .CK(clk), .Q(dataInBuffer_SOUTH[13]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[12]  ( .D(dataIn_SOUTH[12]), .RN(n47), 
        .CK(clk), .Q(dataInBuffer_SOUTH[12]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[11]  ( .D(dataIn_SOUTH[11]), .RN(n35), 
        .CK(clk), .Q(dataInBuffer_SOUTH[11]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[10]  ( .D(dataIn_SOUTH[10]), .RN(n133), 
        .CK(clk), .Q(dataInBuffer_SOUTH[10]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[9]  ( .D(dataIn_SOUTH[9]), .RN(n51), .CK(
        clk), .Q(dataInBuffer_SOUTH[9]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[8]  ( .D(dataIn_SOUTH[8]), .RN(n44), .CK(
        clk), .Q(dataInBuffer_SOUTH[8]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[7]  ( .D(dataIn_SOUTH[7]), .RN(n13), .CK(
        clk), .Q(dataInBuffer_SOUTH[7]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[6]  ( .D(dataIn_SOUTH[6]), .RN(n45), .CK(
        clk), .Q(dataInBuffer_SOUTH[6]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[5]  ( .D(dataIn_SOUTH[5]), .RN(n74), .CK(
        clk), .Q(dataInBuffer_SOUTH[5]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[4]  ( .D(dataIn_SOUTH[4]), .RN(n19), .CK(
        clk), .Q(dataInBuffer_SOUTH[4]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[3]  ( .D(dataIn_SOUTH[3]), .RN(n37), .CK(
        clk), .Q(dataInBuffer_SOUTH[3]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[2]  ( .D(dataIn_SOUTH[2]), .RN(n74), .CK(
        clk), .Q(dataInBuffer_SOUTH[2]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[1]  ( .D(dataIn_SOUTH[1]), .RN(n64), .CK(
        clk), .Q(dataInBuffer_SOUTH[1]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[0]  ( .D(dataIn_SOUTH[0]), .RN(n130), .CK(
        clk), .Q(dataInBuffer_SOUTH[0]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[31]  ( .D(dataIn_NORTH[31]), .RN(n39), 
        .CK(clk), .Q(dataInBuffer_NORTH[31]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[30]  ( .D(dataIn_NORTH[30]), .RN(n61), 
        .CK(clk), .Q(dataInBuffer_NORTH[30]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[29]  ( .D(dataIn_NORTH[29]), .RN(n54), 
        .CK(clk), .Q(dataInBuffer_NORTH[29]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[28]  ( .D(dataIn_NORTH[28]), .RN(n11), 
        .CK(clk), .Q(dataInBuffer_NORTH[28]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[27]  ( .D(dataIn_NORTH[27]), .RN(n34), 
        .CK(clk), .Q(dataInBuffer_NORTH[27]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[26]  ( .D(dataIn_NORTH[26]), .RN(n26), 
        .CK(clk), .Q(dataInBuffer_NORTH[26]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[25]  ( .D(dataIn_NORTH[25]), .RN(n50), 
        .CK(clk), .Q(dataInBuffer_NORTH[25]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[24]  ( .D(dataIn_NORTH[24]), .RN(n43), 
        .CK(clk), .Q(dataInBuffer_NORTH[24]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[23]  ( .D(dataIn_NORTH[23]), .RN(n49), 
        .CK(clk), .Q(dataInBuffer_NORTH[23]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[22]  ( .D(dataIn_NORTH[22]), .RN(n53), 
        .CK(clk), .Q(dataInBuffer_NORTH[22]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[21]  ( .D(dataIn_NORTH[21]), .RN(n31), 
        .CK(clk), .Q(dataInBuffer_NORTH[21]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[20]  ( .D(dataIn_NORTH[20]), .RN(n73), 
        .CK(clk), .Q(dataInBuffer_NORTH[20]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[19]  ( .D(dataIn_NORTH[19]), .RN(n25), 
        .CK(clk), .Q(dataInBuffer_NORTH[19]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[18]  ( .D(dataIn_NORTH[18]), .RN(n138), 
        .CK(clk), .Q(dataInBuffer_NORTH[18]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[17]  ( .D(dataIn_NORTH[17]), .RN(n27), 
        .CK(clk), .Q(dataInBuffer_NORTH[17]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[16]  ( .D(dataIn_NORTH[16]), .RN(n25), 
        .CK(clk), .Q(dataInBuffer_NORTH[16]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[15]  ( .D(dataIn_NORTH[15]), .RN(n42), 
        .CK(clk), .Q(dataInBuffer_NORTH[15]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[14]  ( .D(dataIn_NORTH[14]), .RN(n64), 
        .CK(clk), .Q(dataInBuffer_NORTH[14]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[13]  ( .D(dataIn_NORTH[13]), .RN(n57), 
        .CK(clk), .Q(dataInBuffer_NORTH[13]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[12]  ( .D(dataIn_NORTH[12]), .RN(n49), 
        .CK(clk), .Q(dataInBuffer_NORTH[12]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[11]  ( .D(dataIn_NORTH[11]), .RN(n37), 
        .CK(clk), .Q(dataInBuffer_NORTH[11]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[10]  ( .D(dataIn_NORTH[10]), .RN(n60), 
        .CK(clk), .Q(dataInBuffer_NORTH[10]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[9]  ( .D(dataIn_NORTH[9]), .RN(n53), .CK(
        clk), .Q(dataInBuffer_NORTH[9]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[8]  ( .D(dataIn_NORTH[8]), .RN(n46), .CK(
        clk), .Q(dataInBuffer_NORTH[8]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[7]  ( .D(dataIn_NORTH[7]), .RN(n67), .CK(
        clk), .Q(dataInBuffer_NORTH[7]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[6]  ( .D(dataIn_NORTH[6]), .RN(n138), .CK(
        clk), .Q(dataInBuffer_NORTH[6]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[5]  ( .D(dataIn_NORTH[5]), .RN(n72), .CK(
        clk), .Q(dataInBuffer_NORTH[5]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[4]  ( .D(dataIn_NORTH[4]), .RN(n70), .CK(
        clk), .Q(dataInBuffer_NORTH[4]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[3]  ( .D(dataIn_NORTH[3]), .RN(n19), .CK(
        clk), .Q(dataInBuffer_NORTH[3]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[2]  ( .D(dataIn_NORTH[2]), .RN(n130), .CK(
        clk), .Q(dataInBuffer_NORTH[2]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[1]  ( .D(dataIn_NORTH[1]), .RN(n132), .CK(
        clk), .Q(dataInBuffer_NORTH[1]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[0]  ( .D(dataIn_NORTH[0]), .RN(n24), .CK(
        clk), .Q(dataInBuffer_NORTH[0]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[31]  ( .D(dataIn_EAST[31]), .RN(n41), .CK(
        clk), .Q(dataInBuffer_EAST[31]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[30]  ( .D(dataIn_EAST[30]), .RN(n63), .CK(
        clk), .Q(dataInBuffer_EAST[30]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[29]  ( .D(dataIn_EAST[29]), .RN(n56), .CK(
        clk), .Q(dataInBuffer_EAST[29]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[28]  ( .D(dataIn_EAST[28]), .RN(n48), .CK(
        clk), .Q(dataInBuffer_EAST[28]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[27]  ( .D(dataIn_EAST[27]), .RN(n36), .CK(
        clk), .Q(dataInBuffer_EAST[27]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[26]  ( .D(dataIn_EAST[26]), .RN(n59), .CK(
        clk), .Q(dataInBuffer_EAST[26]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[25]  ( .D(dataIn_EAST[25]), .RN(n52), .CK(
        clk), .Q(dataInBuffer_EAST[25]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[24]  ( .D(dataIn_EAST[24]), .RN(n45), .CK(
        clk), .Q(dataInBuffer_EAST[24]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[23]  ( .D(dataIn_EAST[23]), .RN(n42), .CK(
        clk), .Q(dataInBuffer_EAST[23]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[22]  ( .D(dataIn_EAST[22]), .RN(n59), .CK(
        clk), .Q(dataInBuffer_EAST[22]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[21]  ( .D(dataIn_EAST[21]), .RN(n32), .CK(
        clk), .Q(dataInBuffer_EAST[21]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[20]  ( .D(dataIn_EAST[20]), .RN(n56), .CK(
        clk), .Q(dataInBuffer_EAST[20]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[19]  ( .D(dataIn_EAST[19]), .RN(n48), .CK(
        clk), .Q(dataInBuffer_EAST[19]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[18]  ( .D(dataIn_EAST[18]), .RN(n52), .CK(
        clk), .Q(dataInBuffer_EAST[18]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[17]  ( .D(dataIn_EAST[17]), .RN(n132), .CK(
        clk), .Q(dataInBuffer_EAST[17]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[16]  ( .D(dataIn_EAST[16]), .RN(n31), .CK(
        clk), .Q(dataInBuffer_EAST[16]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[15]  ( .D(dataIn_EAST[15]), .RN(n40), .CK(
        clk), .Q(dataInBuffer_EAST[15]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[14]  ( .D(dataIn_EAST[14]), .RN(n62), .CK(
        clk), .Q(dataInBuffer_EAST[14]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[13]  ( .D(dataIn_EAST[13]), .RN(n55), .CK(
        clk), .Q(dataInBuffer_EAST[13]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[12]  ( .D(dataIn_EAST[12]), .RN(n47), .CK(
        clk), .Q(dataInBuffer_EAST[12]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[11]  ( .D(dataIn_EAST[11]), .RN(n35), .CK(
        clk), .Q(dataInBuffer_EAST[11]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[10]  ( .D(dataIn_EAST[10]), .RN(n133), .CK(
        clk), .Q(dataInBuffer_EAST[10]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[9]  ( .D(dataIn_EAST[9]), .RN(n51), .CK(clk), .Q(dataInBuffer_EAST[9]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[8]  ( .D(dataIn_EAST[8]), .RN(n44), .CK(clk), .Q(dataInBuffer_EAST[8]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[7]  ( .D(dataIn_EAST[7]), .RN(n66), .CK(clk), .Q(dataInBuffer_EAST[7]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[6]  ( .D(dataIn_EAST[6]), .RN(n73), .CK(clk), .Q(dataInBuffer_EAST[6]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[5]  ( .D(dataIn_EAST[5]), .RN(n71), .CK(clk), .Q(dataInBuffer_EAST[5]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[4]  ( .D(dataIn_EAST[4]), .RN(n69), .CK(clk), .Q(dataInBuffer_EAST[4]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[3]  ( .D(dataIn_EAST[3]), .RN(n18), .CK(clk), .Q(dataInBuffer_EAST[3]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[2]  ( .D(dataIn_EAST[2]), .RN(n29), .CK(clk), .Q(dataInBuffer_EAST[2]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[1]  ( .D(dataIn_EAST[1]), .RN(n26), .CK(clk), .Q(dataInBuffer_EAST[1]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[0]  ( .D(dataIn_EAST[0]), .RN(n24), .CK(clk), .Q(dataInBuffer_EAST[0]) );
  DFFTRX2TS \requesterAddressInBuffer_NORTH_reg[1]  ( .D(
        requesterAddressIn_NORTH[1]), .RN(n39), .CK(clk), .Q(
        requesterAddressInBuffer_NORTH[1]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[8]  ( .D(dataIn_WEST[8]), .RN(n61), .CK(clk), .Q(dataInBuffer_WEST[8]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[7]  ( .D(dataIn_WEST[7]), .RN(n54), .CK(clk), .Q(dataInBuffer_WEST[7]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[6]  ( .D(dataIn_WEST[6]), .RN(n71), .CK(clk), .Q(dataInBuffer_WEST[6]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[5]  ( .D(dataIn_WEST[5]), .RN(n34), .CK(clk), .Q(dataInBuffer_WEST[5]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[4]  ( .D(dataIn_WEST[4]), .RN(n131), .CK(
        clk), .Q(dataInBuffer_WEST[4]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[3]  ( .D(dataIn_WEST[3]), .RN(n50), .CK(clk), .Q(dataInBuffer_WEST[3]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[2]  ( .D(dataIn_WEST[2]), .RN(n43), .CK(clk), .Q(dataInBuffer_WEST[2]) );
  INVXLTS U219 ( .A(n4), .Y(n6) );
  INVXLTS U220 ( .A(n3), .Y(n7) );
  INVXLTS U221 ( .A(n30), .Y(n8) );
  INVXLTS U222 ( .A(n8), .Y(n9) );
  INVXLTS U223 ( .A(n23), .Y(n10) );
  INVXLTS U224 ( .A(n17), .Y(n11) );
  INVXLTS U225 ( .A(n32), .Y(n12) );
  INVXLTS U226 ( .A(n12), .Y(n13) );
  INVXLTS U227 ( .A(n65), .Y(n14) );
  INVXLTS U228 ( .A(n14), .Y(n15) );
  INVXLTS U229 ( .A(n14), .Y(n16) );
  INVXLTS U230 ( .A(n67), .Y(n17) );
  INVXLTS U231 ( .A(n17), .Y(n18) );
  INVXLTS U232 ( .A(n17), .Y(n19) );
  INVXLTS U233 ( .A(n68), .Y(n20) );
  INVXLTS U234 ( .A(n20), .Y(n21) );
  INVXLTS U235 ( .A(n20), .Y(n22) );
  INVXLTS U236 ( .A(n70), .Y(n23) );
  INVXLTS U237 ( .A(n23), .Y(n24) );
  INVXLTS U238 ( .A(n23), .Y(n25) );
  INVXLTS U239 ( .A(n8), .Y(n26) );
  INVXLTS U240 ( .A(n15), .Y(n27) );
  INVXLTS U241 ( .A(n68), .Y(n28) );
  INVXLTS U242 ( .A(n16), .Y(n29) );
  CLKBUFX2TS U243 ( .A(n130), .Y(n30) );
  CLKBUFX2TS U244 ( .A(n131), .Y(n31) );
  CLKBUFX2TS U245 ( .A(n133), .Y(n32) );
  INVXLTS U246 ( .A(n66), .Y(n33) );
  INVXLTS U247 ( .A(n33), .Y(n34) );
  INVXLTS U248 ( .A(n33), .Y(n35) );
  INVXLTS U249 ( .A(n33), .Y(n36) );
  INVXLTS U250 ( .A(n33), .Y(n37) );
  INVXLTS U251 ( .A(n9), .Y(n38) );
  INVXLTS U252 ( .A(n38), .Y(n39) );
  INVXLTS U253 ( .A(n38), .Y(n40) );
  INVXLTS U254 ( .A(n38), .Y(n41) );
  INVXLTS U255 ( .A(n38), .Y(n42) );
  INVXLTS U256 ( .A(n65), .Y(n43) );
  INVXLTS U257 ( .A(n68), .Y(n44) );
  INVXLTS U258 ( .A(n65), .Y(n45) );
  INVXLTS U259 ( .A(n15), .Y(n46) );
  INVXLTS U260 ( .A(n21), .Y(n47) );
  INVXLTS U261 ( .A(n21), .Y(n48) );
  INVXLTS U262 ( .A(n22), .Y(n49) );
  INVXLTS U263 ( .A(n16), .Y(n50) );
  INVXLTS U264 ( .A(n23), .Y(n51) );
  INVXLTS U265 ( .A(n22), .Y(n52) );
  INVXLTS U266 ( .A(n16), .Y(n53) );
  INVXLTS U267 ( .A(n8), .Y(n54) );
  INVXLTS U268 ( .A(n8), .Y(n55) );
  INVXLTS U269 ( .A(n58), .Y(n56) );
  INVXLTS U270 ( .A(n15), .Y(n57) );
  INVXLTS U271 ( .A(n13), .Y(n58) );
  INVXLTS U272 ( .A(n58), .Y(n59) );
  INVXLTS U273 ( .A(n58), .Y(n60) );
  INVXLTS U274 ( .A(n12), .Y(n61) );
  INVXLTS U275 ( .A(n58), .Y(n62) );
  INVXLTS U276 ( .A(n12), .Y(n63) );
  INVXLTS U277 ( .A(n12), .Y(n64) );
  INVXLTS U278 ( .A(n130), .Y(n65) );
  INVXLTS U279 ( .A(n15), .Y(n66) );
  INVXLTS U280 ( .A(n16), .Y(n67) );
  INVXLTS U281 ( .A(n131), .Y(n68) );
  INVXLTS U282 ( .A(n21), .Y(n69) );
  INVXLTS U283 ( .A(n22), .Y(n70) );
  INVXLTS U284 ( .A(n22), .Y(n71) );
  INVXLTS U285 ( .A(n21), .Y(n72) );
  INVXLTS U286 ( .A(n17), .Y(n73) );
  INVXLTS U287 ( .A(reset), .Y(n74) );
  INVXLTS U288 ( .A(n74), .Y(n75) );
  INVXLTS U289 ( .A(destinationAddressIn_WEST[8]), .Y(n76) );
  INVXLTS U290 ( .A(n76), .Y(n77) );
  INVXLTS U291 ( .A(destinationAddressIn_EAST[8]), .Y(n78) );
  INVXLTS U292 ( .A(n78), .Y(n79) );
  INVXLTS U293 ( .A(destinationAddressIn_SOUTH[8]), .Y(n80) );
  INVXLTS U294 ( .A(n80), .Y(n81) );
  INVXLTS U295 ( .A(destinationAddressIn_NORTH[8]), .Y(n82) );
  INVXLTS U296 ( .A(n82), .Y(n83) );
  INVXLTS U297 ( .A(localRouterAddress[0]), .Y(n84) );
  INVXLTS U298 ( .A(n84), .Y(n85) );
  INVXLTS U299 ( .A(readIn_WEST), .Y(n86) );
  INVXLTS U300 ( .A(n86), .Y(n87) );
  INVXLTS U301 ( .A(readIn_EAST), .Y(n88) );
  INVXLTS U302 ( .A(n88), .Y(n89) );
  INVXLTS U303 ( .A(readIn_SOUTH), .Y(n90) );
  INVXLTS U304 ( .A(n90), .Y(n91) );
  INVXLTS U305 ( .A(readIn_NORTH), .Y(n92) );
  INVXLTS U306 ( .A(n92), .Y(n93) );
  INVXLTS U307 ( .A(writeIn_WEST), .Y(n94) );
  INVXLTS U308 ( .A(n94), .Y(n95) );
  INVXLTS U309 ( .A(writeIn_EAST), .Y(n96) );
  INVXLTS U310 ( .A(n96), .Y(n97) );
  INVXLTS U311 ( .A(writeIn_SOUTH), .Y(n98) );
  INVXLTS U312 ( .A(n98), .Y(n99) );
  INVXLTS U313 ( .A(writeIn_NORTH), .Y(n100) );
  INVXLTS U314 ( .A(n100), .Y(n101) );
  INVXLTS U315 ( .A(destinationAddressIn_WEST[11]), .Y(n102) );
  INVXLTS U316 ( .A(n102), .Y(n103) );
  INVXLTS U317 ( .A(destinationAddressIn_EAST[11]), .Y(n104) );
  INVXLTS U318 ( .A(n104), .Y(n105) );
  INVXLTS U319 ( .A(destinationAddressIn_SOUTH[11]), .Y(n106) );
  INVXLTS U320 ( .A(n106), .Y(n107) );
  INVXLTS U321 ( .A(destinationAddressIn_NORTH[11]), .Y(n108) );
  INVXLTS U322 ( .A(n108), .Y(n109) );
  INVXLTS U323 ( .A(localRouterAddress[5]), .Y(n110) );
  INVXLTS U324 ( .A(n110), .Y(n111) );
  INVXLTS U325 ( .A(n110), .Y(n112) );
  INVXLTS U326 ( .A(localRouterAddress[1]), .Y(n113) );
  INVXLTS U327 ( .A(n113), .Y(n114) );
  INVXLTS U328 ( .A(n113), .Y(n115) );
  INVXLTS U329 ( .A(localRouterAddress[2]), .Y(n116) );
  INVXLTS U330 ( .A(n116), .Y(n117) );
  INVXLTS U331 ( .A(n116), .Y(n118) );
  INVXLTS U332 ( .A(localRouterAddress[3]), .Y(n119) );
  INVXLTS U333 ( .A(n119), .Y(n120) );
  INVXLTS U334 ( .A(n119), .Y(n121) );
  INVXLTS U335 ( .A(n119), .Y(n122) );
  INVXLTS U336 ( .A(n119), .Y(n123) );
  INVXLTS U337 ( .A(localRouterAddress[4]), .Y(n124) );
  INVXLTS U338 ( .A(n124), .Y(n125) );
  INVXLTS U339 ( .A(n124), .Y(n126) );
  INVXLTS U340 ( .A(n124), .Y(n127) );
  INVXLTS U341 ( .A(n124), .Y(n128) );
  INVXLTS U342 ( .A(n138), .Y(n129) );
  CLKINVX2TS U343 ( .A(n129), .Y(n130) );
  CLKINVX2TS U344 ( .A(n129), .Y(n131) );
  CLKINVX2TS U345 ( .A(n129), .Y(n132) );
  INVX2TS U346 ( .A(n129), .Y(n133) );
  INVX2TS U347 ( .A(n134), .Y(n135) );
  INVX2TS U348 ( .A(n134), .Y(n136) );
  INVX2TS U349 ( .A(n134), .Y(n137) );
  CLKBUFX2TS U350 ( .A(destinationAddressInBuffer_SOUTH[0]), .Y(n297) );
  CLKBUFX2TS U351 ( .A(requesterAddressInBuffer_SOUTH[5]), .Y(n296) );
  CLKBUFX2TS U352 ( .A(requesterAddressInBuffer_SOUTH[4]), .Y(n295) );
  CLKBUFX2TS U353 ( .A(requesterAddressInBuffer_SOUTH[2]), .Y(n293) );
  CLKBUFX2TS U354 ( .A(destinationAddressInBuffer_SOUTH[5]), .Y(n302) );
  CLKBUFX2TS U355 ( .A(destinationAddressInBuffer_SOUTH[3]), .Y(n300) );
  CLKBUFX2TS U356 ( .A(destinationAddressInBuffer_SOUTH[2]), .Y(n299) );
  CLKBUFX2TS U357 ( .A(destinationAddressInBuffer_SOUTH[1]), .Y(n298) );
  CLKBUFX2TS U358 ( .A(dataInBuffer_WEST[31]), .Y(n170) );
  CLKBUFX2TS U359 ( .A(dataInBuffer_SOUTH[30]), .Y(n289) );
  CLKBUFX2TS U360 ( .A(dataInBuffer_WEST[30]), .Y(n169) );
  CLKBUFX2TS U361 ( .A(dataInBuffer_SOUTH[29]), .Y(n288) );
  CLKBUFX2TS U362 ( .A(dataInBuffer_WEST[29]), .Y(n168) );
  CLKBUFX2TS U363 ( .A(dataInBuffer_SOUTH[26]), .Y(n285) );
  CLKBUFX2TS U364 ( .A(dataInBuffer_WEST[26]), .Y(n165) );
  CLKBUFX2TS U365 ( .A(dataInBuffer_WEST[24]), .Y(n163) );
  CLKBUFX2TS U366 ( .A(dataInBuffer_WEST[22]), .Y(n161) );
  CLKBUFX2TS U367 ( .A(dataInBuffer_SOUTH[21]), .Y(n280) );
  CLKBUFX2TS U368 ( .A(dataInBuffer_WEST[21]), .Y(n160) );
  CLKBUFX2TS U369 ( .A(dataInBuffer_SOUTH[19]), .Y(n278) );
  CLKBUFX2TS U370 ( .A(dataInBuffer_WEST[19]), .Y(n158) );
  CLKBUFX2TS U371 ( .A(dataInBuffer_WEST[16]), .Y(n155) );
  CLKBUFX2TS U372 ( .A(dataInBuffer_SOUTH[13]), .Y(n272) );
  CLKBUFX2TS U373 ( .A(dataInBuffer_WEST[13]), .Y(n152) );
  CLKBUFX2TS U374 ( .A(dataInBuffer_SOUTH[12]), .Y(n271) );
  CLKBUFX2TS U375 ( .A(dataInBuffer_WEST[12]), .Y(n151) );
  CLKBUFX2TS U376 ( .A(dataInBuffer_SOUTH[11]), .Y(n270) );
  CLKBUFX2TS U377 ( .A(dataInBuffer_WEST[11]), .Y(n150) );
  CLKBUFX2TS U378 ( .A(dataInBuffer_SOUTH[10]), .Y(n269) );
  CLKBUFX2TS U379 ( .A(dataInBuffer_WEST[10]), .Y(n149) );
  CLKBUFX2TS U380 ( .A(dataInBuffer_SOUTH[8]), .Y(n267) );
  CLKBUFX2TS U381 ( .A(dataInBuffer_WEST[8]), .Y(n147) );
  CLKBUFX2TS U382 ( .A(dataInBuffer_WEST[6]), .Y(n145) );
  CLKBUFX2TS U383 ( .A(requesterAddressInBuffer_SOUTH[3]), .Y(n294) );
  CLKBUFX2TS U384 ( .A(requesterAddressInBuffer_SOUTH[1]), .Y(n292) );
  CLKBUFX2TS U385 ( .A(requesterAddressInBuffer_SOUTH[0]), .Y(n291) );
  CLKBUFX2TS U386 ( .A(dataInBuffer_WEST[28]), .Y(n167) );
  CLKBUFX2TS U387 ( .A(dataInBuffer_SOUTH[28]), .Y(n287) );
  CLKBUFX2TS U388 ( .A(dataInBuffer_WEST[27]), .Y(n166) );
  CLKBUFX2TS U389 ( .A(dataInBuffer_SOUTH[27]), .Y(n286) );
  CLKBUFX2TS U390 ( .A(dataInBuffer_WEST[23]), .Y(n162) );
  CLKBUFX2TS U391 ( .A(dataInBuffer_SOUTH[23]), .Y(n282) );
  CLKBUFX2TS U392 ( .A(dataInBuffer_WEST[20]), .Y(n159) );
  CLKBUFX2TS U393 ( .A(dataInBuffer_SOUTH[20]), .Y(n279) );
  CLKBUFX2TS U394 ( .A(dataInBuffer_WEST[9]), .Y(n148) );
  CLKBUFX2TS U395 ( .A(dataInBuffer_SOUTH[9]), .Y(n268) );
  CLKBUFX2TS U396 ( .A(dataInBuffer_WEST[5]), .Y(n144) );
  CLKBUFX2TS U397 ( .A(dataInBuffer_SOUTH[5]), .Y(n264) );
  CLKBUFX2TS U398 ( .A(dataInBuffer_WEST[2]), .Y(n141) );
  CLKBUFX2TS U399 ( .A(dataInBuffer_WEST[1]), .Y(n140) );
  CLKBUFX2TS U400 ( .A(dataInBuffer_SOUTH[1]), .Y(n260) );
  CLKBUFX2TS U401 ( .A(dataInBuffer_WEST[0]), .Y(n139) );
  CLKBUFX2TS U402 ( .A(dataInBuffer_SOUTH[31]), .Y(n290) );
  CLKBUFX2TS U403 ( .A(dataInBuffer_SOUTH[24]), .Y(n283) );
  CLKBUFX2TS U404 ( .A(dataInBuffer_SOUTH[22]), .Y(n281) );
  CLKBUFX2TS U405 ( .A(dataInBuffer_SOUTH[16]), .Y(n275) );
  CLKBUFX2TS U406 ( .A(dataInBuffer_SOUTH[6]), .Y(n265) );
  CLKBUFX2TS U407 ( .A(dataInBuffer_SOUTH[2]), .Y(n261) );
  CLKBUFX2TS U408 ( .A(dataInBuffer_SOUTH[0]), .Y(n259) );
  CLKBUFX2TS U409 ( .A(dataInBuffer_WEST[7]), .Y(n146) );
  CLKBUFX2TS U410 ( .A(dataInBuffer_SOUTH[7]), .Y(n266) );
  CLKBUFX2TS U411 ( .A(dataInBuffer_WEST[17]), .Y(n156) );
  CLKBUFX2TS U412 ( .A(dataInBuffer_SOUTH[17]), .Y(n276) );
  CLKBUFX2TS U413 ( .A(dataInBuffer_WEST[15]), .Y(n154) );
  CLKBUFX2TS U414 ( .A(dataInBuffer_SOUTH[15]), .Y(n274) );
  CLKBUFX2TS U415 ( .A(dataInBuffer_WEST[14]), .Y(n153) );
  CLKBUFX2TS U416 ( .A(dataInBuffer_SOUTH[14]), .Y(n273) );
  CLKBUFX2TS U417 ( .A(dataInBuffer_WEST[3]), .Y(n142) );
  CLKBUFX2TS U418 ( .A(dataInBuffer_SOUTH[3]), .Y(n262) );
  CLKBUFX2TS U419 ( .A(destinationAddressInBuffer_SOUTH[4]), .Y(n301) );
  CLKBUFX2TS U420 ( .A(dataInBuffer_WEST[25]), .Y(n164) );
  CLKBUFX2TS U421 ( .A(dataInBuffer_SOUTH[25]), .Y(n284) );
  CLKBUFX2TS U422 ( .A(dataInBuffer_WEST[18]), .Y(n157) );
  CLKBUFX2TS U423 ( .A(dataInBuffer_SOUTH[18]), .Y(n277) );
  CLKBUFX2TS U424 ( .A(dataInBuffer_WEST[4]), .Y(n143) );
  CLKBUFX2TS U425 ( .A(dataInBuffer_SOUTH[4]), .Y(n263) );
  CLKBUFX2TS U426 ( .A(dataInBuffer_EAST[31]), .Y(n230) );
  CLKBUFX2TS U427 ( .A(dataInBuffer_EAST[30]), .Y(n229) );
  CLKBUFX2TS U428 ( .A(dataInBuffer_EAST[29]), .Y(n228) );
  CLKBUFX2TS U429 ( .A(dataInBuffer_EAST[26]), .Y(n225) );
  CLKBUFX2TS U430 ( .A(dataInBuffer_EAST[24]), .Y(n223) );
  CLKBUFX2TS U431 ( .A(dataInBuffer_EAST[22]), .Y(n221) );
  CLKBUFX2TS U432 ( .A(dataInBuffer_EAST[21]), .Y(n220) );
  CLKBUFX2TS U433 ( .A(dataInBuffer_EAST[19]), .Y(n218) );
  CLKBUFX2TS U434 ( .A(dataInBuffer_EAST[17]), .Y(n216) );
  CLKBUFX2TS U435 ( .A(dataInBuffer_EAST[16]), .Y(n215) );
  CLKBUFX2TS U436 ( .A(dataInBuffer_EAST[14]), .Y(n213) );
  CLKBUFX2TS U437 ( .A(dataInBuffer_EAST[12]), .Y(n211) );
  CLKBUFX2TS U438 ( .A(dataInBuffer_EAST[11]), .Y(n210) );
  CLKBUFX2TS U439 ( .A(dataInBuffer_EAST[10]), .Y(n209) );
  CLKBUFX2TS U440 ( .A(dataInBuffer_EAST[8]), .Y(n207) );
  CLKBUFX2TS U441 ( .A(dataInBuffer_EAST[6]), .Y(n205) );
  CLKBUFX2TS U442 ( .A(dataInBuffer_EAST[3]), .Y(n202) );
  CLKBUFX2TS U443 ( .A(dataInBuffer_EAST[25]), .Y(n224) );
  CLKBUFX2TS U444 ( .A(dataInBuffer_EAST[18]), .Y(n217) );
  CLKBUFX2TS U445 ( .A(dataInBuffer_EAST[15]), .Y(n214) );
  CLKBUFX2TS U446 ( .A(dataInBuffer_EAST[13]), .Y(n212) );
  CLKBUFX2TS U447 ( .A(dataInBuffer_EAST[4]), .Y(n203) );
  CLKBUFX2TS U448 ( .A(dataInBuffer_EAST[28]), .Y(n227) );
  CLKBUFX2TS U449 ( .A(dataInBuffer_EAST[27]), .Y(n226) );
  CLKBUFX2TS U450 ( .A(dataInBuffer_EAST[23]), .Y(n222) );
  CLKBUFX2TS U451 ( .A(dataInBuffer_EAST[20]), .Y(n219) );
  CLKBUFX2TS U452 ( .A(dataInBuffer_EAST[9]), .Y(n208) );
  CLKBUFX2TS U453 ( .A(dataInBuffer_EAST[5]), .Y(n204) );
  CLKBUFX2TS U454 ( .A(dataInBuffer_EAST[2]), .Y(n201) );
  CLKBUFX2TS U455 ( .A(dataInBuffer_EAST[1]), .Y(n200) );
  CLKBUFX2TS U456 ( .A(dataInBuffer_EAST[0]), .Y(n199) );
  CLKBUFX2TS U457 ( .A(dataInBuffer_EAST[7]), .Y(n206) );
  CLKBUFX2TS U458 ( .A(requesterAddressInBuffer_EAST[3]), .Y(n234) );
  CLKBUFX2TS U459 ( .A(requesterAddressInBuffer_EAST[4]), .Y(n235) );
  CLKBUFX2TS U460 ( .A(n68), .Y(n361) );
  CLKBUFX2TS U461 ( .A(n65), .Y(n362) );
  CLKBUFX2TS U462 ( .A(n366), .Y(n363) );
  CLKBUFX2TS U463 ( .A(n366), .Y(n364) );
  CLKBUFX2TS U464 ( .A(n364), .Y(n365) );
  CLKBUFX2TS U465 ( .A(n75), .Y(n366) );
  CLKBUFX2TS U466 ( .A(requesterAddressInBuffer_EAST[5]), .Y(n236) );
  CLKBUFX2TS U467 ( .A(requesterAddressInBuffer_EAST[2]), .Y(n233) );
  CLKBUFX2TS U468 ( .A(requesterAddressInBuffer_EAST[1]), .Y(n232) );
  CLKBUFX2TS U469 ( .A(requesterAddressInBuffer_EAST[0]), .Y(n231) );
  CLKBUFX2TS U470 ( .A(destinationAddressInBuffer_WEST[0]), .Y(n177) );
  CLKBUFX2TS U471 ( .A(destinationAddressInBuffer_EAST[0]), .Y(n237) );
  CLKBUFX2TS U472 ( .A(destinationAddressInBuffer_WEST[1]), .Y(n178) );
  CLKBUFX2TS U473 ( .A(destinationAddressInBuffer_EAST[1]), .Y(n238) );
  CLKBUFX2TS U474 ( .A(destinationAddressInBuffer_WEST[2]), .Y(n179) );
  CLKBUFX2TS U475 ( .A(destinationAddressInBuffer_EAST[2]), .Y(n239) );
  CLKBUFX2TS U476 ( .A(destinationAddressInBuffer_WEST[3]), .Y(n180) );
  CLKBUFX2TS U477 ( .A(destinationAddressInBuffer_EAST[3]), .Y(n240) );
  CLKBUFX2TS U478 ( .A(destinationAddressInBuffer_WEST[4]), .Y(n181) );
  CLKBUFX2TS U479 ( .A(destinationAddressInBuffer_EAST[4]), .Y(n241) );
  CLKBUFX2TS U480 ( .A(destinationAddressInBuffer_WEST[5]), .Y(n182) );
  CLKBUFX2TS U481 ( .A(destinationAddressInBuffer_EAST[5]), .Y(n242) );
  CLKBUFX2TS U482 ( .A(requesterAddressInBuffer_WEST[0]), .Y(n171) );
  CLKBUFX2TS U483 ( .A(requesterAddressInBuffer_WEST[1]), .Y(n172) );
  CLKBUFX2TS U484 ( .A(requesterAddressInBuffer_WEST[2]), .Y(n173) );
  CLKBUFX2TS U485 ( .A(requesterAddressInBuffer_WEST[3]), .Y(n174) );
  CLKBUFX2TS U486 ( .A(requesterAddressInBuffer_WEST[4]), .Y(n175) );
  CLKBUFX2TS U487 ( .A(requesterAddressInBuffer_WEST[5]), .Y(n176) );
  CLKBUFX2TS U488 ( .A(destinationAddressInBuffer_SOUTH[6]), .Y(n303) );
  CLKBUFX2TS U489 ( .A(destinationAddressInBuffer_SOUTH[7]), .Y(n304) );
  CLKBUFX2TS U490 ( .A(destinationAddressInBuffer_WEST[6]), .Y(n184) );
  CLKBUFX2TS U491 ( .A(destinationAddressInBuffer_EAST[6]), .Y(n244) );
  CLKBUFX2TS U492 ( .A(destinationAddressInBuffer_WEST[7]), .Y(n186) );
  CLKBUFX2TS U493 ( .A(destinationAddressInBuffer_EAST[7]), .Y(n246) );
  CLKBUFX2TS U494 ( .A(destinationAddressInBuffer_WEST[6]), .Y(n183) );
  CLKBUFX2TS U495 ( .A(destinationAddressInBuffer_EAST[6]), .Y(n243) );
  CLKBUFX2TS U496 ( .A(destinationAddressInBuffer_WEST[7]), .Y(n185) );
  CLKBUFX2TS U497 ( .A(destinationAddressInBuffer_EAST[7]), .Y(n245) );
  CLKBUFX2TS U498 ( .A(destinationAddressInBuffer_WEST[12]), .Y(n196) );
  CLKBUFX2TS U499 ( .A(destinationAddressInBuffer_SOUTH[12]), .Y(n314) );
  CLKBUFX2TS U500 ( .A(destinationAddressInBuffer_EAST[12]), .Y(n256) );
  CLKBUFX2TS U501 ( .A(destinationAddressInBuffer_EAST[10]), .Y(n252) );
  CLKBUFX2TS U502 ( .A(destinationAddressInBuffer_SOUTH[10]), .Y(n310) );
  CLKBUFX2TS U503 ( .A(destinationAddressInBuffer_WEST[10]), .Y(n192) );
  CLKBUFX2TS U504 ( .A(destinationAddressInBuffer_EAST[9]), .Y(n250) );
  CLKBUFX2TS U505 ( .A(destinationAddressInBuffer_WEST[9]), .Y(n190) );
  CLKBUFX2TS U506 ( .A(destinationAddressInBuffer_SOUTH[9]), .Y(n308) );
  CLKBUFX2TS U507 ( .A(destinationAddressInBuffer_WEST[13]), .Y(n198) );
  CLKBUFX2TS U508 ( .A(destinationAddressInBuffer_EAST[13]), .Y(n258) );
  CLKBUFX2TS U509 ( .A(destinationAddressInBuffer_SOUTH[13]), .Y(n316) );
  CLKBUFX2TS U510 ( .A(destinationAddressInBuffer_WEST[11]), .Y(n194) );
  CLKBUFX2TS U511 ( .A(destinationAddressInBuffer_EAST[11]), .Y(n254) );
  CLKBUFX2TS U512 ( .A(destinationAddressInBuffer_SOUTH[11]), .Y(n312) );
  CLKBUFX2TS U513 ( .A(destinationAddressInBuffer_WEST[8]), .Y(n188) );
  CLKBUFX2TS U514 ( .A(destinationAddressInBuffer_EAST[8]), .Y(n248) );
  CLKBUFX2TS U515 ( .A(destinationAddressInBuffer_SOUTH[8]), .Y(n306) );
  CLKBUFX2TS U516 ( .A(destinationAddressInBuffer_WEST[12]), .Y(n195) );
  CLKBUFX2TS U517 ( .A(destinationAddressInBuffer_SOUTH[12]), .Y(n313) );
  CLKBUFX2TS U518 ( .A(destinationAddressInBuffer_EAST[12]), .Y(n255) );
  CLKBUFX2TS U519 ( .A(destinationAddressInBuffer_EAST[10]), .Y(n251) );
  CLKBUFX2TS U520 ( .A(destinationAddressInBuffer_SOUTH[10]), .Y(n309) );
  CLKBUFX2TS U521 ( .A(destinationAddressInBuffer_WEST[10]), .Y(n191) );
  CLKBUFX2TS U522 ( .A(destinationAddressInBuffer_EAST[9]), .Y(n249) );
  CLKBUFX2TS U523 ( .A(destinationAddressInBuffer_WEST[9]), .Y(n189) );
  CLKBUFX2TS U524 ( .A(destinationAddressInBuffer_SOUTH[9]), .Y(n307) );
  CLKBUFX2TS U525 ( .A(destinationAddressInBuffer_WEST[13]), .Y(n197) );
  CLKBUFX2TS U526 ( .A(destinationAddressInBuffer_EAST[13]), .Y(n257) );
  CLKBUFX2TS U527 ( .A(destinationAddressInBuffer_SOUTH[13]), .Y(n315) );
  CLKBUFX2TS U528 ( .A(destinationAddressInBuffer_WEST[11]), .Y(n193) );
  CLKBUFX2TS U529 ( .A(destinationAddressInBuffer_EAST[11]), .Y(n253) );
  CLKBUFX2TS U530 ( .A(destinationAddressInBuffer_SOUTH[11]), .Y(n311) );
  CLKBUFX2TS U531 ( .A(destinationAddressInBuffer_WEST[8]), .Y(n187) );
  CLKBUFX2TS U532 ( .A(destinationAddressInBuffer_EAST[8]), .Y(n247) );
  CLKBUFX2TS U533 ( .A(destinationAddressInBuffer_SOUTH[8]), .Y(n305) );
  CLKBUFX2TS U534 ( .A(destinationAddressInBuffer_NORTH[0]), .Y(n355) );
  CLKBUFX2TS U535 ( .A(requesterAddressInBuffer_NORTH[4]), .Y(n353) );
  CLKBUFX2TS U536 ( .A(destinationAddressInBuffer_NORTH[2]), .Y(n357) );
  CLKBUFX2TS U537 ( .A(destinationAddressInBuffer_NORTH[1]), .Y(n356) );
  CLKBUFX2TS U538 ( .A(dataInBuffer_NORTH[30]), .Y(n347) );
  CLKBUFX2TS U539 ( .A(dataInBuffer_NORTH[21]), .Y(n338) );
  CLKBUFX2TS U540 ( .A(dataInBuffer_NORTH[19]), .Y(n336) );
  CLKBUFX2TS U541 ( .A(dataInBuffer_NORTH[13]), .Y(n330) );
  CLKBUFX2TS U542 ( .A(dataInBuffer_NORTH[12]), .Y(n329) );
  CLKBUFX2TS U543 ( .A(dataInBuffer_NORTH[11]), .Y(n328) );
  CLKBUFX2TS U544 ( .A(dataInBuffer_NORTH[10]), .Y(n327) );
  CLKBUFX2TS U545 ( .A(dataInBuffer_NORTH[8]), .Y(n325) );
  CLKBUFX2TS U546 ( .A(requesterAddressInBuffer_NORTH[3]), .Y(n352) );
  CLKBUFX2TS U547 ( .A(requesterAddressInBuffer_NORTH[1]), .Y(n350) );
  CLKBUFX2TS U548 ( .A(requesterAddressInBuffer_NORTH[0]), .Y(n349) );
  CLKBUFX2TS U549 ( .A(dataInBuffer_NORTH[28]), .Y(n345) );
  CLKBUFX2TS U550 ( .A(dataInBuffer_NORTH[27]), .Y(n344) );
  CLKBUFX2TS U551 ( .A(dataInBuffer_NORTH[23]), .Y(n340) );
  CLKBUFX2TS U552 ( .A(dataInBuffer_NORTH[9]), .Y(n326) );
  CLKBUFX2TS U553 ( .A(dataInBuffer_NORTH[1]), .Y(n318) );
  CLKBUFX2TS U554 ( .A(dataInBuffer_NORTH[31]), .Y(n348) );
  CLKBUFX2TS U555 ( .A(dataInBuffer_NORTH[24]), .Y(n341) );
  CLKBUFX2TS U556 ( .A(dataInBuffer_NORTH[22]), .Y(n339) );
  CLKBUFX2TS U557 ( .A(dataInBuffer_NORTH[16]), .Y(n333) );
  CLKBUFX2TS U558 ( .A(dataInBuffer_NORTH[6]), .Y(n323) );
  CLKBUFX2TS U559 ( .A(dataInBuffer_NORTH[2]), .Y(n319) );
  CLKBUFX2TS U560 ( .A(dataInBuffer_NORTH[7]), .Y(n324) );
  CLKBUFX2TS U561 ( .A(dataInBuffer_NORTH[17]), .Y(n334) );
  CLKBUFX2TS U562 ( .A(dataInBuffer_NORTH[15]), .Y(n332) );
  CLKBUFX2TS U563 ( .A(destinationAddressInBuffer_NORTH[4]), .Y(n359) );
  CLKBUFX2TS U564 ( .A(dataInBuffer_NORTH[25]), .Y(n342) );
  CLKBUFX2TS U565 ( .A(dataInBuffer_NORTH[18]), .Y(n335) );
  CLKBUFX2TS U566 ( .A(dataInBuffer_NORTH[4]), .Y(n321) );
  CLKBUFX2TS U567 ( .A(requesterAddressInBuffer_NORTH[5]), .Y(n354) );
  CLKBUFX2TS U568 ( .A(requesterAddressInBuffer_NORTH[2]), .Y(n351) );
  CLKBUFX2TS U569 ( .A(destinationAddressInBuffer_NORTH[5]), .Y(n360) );
  CLKBUFX2TS U570 ( .A(destinationAddressInBuffer_NORTH[3]), .Y(n358) );
  CLKBUFX2TS U571 ( .A(dataInBuffer_NORTH[29]), .Y(n346) );
  CLKBUFX2TS U572 ( .A(dataInBuffer_NORTH[26]), .Y(n343) );
  CLKBUFX2TS U573 ( .A(dataInBuffer_NORTH[20]), .Y(n337) );
  CLKBUFX2TS U574 ( .A(dataInBuffer_NORTH[5]), .Y(n322) );
  CLKBUFX2TS U575 ( .A(dataInBuffer_NORTH[0]), .Y(n317) );
  CLKBUFX2TS U576 ( .A(dataInBuffer_NORTH[14]), .Y(n331) );
  CLKBUFX2TS U577 ( .A(dataInBuffer_NORTH[3]), .Y(n320) );
  INVX2TS U578 ( .A(n364), .Y(n138) );
endmodule

