
module cacheAccessArbiter ( clk, reset, cacheAddressIn_NORTH, 
        requesterAddressIn_NORTH, memRead_NORTH, memWrite_NORTH, dataIn_NORTH, 
        readReady_NORTH, requesterAddressOut_NORTH, cacheDataOut_NORTH, 
        cacheAddressIn_SOUTH, requesterAddressIn_SOUTH, memRead_SOUTH, 
        memWrite_SOUTH, dataIn_SOUTH, readReady_SOUTH, 
        requesterAddressOut_SOUTH, cacheDataOut_SOUTH, cacheAddressIn_EAST, 
        requesterAddressIn_EAST, memRead_EAST, memWrite_EAST, dataIn_EAST, 
        readReady_EAST, requesterAddressOut_EAST, cacheDataOut_EAST, 
        cacheAddressIn_WEST, requesterAddressIn_WEST, memRead_WEST, 
        memWrite_WEST, dataIn_WEST, readReady_WEST, requesterAddressOut_WEST, 
        cacheDataOut_WEST, cacheDataIn_A, cacheAddressIn_A, cacheDataOut_A, 
        memWrite_A, cacheDataIn_B, cacheAddressIn_B, cacheDataOut_B, 
        memWrite_B );
  input [7:0] cacheAddressIn_NORTH;
  input [3:0] requesterAddressIn_NORTH;
  input [5:0] dataIn_NORTH;
  output [3:0] requesterAddressOut_NORTH;
  output [5:0] cacheDataOut_NORTH;
  input [7:0] cacheAddressIn_SOUTH;
  input [3:0] requesterAddressIn_SOUTH;
  input [5:0] dataIn_SOUTH;
  output [3:0] requesterAddressOut_SOUTH;
  output [5:0] cacheDataOut_SOUTH;
  input [7:0] cacheAddressIn_EAST;
  input [3:0] requesterAddressIn_EAST;
  input [5:0] dataIn_EAST;
  output [3:0] requesterAddressOut_EAST;
  output [5:0] cacheDataOut_EAST;
  input [7:0] cacheAddressIn_WEST;
  input [3:0] requesterAddressIn_WEST;
  input [5:0] dataIn_WEST;
  output [3:0] requesterAddressOut_WEST;
  output [5:0] cacheDataOut_WEST;
  output [5:0] cacheDataIn_A;
  output [7:0] cacheAddressIn_A;
  input [5:0] cacheDataOut_A;
  output [5:0] cacheDataIn_B;
  output [7:0] cacheAddressIn_B;
  input [5:0] cacheDataOut_B;
  input clk, reset, memRead_NORTH, memWrite_NORTH, memRead_SOUTH,
         memWrite_SOUTH, memRead_EAST, memWrite_EAST, memRead_WEST,
         memWrite_WEST;
  output readReady_NORTH, readReady_SOUTH, readReady_EAST, readReady_WEST,
         memWrite_A, memWrite_B;
  wire   N741, N742, \dataToWriteBuffer[6][5] , \dataToWriteBuffer[6][4] ,
         \dataToWriteBuffer[6][3] , \dataToWriteBuffer[6][2] ,
         \dataToWriteBuffer[6][1] , \dataToWriteBuffer[6][0] ,
         \dataToWriteBuffer[5][5] , \dataToWriteBuffer[5][4] ,
         \dataToWriteBuffer[5][3] , \dataToWriteBuffer[5][2] ,
         \dataToWriteBuffer[5][1] , \dataToWriteBuffer[5][0] ,
         \dataToWriteBuffer[4][5] , \dataToWriteBuffer[4][4] ,
         \dataToWriteBuffer[4][3] , \dataToWriteBuffer[4][2] ,
         \dataToWriteBuffer[4][1] , \dataToWriteBuffer[4][0] ,
         \dataToWriteBuffer[3][5] , \dataToWriteBuffer[3][4] ,
         \dataToWriteBuffer[3][3] , \dataToWriteBuffer[3][2] ,
         \dataToWriteBuffer[3][1] , \dataToWriteBuffer[3][0] ,
         \dataToWriteBuffer[2][5] , \dataToWriteBuffer[2][4] ,
         \dataToWriteBuffer[2][3] , \dataToWriteBuffer[2][2] ,
         \dataToWriteBuffer[2][1] , \dataToWriteBuffer[2][0] ,
         \dataToWriteBuffer[1][5] , \dataToWriteBuffer[1][4] ,
         \dataToWriteBuffer[1][3] , \dataToWriteBuffer[1][2] ,
         \dataToWriteBuffer[1][1] , \dataToWriteBuffer[1][0] ,
         \dataToWriteBuffer[0][5] , \dataToWriteBuffer[0][4] ,
         \dataToWriteBuffer[0][3] , \dataToWriteBuffer[0][2] ,
         \dataToWriteBuffer[0][1] , \dataToWriteBuffer[0][0] ,
         \addressToWriteBuffer[6][7] , \addressToWriteBuffer[6][6] ,
         \addressToWriteBuffer[6][5] , \addressToWriteBuffer[6][4] ,
         \addressToWriteBuffer[6][3] , \addressToWriteBuffer[6][2] ,
         \addressToWriteBuffer[6][1] , \addressToWriteBuffer[6][0] ,
         \addressToWriteBuffer[5][7] , \addressToWriteBuffer[5][6] ,
         \addressToWriteBuffer[5][5] , \addressToWriteBuffer[5][4] ,
         \addressToWriteBuffer[5][3] , \addressToWriteBuffer[5][2] ,
         \addressToWriteBuffer[5][1] , \addressToWriteBuffer[5][0] ,
         \addressToWriteBuffer[4][7] , \addressToWriteBuffer[4][6] ,
         \addressToWriteBuffer[4][5] , \addressToWriteBuffer[4][4] ,
         \addressToWriteBuffer[4][3] , \addressToWriteBuffer[4][2] ,
         \addressToWriteBuffer[4][1] , \addressToWriteBuffer[4][0] ,
         \addressToWriteBuffer[3][7] , \addressToWriteBuffer[3][6] ,
         \addressToWriteBuffer[3][5] , \addressToWriteBuffer[3][4] ,
         \addressToWriteBuffer[3][3] , \addressToWriteBuffer[3][2] ,
         \addressToWriteBuffer[3][1] , \addressToWriteBuffer[3][0] ,
         \addressToWriteBuffer[2][7] , \addressToWriteBuffer[2][6] ,
         \addressToWriteBuffer[2][5] , \addressToWriteBuffer[2][4] ,
         \addressToWriteBuffer[2][3] , \addressToWriteBuffer[2][2] ,
         \addressToWriteBuffer[2][1] , \addressToWriteBuffer[2][0] ,
         \addressToWriteBuffer[1][7] , \addressToWriteBuffer[1][6] ,
         \addressToWriteBuffer[1][5] , \addressToWriteBuffer[1][4] ,
         \addressToWriteBuffer[1][3] , \addressToWriteBuffer[1][2] ,
         \addressToWriteBuffer[1][1] , \addressToWriteBuffer[1][0] ,
         \addressToWriteBuffer[0][7] , \addressToWriteBuffer[0][6] ,
         \addressToWriteBuffer[0][5] , \addressToWriteBuffer[0][4] ,
         \addressToWriteBuffer[0][3] , \addressToWriteBuffer[0][2] ,
         \addressToWriteBuffer[0][1] , \addressToWriteBuffer[0][0] ,
         \requesterAddressBuffer[1][3] , \requesterAddressBuffer[1][2] ,
         \requesterAddressBuffer[1][1] , \requesterAddressBuffer[1][0] ,
         \requesterAddressBuffer[0][3] , \requesterAddressBuffer[0][2] ,
         \requesterAddressBuffer[0][1] , \requesterAddressBuffer[0][0] ,
         \requesterPortBuffer[5][1] , \requesterPortBuffer[5][0] ,
         \requesterPortBuffer[4][0] , \requesterPortBuffer[3][1] ,
         \requesterPortBuffer[3][0] , \requesterPortBuffer[2][1] ,
         \requesterPortBuffer[2][0] , \requesterPortBuffer[1][1] ,
         \requesterPortBuffer[1][0] , \requesterPortBuffer[0][1] ,
         \requesterPortBuffer[0][0] , \prevRequesterPort_B[1] ,
         \prevRequesterPort_A[0] , prevMemRead_B, prevMemRead_A, N5316, N5324,
         N5332, N5340, N5373, N5374, N5375, N5376, N5377, N5378, N5381, N5382,
         N5383, N5384, N5385, N5386, N5389, N5390, N5391, N5392, N5393, N5394,
         N5397, N5398, N5399, N5400, N5401, N5402, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1214, n1215, n1216, n1217, n1218, n1219, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1272,
         n1273, n1274, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837;
  wire   [7:0] isWrite;
  wire   [3:0] prevRequesterAddress_B;
  wire   [3:0] prevRequesterAddress_A;

  EDFFX1TS \readReady_Concatenated_reg[3]  ( .D(N5340), .E(n837), .CK(clk), 
        .Q(readReady_WEST) );
  EDFFX1TS \readReady_Concatenated_reg[2]  ( .D(N5332), .E(n795), .CK(clk), 
        .Q(readReady_EAST) );
  EDFFX1TS \readReady_Concatenated_reg[1]  ( .D(N5324), .E(n795), .CK(clk), 
        .Q(readReady_SOUTH) );
  EDFFX1TS \readReady_Concatenated_reg[0]  ( .D(N5316), .E(n717), .CK(clk), 
        .Q(readReady_NORTH) );
  DFFNSRX1TS \requesterPortBuffer_reg[4][1]  ( .D(n1274), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n833) );
  DFFNSRX1TS \requesterAddressBuffer_reg[1][3]  ( .D(n1347), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressBuffer[1][3] ) );
  DFFNSRX1TS \requesterAddressBuffer_reg[1][2]  ( .D(n1348), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressBuffer[1][2] ) );
  DFFNSRX1TS \requesterAddressBuffer_reg[1][1]  ( .D(n1349), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressBuffer[1][1] ) );
  DFFNSRX1TS \requesterAddressBuffer_reg[1][0]  ( .D(n1350), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressBuffer[1][0] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[0][5]  ( .D(n1262), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[0][5] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[0][4]  ( .D(n1263), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[0][4] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[0][3]  ( .D(n1264), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[0][3] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[0][2]  ( .D(n1265), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[0][2] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[0][1]  ( .D(n1266), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[0][1] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[0][0]  ( .D(n1267), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[0][0] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[0][7]  ( .D(n1339), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[0][7] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[0][6]  ( .D(n1340), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[0][6] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[0][5]  ( .D(n1341), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[0][5] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[0][4]  ( .D(n1342), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[0][4] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[0][3]  ( .D(n1343), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[0][3] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[0][2]  ( .D(n1344), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[0][2] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[0][1]  ( .D(n1345), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[0][1] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[0][0]  ( .D(n1346), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[0][0] ) );
  DFFNSRX1TS \requesterPortBuffer_reg[0][1]  ( .D(n1282), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[0][1] ) );
  DFFNSRX1TS \requesterPortBuffer_reg[0][0]  ( .D(n1363), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[0][0] ) );
  DFFNSRX1TS \requesterAddressBuffer_reg[0][3]  ( .D(n1351), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressBuffer[0][3] ) );
  DFFNSRX1TS \requesterAddressBuffer_reg[0][2]  ( .D(n1352), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressBuffer[0][2] ) );
  DFFNSRX1TS \requesterAddressBuffer_reg[0][1]  ( .D(n1353), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressBuffer[0][1] ) );
  DFFNSRX1TS \requesterAddressBuffer_reg[0][0]  ( .D(n1354), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressBuffer[0][0] ) );
  DFFNSRX1TS \requesterPortBuffer_reg[1][1]  ( .D(n1280), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[1][1] ) );
  DFFNSRX1TS \requesterPortBuffer_reg[1][0]  ( .D(n1281), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[1][0] ) );
  DFFNSRX1TS \isWrite_reg[3]  ( .D(n1216), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(isWrite[3]) );
  DFFNSRX1TS \requesterPortBuffer_reg[4][0]  ( .D(n827), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[4][0] ) );
  DFFNSRX1TS \isWrite_reg[4]  ( .D(n1215), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(isWrite[4]) );
  DFFNSRX1TS \dataToWriteBuffer_reg[4][5]  ( .D(n1238), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[4][5] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[4][4]  ( .D(n1239), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[4][4] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[4][3]  ( .D(n1240), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[4][3] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[4][2]  ( .D(n1241), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[4][2] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[4][1]  ( .D(n1242), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[4][1] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[4][0]  ( .D(n1243), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[4][0] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[4][7]  ( .D(n1307), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[4][7] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[4][6]  ( .D(n1308), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[4][6] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[4][5]  ( .D(n1309), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[4][5] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[4][4]  ( .D(n1310), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[4][4] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[4][3]  ( .D(n1311), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[4][3] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[4][2]  ( .D(n1312), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[4][2] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[4][1]  ( .D(n1313), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[4][1] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[4][0]  ( .D(n1314), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[4][0] ) );
  DFFNSRX1TS \isWrite_reg[2]  ( .D(n1217), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(isWrite[2]) );
  DFFNSRX1TS \dataToWriteBuffer_reg[1][5]  ( .D(n1256), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[1][5] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[1][4]  ( .D(n1257), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[1][4] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[1][3]  ( .D(n1258), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[1][3] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[1][2]  ( .D(n1259), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[1][2] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[1][1]  ( .D(n1260), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[1][1] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[1][0]  ( .D(n1261), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[1][0] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[1][7]  ( .D(n1331), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[1][7] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[1][6]  ( .D(n1332), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[1][6] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[1][5]  ( .D(n1333), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[1][5] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[1][4]  ( .D(n1334), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[1][4] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[1][3]  ( .D(n1335), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[1][3] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[1][2]  ( .D(n1336), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[1][2] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[1][1]  ( .D(n1337), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[1][1] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[1][0]  ( .D(n1338), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[1][0] ) );
  DFFNSRX1TS \requesterPortBuffer_reg[3][0]  ( .D(n1277), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[3][0] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[3][5]  ( .D(n1244), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[3][5] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[3][4]  ( .D(n1245), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[3][4] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[3][3]  ( .D(n1246), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[3][3] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[3][2]  ( .D(n1247), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[3][2] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[3][1]  ( .D(n1248), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[3][1] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[3][0]  ( .D(n1249), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[3][0] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[3][7]  ( .D(n1315), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[3][7] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[3][6]  ( .D(n1316), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[3][6] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[3][5]  ( .D(n1317), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[3][5] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[3][4]  ( .D(n1318), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[3][4] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[3][3]  ( .D(n1319), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[3][3] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[3][2]  ( .D(n1320), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[3][2] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[3][1]  ( .D(n1321), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[3][1] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[3][0]  ( .D(n1322), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[3][0] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[5][5]  ( .D(n1232), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[5][5] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[5][4]  ( .D(n1233), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[5][4] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[5][3]  ( .D(n1234), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[5][3] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[5][2]  ( .D(n1235), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[5][2] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[5][1]  ( .D(n1236), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[5][1] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[5][0]  ( .D(n1237), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[5][0] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[5][7]  ( .D(n1299), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[5][7] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[5][6]  ( .D(n1300), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[5][6] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[5][5]  ( .D(n1301), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[5][5] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[5][4]  ( .D(n1302), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[5][4] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[5][3]  ( .D(n1303), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[5][3] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[5][2]  ( .D(n1304), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[5][2] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[5][1]  ( .D(n1305), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[5][1] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[5][0]  ( .D(n1306), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[5][0] ) );
  DFFNSRX1TS \requesterPortBuffer_reg[2][0]  ( .D(n1279), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[2][0] ) );
  DFFNSRX1TS \isWrite_reg[0]  ( .D(n1219), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(isWrite[0]) );
  DFFNSRX1TS \dataToWriteBuffer_reg[2][5]  ( .D(n1250), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[2][5] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[2][4]  ( .D(n1251), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[2][4] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[2][3]  ( .D(n1252), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[2][3] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[2][2]  ( .D(n1253), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[2][2] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[2][1]  ( .D(n1254), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[2][1] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[2][0]  ( .D(n1255), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[2][0] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[2][7]  ( .D(n1323), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[2][7] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[2][6]  ( .D(n1324), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[2][6] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[2][5]  ( .D(n1325), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[2][5] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[2][4]  ( .D(n1326), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[2][4] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[2][3]  ( .D(n1327), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[2][3] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[2][2]  ( .D(n1328), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[2][2] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[2][1]  ( .D(n1329), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[2][1] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[2][0]  ( .D(n1330), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[2][0] ) );
  DFFNSRX1TS \requesterPortBuffer_reg[2][1]  ( .D(n1278), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[2][1] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[6][5]  ( .D(n1226), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[6][5] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[6][4]  ( .D(n1227), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[6][4] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[6][3]  ( .D(n1228), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[6][3] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[6][2]  ( .D(n1229), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[6][2] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[6][1]  ( .D(n1230), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[6][1] ) );
  DFFNSRX1TS \dataToWriteBuffer_reg[6][0]  ( .D(n1231), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[6][0] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[6][7]  ( .D(n1291), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[6][7] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[6][6]  ( .D(n1292), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[6][6] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[6][5]  ( .D(n1293), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[6][5] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[6][4]  ( .D(n1294), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[6][4] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[6][3]  ( .D(n1295), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[6][3] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[6][2]  ( .D(n1296), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[6][2] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[6][1]  ( .D(n1297), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[6][1] ) );
  DFFNSRX1TS \addressToWriteBuffer_reg[6][0]  ( .D(n1298), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[6][0] ) );
  DFFNSRX1TS \requesterPortBuffer_reg[3][1]  ( .D(n1276), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[3][1] ) );
  DFFNSRX1TS \requesterPortBuffer_reg[5][0]  ( .D(n1273), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[5][0] ) );
  DFFNSRX1TS \requesterPortBuffer_reg[5][1]  ( .D(n1272), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[5][1] ) );
  DFFNSRX1TS \nextEmptyBuffer_reg[1]  ( .D(n1210), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(N742), .QN(n12) );
  DFFNSRX1TS \nextEmptyBuffer_reg[0]  ( .D(n1211), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(N741) );
  DFFNSRX1TS prevMemRead_B_reg ( .D(n1204), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(prevMemRead_B) );
  DFFNSRX1TS prevMemRead_A_reg ( .D(n1203), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(prevMemRead_A) );
  DFFNSRX1TS \prevRequesterAddress_A_reg[3]  ( .D(n1205), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_A[3]), .QN(n8) );
  DFFNSRX1TS \prevRequesterAddress_A_reg[2]  ( .D(n1206), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_A[2]), .QN(n9) );
  DFFNSRX1TS \prevRequesterAddress_A_reg[1]  ( .D(n1207), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_A[1]), .QN(n10) );
  DFFNSRX1TS \prevRequesterAddress_A_reg[0]  ( .D(n1208), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_A[0]), .QN(n11) );
  TLATXLTS \dataOut_Concatenated_reg[3][5]  ( .G(clk), .D(N5402), .Q(
        cacheDataOut_WEST[5]) );
  TLATXLTS \dataOut_Concatenated_reg[3][4]  ( .G(clk), .D(N5401), .Q(
        cacheDataOut_WEST[4]) );
  TLATXLTS \dataOut_Concatenated_reg[3][3]  ( .G(clk), .D(N5400), .Q(
        cacheDataOut_WEST[3]) );
  TLATXLTS \dataOut_Concatenated_reg[3][2]  ( .G(clk), .D(N5399), .Q(
        cacheDataOut_WEST[2]) );
  TLATXLTS \dataOut_Concatenated_reg[3][1]  ( .G(clk), .D(N5398), .Q(
        cacheDataOut_WEST[1]) );
  TLATXLTS \dataOut_Concatenated_reg[3][0]  ( .G(clk), .D(N5397), .Q(
        cacheDataOut_WEST[0]) );
  TLATXLTS \dataOut_Concatenated_reg[2][5]  ( .G(clk), .D(N5394), .Q(
        cacheDataOut_EAST[5]) );
  TLATXLTS \dataOut_Concatenated_reg[2][4]  ( .G(clk), .D(N5393), .Q(
        cacheDataOut_EAST[4]) );
  TLATXLTS \dataOut_Concatenated_reg[2][3]  ( .G(clk), .D(N5392), .Q(
        cacheDataOut_EAST[3]) );
  TLATXLTS \dataOut_Concatenated_reg[2][2]  ( .G(clk), .D(N5391), .Q(
        cacheDataOut_EAST[2]) );
  TLATXLTS \dataOut_Concatenated_reg[2][1]  ( .G(clk), .D(N5390), .Q(
        cacheDataOut_EAST[1]) );
  TLATXLTS \dataOut_Concatenated_reg[2][0]  ( .G(clk), .D(N5389), .Q(
        cacheDataOut_EAST[0]) );
  TLATXLTS \dataOut_Concatenated_reg[1][5]  ( .G(clk), .D(N5386), .Q(
        cacheDataOut_SOUTH[5]) );
  TLATXLTS \dataOut_Concatenated_reg[1][4]  ( .G(clk), .D(N5385), .Q(
        cacheDataOut_SOUTH[4]) );
  TLATXLTS \dataOut_Concatenated_reg[1][3]  ( .G(clk), .D(N5384), .Q(
        cacheDataOut_SOUTH[3]) );
  TLATXLTS \dataOut_Concatenated_reg[1][2]  ( .G(clk), .D(N5383), .Q(
        cacheDataOut_SOUTH[2]) );
  TLATXLTS \dataOut_Concatenated_reg[1][1]  ( .G(clk), .D(N5382), .Q(
        cacheDataOut_SOUTH[1]) );
  TLATXLTS \dataOut_Concatenated_reg[1][0]  ( .G(clk), .D(N5381), .Q(
        cacheDataOut_SOUTH[0]) );
  TLATXLTS \dataOut_Concatenated_reg[0][5]  ( .G(clk), .D(N5378), .Q(
        cacheDataOut_NORTH[5]) );
  TLATXLTS \dataOut_Concatenated_reg[0][4]  ( .G(clk), .D(N5377), .Q(
        cacheDataOut_NORTH[4]) );
  TLATXLTS \dataOut_Concatenated_reg[0][3]  ( .G(clk), .D(N5376), .Q(
        cacheDataOut_NORTH[3]) );
  TLATXLTS \dataOut_Concatenated_reg[0][2]  ( .G(clk), .D(N5375), .Q(
        cacheDataOut_NORTH[2]) );
  TLATXLTS \dataOut_Concatenated_reg[0][1]  ( .G(clk), .D(N5374), .Q(
        cacheDataOut_NORTH[1]) );
  TLATXLTS \dataOut_Concatenated_reg[0][0]  ( .G(clk), .D(N5373), .Q(
        cacheDataOut_NORTH[0]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[3][3]  ( .D(n1171), .CK(clk), 
        .Q(requesterAddressOut_WEST[3]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[3][2]  ( .D(n1170), .CK(clk), 
        .Q(requesterAddressOut_WEST[2]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[3][1]  ( .D(n1169), .CK(clk), 
        .Q(requesterAddressOut_WEST[1]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[2][3]  ( .D(n1167), .CK(clk), 
        .Q(requesterAddressOut_EAST[3]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[2][2]  ( .D(n1166), .CK(clk), 
        .Q(requesterAddressOut_EAST[2]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[2][1]  ( .D(n1165), .CK(clk), 
        .Q(requesterAddressOut_EAST[1]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[1][3]  ( .D(n1163), .CK(clk), 
        .Q(requesterAddressOut_SOUTH[3]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[1][2]  ( .D(n1162), .CK(clk), 
        .Q(requesterAddressOut_SOUTH[2]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[1][1]  ( .D(n1161), .CK(clk), 
        .Q(requesterAddressOut_SOUTH[1]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[3][0]  ( .D(n1168), .CK(clk), 
        .Q(requesterAddressOut_WEST[0]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[2][0]  ( .D(n1164), .CK(clk), 
        .Q(requesterAddressOut_EAST[0]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[1][0]  ( .D(n1160), .CK(clk), 
        .Q(requesterAddressOut_SOUTH[0]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[0][3]  ( .D(n1159), .CK(clk), 
        .Q(requesterAddressOut_NORTH[3]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[0][2]  ( .D(n1158), .CK(clk), 
        .Q(requesterAddressOut_NORTH[2]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[0][1]  ( .D(n1157), .CK(clk), 
        .Q(requesterAddressOut_NORTH[1]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[0][0]  ( .D(n1156), .CK(clk), 
        .Q(requesterAddressOut_NORTH[0]) );
  DFFNSRX1TS \prevRequesterPort_A_reg[1]  ( .D(n1355), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n4), .QN(n18) );
  DFFNSRX1TS \prevRequesterPort_A_reg[0]  ( .D(n1356), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\prevRequesterPort_A[0] ), .QN(n6) );
  DFFNSRX1TS \prevRequesterPort_B_reg[1]  ( .D(n1357), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\prevRequesterPort_B[1] ), .QN(n5) );
  DFFNSRX1TS \prevRequesterPort_B_reg[0]  ( .D(n1358), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n7), .QN(n20) );
  DFFNSRX1TS memWrite_B_reg ( .D(n1202), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        memWrite_B) );
  DFFNSRX1TS memWrite_A_reg ( .D(n1181), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        memWrite_A) );
  DFFNSRX1TS \cacheDataIn_A_reg[5]  ( .D(n1196), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[5]) );
  DFFNSRX1TS \cacheDataIn_A_reg[4]  ( .D(n1197), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[4]) );
  DFFNSRX1TS \cacheDataIn_A_reg[3]  ( .D(n1198), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[3]) );
  DFFNSRX1TS \cacheDataIn_A_reg[2]  ( .D(n1199), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[2]) );
  DFFNSRX1TS \cacheDataIn_A_reg[1]  ( .D(n1200), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[1]) );
  DFFNSRX1TS \cacheDataIn_A_reg[0]  ( .D(n1201), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[0]) );
  DFFNSRX1TS \cacheAddressIn_B_reg[7]  ( .D(n1195), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_B[7]) );
  DFFNSRX1TS \cacheAddressIn_B_reg[6]  ( .D(n1194), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_B[6]) );
  DFFNSRX1TS \cacheAddressIn_B_reg[5]  ( .D(n1193), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_B[5]) );
  DFFNSRX1TS \cacheAddressIn_B_reg[4]  ( .D(n1192), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_B[4]) );
  DFFNSRX1TS \cacheAddressIn_B_reg[3]  ( .D(n1191), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_B[3]) );
  DFFNSRX1TS \cacheAddressIn_B_reg[2]  ( .D(n1190), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_B[2]) );
  DFFNSRX1TS \cacheAddressIn_B_reg[1]  ( .D(n1189), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_B[1]) );
  DFFNSRX1TS \cacheAddressIn_B_reg[0]  ( .D(n1188), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_B[0]) );
  DFFNSRX1TS \cacheDataIn_B_reg[5]  ( .D(n1187), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[5]) );
  DFFNSRX1TS \cacheDataIn_B_reg[4]  ( .D(n1186), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[4]) );
  DFFNSRX1TS \cacheDataIn_B_reg[3]  ( .D(n1185), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[3]) );
  DFFNSRX1TS \cacheDataIn_B_reg[2]  ( .D(n1184), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[2]) );
  DFFNSRX1TS \cacheDataIn_B_reg[1]  ( .D(n1183), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[1]) );
  DFFNSRX1TS \cacheDataIn_B_reg[0]  ( .D(n1182), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[0]) );
  DFFNSRX1TS \cacheAddressIn_A_reg[7]  ( .D(n1180), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_A[7]) );
  DFFNSRX1TS \cacheAddressIn_A_reg[6]  ( .D(n1179), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_A[6]) );
  DFFNSRX1TS \cacheAddressIn_A_reg[5]  ( .D(n1178), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_A[5]) );
  DFFNSRX1TS \cacheAddressIn_A_reg[4]  ( .D(n1177), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_A[4]) );
  DFFNSRX1TS \cacheAddressIn_A_reg[3]  ( .D(n1176), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_A[3]) );
  DFFNSRX1TS \cacheAddressIn_A_reg[2]  ( .D(n1175), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_A[2]) );
  DFFNSRX1TS \cacheAddressIn_A_reg[1]  ( .D(n1174), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_A[1]) );
  DFFNSRX1TS \cacheAddressIn_A_reg[0]  ( .D(n1173), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_A[0]) );
  DFFNSRX1TS \nextEmptyBuffer_reg[2]  ( .D(n1209), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n836), .QN(n832) );
  DFFNSRX1TS \isWrite_reg[5]  ( .D(n1214), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(isWrite[5]), .QN(n835) );
  DFFNSRX1TS \prevRequesterAddress_B_reg[2]  ( .D(n1360), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_B[2]), .QN(n829) );
  DFFNSRX1TS \prevRequesterAddress_B_reg[1]  ( .D(n1361), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_B[1]), .QN(n830) );
  DFFNSRX1TS \prevRequesterAddress_B_reg[0]  ( .D(n1362), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_B[0]), .QN(n831) );
  DFFNSRX1TS \prevRequesterAddress_B_reg[3]  ( .D(n1359), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_B[3]), .QN(n828) );
  DFFNSRX1TS \isWrite_reg[1]  ( .D(n1218), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(isWrite[1]), .QN(n834) );
  CLKBUFX2TS U3 ( .A(n55), .Y(n536) );
  CLKBUFX2TS U4 ( .A(n34), .Y(n81) );
  INVX2TS U5 ( .A(n15), .Y(n633) );
  NOR2XLTS U6 ( .A(n685), .B(n353), .Y(n354) );
  NOR2XLTS U7 ( .A(n685), .B(n460), .Y(n56) );
  NOR2XLTS U8 ( .A(n52), .B(n836), .Y(n36) );
  NOR2XLTS U9 ( .A(N741), .B(n572), .Y(n40) );
  NOR2XLTS U10 ( .A(n228), .B(n138), .Y(n139) );
  INVX2TS U11 ( .A(memWrite_NORTH), .Y(n674) );
  INVX2TS U12 ( .A(n645), .Y(n632) );
  NOR2XLTS U13 ( .A(memRead_EAST), .B(memWrite_EAST), .Y(n33) );
  CLKBUFX2TS U14 ( .A(n442), .Y(n443) );
  INVX2TS U15 ( .A(n252), .Y(n270) );
  INVX2TS U16 ( .A(n35), .Y(n501) );
  NOR2XLTS U17 ( .A(\prevRequesterPort_A[0] ), .B(n192), .Y(n193) );
  CLKBUFX2TS U18 ( .A(n448), .Y(n556) );
  NAND2X1TS U19 ( .A(n351), .B(n353), .Y(n350) );
  NAND3X1TS U20 ( .A(n608), .B(n671), .C(n574), .Y(n611) );
  CLKBUFX2TS U21 ( .A(n764), .Y(n711) );
  INVX2TS U22 ( .A(n48), .Y(n340) );
  XNOR2X1TS U23 ( .A(n632), .B(n47), .Y(n48) );
  CLKBUFX2TS U24 ( .A(n691), .Y(n724) );
  NOR3BX1TS U25 ( .AN(n574), .B(n441), .C(n307), .Y(n54) );
  NOR3X1TS U26 ( .A(n633), .B(n334), .C(n133), .Y(n134) );
  NOR2X1TS U27 ( .A(n501), .B(n521), .Y(n53) );
  NOR2X1TS U28 ( .A(n512), .B(n578), .Y(n672) );
  NAND3X1TS U29 ( .A(n27), .B(n194), .C(n7), .Y(n3) );
  NOR2X1TS U30 ( .A(memRead_NORTH), .B(memWrite_NORTH), .Y(n34) );
  NOR2X1TS U31 ( .A(n44), .B(n49), .Y(n43) );
  NOR3XLTS U32 ( .A(n133), .B(n440), .C(n516), .Y(n441) );
  XOR2XLTS U33 ( .A(n334), .B(n336), .Y(n343) );
  NAND3XLTS U34 ( .A(n53), .B(n345), .C(n77), .Y(n574) );
  NOR2XLTS U35 ( .A(n44), .B(n77), .Y(n344) );
  NAND3XLTS U36 ( .A(n21), .B(N742), .C(n578), .Y(n338) );
  NOR2XLTS U37 ( .A(n45), .B(n49), .Y(n50) );
  AOI211XLTS U38 ( .A0(n34), .A1(n517), .B0(n673), .C0(n516), .Y(n652) );
  CLKAND2X2TS U39 ( .A(n518), .B(n684), .Y(n16) );
  NOR3XLTS U40 ( .A(n633), .B(n640), .C(n515), .Y(n673) );
  NOR4BXLTS U41 ( .AN(n44), .B(n19), .C(n512), .D(n578), .Y(n438) );
  NOR2X1TS U42 ( .A(memRead_SOUTH), .B(memWrite_SOUTH), .Y(n514) );
  NOR2XLTS U43 ( .A(n133), .B(n80), .Y(n342) );
  AOI211XLTS U44 ( .A0(n81), .A1(n42), .B0(n339), .C0(n338), .Y(n355) );
  NOR2XLTS U45 ( .A(n13), .B(n78), .Y(n345) );
  INVX2TS U46 ( .A(n518), .Y(n513) );
  NAND2X1TS U47 ( .A(n440), .B(n135), .Y(n643) );
  NOR2XLTS U48 ( .A(n640), .B(n639), .Y(n641) );
  INVX2TS U49 ( .A(memWrite_SOUTH), .Y(n676) );
  NAND3XLTS U50 ( .A(n617), .B(n720), .C(n673), .Y(n650) );
  NOR3BXLTS U51 ( .AN(n672), .B(n521), .C(n677), .Y(n522) );
  INVX2TS U52 ( .A(n79), .Y(n440) );
  NAND3XLTS U53 ( .A(n32), .B(n580), .C(n332), .Y(n622) );
  INVX2TS U54 ( .A(cacheAddressIn_EAST[4]), .Y(n487) );
  INVX2TS U55 ( .A(cacheAddressIn_EAST[6]), .Y(n456) );
  INVX2TS U56 ( .A(cacheAddressIn_EAST[7]), .Y(n464) );
  OR2X1TS U57 ( .A(n516), .B(n513), .Y(n252) );
  OAI21XLTS U58 ( .A0(n621), .A1(n55), .B0(n609), .Y(n610) );
  OAI21XLTS U59 ( .A0(n224), .A1(n833), .B0(n223), .Y(n1276) );
  OAI211XLTS U60 ( .A0(n446), .A1(n833), .B0(n445), .C0(n444), .Y(n1278) );
  OAI21XLTS U61 ( .A0(n451), .A1(n450), .B0(n449), .Y(n1279) );
  AOI2BB2XLTS U62 ( .B0(n435), .B1(n42), .A0N(n336), .A1N(n435), .Y(n78) );
  NOR2X1TS U63 ( .A(n35), .B(n672), .Y(n435) );
  CLKAND2X2TS U64 ( .A(n13), .B(n344), .Y(n83) );
  NOR3BXLTS U65 ( .AN(n7), .B(n194), .C(n816), .Y(n29) );
  NOR3BXLTS U66 ( .AN(n194), .B(n7), .C(n23), .Y(n24) );
  INVX2TS U67 ( .A(memWrite_WEST), .Y(n621) );
  AOI31XLTS U68 ( .A0(n32), .A1(n633), .A2(n341), .B0(n719), .Y(n608) );
  NOR2XLTS U69 ( .A(n134), .B(n500), .Y(n243) );
  NAND3XLTS U70 ( .A(n532), .B(n135), .C(n681), .Y(n138) );
  CLKAND2X2TS U71 ( .A(n84), .B(n678), .Y(n85) );
  INVX2TS U72 ( .A(cacheAddressIn_EAST[5]), .Y(n147) );
  OR2X1TS U73 ( .A(n608), .B(n346), .Y(n543) );
  OAI21XLTS U74 ( .A0(n649), .A1(n648), .B0(n646), .Y(n647) );
  OAI32X1TS U75 ( .A0(memRead_EAST), .A1(memRead_SOUTH), .A2(n674), .B0(n676), 
        .B1(memRead_EAST), .Y(n626) );
  NAND3XLTS U76 ( .A(n776), .B(n775), .C(n774), .Y(n1173) );
  NAND3XLTS U77 ( .A(n768), .B(n767), .C(n766), .Y(n1174) );
  NAND3XLTS U78 ( .A(n760), .B(n759), .C(n758), .Y(n1175) );
  NAND3XLTS U79 ( .A(n752), .B(n751), .C(n750), .Y(n1176) );
  NAND3XLTS U80 ( .A(n744), .B(n743), .C(n742), .Y(n1177) );
  NAND3XLTS U81 ( .A(n738), .B(n737), .C(n736), .Y(n1178) );
  NAND3XLTS U82 ( .A(n732), .B(n731), .C(n730), .Y(n1179) );
  NAND3XLTS U83 ( .A(n727), .B(n726), .C(n725), .Y(n1180) );
  NAND3XLTS U84 ( .A(n689), .B(n688), .C(n687), .Y(n1201) );
  NAND3XLTS U85 ( .A(n694), .B(n693), .C(n692), .Y(n1200) );
  NAND3XLTS U86 ( .A(n698), .B(n697), .C(n696), .Y(n1199) );
  NAND3XLTS U87 ( .A(n705), .B(n704), .C(n703), .Y(n1198) );
  NAND3XLTS U88 ( .A(n710), .B(n709), .C(n708), .Y(n1197) );
  NAND3XLTS U89 ( .A(n716), .B(n715), .C(n714), .Y(n1196) );
  AO22XLTS U90 ( .A0(n682), .A1(memWrite_B), .B0(n681), .B1(n680), .Y(n1202)
         );
  OAI211XLTS U91 ( .A0(n501), .A1(n500), .B0(n499), .C0(n498), .Y(n1358) );
  OAI211XLTS U92 ( .A0(n229), .A1(n500), .B0(n496), .C0(n498), .Y(n1357) );
  NAND3BXLTS U93 ( .AN(n724), .B(n520), .C(n650), .Y(n1356) );
  NAND3BXLTS U94 ( .AN(n746), .B(n523), .C(n650), .Y(n1355) );
  NAND3XLTS U95 ( .A(n656), .B(n655), .C(n654), .Y(n1208) );
  NAND3XLTS U96 ( .A(n659), .B(n658), .C(n657), .Y(n1207) );
  NAND3XLTS U97 ( .A(n663), .B(n662), .C(n661), .Y(n1206) );
  NAND3XLTS U98 ( .A(n670), .B(n669), .C(n668), .Y(n1205) );
  AOI211XLTS U99 ( .A0(n440), .A1(n439), .B0(n679), .C0(n677), .Y(n1204) );
  NAND3XLTS U100 ( .A(n622), .B(n582), .C(n581), .Y(n1273) );
  OAI21XLTS U101 ( .A0(n834), .A1(n224), .B0(n222), .Y(n1219) );
  AO21XLTS U102 ( .A0(cacheAddressIn_NORTH[0]), .A1(n426), .B0(n359), .Y(n1306) );
  AO21XLTS U103 ( .A0(n434), .A1(cacheAddressIn_NORTH[1]), .B0(n402), .Y(n1305) );
  OAI211XLTS U104 ( .A0(n432), .A1(n401), .B0(n400), .C0(n399), .Y(n402) );
  AO21XLTS U105 ( .A0(n417), .A1(cacheAddressIn_NORTH[2]), .B0(n416), .Y(n1304) );
  OAI211XLTS U106 ( .A0(n415), .A1(n414), .B0(n413), .C0(n412), .Y(n416) );
  AO21XLTS U107 ( .A0(n409), .A1(cacheAddressIn_NORTH[3]), .B0(n408), .Y(n1303) );
  OAI211XLTS U108 ( .A0(n352), .A1(n407), .B0(n406), .C0(n405), .Y(n408) );
  AO21XLTS U109 ( .A0(n409), .A1(cacheAddressIn_NORTH[4]), .B0(n367), .Y(n1302) );
  AO21XLTS U110 ( .A0(n426), .A1(cacheAddressIn_NORTH[5]), .B0(n378), .Y(n1301) );
  AO21XLTS U111 ( .A0(n417), .A1(cacheAddressIn_NORTH[6]), .B0(n373), .Y(n1300) );
  AO21XLTS U112 ( .A0(n434), .A1(cacheAddressIn_NORTH[7]), .B0(n363), .Y(n1299) );
  AO21XLTS U113 ( .A0(n434), .A1(dataIn_NORTH[0]), .B0(n433), .Y(n1237) );
  OAI211XLTS U114 ( .A0(n432), .A1(n431), .B0(n430), .C0(n429), .Y(n433) );
  AO21XLTS U115 ( .A0(n426), .A1(dataIn_NORTH[1]), .B0(n425), .Y(n1236) );
  OAI211XLTS U116 ( .A0(n424), .A1(n423), .B0(n422), .C0(n421), .Y(n425) );
  AO21XLTS U117 ( .A0(n434), .A1(dataIn_NORTH[2]), .B0(n382), .Y(n1235) );
  AO21XLTS U118 ( .A0(n417), .A1(dataIn_NORTH[3]), .B0(n391), .Y(n1234) );
  OAI211XLTS U119 ( .A0(n415), .A1(n390), .B0(n389), .C0(n388), .Y(n391) );
  AO21XLTS U120 ( .A0(n426), .A1(dataIn_NORTH[4]), .B0(n396), .Y(n1233) );
  OAI211XLTS U121 ( .A0(n424), .A1(n395), .B0(n394), .C0(n393), .Y(n396) );
  AO21XLTS U122 ( .A0(n409), .A1(dataIn_NORTH[5]), .B0(n386), .Y(n1232) );
  OAI211XLTS U123 ( .A0(n352), .A1(n385), .B0(n384), .C0(n383), .Y(n386) );
  OAI211XLTS U124 ( .A0(n468), .A1(n494), .B0(n467), .C0(n466), .Y(n1336) );
  OAI211XLTS U125 ( .A0(n487), .A1(n486), .B0(n485), .C0(n484), .Y(n1334) );
  OAI211XLTS U126 ( .A0(n456), .A1(n472), .B0(n455), .C0(n454), .Y(n1332) );
  OAI211XLTS U127 ( .A0(n464), .A1(n486), .B0(n463), .C0(n462), .Y(n1331) );
  OAI211XLTS U128 ( .A0(n459), .A1(n478), .B0(n458), .C0(n457), .Y(n1261) );
  OAI211XLTS U129 ( .A0(n473), .A1(n472), .B0(n471), .C0(n470), .Y(n1260) );
  OAI211XLTS U130 ( .A0(n479), .A1(n478), .B0(n477), .C0(n476), .Y(n1257) );
  OAI211XLTS U131 ( .A0(n495), .A1(n494), .B0(n493), .C0(n492), .Y(n1256) );
  AO21XLTS U132 ( .A0(n577), .A1(\requesterPortBuffer[1][0] ), .B0(n571), .Y(
        n1281) );
  AO21XLTS U133 ( .A0(n577), .A1(\requesterPortBuffer[1][1] ), .B0(n576), .Y(
        n1280) );
  OAI21XLTS U134 ( .A0(n252), .A1(n833), .B0(n221), .Y(n1274) );
  AO22XLTS U135 ( .A0(n508), .A1(prevMemRead_A), .B0(n504), .B1(prevMemRead_B), 
        .Y(N5316) );
  AO22XLTS U136 ( .A0(n808), .A1(prevMemRead_A), .B0(n804), .B1(prevMemRead_B), 
        .Y(N5324) );
  AO22XLTS U137 ( .A0(n793), .A1(prevMemRead_A), .B0(n791), .B1(prevMemRead_B), 
        .Y(N5332) );
  NOR2BX1TS U138 ( .AN(n519), .B(n4), .Y(n28) );
  NOR2BX1TS U139 ( .AN(n4), .B(n519), .Y(n22) );
  NOR2BX1TS U140 ( .AN(n443), .B(n806), .Y(n546) );
  NOR3BX2TS U141 ( .AN(n347), .B(n350), .C(n355), .Y(n348) );
  NOR2BX1TS U142 ( .AN(n56), .B(n536), .Y(n57) );
  NOR2XLTS U143 ( .A(n81), .B(n514), .Y(n35) );
  INVX2TS U144 ( .A(n228), .Y(n229) );
  OA21XLTS U145 ( .A0(n35), .A1(n50), .B0(n632), .Y(n13) );
  OR2X1TS U146 ( .A(n685), .B(n684), .Y(n14) );
  OA21XLTS U147 ( .A0(n521), .A1(n672), .B0(n501), .Y(n15) );
  NOR4BXLTS U148 ( .AN(n342), .B(n343), .C(n806), .D(n48), .Y(n86) );
  NOR2BX1TS U149 ( .AN(n652), .B(n651), .Y(n653) );
  NAND2X1TS U150 ( .A(n355), .B(n678), .Y(n17) );
  OR2X1TS U151 ( .A(memRead_WEST), .B(memWrite_WEST), .Y(n19) );
  NOR2XLTS U152 ( .A(n537), .B(n451), .Y(n59) );
  OAI21XLTS U153 ( .A0(N741), .A1(n41), .B0(n217), .Y(n42) );
  INVX2TS U154 ( .A(n832), .Y(n21) );
  INVX2TS U162 ( .A(n6), .Y(n519) );
  INVX2TS U163 ( .A(n22), .Y(n25) );
  CLKBUFX2TS U164 ( .A(cacheDataOut_A[5]), .Y(n511) );
  INVX2TS U165 ( .A(n25), .Y(n23) );
  INVX2TS U166 ( .A(n24), .Y(n26) );
  INVX2TS U167 ( .A(n26), .Y(n791) );
  CLKBUFX2TS U168 ( .A(cacheDataOut_B[5]), .Y(n509) );
  AO22X2TS U169 ( .A0(n23), .A1(n511), .B0(n791), .B1(n509), .Y(N5394) );
  INVX2TS U170 ( .A(n25), .Y(n799) );
  CLKBUFX2TS U171 ( .A(cacheDataOut_A[4]), .Y(n507) );
  CLKBUFX2TS U172 ( .A(cacheDataOut_B[4]), .Y(n505) );
  AO22X2TS U173 ( .A0(n799), .A1(n507), .B0(n791), .B1(n505), .Y(N5393) );
  INVX2TS U174 ( .A(n25), .Y(n793) );
  CLKBUFX2TS U175 ( .A(cacheDataOut_A[3]), .Y(n215) );
  INVX2TS U176 ( .A(n26), .Y(n796) );
  CLKBUFX2TS U177 ( .A(cacheDataOut_B[3]), .Y(n214) );
  AO22X2TS U178 ( .A0(n793), .A1(n215), .B0(n796), .B1(n214), .Y(N5392) );
  CLKBUFX2TS U179 ( .A(cacheDataOut_A[2]), .Y(n213) );
  INVX2TS U180 ( .A(n26), .Y(n798) );
  CLKBUFX2TS U181 ( .A(cacheDataOut_B[2]), .Y(n212) );
  AO22X2TS U182 ( .A0(n22), .A1(n213), .B0(n798), .B1(n212), .Y(N5391) );
  CLKBUFX2TS U183 ( .A(cacheDataOut_A[1]), .Y(n211) );
  CLKBUFX2TS U184 ( .A(cacheDataOut_B[1]), .Y(n210) );
  AO22X2TS U185 ( .A0(n793), .A1(n211), .B0(n796), .B1(n210), .Y(N5390) );
  CLKBUFX2TS U186 ( .A(cacheDataOut_A[0]), .Y(n209) );
  CLKBUFX2TS U187 ( .A(cacheDataOut_B[0]), .Y(n208) );
  AO22X2TS U188 ( .A0(n22), .A1(n209), .B0(n798), .B1(n208), .Y(N5389) );
  NAND2X1TS U189 ( .A(n519), .B(n4), .Y(n27) );
  INVX2TS U190 ( .A(n27), .Y(n784) );
  INVX2TS U191 ( .A(n3), .Y(n786) );
  AO22X2TS U192 ( .A0(n784), .A1(n511), .B0(n786), .B1(n509), .Y(N5402) );
  INVX2TS U193 ( .A(n27), .Y(n781) );
  INVX2TS U194 ( .A(n3), .Y(n783) );
  AO22X2TS U195 ( .A0(n781), .A1(n507), .B0(n783), .B1(n505), .Y(N5401) );
  INVX2TS U196 ( .A(n27), .Y(n787) );
  AO22X2TS U197 ( .A0(n787), .A1(n215), .B0(n786), .B1(n214), .Y(N5400) );
  AO22X2TS U198 ( .A0(n784), .A1(n213), .B0(n783), .B1(n212), .Y(N5399) );
  INVX2TS U199 ( .A(n3), .Y(n777) );
  AO22X2TS U200 ( .A0(n781), .A1(n211), .B0(n777), .B1(n210), .Y(N5398) );
  AO22X2TS U201 ( .A0(n787), .A1(n209), .B0(n777), .B1(n208), .Y(N5397) );
  INVX2TS U202 ( .A(n28), .Y(n30) );
  INVX2TS U203 ( .A(n30), .Y(n816) );
  INVX2TS U204 ( .A(n29), .Y(n31) );
  INVX2TS U205 ( .A(n31), .Y(n815) );
  AO22X2TS U206 ( .A0(n816), .A1(n511), .B0(n815), .B1(n509), .Y(N5386) );
  INVX2TS U207 ( .A(n31), .Y(n811) );
  AO22X2TS U208 ( .A0(n808), .A1(n507), .B0(n811), .B1(n505), .Y(N5385) );
  INVX2TS U209 ( .A(n30), .Y(n808) );
  AO22X2TS U210 ( .A0(n808), .A1(n215), .B0(n815), .B1(n214), .Y(N5384) );
  INVX2TS U211 ( .A(n30), .Y(n805) );
  AO22X2TS U212 ( .A0(n805), .A1(n213), .B0(n811), .B1(n212), .Y(N5383) );
  INVX2TS U213 ( .A(n31), .Y(n804) );
  AO22X2TS U214 ( .A0(n816), .A1(n211), .B0(n804), .B1(n210), .Y(N5382) );
  AO22X2TS U215 ( .A0(n805), .A1(n209), .B0(n804), .B1(n208), .Y(N5381) );
  INVX2TS U216 ( .A(n19), .Y(n133) );
  INVX2TS U217 ( .A(n133), .Y(n32) );
  INVX2TS U218 ( .A(n32), .Y(n216) );
  INVX2TS U219 ( .A(n33), .Y(n76) );
  INVX2TS U220 ( .A(n76), .Y(n521) );
  INVX2TS U221 ( .A(n81), .Y(n512) );
  INVX2TS U222 ( .A(n514), .Y(n578) );
  INVX2TS U223 ( .A(n12), .Y(n52) );
  INVX2TS U224 ( .A(n36), .Y(n38) );
  NAND2X1TS U225 ( .A(n36), .B(N741), .Y(n217) );
  INVX2TS U226 ( .A(n217), .Y(n37) );
  INVX2TS U227 ( .A(n37), .Y(n535) );
  INVX2TS U228 ( .A(n535), .Y(n346) );
  NOR2XLTS U229 ( .A(n52), .B(n346), .Y(n645) );
  INVX2TS U230 ( .A(n38), .Y(n537) );
  INVX2TS U231 ( .A(n537), .Y(n39) );
  INVX2TS U232 ( .A(n36), .Y(n572) );
  INVX2TS U233 ( .A(n40), .Y(n137) );
  INVX2TS U234 ( .A(n137), .Y(n41) );
  INVX2TS U235 ( .A(n42), .Y(n51) );
  INVX2TS U236 ( .A(n51), .Y(n45) );
  INVX2TS U237 ( .A(n76), .Y(n44) );
  INVX2TS U238 ( .A(n435), .Y(n49) );
  INVX2TS U239 ( .A(n43), .Y(n227) );
  INVX2TS U240 ( .A(n227), .Y(n228) );
  AOI21X1TS U241 ( .A0(n44), .A1(n49), .B0(n228), .Y(n515) );
  INVX2TS U242 ( .A(n515), .Y(n334) );
  NOR2X1TS U243 ( .A(n45), .B(n334), .Y(n46) );
  INVX2TS U244 ( .A(n15), .Y(n79) );
  INVX2TS U245 ( .A(n53), .Y(n639) );
  OAI22X1TS U246 ( .A0(n46), .A1(n79), .B0(n639), .B1(n45), .Y(n47) );
  INVX2TS U247 ( .A(n41), .Y(n719) );
  INVX2TS U248 ( .A(reset), .Y(n795) );
  CLKBUFX2TS U249 ( .A(n795), .Y(n717) );
  CLKBUFX2TS U250 ( .A(n717), .Y(n197) );
  INVX2TS U251 ( .A(n197), .Y(n685) );
  INVX2TS U252 ( .A(n51), .Y(n336) );
  OAI21XLTS U253 ( .A0(n52), .A1(n35), .B0(n836), .Y(n77) );
  INVX2TS U254 ( .A(n40), .Y(n516) );
  CLKBUFX2TS U255 ( .A(n795), .Y(n196) );
  CLKBUFX2TS U256 ( .A(n196), .Y(n518) );
  CLKBUFX2TS U257 ( .A(n252), .Y(n230) );
  CLKBUFX2TS U258 ( .A(n230), .Y(n307) );
  INVX2TS U259 ( .A(n54), .Y(n73) );
  INVX2TS U260 ( .A(n73), .Y(n460) );
  CLKAND2X2TS U261 ( .A(n608), .B(n56), .Y(n68) );
  INVX2TS U262 ( .A(n68), .Y(n486) );
  INVX2TS U263 ( .A(cacheAddressIn_WEST[5]), .Y(n377) );
  INVX2TS U264 ( .A(n377), .Y(n734) );
  NAND2X1TS U265 ( .A(n343), .B(n41), .Y(n55) );
  INVX2TS U266 ( .A(n57), .Y(n452) );
  INVX2TS U267 ( .A(n73), .Y(n488) );
  AOI22X1TS U268 ( .A0(n734), .A1(n57), .B0(n488), .B1(
        \addressToWriteBuffer[1][5] ), .Y(n61) );
  OR2X1TS U269 ( .A(n685), .B(n217), .Y(n58) );
  INVX2TS U270 ( .A(n58), .Y(n62) );
  INVX2TS U271 ( .A(n65), .Y(n469) );
  CLKBUFX2TS U272 ( .A(n717), .Y(n678) );
  INVX2TS U273 ( .A(n678), .Y(n451) );
  INVX2TS U274 ( .A(n59), .Y(n453) );
  AOI22X1TS U275 ( .A0(n469), .A1(\addressToWriteBuffer[2][5] ), .B0(n59), 
        .B1(\addressToWriteBuffer[3][5] ), .Y(n60) );
  OAI211XLTS U276 ( .A0(n147), .A1(n486), .B0(n61), .C0(n60), .Y(n1333) );
  INVX2TS U277 ( .A(cacheAddressIn_EAST[1]), .Y(n144) );
  INVX2TS U278 ( .A(n68), .Y(n494) );
  INVX2TS U279 ( .A(cacheAddressIn_WEST[1]), .Y(n401) );
  INVX2TS U280 ( .A(n401), .Y(n765) );
  INVX2TS U281 ( .A(n452), .Y(n474) );
  AOI22X1TS U282 ( .A0(n765), .A1(n474), .B0(n488), .B1(
        \addressToWriteBuffer[1][1] ), .Y(n64) );
  INVX2TS U283 ( .A(n62), .Y(n65) );
  INVX2TS U284 ( .A(n453), .Y(n475) );
  AOI22X1TS U285 ( .A0(n62), .A1(\addressToWriteBuffer[2][1] ), .B0(n475), 
        .B1(\addressToWriteBuffer[3][1] ), .Y(n63) );
  OAI211XLTS U286 ( .A0(n144), .A1(n494), .B0(n64), .C0(n63), .Y(n1337) );
  INVX2TS U287 ( .A(cacheAddressIn_EAST[0]), .Y(n191) );
  INVX2TS U288 ( .A(n68), .Y(n472) );
  INVX2TS U289 ( .A(cacheAddressIn_WEST[0]), .Y(n358) );
  INVX2TS U290 ( .A(n358), .Y(n771) );
  INVX2TS U291 ( .A(n73), .Y(n480) );
  AOI22X1TS U292 ( .A0(n771), .A1(n57), .B0(n480), .B1(
        \addressToWriteBuffer[1][0] ), .Y(n67) );
  INVX2TS U293 ( .A(n65), .Y(n461) );
  INVX2TS U294 ( .A(n58), .Y(n483) );
  AOI22X1TS U295 ( .A0(n483), .A1(\addressToWriteBuffer[2][0] ), .B0(n59), 
        .B1(\addressToWriteBuffer[3][0] ), .Y(n66) );
  OAI211XLTS U296 ( .A0(n191), .A1(n472), .B0(n67), .C0(n66), .Y(n1338) );
  INVX2TS U297 ( .A(cacheAddressIn_EAST[3]), .Y(n166) );
  INVX2TS U298 ( .A(n68), .Y(n478) );
  INVX2TS U299 ( .A(cacheAddressIn_WEST[3]), .Y(n407) );
  INVX2TS U300 ( .A(n407), .Y(n748) );
  INVX2TS U301 ( .A(n452), .Y(n489) );
  AOI22X1TS U302 ( .A0(n748), .A1(n489), .B0(n460), .B1(
        \addressToWriteBuffer[1][3] ), .Y(n70) );
  INVX2TS U303 ( .A(n65), .Y(n398) );
  INVX2TS U304 ( .A(n453), .Y(n490) );
  AOI22X1TS U305 ( .A0(n398), .A1(\addressToWriteBuffer[2][3] ), .B0(n490), 
        .B1(\addressToWriteBuffer[3][3] ), .Y(n69) );
  OAI211XLTS U306 ( .A0(n166), .A1(n478), .B0(n70), .C0(n69), .Y(n1335) );
  INVX2TS U307 ( .A(dataIn_EAST[3]), .Y(n183) );
  INVX2TS U308 ( .A(dataIn_WEST[3]), .Y(n390) );
  INVX2TS U309 ( .A(n390), .Y(n701) );
  AOI22X1TS U310 ( .A0(n701), .A1(n489), .B0(n460), .B1(
        \dataToWriteBuffer[1][3] ), .Y(n72) );
  AOI22X1TS U311 ( .A0(n461), .A1(\dataToWriteBuffer[2][3] ), .B0(n490), .B1(
        \dataToWriteBuffer[3][3] ), .Y(n71) );
  OAI211XLTS U312 ( .A0(n183), .A1(n486), .B0(n72), .C0(n71), .Y(n1258) );
  INVX2TS U313 ( .A(dataIn_EAST[2]), .Y(n154) );
  INVX2TS U314 ( .A(dataIn_WEST[2]), .Y(n381) );
  INVX2TS U315 ( .A(n381), .Y(n695) );
  AOI22X1TS U316 ( .A0(n695), .A1(n474), .B0(n54), .B1(
        \dataToWriteBuffer[1][2] ), .Y(n75) );
  INVX2TS U317 ( .A(n58), .Y(n465) );
  AOI22X1TS U318 ( .A0(n465), .A1(\dataToWriteBuffer[2][2] ), .B0(n475), .B1(
        \dataToWriteBuffer[3][2] ), .Y(n74) );
  OAI211XLTS U319 ( .A0(n154), .A1(n494), .B0(n75), .C0(n74), .Y(n1259) );
  CLKBUFX2TS U320 ( .A(n197), .Y(n837) );
  AND4X1TS U321 ( .A(n344), .B(n13), .C(n78), .D(n837), .Y(n93) );
  INVX2TS U322 ( .A(n93), .Y(n126) );
  INVX2TS U323 ( .A(dataIn_EAST[1]), .Y(n473) );
  CLKBUFX2TS U324 ( .A(n196), .Y(n538) );
  INVX2TS U325 ( .A(n538), .Y(n780) );
  OAI21XLTS U326 ( .A0(n79), .A1(N742), .B0(n836), .Y(n80) );
  NOR2BX1TS U327 ( .AN(n342), .B(n48), .Y(n82) );
  NOR2XLTS U328 ( .A(n81), .B(n336), .Y(n339) );
  NOR2BX1TS U329 ( .AN(n339), .B(n338), .Y(n84) );
  OR4X2TS U330 ( .A(n780), .B(n83), .C(n82), .D(n84), .Y(n96) );
  INVX2TS U331 ( .A(n96), .Y(n117) );
  INVX2TS U332 ( .A(n85), .Y(n100) );
  AOI22X1TS U333 ( .A0(\dataToWriteBuffer[6][1] ), .A1(n117), .B0(
        dataIn_SOUTH[1]), .B1(n116), .Y(n88) );
  INVX2TS U334 ( .A(n197), .Y(n806) );
  INVX2TS U335 ( .A(n86), .Y(n97) );
  INVX2TS U336 ( .A(n97), .Y(n118) );
  NAND2X1TS U337 ( .A(dataIn_WEST[1]), .B(n118), .Y(n87) );
  OAI211XLTS U338 ( .A0(n126), .A1(n473), .B0(n88), .C0(n87), .Y(n1230) );
  INVX2TS U339 ( .A(n93), .Y(n132) );
  INVX2TS U340 ( .A(n96), .Y(n128) );
  INVX2TS U341 ( .A(n100), .Y(n116) );
  AOI22X1TS U342 ( .A0(\dataToWriteBuffer[6][3] ), .A1(n128), .B0(
        dataIn_SOUTH[3]), .B1(n116), .Y(n90) );
  INVX2TS U343 ( .A(n97), .Y(n129) );
  NAND2X1TS U344 ( .A(dataIn_WEST[3]), .B(n129), .Y(n89) );
  OAI211XLTS U345 ( .A0(n132), .A1(n183), .B0(n90), .C0(n89), .Y(n1228) );
  INVX2TS U346 ( .A(n93), .Y(n115) );
  INVX2TS U347 ( .A(n96), .Y(n112) );
  INVX2TS U348 ( .A(n100), .Y(n127) );
  AOI22X1TS U349 ( .A0(\dataToWriteBuffer[6][2] ), .A1(n112), .B0(
        dataIn_SOUTH[2]), .B1(n127), .Y(n92) );
  NAND2X1TS U350 ( .A(dataIn_WEST[2]), .B(n129), .Y(n91) );
  OAI211XLTS U351 ( .A0(n115), .A1(n154), .B0(n92), .C0(n91), .Y(n1229) );
  INVX2TS U352 ( .A(n93), .Y(n121) );
  INVX2TS U353 ( .A(dataIn_EAST[5]), .Y(n495) );
  AOI22X1TS U354 ( .A0(\dataToWriteBuffer[6][5] ), .A1(n117), .B0(
        dataIn_SOUTH[5]), .B1(n127), .Y(n95) );
  NAND2X1TS U355 ( .A(dataIn_WEST[5]), .B(n118), .Y(n94) );
  OAI211XLTS U356 ( .A0(n121), .A1(n495), .B0(n95), .C0(n94), .Y(n1226) );
  INVX2TS U357 ( .A(dataIn_EAST[4]), .Y(n479) );
  INVX2TS U358 ( .A(n96), .Y(n122) );
  AOI22X1TS U359 ( .A0(\dataToWriteBuffer[6][4] ), .A1(n122), .B0(
        dataIn_SOUTH[4]), .B1(n85), .Y(n99) );
  INVX2TS U360 ( .A(n97), .Y(n123) );
  NAND2X1TS U361 ( .A(dataIn_WEST[4]), .B(n123), .Y(n98) );
  OAI211XLTS U362 ( .A0(n126), .A1(n479), .B0(n99), .C0(n98), .Y(n1227) );
  INVX2TS U363 ( .A(n100), .Y(n107) );
  AOI22X1TS U364 ( .A0(\addressToWriteBuffer[6][3] ), .A1(n128), .B0(
        cacheAddressIn_SOUTH[3]), .B1(n107), .Y(n102) );
  NAND2X1TS U365 ( .A(cacheAddressIn_WEST[3]), .B(n129), .Y(n101) );
  OAI211XLTS U366 ( .A0(n132), .A1(n166), .B0(n102), .C0(n101), .Y(n1295) );
  INVX2TS U367 ( .A(cacheAddressIn_EAST[2]), .Y(n468) );
  AOI22X1TS U368 ( .A0(\addressToWriteBuffer[6][2] ), .A1(n112), .B0(
        cacheAddressIn_SOUTH[2]), .B1(n107), .Y(n104) );
  NAND2X1TS U369 ( .A(cacheAddressIn_WEST[2]), .B(n86), .Y(n103) );
  OAI211XLTS U370 ( .A0(n115), .A1(n468), .B0(n104), .C0(n103), .Y(n1296) );
  AOI22X1TS U371 ( .A0(\addressToWriteBuffer[6][1] ), .A1(n117), .B0(
        cacheAddressIn_SOUTH[1]), .B1(n107), .Y(n106) );
  NAND2X1TS U372 ( .A(cacheAddressIn_WEST[1]), .B(n118), .Y(n105) );
  OAI211XLTS U373 ( .A0(n121), .A1(n144), .B0(n106), .C0(n105), .Y(n1297) );
  AOI22X1TS U374 ( .A0(\addressToWriteBuffer[6][0] ), .A1(n122), .B0(
        cacheAddressIn_SOUTH[0]), .B1(n107), .Y(n109) );
  NAND2X1TS U375 ( .A(cacheAddressIn_WEST[0]), .B(n123), .Y(n108) );
  OAI211XLTS U376 ( .A0(n126), .A1(n191), .B0(n109), .C0(n108), .Y(n1298) );
  INVX2TS U377 ( .A(dataIn_EAST[0]), .Y(n459) );
  AOI22X1TS U378 ( .A0(\dataToWriteBuffer[6][0] ), .A1(n122), .B0(
        dataIn_SOUTH[0]), .B1(n116), .Y(n111) );
  NAND2X1TS U379 ( .A(dataIn_WEST[0]), .B(n123), .Y(n110) );
  OAI211XLTS U380 ( .A0(n132), .A1(n459), .B0(n111), .C0(n110), .Y(n1231) );
  AOI22X1TS U381 ( .A0(\addressToWriteBuffer[6][6] ), .A1(n112), .B0(
        cacheAddressIn_SOUTH[6]), .B1(n85), .Y(n114) );
  NAND2X1TS U382 ( .A(cacheAddressIn_WEST[6]), .B(n86), .Y(n113) );
  OAI211XLTS U383 ( .A0(n115), .A1(n456), .B0(n114), .C0(n113), .Y(n1292) );
  AOI22X1TS U384 ( .A0(\addressToWriteBuffer[6][5] ), .A1(n117), .B0(
        cacheAddressIn_SOUTH[5]), .B1(n116), .Y(n120) );
  NAND2X1TS U385 ( .A(cacheAddressIn_WEST[5]), .B(n118), .Y(n119) );
  OAI211XLTS U386 ( .A0(n121), .A1(n147), .B0(n120), .C0(n119), .Y(n1293) );
  AOI22X1TS U387 ( .A0(\addressToWriteBuffer[6][4] ), .A1(n122), .B0(
        cacheAddressIn_SOUTH[4]), .B1(n127), .Y(n125) );
  NAND2X1TS U388 ( .A(cacheAddressIn_WEST[4]), .B(n123), .Y(n124) );
  OAI211XLTS U389 ( .A0(n126), .A1(n487), .B0(n125), .C0(n124), .Y(n1294) );
  AOI22X1TS U390 ( .A0(\addressToWriteBuffer[6][7] ), .A1(n128), .B0(
        cacheAddressIn_SOUTH[7]), .B1(n127), .Y(n131) );
  NAND2X1TS U391 ( .A(cacheAddressIn_WEST[7]), .B(n129), .Y(n130) );
  OAI211XLTS U392 ( .A0(n132), .A1(n464), .B0(n131), .C0(n130), .Y(n1291) );
  INVX2TS U393 ( .A(n230), .Y(n528) );
  CLKAND2X2TS U394 ( .A(n228), .B(n528), .Y(n148) );
  INVX2TS U395 ( .A(n148), .Y(n182) );
  INVX2TS U396 ( .A(dataIn_WEST[4]), .Y(n395) );
  INVX2TS U397 ( .A(n395), .Y(n707) );
  CLKBUFX2TS U398 ( .A(n252), .Y(n262) );
  CLKBUFX2TS U399 ( .A(n262), .Y(n615) );
  INVX2TS U400 ( .A(n615), .Y(n503) );
  INVX2TS U401 ( .A(n134), .Y(n135) );
  NAND2X1TS U402 ( .A(n503), .B(n136), .Y(n498) );
  CLKBUFX2TS U403 ( .A(n498), .Y(n151) );
  INVX2TS U404 ( .A(n151), .Y(n185) );
  INVX2TS U405 ( .A(n151), .Y(n226) );
  CLKBUFX2TS U406 ( .A(n196), .Y(n671) );
  NAND2X1TS U407 ( .A(n572), .B(n671), .Y(n446) );
  INVX2TS U408 ( .A(n446), .Y(n534) );
  CLKBUFX2TS U409 ( .A(n534), .Y(n530) );
  CLKBUFX2TS U410 ( .A(n530), .Y(n273) );
  CLKBUFX2TS U411 ( .A(n273), .Y(n289) );
  CLKBUFX2TS U412 ( .A(n289), .Y(n234) );
  AOI22X1TS U413 ( .A0(n707), .A1(n226), .B0(\dataToWriteBuffer[1][4] ), .B1(
        n234), .Y(n141) );
  INVX2TS U414 ( .A(n230), .Y(n532) );
  INVX2TS U415 ( .A(n135), .Y(n136) );
  INVX2TS U416 ( .A(n137), .Y(n720) );
  AOI21X1TS U417 ( .A0(n720), .A1(n643), .B0(n572), .Y(n225) );
  NAND2X1TS U418 ( .A(n538), .B(n225), .Y(n681) );
  INVX2TS U419 ( .A(n139), .Y(n159) );
  CLKBUFX2TS U420 ( .A(n681), .Y(n155) );
  INVX2TS U421 ( .A(n155), .Y(n167) );
  AOI22X1TS U422 ( .A0(dataIn_SOUTH[4]), .A1(n170), .B0(n167), .B1(
        cacheDataIn_B[4]), .Y(n140) );
  OAI211XLTS U423 ( .A0(n479), .A1(n182), .B0(n141), .C0(n140), .Y(n1186) );
  INVX2TS U424 ( .A(n148), .Y(n190) );
  INVX2TS U425 ( .A(n151), .Y(n235) );
  CLKBUFX2TS U426 ( .A(n289), .Y(n174) );
  AOI22X1TS U427 ( .A0(n765), .A1(n235), .B0(\addressToWriteBuffer[1][1] ), 
        .B1(n174), .Y(n143) );
  INVX2TS U428 ( .A(n155), .Y(n682) );
  AOI22X1TS U429 ( .A0(cacheAddressIn_SOUTH[1]), .A1(n139), .B0(n682), .B1(
        cacheAddressIn_B[1]), .Y(n142) );
  OAI211XLTS U430 ( .A0(n144), .A1(n190), .B0(n143), .C0(n142), .Y(n1189) );
  INVX2TS U431 ( .A(n148), .Y(n173) );
  CLKBUFX2TS U432 ( .A(n530), .Y(n305) );
  CLKBUFX2TS U433 ( .A(n305), .Y(n238) );
  AOI22X1TS U434 ( .A0(n734), .A1(n242), .B0(\addressToWriteBuffer[1][5] ), 
        .B1(n238), .Y(n146) );
  INVX2TS U435 ( .A(n159), .Y(n176) );
  AOI22X1TS U436 ( .A0(cacheAddressIn_SOUTH[5]), .A1(n176), .B0(n682), .B1(
        cacheAddressIn_B[5]), .Y(n145) );
  OAI211XLTS U437 ( .A0(n147), .A1(n173), .B0(n146), .C0(n145), .Y(n1193) );
  INVX2TS U438 ( .A(n148), .Y(n179) );
  INVX2TS U439 ( .A(cacheAddressIn_WEST[6]), .Y(n372) );
  INVX2TS U440 ( .A(n372), .Y(n729) );
  INVX2TS U441 ( .A(n498), .Y(n158) );
  AOI22X1TS U442 ( .A0(n729), .A1(n158), .B0(\addressToWriteBuffer[1][6] ), 
        .B1(n238), .Y(n150) );
  AOI22X1TS U443 ( .A0(cacheAddressIn_SOUTH[6]), .A1(n176), .B0(n167), .B1(
        cacheAddressIn_B[6]), .Y(n149) );
  OAI211XLTS U444 ( .A0(n456), .A1(n179), .B0(n150), .C0(n149), .Y(n1194) );
  INVX2TS U445 ( .A(n151), .Y(n242) );
  CLKBUFX2TS U446 ( .A(n305), .Y(n184) );
  AOI22X1TS U447 ( .A0(n695), .A1(n242), .B0(\dataToWriteBuffer[1][2] ), .B1(
        n184), .Y(n153) );
  INVX2TS U448 ( .A(n159), .Y(n170) );
  INVX2TS U449 ( .A(n155), .Y(n186) );
  AOI22X1TS U450 ( .A0(dataIn_SOUTH[2]), .A1(n170), .B0(n186), .B1(
        cacheDataIn_B[2]), .Y(n152) );
  OAI211XLTS U451 ( .A0(n154), .A1(n182), .B0(n153), .C0(n152), .Y(n1184) );
  INVX2TS U452 ( .A(dataIn_WEST[1]), .Y(n423) );
  INVX2TS U453 ( .A(n423), .Y(n690) );
  AOI22X1TS U454 ( .A0(n690), .A1(n158), .B0(\dataToWriteBuffer[1][1] ), .B1(
        n234), .Y(n157) );
  INVX2TS U455 ( .A(n155), .Y(n175) );
  AOI22X1TS U456 ( .A0(dataIn_SOUTH[1]), .A1(n139), .B0(n175), .B1(
        cacheDataIn_B[1]), .Y(n156) );
  OAI211XLTS U457 ( .A0(n473), .A1(n190), .B0(n157), .C0(n156), .Y(n1183) );
  INVX2TS U458 ( .A(dataIn_WEST[0]), .Y(n431) );
  INVX2TS U459 ( .A(n431), .Y(n686) );
  CLKBUFX2TS U460 ( .A(n305), .Y(n589) );
  AOI22X1TS U461 ( .A0(n686), .A1(n158), .B0(\dataToWriteBuffer[1][0] ), .B1(
        n589), .Y(n161) );
  INVX2TS U462 ( .A(n159), .Y(n187) );
  AOI22X1TS U463 ( .A0(dataIn_SOUTH[0]), .A1(n187), .B0(n167), .B1(
        cacheDataIn_B[0]), .Y(n160) );
  OAI211XLTS U464 ( .A0(n459), .A1(n173), .B0(n161), .C0(n160), .Y(n1182) );
  INVX2TS U465 ( .A(cacheAddressIn_WEST[4]), .Y(n366) );
  INVX2TS U466 ( .A(n366), .Y(n740) );
  AOI22X1TS U467 ( .A0(n740), .A1(n235), .B0(\addressToWriteBuffer[1][4] ), 
        .B1(n174), .Y(n163) );
  AOI22X1TS U468 ( .A0(cacheAddressIn_SOUTH[4]), .A1(n176), .B0(n186), .B1(
        cacheAddressIn_B[4]), .Y(n162) );
  OAI211XLTS U469 ( .A0(n487), .A1(n179), .B0(n163), .C0(n162), .Y(n1192) );
  AOI22X1TS U470 ( .A0(n748), .A1(n185), .B0(\addressToWriteBuffer[1][3] ), 
        .B1(n238), .Y(n165) );
  AOI22X1TS U471 ( .A0(cacheAddressIn_SOUTH[3]), .A1(n187), .B0(n175), .B1(
        cacheAddressIn_B[3]), .Y(n164) );
  OAI211XLTS U472 ( .A0(n166), .A1(n182), .B0(n165), .C0(n164), .Y(n1191) );
  INVX2TS U473 ( .A(cacheAddressIn_WEST[2]), .Y(n414) );
  INVX2TS U474 ( .A(n414), .Y(n756) );
  AOI22X1TS U475 ( .A0(n756), .A1(n226), .B0(\addressToWriteBuffer[1][2] ), 
        .B1(n184), .Y(n169) );
  AOI22X1TS U476 ( .A0(cacheAddressIn_SOUTH[2]), .A1(n170), .B0(n167), .B1(
        cacheAddressIn_B[2]), .Y(n168) );
  OAI211XLTS U477 ( .A0(n468), .A1(n190), .B0(n169), .C0(n168), .Y(n1190) );
  INVX2TS U478 ( .A(dataIn_WEST[5]), .Y(n385) );
  INVX2TS U479 ( .A(n385), .Y(n712) );
  AOI22X1TS U480 ( .A0(n712), .A1(n242), .B0(\dataToWriteBuffer[1][5] ), .B1(
        n174), .Y(n172) );
  AOI22X1TS U481 ( .A0(dataIn_SOUTH[5]), .A1(n170), .B0(n175), .B1(
        cacheDataIn_B[5]), .Y(n171) );
  OAI211XLTS U482 ( .A0(n495), .A1(n173), .B0(n172), .C0(n171), .Y(n1187) );
  INVX2TS U483 ( .A(cacheAddressIn_WEST[7]), .Y(n362) );
  INVX2TS U484 ( .A(n362), .Y(n723) );
  AOI22X1TS U485 ( .A0(n723), .A1(n235), .B0(\addressToWriteBuffer[1][7] ), 
        .B1(n174), .Y(n178) );
  AOI22X1TS U486 ( .A0(cacheAddressIn_SOUTH[7]), .A1(n176), .B0(n175), .B1(
        cacheAddressIn_B[7]), .Y(n177) );
  OAI211XLTS U487 ( .A0(n464), .A1(n179), .B0(n178), .C0(n177), .Y(n1195) );
  AOI22X1TS U488 ( .A0(n701), .A1(n185), .B0(\dataToWriteBuffer[1][3] ), .B1(
        n184), .Y(n181) );
  AOI22X1TS U489 ( .A0(dataIn_SOUTH[3]), .A1(n187), .B0(n682), .B1(
        cacheDataIn_B[3]), .Y(n180) );
  OAI211XLTS U490 ( .A0(n183), .A1(n182), .B0(n181), .C0(n180), .Y(n1185) );
  AOI22X1TS U491 ( .A0(n771), .A1(n185), .B0(\addressToWriteBuffer[1][0] ), 
        .B1(n184), .Y(n189) );
  AOI22X1TS U492 ( .A0(cacheAddressIn_SOUTH[0]), .A1(n187), .B0(n186), .B1(
        cacheAddressIn_B[0]), .Y(n188) );
  OAI211XLTS U493 ( .A0(n191), .A1(n190), .B0(n189), .C0(n188), .Y(n1188) );
  INVX2TS U494 ( .A(n20), .Y(n195) );
  INVX2TS U495 ( .A(n5), .Y(n194) );
  INVX2TS U496 ( .A(n18), .Y(n192) );
  INVX2TS U497 ( .A(n193), .Y(n206) );
  INVX2TS U498 ( .A(n206), .Y(n198) );
  OR3X1TS U499 ( .A(n195), .B(n194), .C(n198), .Y(n207) );
  INVX2TS U500 ( .A(n207), .Y(n506) );
  CLKBUFX2TS U501 ( .A(n196), .Y(n617) );
  NAND2X1TS U502 ( .A(n506), .B(n617), .Y(n205) );
  INVX2TS U503 ( .A(n8), .Y(n803) );
  NOR2BX1TS U504 ( .AN(n198), .B(n513), .Y(n203) );
  INVX2TS U505 ( .A(n197), .Y(n778) );
  INVX2TS U506 ( .A(n207), .Y(n510) );
  NOR3XLTS U507 ( .A(n778), .B(n198), .C(n510), .Y(n202) );
  AOI22X1TS U508 ( .A0(n803), .A1(n203), .B0(n202), .B1(
        requesterAddressOut_NORTH[3]), .Y(n199) );
  OAI21XLTS U509 ( .A0(n828), .A1(n205), .B0(n199), .Y(n1159) );
  INVX2TS U510 ( .A(n9), .Y(n809) );
  AOI22X1TS U511 ( .A0(n809), .A1(n203), .B0(n202), .B1(
        requesterAddressOut_NORTH[2]), .Y(n200) );
  OAI21XLTS U512 ( .A0(n829), .A1(n205), .B0(n200), .Y(n1158) );
  INVX2TS U513 ( .A(n10), .Y(n812) );
  AOI22X1TS U514 ( .A0(n812), .A1(n203), .B0(n202), .B1(
        requesterAddressOut_NORTH[1]), .Y(n201) );
  OAI21XLTS U515 ( .A0(n830), .A1(n205), .B0(n201), .Y(n1157) );
  INVX2TS U516 ( .A(n11), .Y(n817) );
  AOI22X1TS U517 ( .A0(n817), .A1(n203), .B0(n202), .B1(
        requesterAddressOut_NORTH[0]), .Y(n204) );
  OAI21XLTS U518 ( .A0(n831), .A1(n205), .B0(n204), .Y(n1156) );
  INVX2TS U519 ( .A(n206), .Y(n508) );
  INVX2TS U520 ( .A(n207), .Y(n504) );
  AO22X2TS U521 ( .A0(n508), .A1(n209), .B0(n504), .B1(n208), .Y(N5373) );
  AO22X2TS U522 ( .A0(n193), .A1(n211), .B0(n506), .B1(n210), .Y(N5374) );
  AO22X2TS U523 ( .A0(n193), .A1(n213), .B0(n510), .B1(n212), .Y(N5375) );
  AO22X2TS U524 ( .A0(n508), .A1(n215), .B0(n504), .B1(n214), .Y(N5376) );
  NAND3XLTS U525 ( .A(n52), .B(n836), .C(N741), .Y(n218) );
  INVX2TS U526 ( .A(n218), .Y(n580) );
  CLKBUFX2TS U527 ( .A(n289), .Y(n332) );
  NAND2X1TS U528 ( .A(n580), .B(n332), .Y(n220) );
  OAI211XLTS U529 ( .A0(n438), .A1(n218), .B0(n217), .C0(n837), .Y(n630) );
  INVX2TS U530 ( .A(n630), .Y(n628) );
  NAND2X1TS U531 ( .A(n628), .B(\requesterPortBuffer[5][1] ), .Y(n219) );
  OAI211XLTS U532 ( .A0(n521), .A1(n220), .B0(n219), .C0(n622), .Y(n1272) );
  NAND2X1TS U533 ( .A(n538), .B(n346), .Y(n224) );
  INVX2TS U534 ( .A(n224), .Y(n282) );
  CLKBUFX2TS U535 ( .A(n282), .Y(n563) );
  CLKBUFX2TS U536 ( .A(n563), .Y(n555) );
  CLKBUFX2TS U537 ( .A(n555), .Y(n527) );
  NAND2X1TS U538 ( .A(n527), .B(\requesterPortBuffer[5][1] ), .Y(n221) );
  CLKBUFX2TS U539 ( .A(n534), .Y(n554) );
  CLKBUFX2TS U540 ( .A(n554), .Y(n602) );
  AOI22X1TS U541 ( .A0(n532), .A1(isWrite[0]), .B0(n602), .B1(isWrite[2]), .Y(
        n222) );
  AOI22X1TS U542 ( .A0(n532), .A1(\requesterPortBuffer[3][1] ), .B0(n589), 
        .B1(\requesterPortBuffer[5][1] ), .Y(n223) );
  NOR2XLTS U543 ( .A(n778), .B(n225), .Y(n246) );
  INVX2TS U544 ( .A(n246), .Y(n497) );
  INVX2TS U545 ( .A(n497), .Y(n233) );
  AOI22X1TS U546 ( .A0(requesterAddressIn_WEST[3]), .A1(n226), .B0(
        \requesterAddressBuffer[1][3] ), .B1(n234), .Y(n232) );
  INVX2TS U547 ( .A(n229), .Y(n239) );
  INVX2TS U548 ( .A(n230), .Y(n319) );
  NAND2X1TS U549 ( .A(n319), .B(n643), .Y(n500) );
  OAI221XLTS U550 ( .A0(n43), .A1(requesterAddressIn_SOUTH[3]), .B0(n229), 
        .B1(requesterAddressIn_EAST[3]), .C0(n243), .Y(n231) );
  OAI211XLTS U551 ( .A0(n233), .A1(n828), .B0(n232), .C0(n231), .Y(n1359) );
  AOI22X1TS U552 ( .A0(requesterAddressIn_WEST[2]), .A1(n235), .B0(
        \requesterAddressBuffer[1][2] ), .B1(n234), .Y(n237) );
  OAI221XLTS U553 ( .A0(n239), .A1(requesterAddressIn_SOUTH[2]), .B0(n227), 
        .B1(requesterAddressIn_EAST[2]), .C0(n243), .Y(n236) );
  OAI211XLTS U554 ( .A0(n246), .A1(n829), .B0(n237), .C0(n236), .Y(n1360) );
  AOI22X1TS U555 ( .A0(requesterAddressIn_WEST[0]), .A1(n226), .B0(
        \requesterAddressBuffer[1][0] ), .B1(n238), .Y(n241) );
  OAI221XLTS U556 ( .A0(n43), .A1(requesterAddressIn_SOUTH[0]), .B0(n227), 
        .B1(requesterAddressIn_EAST[0]), .C0(n243), .Y(n240) );
  OAI211XLTS U557 ( .A0(n246), .A1(n831), .B0(n241), .C0(n240), .Y(n1362) );
  AOI22X1TS U558 ( .A0(requesterAddressIn_WEST[1]), .A1(n242), .B0(
        \requesterAddressBuffer[1][1] ), .B1(n589), .Y(n245) );
  OAI221XLTS U559 ( .A0(n239), .A1(requesterAddressIn_SOUTH[1]), .B0(n227), 
        .B1(requesterAddressIn_EAST[1]), .C0(n243), .Y(n244) );
  OAI211XLTS U560 ( .A0(n246), .A1(n830), .B0(n245), .C0(n244), .Y(n1361) );
  CLKBUFX2TS U561 ( .A(n332), .Y(n250) );
  CLKBUFX2TS U562 ( .A(n282), .Y(n260) );
  INVX2TS U563 ( .A(n262), .Y(n259) );
  AOI222XLTS U564 ( .A0(\addressToWriteBuffer[6][5] ), .A1(n250), .B0(
        \addressToWriteBuffer[5][5] ), .B1(n260), .C0(n259), .C1(
        \addressToWriteBuffer[4][5] ), .Y(n247) );
  INVX2TS U565 ( .A(n247), .Y(n1309) );
  INVX2TS U566 ( .A(n262), .Y(n256) );
  AOI222XLTS U567 ( .A0(\addressToWriteBuffer[6][3] ), .A1(n250), .B0(
        \addressToWriteBuffer[5][3] ), .B1(n260), .C0(n256), .C1(
        \addressToWriteBuffer[4][3] ), .Y(n248) );
  INVX2TS U568 ( .A(n248), .Y(n1311) );
  CLKBUFX2TS U569 ( .A(n282), .Y(n263) );
  CLKBUFX2TS U570 ( .A(n263), .Y(n309) );
  CLKBUFX2TS U571 ( .A(n309), .Y(n301) );
  AOI222XLTS U572 ( .A0(\addressToWriteBuffer[6][4] ), .A1(n250), .B0(
        \addressToWriteBuffer[5][4] ), .B1(n301), .C0(n256), .C1(
        \addressToWriteBuffer[4][4] ), .Y(n249) );
  INVX2TS U573 ( .A(n249), .Y(n1310) );
  AOI222XLTS U574 ( .A0(\addressToWriteBuffer[6][2] ), .A1(n250), .B0(
        \addressToWriteBuffer[5][2] ), .B1(n260), .C0(n256), .C1(
        \addressToWriteBuffer[4][2] ), .Y(n251) );
  INVX2TS U575 ( .A(n251), .Y(n1312) );
  CLKBUFX2TS U576 ( .A(n530), .Y(n280) );
  CLKBUFX2TS U577 ( .A(n263), .Y(n271) );
  AOI222XLTS U578 ( .A0(\dataToWriteBuffer[6][0] ), .A1(n280), .B0(
        \dataToWriteBuffer[5][0] ), .B1(n271), .C0(n270), .C1(
        \dataToWriteBuffer[4][0] ), .Y(n253) );
  INVX2TS U579 ( .A(n253), .Y(n1243) );
  CLKBUFX2TS U580 ( .A(n263), .Y(n274) );
  AOI222XLTS U581 ( .A0(\dataToWriteBuffer[6][2] ), .A1(n280), .B0(
        \dataToWriteBuffer[5][2] ), .B1(n274), .C0(n270), .C1(
        \dataToWriteBuffer[4][2] ), .Y(n254) );
  INVX2TS U582 ( .A(n254), .Y(n1241) );
  CLKBUFX2TS U583 ( .A(n273), .Y(n299) );
  AOI222XLTS U584 ( .A0(\dataToWriteBuffer[6][3] ), .A1(n299), .B0(
        \dataToWriteBuffer[5][3] ), .B1(n271), .C0(n259), .C1(
        \dataToWriteBuffer[4][3] ), .Y(n255) );
  INVX2TS U585 ( .A(n255), .Y(n1240) );
  CLKBUFX2TS U586 ( .A(n273), .Y(n277) );
  AOI222XLTS U587 ( .A0(\addressToWriteBuffer[6][0] ), .A1(n277), .B0(
        \addressToWriteBuffer[5][0] ), .B1(n274), .C0(n256), .C1(
        \addressToWriteBuffer[4][0] ), .Y(n257) );
  INVX2TS U588 ( .A(n257), .Y(n1314) );
  AOI222XLTS U589 ( .A0(\dataToWriteBuffer[6][1] ), .A1(n280), .B0(
        \dataToWriteBuffer[5][1] ), .B1(n271), .C0(n259), .C1(
        \dataToWriteBuffer[4][1] ), .Y(n258) );
  INVX2TS U590 ( .A(n258), .Y(n1242) );
  AOI222XLTS U591 ( .A0(\addressToWriteBuffer[6][1] ), .A1(n277), .B0(
        \addressToWriteBuffer[5][1] ), .B1(n260), .C0(n259), .C1(
        \addressToWriteBuffer[4][1] ), .Y(n261) );
  INVX2TS U592 ( .A(n261), .Y(n1313) );
  CLKBUFX2TS U593 ( .A(n262), .Y(n437) );
  INVX2TS U594 ( .A(n437), .Y(n302) );
  CLKBUFX2TS U595 ( .A(n263), .Y(n268) );
  AOI222XLTS U596 ( .A0(\addressToWriteBuffer[5][6] ), .A1(n299), .B0(n302), 
        .B1(\addressToWriteBuffer[3][6] ), .C0(n268), .C1(
        \addressToWriteBuffer[4][6] ), .Y(n264) );
  INVX2TS U597 ( .A(n264), .Y(n1316) );
  CLKBUFX2TS U598 ( .A(n554), .Y(n447) );
  CLKBUFX2TS U599 ( .A(n447), .Y(n287) );
  INVX2TS U600 ( .A(n437), .Y(n291) );
  AOI222XLTS U601 ( .A0(\addressToWriteBuffer[5][1] ), .A1(n287), .B0(n291), 
        .B1(\addressToWriteBuffer[3][1] ), .C0(n268), .C1(
        \addressToWriteBuffer[4][1] ), .Y(n265) );
  INVX2TS U602 ( .A(n265), .Y(n1321) );
  AOI222XLTS U603 ( .A0(\addressToWriteBuffer[5][0] ), .A1(n287), .B0(n291), 
        .B1(\addressToWriteBuffer[3][0] ), .C0(n268), .C1(
        \addressToWriteBuffer[4][0] ), .Y(n266) );
  INVX2TS U604 ( .A(n266), .Y(n1322) );
  CLKBUFX2TS U605 ( .A(n447), .Y(n303) );
  AOI222XLTS U606 ( .A0(\dataToWriteBuffer[6][5] ), .A1(n303), .B0(
        \dataToWriteBuffer[5][5] ), .B1(n274), .C0(n270), .C1(
        \dataToWriteBuffer[4][5] ), .Y(n267) );
  INVX2TS U607 ( .A(n267), .Y(n1238) );
  INVX2TS U608 ( .A(n437), .Y(n297) );
  AOI222XLTS U609 ( .A0(\addressToWriteBuffer[5][2] ), .A1(n303), .B0(n297), 
        .B1(\addressToWriteBuffer[3][2] ), .C0(n268), .C1(
        \addressToWriteBuffer[4][2] ), .Y(n269) );
  INVX2TS U610 ( .A(n269), .Y(n1320) );
  AOI222XLTS U611 ( .A0(\dataToWriteBuffer[6][4] ), .A1(n303), .B0(
        \dataToWriteBuffer[5][4] ), .B1(n271), .C0(n270), .C1(
        \dataToWriteBuffer[4][4] ), .Y(n272) );
  INVX2TS U612 ( .A(n272), .Y(n1239) );
  CLKBUFX2TS U613 ( .A(n273), .Y(n314) );
  AOI222XLTS U614 ( .A0(\addressToWriteBuffer[6][6] ), .A1(n314), .B0(
        \addressToWriteBuffer[5][6] ), .B1(n274), .C0(n297), .C1(
        \addressToWriteBuffer[4][6] ), .Y(n275) );
  INVX2TS U615 ( .A(n275), .Y(n1308) );
  INVX2TS U616 ( .A(n615), .Y(n294) );
  CLKBUFX2TS U617 ( .A(n563), .Y(n559) );
  CLKBUFX2TS U618 ( .A(n559), .Y(n331) );
  AOI222XLTS U619 ( .A0(\dataToWriteBuffer[5][0] ), .A1(n277), .B0(n294), .B1(
        \dataToWriteBuffer[3][0] ), .C0(n331), .C1(\dataToWriteBuffer[4][0] ), 
        .Y(n276) );
  INVX2TS U620 ( .A(n276), .Y(n1249) );
  AOI222XLTS U621 ( .A0(\addressToWriteBuffer[5][7] ), .A1(n277), .B0(n302), 
        .B1(\addressToWriteBuffer[3][7] ), .C0(n331), .C1(
        \addressToWriteBuffer[4][7] ), .Y(n278) );
  INVX2TS U622 ( .A(n278), .Y(n1315) );
  AOI222XLTS U623 ( .A0(\addressToWriteBuffer[5][4] ), .A1(n299), .B0(n297), 
        .B1(\addressToWriteBuffer[3][4] ), .C0(n331), .C1(
        \addressToWriteBuffer[4][4] ), .Y(n279) );
  INVX2TS U624 ( .A(n279), .Y(n1318) );
  CLKBUFX2TS U625 ( .A(n559), .Y(n531) );
  AOI222XLTS U626 ( .A0(\dataToWriteBuffer[5][5] ), .A1(n280), .B0(n291), .B1(
        \dataToWriteBuffer[3][5] ), .C0(n531), .C1(\dataToWriteBuffer[4][5] ), 
        .Y(n281) );
  INVX2TS U627 ( .A(n281), .Y(n1244) );
  INVX2TS U628 ( .A(n307), .Y(n329) );
  CLKBUFX2TS U629 ( .A(n447), .Y(n325) );
  CLKBUFX2TS U630 ( .A(n282), .Y(n286) );
  AOI222XLTS U631 ( .A0(n329), .A1(\dataToWriteBuffer[0][4] ), .B0(
        \dataToWriteBuffer[2][4] ), .B1(n325), .C0(\dataToWriteBuffer[1][4] ), 
        .C1(n286), .Y(n283) );
  INVX2TS U632 ( .A(n283), .Y(n1263) );
  INVX2TS U633 ( .A(n307), .Y(n315) );
  AOI222XLTS U634 ( .A0(n315), .A1(\dataToWriteBuffer[0][3] ), .B0(
        \dataToWriteBuffer[2][3] ), .B1(n325), .C0(\dataToWriteBuffer[1][3] ), 
        .C1(n286), .Y(n284) );
  INVX2TS U635 ( .A(n284), .Y(n1264) );
  AOI222XLTS U636 ( .A0(n315), .A1(\dataToWriteBuffer[0][0] ), .B0(
        \dataToWriteBuffer[2][0] ), .B1(n287), .C0(\dataToWriteBuffer[1][0] ), 
        .C1(n286), .Y(n285) );
  INVX2TS U637 ( .A(n285), .Y(n1267) );
  AOI222XLTS U638 ( .A0(n503), .A1(\dataToWriteBuffer[0][1] ), .B0(
        \dataToWriteBuffer[2][1] ), .B1(n287), .C0(\dataToWriteBuffer[1][1] ), 
        .C1(n286), .Y(n288) );
  INVX2TS U639 ( .A(n288), .Y(n1266) );
  CLKBUFX2TS U640 ( .A(n289), .Y(n295) );
  AOI222XLTS U641 ( .A0(\dataToWriteBuffer[5][3] ), .A1(n295), .B0(n294), .B1(
        \dataToWriteBuffer[3][3] ), .C0(n531), .C1(\dataToWriteBuffer[4][3] ), 
        .Y(n290) );
  INVX2TS U642 ( .A(n290), .Y(n1246) );
  CLKBUFX2TS U643 ( .A(n559), .Y(n502) );
  AOI222XLTS U644 ( .A0(\dataToWriteBuffer[5][2] ), .A1(n295), .B0(n291), .B1(
        \dataToWriteBuffer[3][2] ), .C0(n502), .C1(\dataToWriteBuffer[4][2] ), 
        .Y(n292) );
  INVX2TS U645 ( .A(n292), .Y(n1247) );
  AOI222XLTS U646 ( .A0(\dataToWriteBuffer[5][4] ), .A1(n295), .B0(n294), .B1(
        \dataToWriteBuffer[3][4] ), .C0(n502), .C1(\dataToWriteBuffer[4][4] ), 
        .Y(n293) );
  INVX2TS U647 ( .A(n293), .Y(n1245) );
  AOI222XLTS U648 ( .A0(\dataToWriteBuffer[5][1] ), .A1(n295), .B0(n294), .B1(
        \dataToWriteBuffer[3][1] ), .C0(n502), .C1(\dataToWriteBuffer[4][1] ), 
        .Y(n296) );
  INVX2TS U649 ( .A(n296), .Y(n1248) );
  AOI222XLTS U650 ( .A0(\addressToWriteBuffer[6][7] ), .A1(n314), .B0(
        \addressToWriteBuffer[5][7] ), .B1(n301), .C0(n297), .C1(
        \addressToWriteBuffer[4][7] ), .Y(n298) );
  INVX2TS U651 ( .A(n298), .Y(n1307) );
  AOI222XLTS U652 ( .A0(\addressToWriteBuffer[5][5] ), .A1(n299), .B0(n302), 
        .B1(\addressToWriteBuffer[3][5] ), .C0(n301), .C1(
        \addressToWriteBuffer[4][5] ), .Y(n300) );
  INVX2TS U653 ( .A(n300), .Y(n1317) );
  AOI222XLTS U654 ( .A0(\addressToWriteBuffer[5][3] ), .A1(n303), .B0(n302), 
        .B1(\addressToWriteBuffer[3][3] ), .C0(n301), .C1(
        \addressToWriteBuffer[4][3] ), .Y(n304) );
  INVX2TS U655 ( .A(n304), .Y(n1319) );
  CLKBUFX2TS U656 ( .A(n305), .Y(n526) );
  CLKBUFX2TS U657 ( .A(n526), .Y(n322) );
  CLKBUFX2TS U658 ( .A(n309), .Y(n321) );
  AOI222XLTS U659 ( .A0(n319), .A1(\addressToWriteBuffer[0][0] ), .B0(
        \addressToWriteBuffer[2][0] ), .B1(n322), .C0(
        \addressToWriteBuffer[1][0] ), .C1(n321), .Y(n306) );
  INVX2TS U660 ( .A(n306), .Y(n1346) );
  INVX2TS U661 ( .A(n307), .Y(n323) );
  CLKBUFX2TS U662 ( .A(n526), .Y(n328) );
  CLKBUFX2TS U663 ( .A(n309), .Y(n317) );
  AOI222XLTS U664 ( .A0(n323), .A1(\addressToWriteBuffer[0][6] ), .B0(
        \addressToWriteBuffer[2][6] ), .B1(n328), .C0(
        \addressToWriteBuffer[1][6] ), .C1(n317), .Y(n308) );
  INVX2TS U665 ( .A(n308), .Y(n1340) );
  CLKBUFX2TS U666 ( .A(n309), .Y(n327) );
  AOI222XLTS U667 ( .A0(n315), .A1(\dataToWriteBuffer[0][5] ), .B0(
        \dataToWriteBuffer[2][5] ), .B1(n325), .C0(\dataToWriteBuffer[1][5] ), 
        .C1(n327), .Y(n310) );
  INVX2TS U668 ( .A(n310), .Y(n1262) );
  AOI222XLTS U669 ( .A0(n319), .A1(\requesterPortBuffer[0][0] ), .B0(n314), 
        .B1(\requesterPortBuffer[2][0] ), .C0(\requesterPortBuffer[1][0] ), 
        .C1(n321), .Y(n311) );
  INVX2TS U670 ( .A(n311), .Y(n1363) );
  AOI222XLTS U671 ( .A0(n323), .A1(\addressToWriteBuffer[0][4] ), .B0(
        \addressToWriteBuffer[2][4] ), .B1(n328), .C0(
        \addressToWriteBuffer[1][4] ), .C1(n317), .Y(n312) );
  INVX2TS U672 ( .A(n312), .Y(n1342) );
  AOI222XLTS U673 ( .A0(n329), .A1(\addressToWriteBuffer[0][2] ), .B0(
        \addressToWriteBuffer[2][2] ), .B1(n322), .C0(
        \addressToWriteBuffer[1][2] ), .C1(n317), .Y(n313) );
  INVX2TS U674 ( .A(n313), .Y(n1344) );
  AOI222XLTS U675 ( .A0(n315), .A1(\requesterPortBuffer[0][1] ), .B0(n314), 
        .B1(\requesterPortBuffer[2][1] ), .C0(\requesterPortBuffer[1][1] ), 
        .C1(n327), .Y(n316) );
  INVX2TS U676 ( .A(n316), .Y(n1282) );
  AOI222XLTS U677 ( .A0(n323), .A1(\addressToWriteBuffer[0][5] ), .B0(
        \addressToWriteBuffer[2][5] ), .B1(n328), .C0(
        \addressToWriteBuffer[1][5] ), .C1(n317), .Y(n318) );
  INVX2TS U678 ( .A(n318), .Y(n1341) );
  AOI222XLTS U679 ( .A0(n319), .A1(\addressToWriteBuffer[0][1] ), .B0(
        \addressToWriteBuffer[2][1] ), .B1(n322), .C0(
        \addressToWriteBuffer[1][1] ), .C1(n321), .Y(n320) );
  INVX2TS U680 ( .A(n320), .Y(n1345) );
  AOI222XLTS U681 ( .A0(n323), .A1(\addressToWriteBuffer[0][3] ), .B0(
        \addressToWriteBuffer[2][3] ), .B1(n322), .C0(
        \addressToWriteBuffer[1][3] ), .C1(n321), .Y(n324) );
  INVX2TS U682 ( .A(n324), .Y(n1343) );
  AOI222XLTS U683 ( .A0(n329), .A1(\dataToWriteBuffer[0][2] ), .B0(
        \dataToWriteBuffer[2][2] ), .B1(n325), .C0(\dataToWriteBuffer[1][2] ), 
        .C1(n327), .Y(n326) );
  INVX2TS U684 ( .A(n326), .Y(n1265) );
  AOI222XLTS U685 ( .A0(n329), .A1(\addressToWriteBuffer[0][7] ), .B0(
        \addressToWriteBuffer[2][7] ), .B1(n328), .C0(
        \addressToWriteBuffer[1][7] ), .C1(n327), .Y(n330) );
  INVX2TS U686 ( .A(n330), .Y(n1339) );
  AOI222XLTS U687 ( .A0(n503), .A1(\requesterPortBuffer[3][0] ), .B0(n332), 
        .B1(\requesterPortBuffer[5][0] ), .C0(n331), .C1(
        \requesterPortBuffer[4][0] ), .Y(n333) );
  INVX2TS U688 ( .A(n333), .Y(n1277) );
  INVX2TS U689 ( .A(n19), .Y(n640) );
  OAI22X1TS U690 ( .A0(n32), .A1(n334), .B0(n515), .B1(n640), .Y(n439) );
  INVX2TS U691 ( .A(n439), .Y(n337) );
  NOR2XLTS U692 ( .A(n337), .B(n42), .Y(n638) );
  AOI21X1TS U693 ( .A0(n40), .A1(n438), .B0(n451), .Y(n646) );
  INVX2TS U694 ( .A(n646), .Y(n335) );
  AOI211XLTS U695 ( .A0(n337), .A1(n336), .B0(n638), .C0(n335), .Y(n1211) );
  INVX2TS U696 ( .A(n340), .Y(n341) );
  NAND3X1TS U697 ( .A(n343), .B(n342), .C(n341), .Y(n351) );
  NAND2X1TS U698 ( .A(n345), .B(n344), .Y(n353) );
  AOI211XLTS U699 ( .A0(n580), .A1(n512), .B0(n346), .C0(n778), .Y(n347) );
  INVX2TS U700 ( .A(n348), .Y(n374) );
  INVX2TS U701 ( .A(n374), .Y(n410) );
  NAND2BX1TS U702 ( .AN(n410), .B(n518), .Y(n349) );
  OR4X2TS U703 ( .A(n537), .B(n355), .C(n350), .D(n349), .Y(n368) );
  INVX2TS U704 ( .A(n368), .Y(n426) );
  NAND2BX1TS U705 ( .AN(n351), .B(n518), .Y(n352) );
  INVX2TS U706 ( .A(n352), .Y(n369) );
  INVX2TS U707 ( .A(n369), .Y(n424) );
  INVX2TS U708 ( .A(n374), .Y(n419) );
  INVX2TS U709 ( .A(n354), .Y(n397) );
  INVX2TS U710 ( .A(n397), .Y(n418) );
  AOI22X1TS U711 ( .A0(n419), .A1(\addressToWriteBuffer[5][0] ), .B0(
        cacheAddressIn_EAST[0]), .B1(n418), .Y(n357) );
  INVX2TS U712 ( .A(n17), .Y(n387) );
  AOI22X1TS U713 ( .A0(n469), .A1(\addressToWriteBuffer[6][0] ), .B0(
        cacheAddressIn_SOUTH[0]), .B1(n387), .Y(n356) );
  OAI211XLTS U714 ( .A0(n358), .A1(n424), .B0(n357), .C0(n356), .Y(n359) );
  INVX2TS U715 ( .A(n368), .Y(n434) );
  INVX2TS U716 ( .A(n369), .Y(n432) );
  INVX2TS U717 ( .A(n374), .Y(n403) );
  AOI22X1TS U718 ( .A0(n403), .A1(\addressToWriteBuffer[5][7] ), .B0(n354), 
        .B1(cacheAddressIn_EAST[7]), .Y(n361) );
  AOI22X1TS U719 ( .A0(n465), .A1(\addressToWriteBuffer[6][7] ), .B0(n387), 
        .B1(cacheAddressIn_SOUTH[7]), .Y(n360) );
  OAI211XLTS U720 ( .A0(n432), .A1(n362), .B0(n361), .C0(n360), .Y(n363) );
  INVX2TS U721 ( .A(n368), .Y(n409) );
  AOI22X1TS U722 ( .A0(n403), .A1(\addressToWriteBuffer[5][4] ), .B0(n354), 
        .B1(cacheAddressIn_EAST[4]), .Y(n365) );
  AOI22X1TS U723 ( .A0(n491), .A1(\addressToWriteBuffer[6][4] ), .B0(n387), 
        .B1(cacheAddressIn_SOUTH[4]), .Y(n364) );
  OAI211XLTS U724 ( .A0(n415), .A1(n366), .B0(n365), .C0(n364), .Y(n367) );
  INVX2TS U725 ( .A(n368), .Y(n417) );
  INVX2TS U726 ( .A(n369), .Y(n415) );
  AOI22X1TS U727 ( .A0(n419), .A1(\addressToWriteBuffer[5][6] ), .B0(n418), 
        .B1(cacheAddressIn_EAST[6]), .Y(n371) );
  INVX2TS U728 ( .A(n65), .Y(n404) );
  INVX2TS U729 ( .A(n17), .Y(n420) );
  AOI22X1TS U730 ( .A0(n404), .A1(\addressToWriteBuffer[6][6] ), .B0(n420), 
        .B1(cacheAddressIn_SOUTH[6]), .Y(n370) );
  OAI211XLTS U731 ( .A0(n415), .A1(n372), .B0(n371), .C0(n370), .Y(n373) );
  INVX2TS U732 ( .A(n397), .Y(n392) );
  AOI22X1TS U733 ( .A0(n348), .A1(\addressToWriteBuffer[5][5] ), .B0(n392), 
        .B1(cacheAddressIn_EAST[5]), .Y(n376) );
  INVX2TS U734 ( .A(n58), .Y(n491) );
  INVX2TS U735 ( .A(n17), .Y(n428) );
  AOI22X1TS U736 ( .A0(n491), .A1(\addressToWriteBuffer[6][5] ), .B0(n428), 
        .B1(cacheAddressIn_SOUTH[5]), .Y(n375) );
  OAI211XLTS U737 ( .A0(n424), .A1(n377), .B0(n376), .C0(n375), .Y(n378) );
  AOI22X1TS U738 ( .A0(n348), .A1(\dataToWriteBuffer[5][2] ), .B0(n392), .B1(
        dataIn_EAST[2]), .Y(n380) );
  AOI22X1TS U739 ( .A0(n398), .A1(\dataToWriteBuffer[6][2] ), .B0(n428), .B1(
        dataIn_SOUTH[2]), .Y(n379) );
  OAI211XLTS U740 ( .A0(n432), .A1(n381), .B0(n380), .C0(n379), .Y(n382) );
  AOI22X1TS U741 ( .A0(n419), .A1(\dataToWriteBuffer[5][5] ), .B0(n418), .B1(
        dataIn_EAST[5]), .Y(n384) );
  AOI22X1TS U742 ( .A0(n469), .A1(\dataToWriteBuffer[6][5] ), .B0(n420), .B1(
        dataIn_SOUTH[5]), .Y(n383) );
  AOI22X1TS U743 ( .A0(n403), .A1(\dataToWriteBuffer[5][3] ), .B0(n392), .B1(
        dataIn_EAST[3]), .Y(n389) );
  AOI22X1TS U744 ( .A0(n404), .A1(\dataToWriteBuffer[6][3] ), .B0(n387), .B1(
        dataIn_SOUTH[3]), .Y(n388) );
  AOI22X1TS U745 ( .A0(n410), .A1(\dataToWriteBuffer[5][4] ), .B0(n392), .B1(
        dataIn_EAST[4]), .Y(n394) );
  AOI22X1TS U746 ( .A0(n465), .A1(\dataToWriteBuffer[6][4] ), .B0(n428), .B1(
        dataIn_SOUTH[4]), .Y(n393) );
  INVX2TS U747 ( .A(n397), .Y(n427) );
  AOI22X1TS U748 ( .A0(n410), .A1(\addressToWriteBuffer[5][1] ), .B0(n427), 
        .B1(cacheAddressIn_EAST[1]), .Y(n400) );
  INVX2TS U749 ( .A(n17), .Y(n411) );
  AOI22X1TS U750 ( .A0(n398), .A1(\addressToWriteBuffer[6][1] ), .B0(n411), 
        .B1(cacheAddressIn_SOUTH[1]), .Y(n399) );
  AOI22X1TS U751 ( .A0(n403), .A1(\addressToWriteBuffer[5][3] ), .B0(n427), 
        .B1(cacheAddressIn_EAST[3]), .Y(n406) );
  AOI22X1TS U752 ( .A0(n404), .A1(\addressToWriteBuffer[6][3] ), .B0(n411), 
        .B1(cacheAddressIn_SOUTH[3]), .Y(n405) );
  AOI22X1TS U753 ( .A0(n410), .A1(\addressToWriteBuffer[5][2] ), .B0(n427), 
        .B1(cacheAddressIn_EAST[2]), .Y(n413) );
  AOI22X1TS U754 ( .A0(n461), .A1(\addressToWriteBuffer[6][2] ), .B0(n411), 
        .B1(cacheAddressIn_SOUTH[2]), .Y(n412) );
  AOI22X1TS U755 ( .A0(n419), .A1(\dataToWriteBuffer[5][1] ), .B0(n418), .B1(
        dataIn_EAST[1]), .Y(n422) );
  AOI22X1TS U756 ( .A0(n491), .A1(\dataToWriteBuffer[6][1] ), .B0(n420), .B1(
        dataIn_SOUTH[1]), .Y(n421) );
  AOI22X1TS U757 ( .A0(n348), .A1(\dataToWriteBuffer[5][0] ), .B0(n427), .B1(
        dataIn_EAST[0]), .Y(n430) );
  AOI22X1TS U758 ( .A0(n398), .A1(\dataToWriteBuffer[6][0] ), .B0(n428), .B1(
        dataIn_SOUTH[0]), .Y(n429) );
  AOI22X1TS U759 ( .A0(memWrite_EAST), .A1(n435), .B0(memWrite_SOUTH), .B1(
        n229), .Y(n436) );
  AOI22X1TS U760 ( .A0(n136), .A1(n621), .B0(n436), .B1(n135), .Y(n679) );
  OR2X1TS U761 ( .A(n438), .B(n437), .Y(n677) );
  NOR2BX1TS U762 ( .AN(n441), .B(n341), .Y(n442) );
  OR2X1TS U763 ( .A(n443), .B(n615), .Y(n549) );
  INVX2TS U764 ( .A(n549), .Y(n590) );
  AOI22X1TS U765 ( .A0(\requesterPortBuffer[2][1] ), .A1(n590), .B0(
        \requesterPortBuffer[3][1] ), .B1(n531), .Y(n445) );
  NAND2X1TS U766 ( .A(n442), .B(n617), .Y(n444) );
  INVX2TS U767 ( .A(n535), .Y(n618) );
  AOI21X1TS U768 ( .A0(\requesterPortBuffer[3][0] ), .A1(n618), .B0(n443), .Y(
        n450) );
  CLKBUFX2TS U769 ( .A(n447), .Y(n579) );
  CLKBUFX2TS U770 ( .A(n579), .Y(n625) );
  INVX2TS U771 ( .A(n549), .Y(n448) );
  AOI22X1TS U772 ( .A0(n625), .A1(\requesterPortBuffer[4][0] ), .B0(
        \requesterPortBuffer[2][0] ), .B1(n556), .Y(n449) );
  INVX2TS U773 ( .A(n452), .Y(n481) );
  AOI22X1TS U774 ( .A0(n729), .A1(n481), .B0(n54), .B1(
        \addressToWriteBuffer[1][6] ), .Y(n455) );
  INVX2TS U775 ( .A(n453), .Y(n482) );
  AOI22X1TS U776 ( .A0(n62), .A1(\addressToWriteBuffer[2][6] ), .B0(n482), 
        .B1(\addressToWriteBuffer[3][6] ), .Y(n454) );
  AOI22X1TS U777 ( .A0(n686), .A1(n489), .B0(n480), .B1(
        \dataToWriteBuffer[1][0] ), .Y(n458) );
  AOI22X1TS U778 ( .A0(n483), .A1(\dataToWriteBuffer[2][0] ), .B0(n490), .B1(
        \dataToWriteBuffer[3][0] ), .Y(n457) );
  AOI22X1TS U779 ( .A0(n723), .A1(n481), .B0(n460), .B1(
        \addressToWriteBuffer[1][7] ), .Y(n463) );
  AOI22X1TS U780 ( .A0(n461), .A1(\addressToWriteBuffer[2][7] ), .B0(n475), 
        .B1(\addressToWriteBuffer[3][7] ), .Y(n462) );
  AOI22X1TS U781 ( .A0(n756), .A1(n481), .B0(n54), .B1(
        \addressToWriteBuffer[1][2] ), .Y(n467) );
  AOI22X1TS U782 ( .A0(n465), .A1(\addressToWriteBuffer[2][2] ), .B0(n482), 
        .B1(\addressToWriteBuffer[3][2] ), .Y(n466) );
  AOI22X1TS U783 ( .A0(n690), .A1(n474), .B0(n488), .B1(
        \dataToWriteBuffer[1][1] ), .Y(n471) );
  AOI22X1TS U784 ( .A0(n469), .A1(\dataToWriteBuffer[2][1] ), .B0(n482), .B1(
        \dataToWriteBuffer[3][1] ), .Y(n470) );
  AOI22X1TS U785 ( .A0(n707), .A1(n474), .B0(n480), .B1(
        \dataToWriteBuffer[1][4] ), .Y(n477) );
  AOI22X1TS U786 ( .A0(n483), .A1(\dataToWriteBuffer[2][4] ), .B0(n475), .B1(
        \dataToWriteBuffer[3][4] ), .Y(n476) );
  AOI22X1TS U787 ( .A0(n740), .A1(n481), .B0(n480), .B1(
        \addressToWriteBuffer[1][4] ), .Y(n485) );
  AOI22X1TS U788 ( .A0(n483), .A1(\addressToWriteBuffer[2][4] ), .B0(n482), 
        .B1(\addressToWriteBuffer[3][4] ), .Y(n484) );
  AOI22X1TS U789 ( .A0(n712), .A1(n489), .B0(n488), .B1(
        \dataToWriteBuffer[1][5] ), .Y(n493) );
  AOI22X1TS U790 ( .A0(n491), .A1(\dataToWriteBuffer[2][5] ), .B0(n490), .B1(
        \dataToWriteBuffer[3][5] ), .Y(n492) );
  AOI22X1TS U791 ( .A0(n625), .A1(\requesterPortBuffer[1][1] ), .B0(
        \prevRequesterPort_B[1] ), .B1(n497), .Y(n496) );
  AOI22X1TS U792 ( .A0(n625), .A1(\requesterPortBuffer[1][0] ), .B0(n7), .B1(
        n497), .Y(n499) );
  AO22XLTS U793 ( .A0(n503), .A1(\requesterPortBuffer[4][0] ), .B0(n502), .B1(
        \requesterPortBuffer[5][0] ), .Y(n827) );
  AO22XLTS U794 ( .A0(n784), .A1(prevMemRead_A), .B0(n777), .B1(prevMemRead_B), 
        .Y(N5340) );
  AO22X1TS U795 ( .A0(n508), .A1(n507), .B0(n506), .B1(n505), .Y(N5377) );
  AO22X1TS U796 ( .A0(n198), .A1(n511), .B0(n510), .B1(n509), .Y(N5378) );
  OR3X1TS U797 ( .A(n514), .B(n512), .C(n677), .Y(n702) );
  INVX2TS U798 ( .A(n702), .Y(n691) );
  NOR2XLTS U799 ( .A(n41), .B(n513), .Y(n660) );
  CLKBUFX2TS U800 ( .A(n660), .Y(n666) );
  NAND2X1TS U801 ( .A(n33), .B(n514), .Y(n517) );
  NAND2X1TS U802 ( .A(n34), .B(n652), .Y(n684) );
  INVX2TS U803 ( .A(n16), .Y(n651) );
  AOI22X1TS U804 ( .A0(\requesterPortBuffer[0][0] ), .A1(n666), .B0(n519), 
        .B1(n651), .Y(n520) );
  INVX2TS U805 ( .A(n522), .Y(n665) );
  INVX2TS U806 ( .A(n665), .Y(n746) );
  AOI22X1TS U807 ( .A0(\requesterPortBuffer[0][1] ), .A1(n666), .B0(n4), .B1(
        n651), .Y(n523) );
  AOI22X1TS U808 ( .A0(n528), .A1(\requesterAddressBuffer[0][0] ), .B0(
        requesterAddressIn_SOUTH[0]), .B1(n527), .Y(n524) );
  OAI2BB1X1TS U809 ( .A0N(requesterAddressIn_EAST[0]), .A1N(n526), .B0(n524), 
        .Y(n1354) );
  AOI22X1TS U810 ( .A0(n528), .A1(\requesterAddressBuffer[0][1] ), .B0(
        requesterAddressIn_SOUTH[1]), .B1(n527), .Y(n525) );
  OAI2BB1X1TS U811 ( .A0N(requesterAddressIn_EAST[1]), .A1N(n526), .B0(n525), 
        .Y(n1353) );
  AOI22X1TS U812 ( .A0(n528), .A1(\requesterAddressBuffer[0][2] ), .B0(
        requesterAddressIn_SOUTH[2]), .B1(n527), .Y(n529) );
  OAI2BB1X1TS U813 ( .A0N(requesterAddressIn_EAST[2]), .A1N(n530), .B0(n529), 
        .Y(n1352) );
  AOI22X1TS U814 ( .A0(n532), .A1(\requesterAddressBuffer[0][3] ), .B0(
        requesterAddressIn_SOUTH[3]), .B1(n531), .Y(n533) );
  OAI2BB1X1TS U815 ( .A0N(requesterAddressIn_EAST[3]), .A1N(n534), .B0(n533), 
        .Y(n1351) );
  NAND2X1TS U816 ( .A(n537), .B(n536), .Y(n544) );
  AOI22X1TS U817 ( .A0(requesterAddressIn_EAST[0]), .A1(n543), .B0(
        requesterAddressIn_WEST[0]), .B1(n544), .Y(n540) );
  NAND2X1TS U818 ( .A(n538), .B(n611), .Y(n573) );
  INVX2TS U819 ( .A(n611), .Y(n539) );
  OAI2BB2XLTS U820 ( .B0(n540), .B1(n573), .A0N(n577), .A1N(
        \requesterAddressBuffer[1][0] ), .Y(n1350) );
  AOI22X1TS U821 ( .A0(requesterAddressIn_WEST[1]), .A1(n544), .B0(
        requesterAddressIn_EAST[1]), .B1(n543), .Y(n541) );
  CLKBUFX2TS U822 ( .A(n573), .Y(n612) );
  OAI2BB2XLTS U823 ( .B0(n541), .B1(n612), .A0N(n539), .A1N(
        \requesterAddressBuffer[1][1] ), .Y(n1349) );
  AOI22X1TS U824 ( .A0(requesterAddressIn_WEST[2]), .A1(n544), .B0(
        requesterAddressIn_EAST[2]), .B1(n543), .Y(n542) );
  OAI2BB2XLTS U825 ( .B0(n542), .B1(n612), .A0N(n539), .A1N(
        \requesterAddressBuffer[1][2] ), .Y(n1348) );
  AOI22X1TS U826 ( .A0(requesterAddressIn_WEST[3]), .A1(n544), .B0(
        requesterAddressIn_EAST[3]), .B1(n543), .Y(n545) );
  OAI2BB2XLTS U827 ( .B0(n545), .B1(n612), .A0N(n539), .A1N(
        \requesterAddressBuffer[1][3] ), .Y(n1347) );
  CLKBUFX2TS U828 ( .A(n555), .Y(n603) );
  AOI22X1TS U829 ( .A0(\addressToWriteBuffer[3][0] ), .A1(n603), .B0(n579), 
        .B1(\addressToWriteBuffer[4][0] ), .Y(n548) );
  INVX2TS U830 ( .A(n546), .Y(n560) );
  INVX2TS U831 ( .A(n549), .Y(n599) );
  AOI22X1TS U832 ( .A0(n771), .A1(n591), .B0(\addressToWriteBuffer[2][0] ), 
        .B1(n599), .Y(n547) );
  NAND2X1TS U833 ( .A(n548), .B(n547), .Y(n1330) );
  CLKBUFX2TS U834 ( .A(n554), .Y(n585) );
  AOI22X1TS U835 ( .A0(\addressToWriteBuffer[3][1] ), .A1(n555), .B0(n585), 
        .B1(\addressToWriteBuffer[4][1] ), .Y(n551) );
  INVX2TS U836 ( .A(n560), .Y(n605) );
  INVX2TS U837 ( .A(n549), .Y(n604) );
  AOI22X1TS U838 ( .A0(n765), .A1(n605), .B0(\addressToWriteBuffer[2][1] ), 
        .B1(n604), .Y(n550) );
  NAND2X1TS U839 ( .A(n551), .B(n550), .Y(n1329) );
  AOI22X1TS U840 ( .A0(\addressToWriteBuffer[3][2] ), .A1(n603), .B0(n585), 
        .B1(\addressToWriteBuffer[4][2] ), .Y(n553) );
  INVX2TS U841 ( .A(n560), .Y(n595) );
  AOI22X1TS U842 ( .A0(n756), .A1(n595), .B0(\addressToWriteBuffer[2][2] ), 
        .B1(n590), .Y(n552) );
  NAND2X1TS U843 ( .A(n553), .B(n552), .Y(n1328) );
  CLKBUFX2TS U844 ( .A(n554), .Y(n598) );
  AOI22X1TS U845 ( .A0(\addressToWriteBuffer[3][3] ), .A1(n555), .B0(n598), 
        .B1(\addressToWriteBuffer[4][3] ), .Y(n558) );
  AOI22X1TS U846 ( .A0(n748), .A1(n595), .B0(\addressToWriteBuffer[2][3] ), 
        .B1(n556), .Y(n557) );
  NAND2X1TS U847 ( .A(n558), .B(n557), .Y(n1327) );
  CLKBUFX2TS U848 ( .A(n559), .Y(n594) );
  AOI22X1TS U849 ( .A0(\addressToWriteBuffer[3][4] ), .A1(n594), .B0(n585), 
        .B1(\addressToWriteBuffer[4][4] ), .Y(n562) );
  INVX2TS U850 ( .A(n560), .Y(n591) );
  AOI22X1TS U851 ( .A0(n740), .A1(n591), .B0(\addressToWriteBuffer[2][4] ), 
        .B1(n599), .Y(n561) );
  NAND2X1TS U852 ( .A(n562), .B(n561), .Y(n1326) );
  CLKBUFX2TS U853 ( .A(n563), .Y(n586) );
  AOI22X1TS U854 ( .A0(\addressToWriteBuffer[3][5] ), .A1(n586), .B0(n579), 
        .B1(\addressToWriteBuffer[4][5] ), .Y(n565) );
  AOI22X1TS U855 ( .A0(n734), .A1(n546), .B0(\addressToWriteBuffer[2][5] ), 
        .B1(n604), .Y(n564) );
  NAND2X1TS U856 ( .A(n565), .B(n564), .Y(n1325) );
  AOI22X1TS U857 ( .A0(\addressToWriteBuffer[3][6] ), .A1(n594), .B0(n598), 
        .B1(\addressToWriteBuffer[4][6] ), .Y(n567) );
  AOI22X1TS U858 ( .A0(n729), .A1(n605), .B0(\addressToWriteBuffer[2][6] ), 
        .B1(n590), .Y(n566) );
  NAND2X1TS U859 ( .A(n567), .B(n566), .Y(n1324) );
  AOI22X1TS U860 ( .A0(\addressToWriteBuffer[3][7] ), .A1(n586), .B0(n602), 
        .B1(\addressToWriteBuffer[4][7] ), .Y(n569) );
  AOI22X1TS U861 ( .A0(n723), .A1(n595), .B0(\addressToWriteBuffer[2][7] ), 
        .B1(n556), .Y(n568) );
  NAND2X1TS U862 ( .A(n569), .B(n568), .Y(n1323) );
  INVX2TS U863 ( .A(n611), .Y(n577) );
  AOI22X1TS U864 ( .A0(\requesterPortBuffer[2][0] ), .A1(n618), .B0(
        \requesterPortBuffer[3][0] ), .B1(n39), .Y(n570) );
  AOI21X1TS U865 ( .A0(n570), .A1(n55), .B0(n573), .Y(n571) );
  AOI22X1TS U866 ( .A0(\requesterPortBuffer[2][1] ), .A1(n37), .B0(
        \requesterPortBuffer[3][1] ), .B1(n572), .Y(n575) );
  AOI31XLTS U867 ( .A0(n575), .A1(n574), .A2(n536), .B0(n573), .Y(n576) );
  NAND2X1TS U868 ( .A(n628), .B(\requesterPortBuffer[5][0] ), .Y(n582) );
  NAND4XLTS U869 ( .A(n33), .B(n580), .C(n579), .D(n578), .Y(n581) );
  AOI22X1TS U870 ( .A0(\dataToWriteBuffer[3][0] ), .A1(n586), .B0(n598), .B1(
        \dataToWriteBuffer[4][0] ), .Y(n584) );
  AOI22X1TS U871 ( .A0(n686), .A1(n605), .B0(\dataToWriteBuffer[2][0] ), .B1(
        n599), .Y(n583) );
  NAND2X1TS U872 ( .A(n584), .B(n583), .Y(n1255) );
  AOI22X1TS U873 ( .A0(\dataToWriteBuffer[3][1] ), .A1(n586), .B0(n585), .B1(
        \dataToWriteBuffer[4][1] ), .Y(n588) );
  AOI22X1TS U874 ( .A0(n690), .A1(n591), .B0(\dataToWriteBuffer[2][1] ), .B1(
        n604), .Y(n587) );
  NAND2X1TS U875 ( .A(n588), .B(n587), .Y(n1254) );
  AOI22X1TS U876 ( .A0(\dataToWriteBuffer[3][2] ), .A1(n594), .B0(n589), .B1(
        \dataToWriteBuffer[4][2] ), .Y(n593) );
  AOI22X1TS U877 ( .A0(n695), .A1(n591), .B0(\dataToWriteBuffer[2][2] ), .B1(
        n590), .Y(n592) );
  NAND2X1TS U878 ( .A(n593), .B(n592), .Y(n1253) );
  AOI22X1TS U879 ( .A0(\dataToWriteBuffer[3][3] ), .A1(n594), .B0(n602), .B1(
        \dataToWriteBuffer[4][3] ), .Y(n597) );
  AOI22X1TS U880 ( .A0(n701), .A1(n595), .B0(\dataToWriteBuffer[2][3] ), .B1(
        n448), .Y(n596) );
  NAND2X1TS U881 ( .A(n597), .B(n596), .Y(n1252) );
  AOI22X1TS U882 ( .A0(\dataToWriteBuffer[3][4] ), .A1(n603), .B0(n598), .B1(
        \dataToWriteBuffer[4][4] ), .Y(n601) );
  AOI22X1TS U883 ( .A0(n707), .A1(n546), .B0(\dataToWriteBuffer[2][4] ), .B1(
        n599), .Y(n600) );
  NAND2X1TS U884 ( .A(n601), .B(n600), .Y(n1251) );
  AOI22X1TS U885 ( .A0(\dataToWriteBuffer[3][5] ), .A1(n603), .B0(n602), .B1(
        \dataToWriteBuffer[4][5] ), .Y(n607) );
  AOI22X1TS U886 ( .A0(n712), .A1(n605), .B0(\dataToWriteBuffer[2][5] ), .B1(
        n604), .Y(n606) );
  NAND2X1TS U887 ( .A(n607), .B(n606), .Y(n1250) );
  CLKBUFX2TS U888 ( .A(memWrite_EAST), .Y(n627) );
  AOI22X1TS U889 ( .A0(n608), .A1(n627), .B0(isWrite[3]), .B1(n39), .Y(n609)
         );
  AOI21X1TS U890 ( .A0(n37), .A1(isWrite[2]), .B0(n610), .Y(n613) );
  OAI22X1TS U891 ( .A0(n613), .A1(n612), .B0(n611), .B1(n834), .Y(n1218) );
  INVX2TS U892 ( .A(n837), .Y(n814) );
  AOI222XLTS U893 ( .A0(n39), .A1(isWrite[4]), .B0(isWrite[3]), .B1(n618), 
        .C0(memWrite_WEST), .C1(n443), .Y(n614) );
  OAI2BB2XLTS U894 ( .B0(n814), .B1(n614), .A0N(n556), .A1N(isWrite[2]), .Y(
        n1217) );
  INVX2TS U895 ( .A(n671), .Y(n790) );
  AOI22X1TS U896 ( .A0(isWrite[4]), .A1(n37), .B0(isWrite[5]), .B1(n38), .Y(
        n616) );
  INVX2TS U897 ( .A(n615), .Y(n619) );
  OAI2BB2XLTS U898 ( .B0(n790), .B1(n616), .A0N(isWrite[3]), .A1N(n619), .Y(
        n1216) );
  INVX2TS U899 ( .A(n617), .Y(n802) );
  NAND2X1TS U900 ( .A(isWrite[5]), .B(n618), .Y(n620) );
  OAI2BB2XLTS U901 ( .B0(n802), .B1(n620), .A0N(isWrite[4]), .A1N(n619), .Y(
        n1215) );
  INVX2TS U902 ( .A(n621), .Y(n624) );
  INVX2TS U903 ( .A(n622), .Y(n623) );
  NAND2X1TS U904 ( .A(n624), .B(n623), .Y(n631) );
  OAI211XLTS U905 ( .A0(n627), .A1(n626), .B0(n625), .C0(n216), .Y(n629) );
  AOI32X1TS U906 ( .A0(n631), .A1(n630), .A2(n629), .B0(n628), .B1(n835), .Y(
        n1214) );
  INVX2TS U907 ( .A(n632), .Y(n637) );
  OAI22X1TS U908 ( .A0(n640), .A1(n639), .B0(n134), .B1(n633), .Y(n634) );
  XNOR2X1TS U909 ( .A(n638), .B(n634), .Y(n636) );
  OAI21XLTS U910 ( .A0(n637), .A1(n636), .B0(n646), .Y(n635) );
  AOI21X1TS U911 ( .A0(n637), .A1(n636), .B0(n635), .Y(n1210) );
  OA21XLTS U912 ( .A0(n643), .A1(n645), .B0(n638), .Y(n642) );
  AOI211XLTS U913 ( .A0(n645), .A1(n643), .B0(n642), .C0(n641), .Y(n649) );
  OR2X1TS U914 ( .A(N742), .B(n832), .Y(n644) );
  OAI21XLTS U915 ( .A0(n21), .A1(n645), .B0(n644), .Y(n648) );
  AOI21X1TS U916 ( .A0(n649), .A1(n648), .B0(n647), .Y(n1209) );
  CLKBUFX2TS U917 ( .A(n650), .Y(n706) );
  INVX2TS U918 ( .A(n706), .Y(n764) );
  INVX2TS U919 ( .A(n16), .Y(n664) );
  AOI22X1TS U920 ( .A0(requesterAddressIn_WEST[0]), .A1(n764), .B0(n817), .B1(
        n664), .Y(n656) );
  INVX2TS U921 ( .A(n665), .Y(n763) );
  AOI22X1TS U922 ( .A0(requesterAddressIn_EAST[0]), .A1(n763), .B0(n660), .B1(
        \requesterAddressBuffer[0][0] ), .Y(n655) );
  INVX2TS U923 ( .A(n653), .Y(n667) );
  INVX2TS U924 ( .A(n667), .Y(n749) );
  AOI22X1TS U925 ( .A0(n724), .A1(requesterAddressIn_SOUTH[0]), .B0(n749), 
        .B1(requesterAddressIn_NORTH[0]), .Y(n654) );
  INVX2TS U926 ( .A(n706), .Y(n733) );
  AOI22X1TS U927 ( .A0(requesterAddressIn_WEST[1]), .A1(n733), .B0(n812), .B1(
        n664), .Y(n659) );
  INVX2TS U928 ( .A(n665), .Y(n739) );
  AOI22X1TS U929 ( .A0(requesterAddressIn_EAST[1]), .A1(n739), .B0(n660), .B1(
        \requesterAddressBuffer[0][1] ), .Y(n658) );
  INVX2TS U930 ( .A(n702), .Y(n741) );
  INVX2TS U931 ( .A(n667), .Y(n773) );
  AOI22X1TS U932 ( .A0(n741), .A1(requesterAddressIn_SOUTH[1]), .B0(n773), 
        .B1(requesterAddressIn_NORTH[1]), .Y(n657) );
  INVX2TS U933 ( .A(n706), .Y(n755) );
  AOI22X1TS U934 ( .A0(requesterAddressIn_WEST[2]), .A1(n755), .B0(n809), .B1(
        n664), .Y(n663) );
  AOI22X1TS U935 ( .A0(requesterAddressIn_EAST[2]), .A1(n522), .B0(n660), .B1(
        \requesterAddressBuffer[0][2] ), .Y(n662) );
  INVX2TS U936 ( .A(n702), .Y(n772) );
  INVX2TS U937 ( .A(n667), .Y(n735) );
  AOI22X1TS U938 ( .A0(n772), .A1(requesterAddressIn_SOUTH[2]), .B0(n735), 
        .B1(requesterAddressIn_NORTH[2]), .Y(n661) );
  AOI22X1TS U939 ( .A0(requesterAddressIn_WEST[3]), .A1(n755), .B0(n803), .B1(
        n664), .Y(n670) );
  INVX2TS U940 ( .A(n665), .Y(n728) );
  AOI22X1TS U941 ( .A0(requesterAddressIn_EAST[3]), .A1(n728), .B0(n666), .B1(
        \requesterAddressBuffer[0][3] ), .Y(n669) );
  INVX2TS U942 ( .A(n667), .Y(n757) );
  AOI22X1TS U943 ( .A0(n691), .A1(requesterAddressIn_SOUTH[3]), .B0(n757), 
        .B1(requesterAddressIn_NORTH[3]), .Y(n668) );
  NAND2X1TS U944 ( .A(n719), .B(n671), .Y(n683) );
  AOI22X1TS U945 ( .A0(memWrite_WEST), .A1(n673), .B0(memWrite_EAST), .B1(n672), .Y(n675) );
  OAI211XLTS U946 ( .A0(memRead_NORTH), .A1(n676), .B0(n675), .C0(n674), .Y(
        n718) );
  OAI22X1TS U947 ( .A0(isWrite[0]), .A1(n683), .B0(n718), .B1(n677), .Y(n1203)
         );
  OAI221XLTS U948 ( .A0(n720), .A1(isWrite[1]), .B0(n719), .B1(n679), .C0(n678), .Y(n680) );
  CLKBUFX2TS U949 ( .A(n683), .Y(n699) );
  INVX2TS U950 ( .A(n699), .Y(n762) );
  INVX2TS U951 ( .A(n14), .Y(n700) );
  AOI22X1TS U952 ( .A0(n762), .A1(\dataToWriteBuffer[0][0] ), .B0(n700), .B1(
        cacheDataIn_A[0]), .Y(n689) );
  AOI22X1TS U953 ( .A0(n686), .A1(n755), .B0(dataIn_EAST[0]), .B1(n728), .Y(
        n688) );
  AOI22X1TS U954 ( .A0(dataIn_NORTH[0]), .A1(n749), .B0(dataIn_SOUTH[0]), .B1(
        n691), .Y(n687) );
  INVX2TS U955 ( .A(n699), .Y(n770) );
  AOI22X1TS U956 ( .A0(n770), .A1(\dataToWriteBuffer[0][1] ), .B0(n700), .B1(
        cacheDataIn_A[1]), .Y(n694) );
  AOI22X1TS U957 ( .A0(n690), .A1(n747), .B0(dataIn_EAST[1]), .B1(n746), .Y(
        n693) );
  AOI22X1TS U958 ( .A0(dataIn_NORTH[1]), .A1(n735), .B0(dataIn_SOUTH[1]), .B1(
        n691), .Y(n692) );
  INVX2TS U959 ( .A(n699), .Y(n745) );
  AOI22X1TS U960 ( .A0(n745), .A1(\dataToWriteBuffer[0][2] ), .B0(n700), .B1(
        cacheDataIn_A[2]), .Y(n698) );
  AOI22X1TS U961 ( .A0(n695), .A1(n764), .B0(dataIn_EAST[2]), .B1(n739), .Y(
        n697) );
  AOI22X1TS U962 ( .A0(dataIn_NORTH[2]), .A1(n749), .B0(dataIn_SOUTH[2]), .B1(
        n724), .Y(n696) );
  INVX2TS U963 ( .A(n699), .Y(n754) );
  AOI22X1TS U964 ( .A0(n754), .A1(\dataToWriteBuffer[0][3] ), .B0(n700), .B1(
        cacheDataIn_A[3]), .Y(n705) );
  AOI22X1TS U965 ( .A0(n701), .A1(n733), .B0(dataIn_EAST[3]), .B1(n763), .Y(
        n704) );
  INVX2TS U966 ( .A(n702), .Y(n713) );
  AOI22X1TS U967 ( .A0(dataIn_NORTH[3]), .A1(n735), .B0(dataIn_SOUTH[3]), .B1(
        n713), .Y(n703) );
  INVX2TS U968 ( .A(n14), .Y(n769) );
  AOI22X1TS U969 ( .A0(n762), .A1(\dataToWriteBuffer[0][4] ), .B0(n769), .B1(
        cacheDataIn_A[4]), .Y(n710) );
  INVX2TS U970 ( .A(n706), .Y(n747) );
  AOI22X1TS U971 ( .A0(n707), .A1(n747), .B0(dataIn_EAST[4]), .B1(n728), .Y(
        n709) );
  AOI22X1TS U972 ( .A0(dataIn_NORTH[4]), .A1(n757), .B0(dataIn_SOUTH[4]), .B1(
        n713), .Y(n708) );
  INVX2TS U973 ( .A(n14), .Y(n753) );
  AOI22X1TS U974 ( .A0(n770), .A1(\dataToWriteBuffer[0][5] ), .B0(n753), .B1(
        cacheDataIn_A[5]), .Y(n716) );
  AOI22X1TS U975 ( .A0(n712), .A1(n711), .B0(dataIn_EAST[5]), .B1(n739), .Y(
        n715) );
  AOI22X1TS U976 ( .A0(dataIn_NORTH[5]), .A1(n773), .B0(dataIn_SOUTH[5]), .B1(
        n713), .Y(n714) );
  OAI221XLTS U977 ( .A0(n720), .A1(isWrite[0]), .B0(n719), .B1(n718), .C0(n717), .Y(n721) );
  INVX2TS U978 ( .A(n721), .Y(n722) );
  INVX2TS U979 ( .A(n14), .Y(n761) );
  OAI2BB2XLTS U980 ( .B0(n753), .B1(n722), .A0N(n761), .A1N(memWrite_A), .Y(
        n1181) );
  AOI22X1TS U981 ( .A0(n745), .A1(\addressToWriteBuffer[0][7] ), .B0(n761), 
        .B1(cacheAddressIn_A[7]), .Y(n727) );
  AOI22X1TS U982 ( .A0(n723), .A1(n733), .B0(cacheAddressIn_EAST[7]), .B1(n746), .Y(n726) );
  AOI22X1TS U983 ( .A0(cacheAddressIn_NORTH[7]), .A1(n773), .B0(
        cacheAddressIn_SOUTH[7]), .B1(n713), .Y(n725) );
  AOI22X1TS U984 ( .A0(n754), .A1(\addressToWriteBuffer[0][6] ), .B0(n769), 
        .B1(cacheAddressIn_A[6]), .Y(n732) );
  AOI22X1TS U985 ( .A0(n729), .A1(n747), .B0(cacheAddressIn_EAST[6]), .B1(n728), .Y(n731) );
  AOI22X1TS U986 ( .A0(cacheAddressIn_NORTH[6]), .A1(n757), .B0(
        cacheAddressIn_SOUTH[6]), .B1(n741), .Y(n730) );
  AOI22X1TS U987 ( .A0(n762), .A1(\addressToWriteBuffer[0][5] ), .B0(n753), 
        .B1(cacheAddressIn_A[5]), .Y(n738) );
  AOI22X1TS U988 ( .A0(n734), .A1(n733), .B0(cacheAddressIn_EAST[5]), .B1(n763), .Y(n737) );
  AOI22X1TS U989 ( .A0(cacheAddressIn_NORTH[5]), .A1(n735), .B0(
        cacheAddressIn_SOUTH[5]), .B1(n741), .Y(n736) );
  AOI22X1TS U990 ( .A0(n770), .A1(\addressToWriteBuffer[0][4] ), .B0(n761), 
        .B1(cacheAddressIn_A[4]), .Y(n744) );
  AOI22X1TS U991 ( .A0(n740), .A1(n711), .B0(cacheAddressIn_EAST[4]), .B1(n739), .Y(n743) );
  AOI22X1TS U992 ( .A0(cacheAddressIn_NORTH[4]), .A1(n653), .B0(
        cacheAddressIn_SOUTH[4]), .B1(n741), .Y(n742) );
  AOI22X1TS U993 ( .A0(n745), .A1(\addressToWriteBuffer[0][3] ), .B0(n769), 
        .B1(cacheAddressIn_A[3]), .Y(n752) );
  AOI22X1TS U994 ( .A0(n748), .A1(n747), .B0(cacheAddressIn_EAST[3]), .B1(n746), .Y(n751) );
  AOI22X1TS U995 ( .A0(cacheAddressIn_NORTH[3]), .A1(n749), .B0(
        cacheAddressIn_SOUTH[3]), .B1(n724), .Y(n750) );
  AOI22X1TS U996 ( .A0(n754), .A1(\addressToWriteBuffer[0][2] ), .B0(n753), 
        .B1(cacheAddressIn_A[2]), .Y(n760) );
  AOI22X1TS U997 ( .A0(n756), .A1(n755), .B0(cacheAddressIn_EAST[2]), .B1(n522), .Y(n759) );
  AOI22X1TS U998 ( .A0(cacheAddressIn_NORTH[2]), .A1(n757), .B0(
        cacheAddressIn_SOUTH[2]), .B1(n772), .Y(n758) );
  AOI22X1TS U999 ( .A0(n762), .A1(\addressToWriteBuffer[0][1] ), .B0(n761), 
        .B1(cacheAddressIn_A[1]), .Y(n768) );
  AOI22X1TS U1000 ( .A0(n765), .A1(n764), .B0(cacheAddressIn_EAST[1]), .B1(
        n763), .Y(n767) );
  AOI22X1TS U1001 ( .A0(cacheAddressIn_NORTH[1]), .A1(n653), .B0(
        cacheAddressIn_SOUTH[1]), .B1(n772), .Y(n766) );
  AOI22X1TS U1002 ( .A0(n770), .A1(\addressToWriteBuffer[0][0] ), .B0(n769), 
        .B1(cacheAddressIn_A[0]), .Y(n776) );
  AOI22X1TS U1003 ( .A0(n771), .A1(n711), .B0(cacheAddressIn_EAST[0]), .B1(
        n522), .Y(n775) );
  AOI22X1TS U1004 ( .A0(cacheAddressIn_NORTH[0]), .A1(n773), .B0(
        cacheAddressIn_SOUTH[0]), .B1(n772), .Y(n774) );
  AOI22X1TS U1005 ( .A0(n803), .A1(n787), .B0(prevRequesterAddress_B[3]), .B1(
        n783), .Y(n779) );
  NOR3XLTS U1006 ( .A(n778), .B(n781), .C(n777), .Y(n788) );
  OAI2BB2XLTS U1007 ( .B0(n780), .B1(n779), .A0N(requesterAddressOut_WEST[3]), 
        .A1N(n788), .Y(n1171) );
  AOI22X1TS U1008 ( .A0(n809), .A1(n781), .B0(prevRequesterAddress_B[2]), .B1(
        n786), .Y(n782) );
  OAI2BB2XLTS U1009 ( .B0(n790), .B1(n782), .A0N(requesterAddressOut_WEST[2]), 
        .A1N(n788), .Y(n1170) );
  AOI22X1TS U1010 ( .A0(n812), .A1(n784), .B0(prevRequesterAddress_B[1]), .B1(
        n783), .Y(n785) );
  OAI2BB2XLTS U1011 ( .B0(n790), .B1(n785), .A0N(requesterAddressOut_WEST[1]), 
        .A1N(n788), .Y(n1169) );
  AOI22X1TS U1012 ( .A0(n817), .A1(n787), .B0(prevRequesterAddress_B[0]), .B1(
        n786), .Y(n789) );
  OAI2BB2XLTS U1013 ( .B0(n790), .B1(n789), .A0N(requesterAddressOut_WEST[0]), 
        .A1N(n788), .Y(n1168) );
  AOI22X1TS U1014 ( .A0(prevRequesterAddress_A[3]), .A1(n799), .B0(
        prevRequesterAddress_B[3]), .B1(n796), .Y(n792) );
  NOR3XLTS U1015 ( .A(n806), .B(n799), .C(n791), .Y(n800) );
  OAI2BB2XLTS U1016 ( .B0(n802), .B1(n792), .A0N(requesterAddressOut_EAST[3]), 
        .A1N(n800), .Y(n1167) );
  AOI22X1TS U1017 ( .A0(prevRequesterAddress_A[2]), .A1(n793), .B0(
        prevRequesterAddress_B[2]), .B1(n798), .Y(n794) );
  OAI2BB2XLTS U1018 ( .B0(n802), .B1(n794), .A0N(requesterAddressOut_EAST[2]), 
        .A1N(n800), .Y(n1166) );
  AOI22X1TS U1019 ( .A0(prevRequesterAddress_A[1]), .A1(n22), .B0(
        prevRequesterAddress_B[1]), .B1(n796), .Y(n797) );
  OAI2BB2XLTS U1020 ( .B0(n780), .B1(n797), .A0N(requesterAddressOut_EAST[1]), 
        .A1N(n800), .Y(n1165) );
  AOI22X1TS U1021 ( .A0(prevRequesterAddress_A[0]), .A1(n799), .B0(
        prevRequesterAddress_B[0]), .B1(n798), .Y(n801) );
  OAI2BB2XLTS U1022 ( .B0(n802), .B1(n801), .A0N(requesterAddressOut_EAST[0]), 
        .A1N(n800), .Y(n1164) );
  AOI22X1TS U1023 ( .A0(n803), .A1(n805), .B0(prevRequesterAddress_B[3]), .B1(
        n811), .Y(n807) );
  NOR3XLTS U1024 ( .A(n806), .B(n805), .C(n804), .Y(n818) );
  OAI2BB2XLTS U1025 ( .B0(n814), .B1(n807), .A0N(requesterAddressOut_SOUTH[3]), 
        .A1N(n818), .Y(n1163) );
  AOI22X1TS U1026 ( .A0(n809), .A1(n808), .B0(prevRequesterAddress_B[2]), .B1(
        n815), .Y(n810) );
  OAI2BB2XLTS U1027 ( .B0(n814), .B1(n810), .A0N(requesterAddressOut_SOUTH[2]), 
        .A1N(n818), .Y(n1162) );
  AOI22X1TS U1028 ( .A0(n812), .A1(n28), .B0(prevRequesterAddress_B[1]), .B1(
        n811), .Y(n813) );
  OAI2BB2XLTS U1029 ( .B0(n814), .B1(n813), .A0N(requesterAddressOut_SOUTH[1]), 
        .A1N(n818), .Y(n1161) );
  AOI22X1TS U1030 ( .A0(n817), .A1(n816), .B0(prevRequesterAddress_B[0]), .B1(
        n815), .Y(n819) );
  OAI2BB2XLTS U1031 ( .B0(n780), .B1(n819), .A0N(requesterAddressOut_SOUTH[0]), 
        .A1N(n818), .Y(n1160) );
endmodule


module outputPortArbiter_0 ( clk, reset, selectBit_NORTH, 
        destinationAddressIn_NORTH, requesterAddressIn_NORTH, readIn_NORTH, 
        writeIn_NORTH, dataIn_NORTH, selectBit_SOUTH, 
        destinationAddressIn_SOUTH, requesterAddressIn_SOUTH, readIn_SOUTH, 
        writeIn_SOUTH, dataIn_SOUTH, selectBit_EAST, destinationAddressIn_EAST, 
        requesterAddressIn_EAST, readIn_EAST, writeIn_EAST, dataIn_EAST, 
        selectBit_WEST, destinationAddressIn_WEST, requesterAddressIn_WEST, 
        readIn_WEST, writeIn_WEST, dataIn_WEST, readReady, 
        readRequesterAddress, cacheDataOut, destinationAddressOut, 
        requesterAddressOut, readOut, writeOut, dataOut );
  input [11:0] destinationAddressIn_NORTH;
  input [3:0] requesterAddressIn_NORTH;
  input [5:0] dataIn_NORTH;
  input [11:0] destinationAddressIn_SOUTH;
  input [3:0] requesterAddressIn_SOUTH;
  input [5:0] dataIn_SOUTH;
  input [11:0] destinationAddressIn_EAST;
  input [3:0] requesterAddressIn_EAST;
  input [5:0] dataIn_EAST;
  input [11:0] destinationAddressIn_WEST;
  input [3:0] requesterAddressIn_WEST;
  input [5:0] dataIn_WEST;
  input [3:0] readRequesterAddress;
  input [5:0] cacheDataOut;
  output [11:0] destinationAddressOut;
  output [3:0] requesterAddressOut;
  output [5:0] dataOut;
  input clk, reset, selectBit_NORTH, readIn_NORTH, writeIn_NORTH,
         selectBit_SOUTH, readIn_SOUTH, writeIn_SOUTH, selectBit_EAST,
         readIn_EAST, writeIn_EAST, selectBit_WEST, readIn_WEST, writeIn_WEST,
         readReady;
  output readOut, writeOut;
  wire   \requesterAddressbuffer[0][3] , \requesterAddressbuffer[0][2] ,
         \requesterAddressbuffer[0][1] , \requesterAddressbuffer[0][0] ,
         \requesterAddressbuffer[1][3] , \requesterAddressbuffer[1][2] ,
         \requesterAddressbuffer[1][1] , \requesterAddressbuffer[1][0] ,
         \requesterAddressbuffer[2][3] , \requesterAddressbuffer[2][2] ,
         \requesterAddressbuffer[2][1] , \requesterAddressbuffer[2][0] ,
         \requesterAddressbuffer[3][3] , \requesterAddressbuffer[3][2] ,
         \requesterAddressbuffer[3][1] , \requesterAddressbuffer[3][0] ,
         \requesterAddressbuffer[4][3] , \requesterAddressbuffer[4][2] ,
         \requesterAddressbuffer[4][1] , \requesterAddressbuffer[4][0] ,
         \requesterAddressbuffer[5][3] , \requesterAddressbuffer[5][2] ,
         \requesterAddressbuffer[5][1] , \requesterAddressbuffer[5][0] ,
         \requesterAddressbuffer[6][3] , \requesterAddressbuffer[6][2] ,
         \requesterAddressbuffer[6][1] , \requesterAddressbuffer[6][0] ,
         \requesterAddressbuffer[7][3] , \requesterAddressbuffer[7][2] ,
         \requesterAddressbuffer[7][1] , \requesterAddressbuffer[7][0] ,
         \destinationAddressbuffer[0][11] , \destinationAddressbuffer[0][10] ,
         \destinationAddressbuffer[0][9] , \destinationAddressbuffer[0][8] ,
         \destinationAddressbuffer[0][7] , \destinationAddressbuffer[0][6] ,
         \destinationAddressbuffer[0][5] , \destinationAddressbuffer[0][4] ,
         \destinationAddressbuffer[0][3] , \destinationAddressbuffer[0][2] ,
         \destinationAddressbuffer[0][1] , \destinationAddressbuffer[0][0] ,
         \destinationAddressbuffer[1][11] , \destinationAddressbuffer[1][10] ,
         \destinationAddressbuffer[1][9] , \destinationAddressbuffer[1][8] ,
         \destinationAddressbuffer[1][7] , \destinationAddressbuffer[1][6] ,
         \destinationAddressbuffer[1][5] , \destinationAddressbuffer[1][4] ,
         \destinationAddressbuffer[1][3] , \destinationAddressbuffer[1][2] ,
         \destinationAddressbuffer[1][1] , \destinationAddressbuffer[1][0] ,
         \destinationAddressbuffer[2][11] , \destinationAddressbuffer[2][10] ,
         \destinationAddressbuffer[2][9] , \destinationAddressbuffer[2][8] ,
         \destinationAddressbuffer[2][7] , \destinationAddressbuffer[2][6] ,
         \destinationAddressbuffer[2][5] , \destinationAddressbuffer[2][4] ,
         \destinationAddressbuffer[2][3] , \destinationAddressbuffer[2][2] ,
         \destinationAddressbuffer[2][1] , \destinationAddressbuffer[2][0] ,
         \destinationAddressbuffer[3][11] , \destinationAddressbuffer[3][10] ,
         \destinationAddressbuffer[3][9] , \destinationAddressbuffer[3][8] ,
         \destinationAddressbuffer[3][7] , \destinationAddressbuffer[3][6] ,
         \destinationAddressbuffer[3][5] , \destinationAddressbuffer[3][4] ,
         \destinationAddressbuffer[3][3] , \destinationAddressbuffer[3][2] ,
         \destinationAddressbuffer[3][1] , \destinationAddressbuffer[3][0] ,
         \destinationAddressbuffer[4][11] , \destinationAddressbuffer[4][10] ,
         \destinationAddressbuffer[4][9] , \destinationAddressbuffer[4][8] ,
         \destinationAddressbuffer[4][7] , \destinationAddressbuffer[4][6] ,
         \destinationAddressbuffer[4][5] , \destinationAddressbuffer[4][4] ,
         \destinationAddressbuffer[4][3] , \destinationAddressbuffer[4][2] ,
         \destinationAddressbuffer[4][1] , \destinationAddressbuffer[4][0] ,
         \destinationAddressbuffer[5][11] , \destinationAddressbuffer[5][10] ,
         \destinationAddressbuffer[5][9] , \destinationAddressbuffer[5][8] ,
         \destinationAddressbuffer[5][7] , \destinationAddressbuffer[5][6] ,
         \destinationAddressbuffer[5][5] , \destinationAddressbuffer[5][4] ,
         \destinationAddressbuffer[5][3] , \destinationAddressbuffer[5][2] ,
         \destinationAddressbuffer[5][1] , \destinationAddressbuffer[5][0] ,
         \destinationAddressbuffer[6][11] , \destinationAddressbuffer[6][10] ,
         \destinationAddressbuffer[6][9] , \destinationAddressbuffer[6][8] ,
         \destinationAddressbuffer[6][7] , \destinationAddressbuffer[6][6] ,
         \destinationAddressbuffer[6][5] , \destinationAddressbuffer[6][4] ,
         \destinationAddressbuffer[6][3] , \destinationAddressbuffer[6][2] ,
         \destinationAddressbuffer[6][1] , \destinationAddressbuffer[6][0] ,
         \destinationAddressbuffer[7][11] , \destinationAddressbuffer[7][10] ,
         \destinationAddressbuffer[7][9] , \destinationAddressbuffer[7][8] ,
         \destinationAddressbuffer[7][7] , \destinationAddressbuffer[7][6] ,
         \destinationAddressbuffer[7][5] , \destinationAddressbuffer[7][4] ,
         \destinationAddressbuffer[7][3] , \destinationAddressbuffer[7][2] ,
         \destinationAddressbuffer[7][1] , \destinationAddressbuffer[7][0] ,
         \dataoutbuffer[7][5] , \dataoutbuffer[7][4] , \dataoutbuffer[7][3] ,
         \dataoutbuffer[7][2] , \dataoutbuffer[7][1] , \dataoutbuffer[7][0] ,
         \dataoutbuffer[6][5] , \dataoutbuffer[6][4] , \dataoutbuffer[6][3] ,
         \dataoutbuffer[6][2] , \dataoutbuffer[6][1] , \dataoutbuffer[6][0] ,
         \dataoutbuffer[5][5] , \dataoutbuffer[5][4] , \dataoutbuffer[5][3] ,
         \dataoutbuffer[5][2] , \dataoutbuffer[5][1] , \dataoutbuffer[5][0] ,
         \dataoutbuffer[4][5] , \dataoutbuffer[4][4] , \dataoutbuffer[4][3] ,
         \dataoutbuffer[4][2] , \dataoutbuffer[4][1] , \dataoutbuffer[4][0] ,
         \dataoutbuffer[3][5] , \dataoutbuffer[3][4] , \dataoutbuffer[3][3] ,
         \dataoutbuffer[3][2] , \dataoutbuffer[3][1] , \dataoutbuffer[3][0] ,
         \dataoutbuffer[2][5] , \dataoutbuffer[2][4] , \dataoutbuffer[2][3] ,
         \dataoutbuffer[2][2] , \dataoutbuffer[2][1] , \dataoutbuffer[2][0] ,
         \dataoutbuffer[1][5] , \dataoutbuffer[1][4] , \dataoutbuffer[1][3] ,
         \dataoutbuffer[1][2] , \dataoutbuffer[1][1] , \dataoutbuffer[1][0] ,
         \dataoutbuffer[0][5] , \dataoutbuffer[0][4] , \dataoutbuffer[0][3] ,
         \dataoutbuffer[0][2] , \dataoutbuffer[0][1] , \dataoutbuffer[0][0] ,
         N2624, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
         n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
         n1967, n1968, n1969, n1970, n1971;
  wire   [0:7] writeOutbuffer;
  wire   [0:7] readOutbuffer;

  DFFNSRX1TS full_reg_reg ( .D(N2624), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(
        n1963) );
  DFFNSRX1TS \requesterAddressbuffer_reg[2][0]  ( .D(n1285), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[2][1]  ( .D(n1284), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[2][2]  ( .D(n1283), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[2][3]  ( .D(n1282), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][0]  ( .D(n1149), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][1]  ( .D(n1148), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][2]  ( .D(n1147), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][3]  ( .D(n1146), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][0]  ( .D(n1273), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][1]  ( .D(n1272), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][2]  ( .D(n1271), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][3]  ( .D(n1270), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][4]  ( .D(n1269), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][5]  ( .D(n1268), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][5] ) );
  DFFNSRX1TS \writeOutbuffer_reg[7]  ( .D(n1225), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[7]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][4]  ( .D(n1205), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][5]  ( .D(n1204), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][6]  ( .D(n1203), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][7]  ( .D(n1202), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][8]  ( .D(n1201), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][9]  ( .D(n1200), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][11]  ( .D(n1198), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[6]  ( .D(n1224), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[6]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][4]  ( .D(n1193), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][5]  ( .D(n1192), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][6]  ( .D(n1191), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][7]  ( .D(n1190), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][8]  ( .D(n1189), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][9]  ( .D(n1188), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][10]  ( .D(n1187), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][11]  ( .D(n1186), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[3]  ( .D(n1221), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[3]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][4]  ( .D(n1157), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][5]  ( .D(n1156), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][6]  ( .D(n1155), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][7]  ( .D(n1154), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][8]  ( .D(n1153), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][9]  ( .D(n1152), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][10]  ( .D(n1151), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][11]  ( .D(n1150), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[2]  ( .D(n1220), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[2]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][4]  ( .D(n1145), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][5]  ( .D(n1144), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][6]  ( .D(n1143), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][7]  ( .D(n1142), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][8]  ( .D(n1141), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][9]  ( .D(n1140), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][10]  ( .D(n1139), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][11]  ( .D(n1138), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][11] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][0]  ( .D(n1231), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][1]  ( .D(n1230), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][2]  ( .D(n1229), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][3]  ( .D(n1228), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][4]  ( .D(n1227), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][5]  ( .D(n1226), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][0]  ( .D(n1237), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][1]  ( .D(n1236), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][2]  ( .D(n1235), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][3]  ( .D(n1234), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][4]  ( .D(n1233), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][5]  ( .D(n1232), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][5] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[5][0]  ( .D(n1297), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[5][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[5][1]  ( .D(n1296), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[5][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[5][2]  ( .D(n1295), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[5][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[5][3]  ( .D(n1294), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[5][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][0]  ( .D(n1185), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][1]  ( .D(n1184), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][2]  ( .D(n1183), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][3]  ( .D(n1182), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[4][0]  ( .D(n1293), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[4][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[4][1]  ( .D(n1292), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[4][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[4][2]  ( .D(n1291), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[4][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[4][3]  ( .D(n1290), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[4][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][0]  ( .D(n1173), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][1]  ( .D(n1172), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][2]  ( .D(n1171), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][3]  ( .D(n1170), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][0]  ( .D(n1255), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][1]  ( .D(n1254), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][2]  ( .D(n1253), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][3]  ( .D(n1252), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][4]  ( .D(n1251), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][5]  ( .D(n1250), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][0]  ( .D(n1261), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][1]  ( .D(n1260), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][2]  ( .D(n1259), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][3]  ( .D(n1258), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][4]  ( .D(n1257), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][5]  ( .D(n1256), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][5] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[1][0]  ( .D(n1281), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[1][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[1][1]  ( .D(n1280), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[1][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[1][2]  ( .D(n1279), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[1][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[1][3]  ( .D(n1278), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[1][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][0]  ( .D(n1137), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][1]  ( .D(n1136), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][2]  ( .D(n1135), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][3]  ( .D(n1134), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[0][0]  ( .D(n1277), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[0][1]  ( .D(n1276), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[0][2]  ( .D(n1275), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[0][3]  ( .D(n1274), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][0]  ( .D(n1125), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][1]  ( .D(n1124), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][2]  ( .D(n1123), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][3]  ( .D(n1122), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[7][0]  ( .D(n1305), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[7][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[7][1]  ( .D(n1304), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[7][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[7][2]  ( .D(n1303), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[7][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[7][3]  ( .D(n1302), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[7][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][0]  ( .D(n1209), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][1]  ( .D(n1208), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][2]  ( .D(n1207), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][3]  ( .D(n1206), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[6][0]  ( .D(n1301), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[6][1]  ( .D(n1300), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[6][2]  ( .D(n1299), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[6][3]  ( .D(n1298), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][0]  ( .D(n1197), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][1]  ( .D(n1196), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][2]  ( .D(n1195), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][3]  ( .D(n1194), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][0]  ( .D(n1243), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][1]  ( .D(n1242), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][2]  ( .D(n1241), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][3]  ( .D(n1240), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][4]  ( .D(n1239), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][5]  ( .D(n1238), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][0]  ( .D(n1249), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][1]  ( .D(n1248), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][2]  ( .D(n1247), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][3]  ( .D(n1246), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][4]  ( .D(n1245), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][5]  ( .D(n1244), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][5] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[3][0]  ( .D(n1289), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[3][1]  ( .D(n1288), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[3][2]  ( .D(n1287), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[3][3]  ( .D(n1286), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][0]  ( .D(n1161), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][1]  ( .D(n1160), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][2]  ( .D(n1159), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][3]  ( .D(n1158), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][0]  ( .D(n1267), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][1]  ( .D(n1266), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][2]  ( .D(n1265), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][3]  ( .D(n1264), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][4]  ( .D(n1263), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][5]  ( .D(n1262), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][5] ) );
  DFFNSRX1TS \writeOutbuffer_reg[5]  ( .D(n1223), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[5]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][4]  ( .D(n1181), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][5]  ( .D(n1180), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][6]  ( .D(n1179), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][7]  ( .D(n1178), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][8]  ( .D(n1177), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][9]  ( .D(n1176), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][10]  ( .D(n1175), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][11]  ( .D(n1174), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[4]  ( .D(n1222), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[4]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][4]  ( .D(n1169), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][5]  ( .D(n1168), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][6]  ( .D(n1167), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][7]  ( .D(n1166), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][8]  ( .D(n1165), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][9]  ( .D(n1164), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][10]  ( .D(n1163), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][11]  ( .D(n1162), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[1]  ( .D(n1219), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[1]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][4]  ( .D(n1133), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][5]  ( .D(n1132), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][6]  ( .D(n1131), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][7]  ( .D(n1130), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][8]  ( .D(n1129), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][9]  ( .D(n1128), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][10]  ( .D(n1127), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][11]  ( .D(n1126), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[0]  ( .D(n1218), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[0]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][4]  ( .D(n1121), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][5]  ( .D(n1120), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][6]  ( .D(n1119), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][7]  ( .D(n1118), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][8]  ( .D(n1117), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][9]  ( .D(n1116), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][10]  ( .D(n1115), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][11]  ( .D(n1114), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][11] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][10]  ( .D(n1199), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][10] ) );
  DFFNSRX1TS writeOut_reg ( .D(n1328), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        writeOut) );
  DFFNSRX1TS \destinationAddressOut_reg[4]  ( .D(n1319), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[4]) );
  DFFNSRX1TS \destinationAddressOut_reg[5]  ( .D(n1318), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[5]) );
  DFFNSRX1TS \destinationAddressOut_reg[6]  ( .D(n1317), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[6]) );
  DFFNSRX1TS \destinationAddressOut_reg[7]  ( .D(n1316), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[7]) );
  DFFNSRX1TS \destinationAddressOut_reg[8]  ( .D(n1315), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[8]) );
  DFFNSRX1TS \destinationAddressOut_reg[9]  ( .D(n1314), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[9]) );
  DFFNSRX1TS \destinationAddressOut_reg[10]  ( .D(n1313), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[10]) );
  DFFNSRX1TS \destinationAddressOut_reg[11]  ( .D(n1312), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[11]) );
  DFFNSRX1TS readOut_reg ( .D(n1329), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        readOut) );
  DFFNSRX1TS \requesterAddressOut_reg[0]  ( .D(n1327), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[0]) );
  DFFNSRX1TS \requesterAddressOut_reg[1]  ( .D(n1326), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[1]) );
  DFFNSRX1TS \requesterAddressOut_reg[2]  ( .D(n1325), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[2]) );
  DFFNSRX1TS \requesterAddressOut_reg[3]  ( .D(n1324), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[3]) );
  DFFNSRX1TS \destinationAddressOut_reg[0]  ( .D(n1323), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[0]) );
  DFFNSRX1TS \destinationAddressOut_reg[1]  ( .D(n1322), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[1]) );
  DFFNSRX1TS \destinationAddressOut_reg[2]  ( .D(n1321), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[2]) );
  DFFNSRX1TS \destinationAddressOut_reg[3]  ( .D(n1320), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[3]) );
  DFFNSRX1TS \dataOut_reg[0]  ( .D(n1311), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[0]) );
  DFFNSRX1TS \dataOut_reg[1]  ( .D(n1310), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[1]) );
  DFFNSRX1TS \dataOut_reg[2]  ( .D(n1309), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[2]) );
  DFFNSRX1TS \dataOut_reg[3]  ( .D(n1308), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[3]) );
  DFFNSRX1TS \dataOut_reg[4]  ( .D(n1307), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[4]) );
  DFFNSRX1TS \dataOut_reg[5]  ( .D(n1306), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[5]) );
  DFFNSRX1TS \read_reg_reg[1]  ( .D(n1330), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1956), .QN(n1955) );
  DFFNSRX1TS \write_reg_reg[0]  ( .D(n1335), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1954), .QN(n1958) );
  DFFNSRX1TS \write_reg_reg[2]  ( .D(n1333), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1959), .QN(n1960) );
  DFFNSRX1TS \read_reg_reg[0]  ( .D(n1336), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1949), .QN(n1961) );
  DFFNSRX1TS \read_reg_reg[2]  ( .D(n1331), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1952), .QN(n1953) );
  DFFNSRX1TS empty_reg_reg ( .D(n1332), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        n1951), .QN(n1950) );
  DFFNSRX1TS \readOutbuffer_reg[7]  ( .D(n1217), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[7]), .QN(n1964) );
  DFFNSRX1TS \readOutbuffer_reg[4]  ( .D(n1214), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[4]), .QN(n1967) );
  DFFNSRX1TS \readOutbuffer_reg[6]  ( .D(n1216), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[6]), .QN(n1965) );
  DFFNSRX1TS \readOutbuffer_reg[5]  ( .D(n1215), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[5]), .QN(n1966) );
  DFFNSRX1TS \readOutbuffer_reg[1]  ( .D(n1211), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[1]), .QN(n1970) );
  DFFNSRX1TS \readOutbuffer_reg[2]  ( .D(n1212), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[2]), .QN(n1969) );
  DFFNSRX1TS \readOutbuffer_reg[0]  ( .D(n1210), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[0]), .QN(n1971) );
  DFFNSRX1TS \readOutbuffer_reg[3]  ( .D(n1213), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[3]), .QN(n1968) );
  DFFNSRX1TS \write_reg_reg[1]  ( .D(n1334), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1957), .QN(n1962) );
  CMPR32X2TS U3 ( .A(n488), .B(n487), .C(n486), .CO(n481), .S(n496) );
  CLKBUFX2TS U4 ( .A(n14), .Y(n79) );
  CMPR32X2TS U5 ( .A(n466), .B(n497), .C(n16), .CO(n17), .S(n14) );
  CMPR32X2TS U6 ( .A(n532), .B(n464), .C(n463), .CO(n455), .S(n469) );
  CMPR32X2TS U7 ( .A(n462), .B(n516), .C(n461), .CO(n465), .S(n478) );
  NOR2X1TS U8 ( .A(n460), .B(n506), .Y(n18) );
  INVX2TS U9 ( .A(selectBit_NORTH), .Y(n506) );
  CLKBUFX2TS U10 ( .A(n20), .Y(n81) );
  NOR2XLTS U11 ( .A(n1613), .B(n279), .Y(n292) );
  NOR2XLTS U12 ( .A(n1578), .B(n38), .Y(n43) );
  ADDHXLTS U13 ( .A(n448), .B(n461), .CO(n16), .S(n15) );
  INVX2TS U14 ( .A(n1617), .Y(n1615) );
  INVX2TS U15 ( .A(n1593), .Y(n1591) );
  INVX2TS U16 ( .A(n1582), .Y(n1580) );
  INVX2TS U17 ( .A(n1656), .Y(n1653) );
  INVX2TS U18 ( .A(n1621), .Y(n1618) );
  NOR2XLTS U19 ( .A(selectBit_NORTH), .B(n507), .Y(n540) );
  NOR2XLTS U20 ( .A(n1646), .B(n325), .Y(n326) );
  NOR2XLTS U21 ( .A(n1628), .B(n134), .Y(n135) );
  NOR2XLTS U22 ( .A(n318), .B(n1657), .Y(n319) );
  NOR2XLTS U23 ( .A(n318), .B(n1631), .Y(n131) );
  NOR2XLTS U24 ( .A(n452), .B(n1610), .Y(n225) );
  NOR2XLTS U25 ( .A(n1586), .B(n30), .Y(n34) );
  NOR2XLTS U26 ( .A(n1634), .B(n189), .Y(n190) );
  NOR2X1TS U27 ( .A(n1635), .B(n189), .Y(n193) );
  NOR2X1TS U28 ( .A(n1590), .B(n90), .Y(n102) );
  NAND2BXLTS U29 ( .AN(n323), .B(n322), .Y(n325) );
  NAND2BXLTS U30 ( .AN(n399), .B(n398), .Y(n400) );
  NAND2BXLTS U31 ( .AN(n278), .B(n277), .Y(n279) );
  NAND2BXLTS U32 ( .AN(n89), .B(n88), .Y(n90) );
  NAND2BXLTS U33 ( .AN(n188), .B(n187), .Y(n189) );
  NOR2X1TS U34 ( .A(n125), .B(n386), .Y(n1627) );
  NAND2BX1TS U35 ( .AN(n124), .B(selectBit_EAST), .Y(n386) );
  NAND2X1TS U36 ( .A(n512), .B(n124), .Y(n270) );
  NAND3X1TS U37 ( .A(n83), .B(n29), .C(n222), .Y(n1578) );
  NAND3X1TS U38 ( .A(n29), .B(n222), .C(n271), .Y(n1600) );
  NOR2X1TS U39 ( .A(n222), .B(n80), .Y(n314) );
  INVX1TS U40 ( .A(n1642), .Y(n1640) );
  INVX1TS U41 ( .A(n1596), .Y(n1594) );
  INVX1TS U42 ( .A(n1670), .Y(n1667) );
  NOR2X1TS U43 ( .A(n8), .B(n80), .Y(n28) );
  AND2X2TS U44 ( .A(n525), .B(n1963), .Y(n130) );
  BUFX3TS U45 ( .A(n18), .Y(n19) );
  CLKBUFX2TS U46 ( .A(n55), .Y(n295) );
  CLKBUFX2TS U47 ( .A(readIn_EAST), .Y(n1577) );
  INVX1TS U48 ( .A(n1960), .Y(n482) );
  NAND2BX1TS U49 ( .AN(n123), .B(n462), .Y(n384) );
  OAI21X2TS U50 ( .A0(n28), .A1(n25), .B0(n27), .Y(n124) );
  NOR2XLTS U51 ( .A(n1609), .B(n1606), .Y(n228) );
  NOR3BXLTS U52 ( .AN(n514), .B(n513), .C(n512), .Y(n539) );
  NAND2BXLTS U53 ( .AN(n134), .B(n128), .Y(n133) );
  NAND2X1TS U54 ( .A(n132), .B(n1631), .Y(n134) );
  OR2X1TS U55 ( .A(n276), .B(n930), .Y(n1425) );
  OR2X1TS U56 ( .A(n226), .B(n913), .Y(n1456) );
  OR2X1TS U57 ( .A(n185), .B(n978), .Y(n1357) );
  OR2X1TS U58 ( .A(n132), .B(n956), .Y(n1392) );
  OR2X1TS U59 ( .A(n86), .B(n895), .Y(n1493) );
  OR2X1TS U60 ( .A(n35), .B(n1673), .Y(n1542) );
  XOR2X1TS U61 ( .A(n484), .B(n483), .Y(n498) );
  XNOR2X1TS U62 ( .A(n482), .B(n481), .Y(n483) );
  NAND4XLTS U63 ( .A(n458), .B(n1954), .C(readReady), .D(n444), .Y(n1631) );
  INVX2TS U64 ( .A(n1630), .Y(n1628) );
  CLKBUFX2TS U65 ( .A(n1392), .Y(n1632) );
  NOR3XLTS U66 ( .A(n79), .B(n122), .C(n384), .Y(n1670) );
  INVX2TS U67 ( .A(n1666), .Y(n1663) );
  NOR3XLTS U68 ( .A(n15), .B(n181), .C(n384), .Y(n1642) );
  INVX2TS U69 ( .A(n1639), .Y(n1636) );
  CLKBUFX2TS U70 ( .A(n1357), .Y(n1644) );
  NAND4XLTS U71 ( .A(n449), .B(readReady), .C(n446), .D(n392), .Y(n1657) );
  NOR3XLTS U72 ( .A(n79), .B(n78), .C(n384), .Y(n1656) );
  INVX2TS U73 ( .A(n1652), .Y(n1650) );
  NAND4XLTS U74 ( .A(n448), .B(n273), .C(readReady), .D(n389), .Y(n1610) );
  NOR3X1TS U75 ( .A(n14), .B(n78), .C(n268), .Y(n1609) );
  CLKBUFX2TS U76 ( .A(n1456), .Y(n1611) );
  NOR3XLTS U77 ( .A(n15), .B(n181), .C(n268), .Y(n1596) );
  CLKBUFX2TS U78 ( .A(n1493), .Y(n1598) );
  NOR3XLTS U79 ( .A(n79), .B(n15), .C(n268), .Y(n1621) );
  CLKBUFX2TS U80 ( .A(n1425), .Y(n1623) );
  NAND4XLTS U81 ( .A(n449), .B(n497), .C(n273), .D(n514), .Y(n1586) );
  CLKBUFX2TS U82 ( .A(n1542), .Y(n1587) );
  NAND3XLTS U83 ( .A(n540), .B(n1951), .C(n539), .Y(n561) );
  CLKAND2X2TS U84 ( .A(n525), .B(n523), .Y(n552) );
  CLKAND2X2TS U85 ( .A(n480), .B(n478), .Y(n485) );
  NOR2XLTS U86 ( .A(n1621), .B(n1617), .Y(n277) );
  NOR2XLTS U87 ( .A(n1596), .B(n1593), .Y(n88) );
  NOR2XLTS U88 ( .A(n1585), .B(n1582), .Y(n36) );
  NOR2XLTS U89 ( .A(n1670), .B(n1666), .Y(n398) );
  AO21X1TS U90 ( .A0(n460), .A1(n506), .B0(n19), .Y(n21) );
  NAND3XLTS U91 ( .A(selectBit_NORTH), .B(n509), .C(n508), .Y(n520) );
  NAND3XLTS U92 ( .A(n507), .B(n509), .C(n506), .Y(n519) );
  NOR2XLTS U93 ( .A(n1656), .B(n1652), .Y(n322) );
  NOR2XLTS U94 ( .A(n1630), .B(n1627), .Y(n128) );
  NAND2BXLTS U95 ( .AN(n229), .B(n228), .Y(n230) );
  NAND3XLTS U96 ( .A(n19), .B(n482), .C(n392), .Y(n223) );
  NAND2BXLTS U97 ( .AN(n37), .B(n36), .Y(n38) );
  XOR2XLTS U98 ( .A(n455), .B(n457), .Y(n475) );
  OAI21XLTS U99 ( .A0(n458), .A1(n1955), .B0(n457), .Y(n459) );
  INVX2TS U100 ( .A(n7), .Y(n271) );
  INVX2TS U101 ( .A(n271), .Y(n388) );
  XOR2X1TS U102 ( .A(n482), .B(n17), .Y(n123) );
  CLKAND2X2TS U103 ( .A(n480), .B(n479), .Y(n486) );
  NOR2XLTS U104 ( .A(n85), .B(reset), .Y(n500) );
  NOR3X1TS U105 ( .A(n181), .B(n78), .C(n384), .Y(n1630) );
  INVX2TS U106 ( .A(n1627), .Y(n1625) );
  NAND4XLTS U107 ( .A(n511), .B(n393), .C(n392), .D(n444), .Y(n1671) );
  NOR3XLTS U108 ( .A(n24), .B(n388), .C(n20), .Y(n1662) );
  INVX2TS U109 ( .A(n1662), .Y(n1659) );
  NOR3BXLTS U110 ( .AN(n387), .B(n386), .C(n385), .Y(n1666) );
  NAND4XLTS U111 ( .A(n487), .B(n511), .C(n393), .D(n446), .Y(n1643) );
  NOR3XLTS U112 ( .A(n29), .B(n81), .C(n271), .Y(n1635) );
  INVX2TS U113 ( .A(n1635), .Y(n1634) );
  NOR3XLTS U114 ( .A(n29), .B(n388), .C(n8), .Y(n1649) );
  INVX2TS U115 ( .A(n1649), .Y(n1646) );
  NOR3XLTS U116 ( .A(n315), .B(n314), .C(n386), .Y(n1652) );
  INVX2TS U117 ( .A(n1609), .Y(n1607) );
  NOR3XLTS U118 ( .A(n315), .B(n314), .C(n270), .Y(n1606) );
  NAND4XLTS U119 ( .A(n83), .B(n454), .C(n514), .D(n393), .Y(n1597) );
  INVX2TS U120 ( .A(n1590), .Y(n1589) );
  NAND4XLTS U121 ( .A(n273), .B(n511), .C(n393), .D(n389), .Y(n1622) );
  NOR3XLTS U122 ( .A(n388), .B(n20), .C(n23), .Y(n1614) );
  INVX2TS U123 ( .A(n1614), .Y(n1613) );
  NOR3BXLTS U124 ( .AN(n387), .B(n270), .C(n269), .Y(n1617) );
  NAND4XLTS U125 ( .A(n14), .B(n122), .C(n123), .D(n462), .Y(n1583) );
  INVX2TS U126 ( .A(n1578), .Y(n1579) );
  NOR2XLTS U127 ( .A(n125), .B(n270), .Y(n1582) );
  INVX2TS U128 ( .A(destinationAddressIn_SOUTH[11]), .Y(n142) );
  INVX2TS U129 ( .A(destinationAddressIn_SOUTH[10]), .Y(n138) );
  INVX2TS U130 ( .A(destinationAddressIn_SOUTH[9]), .Y(n151) );
  INVX2TS U131 ( .A(destinationAddressIn_SOUTH[8]), .Y(n146) );
  AO22XLTS U132 ( .A0(n1959), .A1(n500), .B0(n499), .B1(n498), .Y(n1333) );
  AO22XLTS U133 ( .A0(n1954), .A1(n500), .B0(n499), .B1(n495), .Y(n1335) );
  AO22XLTS U134 ( .A0(n497), .A1(n500), .B0(n499), .B1(n496), .Y(n1334) );
  OAI21XLTS U135 ( .A0(n85), .A1(n451), .B0(n494), .Y(n1332) );
  NAND4XLTS U136 ( .A(n874), .B(n873), .C(n872), .D(n871), .Y(n1306) );
  NAND4XLTS U137 ( .A(n850), .B(n849), .C(n848), .D(n847), .Y(n1307) );
  NAND4XLTS U138 ( .A(n838), .B(n837), .C(n836), .D(n835), .Y(n1308) );
  NAND4XLTS U139 ( .A(n826), .B(n825), .C(n824), .D(n823), .Y(n1309) );
  NAND4XLTS U140 ( .A(n807), .B(n806), .C(n805), .D(n804), .Y(n1310) );
  NAND4XLTS U141 ( .A(n787), .B(n786), .C(n785), .D(n784), .Y(n1311) );
  NAND4XLTS U142 ( .A(n658), .B(n657), .C(n656), .D(n655), .Y(n1320) );
  NAND4XLTS U143 ( .A(n646), .B(n645), .C(n644), .D(n643), .Y(n1321) );
  NAND4XLTS U144 ( .A(n626), .B(n625), .C(n624), .D(n623), .Y(n1322) );
  NAND4XLTS U145 ( .A(n611), .B(n610), .C(n609), .D(n608), .Y(n1323) );
  NAND4XLTS U146 ( .A(n600), .B(n599), .C(n598), .D(n655), .Y(n1324) );
  NAND4XLTS U147 ( .A(n589), .B(n588), .C(n587), .D(n643), .Y(n1325) );
  NAND4XLTS U148 ( .A(n581), .B(n580), .C(n579), .D(n623), .Y(n1326) );
  NAND4XLTS U149 ( .A(n564), .B(n563), .C(n562), .D(n608), .Y(n1327) );
  NAND4XLTS U150 ( .A(n543), .B(n542), .C(n541), .D(n561), .Y(n1329) );
  NAND3XLTS U151 ( .A(n777), .B(n776), .C(n775), .Y(n1312) );
  NAND3XLTS U152 ( .A(n763), .B(n762), .C(n761), .Y(n1313) );
  NAND3XLTS U153 ( .A(n748), .B(n747), .C(n746), .Y(n1314) );
  NAND3XLTS U154 ( .A(n730), .B(n729), .C(n728), .Y(n1315) );
  NAND3XLTS U155 ( .A(n716), .B(n715), .C(n714), .Y(n1316) );
  NAND3XLTS U156 ( .A(n705), .B(n704), .C(n703), .Y(n1317) );
  NAND3XLTS U157 ( .A(n690), .B(n689), .C(n688), .Y(n1318) );
  NAND3XLTS U158 ( .A(n669), .B(n668), .C(n667), .Y(n1319) );
  NAND3XLTS U159 ( .A(n555), .B(n554), .C(n553), .Y(n1328) );
  NAND3XLTS U160 ( .A(n1345), .B(n1344), .C(n1343), .Y(n1262) );
  NAND3XLTS U161 ( .A(n1339), .B(n1338), .C(n1337), .Y(n1263) );
  NAND3XLTS U162 ( .A(n1110), .B(n1109), .C(n1108), .Y(n1264) );
  NAND3XLTS U163 ( .A(n1105), .B(n1104), .C(n1103), .Y(n1265) );
  NAND3XLTS U164 ( .A(n1097), .B(n1096), .C(n1095), .Y(n1266) );
  NAND3XLTS U165 ( .A(n1091), .B(n1090), .C(n1089), .Y(n1267) );
  NAND3XLTS U166 ( .A(n1825), .B(n1824), .C(n1823), .Y(n1158) );
  NAND3XLTS U167 ( .A(n1815), .B(n1814), .C(n1813), .Y(n1159) );
  NAND3XLTS U168 ( .A(n1808), .B(n1807), .C(n1806), .Y(n1160) );
  NAND3XLTS U169 ( .A(n1800), .B(n1799), .C(n1798), .Y(n1161) );
  NAND3XLTS U170 ( .A(n973), .B(n972), .C(n971), .Y(n1286) );
  NAND3XLTS U171 ( .A(n968), .B(n967), .C(n966), .Y(n1287) );
  NAND3XLTS U172 ( .A(n961), .B(n960), .C(n959), .Y(n1288) );
  NAND3XLTS U173 ( .A(n954), .B(n953), .C(n952), .Y(n1289) );
  NAND3XLTS U174 ( .A(n1444), .B(n1443), .C(n1442), .Y(n1244) );
  NAND3XLTS U175 ( .A(n1439), .B(n1438), .C(n1437), .Y(n1245) );
  NAND3XLTS U176 ( .A(n1434), .B(n1433), .C(n1432), .Y(n1246) );
  NAND3XLTS U177 ( .A(n1430), .B(n1429), .C(n1428), .Y(n1247) );
  NAND3XLTS U178 ( .A(n1424), .B(n1423), .C(n1422), .Y(n1248) );
  NAND3XLTS U179 ( .A(n1417), .B(n1416), .C(n1415), .Y(n1249) );
  NAND3XLTS U180 ( .A(n1475), .B(n1474), .C(n1473), .Y(n1238) );
  NAND3XLTS U181 ( .A(n1471), .B(n1470), .C(n1469), .Y(n1239) );
  NAND3XLTS U182 ( .A(n1466), .B(n1465), .C(n1464), .Y(n1240) );
  NAND3XLTS U183 ( .A(n1461), .B(n1460), .C(n1459), .Y(n1241) );
  NAND3XLTS U184 ( .A(n1455), .B(n1454), .C(n1453), .Y(n1242) );
  NAND3XLTS U185 ( .A(n1449), .B(n1448), .C(n1447), .Y(n1243) );
  NAND3XLTS U186 ( .A(n1733), .B(n1732), .C(n1731), .Y(n1194) );
  NAND3XLTS U187 ( .A(n1724), .B(n1723), .C(n1722), .Y(n1195) );
  NAND3XLTS U188 ( .A(n1715), .B(n1714), .C(n1713), .Y(n1196) );
  NAND3XLTS U189 ( .A(n1706), .B(n1705), .C(n1704), .Y(n1197) );
  NAND3XLTS U190 ( .A(n908), .B(n907), .C(n906), .Y(n1298) );
  NAND3XLTS U191 ( .A(n904), .B(n903), .C(n902), .Y(n1299) );
  NAND3XLTS U192 ( .A(n900), .B(n899), .C(n898), .Y(n1300) );
  NAND3XLTS U193 ( .A(n894), .B(n893), .C(n892), .Y(n1301) );
  NAND3XLTS U194 ( .A(n1701), .B(n1700), .C(n1699), .Y(n1206) );
  NAND3XLTS U195 ( .A(n1693), .B(n1692), .C(n1691), .Y(n1207) );
  NAND3XLTS U196 ( .A(n1684), .B(n1683), .C(n1682), .Y(n1208) );
  NAND3XLTS U197 ( .A(n1676), .B(n1675), .C(n1674), .Y(n1209) );
  NAND3XLTS U198 ( .A(n891), .B(n890), .C(n889), .Y(n1302) );
  NAND3XLTS U199 ( .A(n885), .B(n884), .C(n883), .Y(n1303) );
  NAND3XLTS U200 ( .A(n882), .B(n881), .C(n880), .Y(n1304) );
  NAND3XLTS U201 ( .A(n878), .B(n877), .C(n876), .Y(n1305) );
  NAND3XLTS U202 ( .A(n1933), .B(n1932), .C(n1931), .Y(n1122) );
  NAND3XLTS U203 ( .A(n1922), .B(n1921), .C(n1920), .Y(n1123) );
  NAND3XLTS U204 ( .A(n1910), .B(n1909), .C(n1908), .Y(n1124) );
  NAND3XLTS U205 ( .A(n1899), .B(n1898), .C(n1897), .Y(n1125) );
  NAND3XLTS U206 ( .A(n1051), .B(n1050), .C(n1049), .Y(n1274) );
  NAND3XLTS U207 ( .A(n1042), .B(n1041), .C(n1040), .Y(n1275) );
  NAND3XLTS U208 ( .A(n1036), .B(n1035), .C(n1034), .Y(n1276) );
  NAND3XLTS U209 ( .A(n1029), .B(n1028), .C(n1027), .Y(n1277) );
  NAND3XLTS U210 ( .A(n1891), .B(n1890), .C(n1889), .Y(n1134) );
  NAND3XLTS U211 ( .A(n1881), .B(n1880), .C(n1879), .Y(n1135) );
  NAND3XLTS U212 ( .A(n1869), .B(n1868), .C(n1867), .Y(n1136) );
  NAND3XLTS U213 ( .A(n1859), .B(n1858), .C(n1857), .Y(n1137) );
  NAND3XLTS U214 ( .A(n1022), .B(n1021), .C(n1020), .Y(n1278) );
  NAND3XLTS U215 ( .A(n1013), .B(n1012), .C(n1011), .Y(n1279) );
  NAND3XLTS U216 ( .A(n1005), .B(n1004), .C(n1003), .Y(n1280) );
  NAND3XLTS U217 ( .A(n997), .B(n996), .C(n995), .Y(n1281) );
  NAND3XLTS U218 ( .A(n1381), .B(n1380), .C(n1379), .Y(n1256) );
  NAND3XLTS U219 ( .A(n1374), .B(n1373), .C(n1372), .Y(n1257) );
  NAND3XLTS U220 ( .A(n1367), .B(n1366), .C(n1365), .Y(n1258) );
  NAND3XLTS U221 ( .A(n1363), .B(n1362), .C(n1361), .Y(n1259) );
  NAND3XLTS U222 ( .A(n1356), .B(n1355), .C(n1354), .Y(n1260) );
  NAND3XLTS U223 ( .A(n1350), .B(n1349), .C(n1348), .Y(n1261) );
  NAND3XLTS U224 ( .A(n1412), .B(n1411), .C(n1410), .Y(n1250) );
  NAND3XLTS U225 ( .A(n1405), .B(n1404), .C(n1403), .Y(n1251) );
  NAND3XLTS U226 ( .A(n1400), .B(n1399), .C(n1398), .Y(n1252) );
  NAND3XLTS U227 ( .A(n1396), .B(n1395), .C(n1394), .Y(n1253) );
  NAND3XLTS U228 ( .A(n1391), .B(n1390), .C(n1389), .Y(n1254) );
  NAND3XLTS U229 ( .A(n1386), .B(n1385), .C(n1384), .Y(n1255) );
  NAND3XLTS U230 ( .A(n1795), .B(n1794), .C(n1793), .Y(n1170) );
  NAND3XLTS U231 ( .A(n1787), .B(n1786), .C(n1785), .Y(n1171) );
  NAND3XLTS U232 ( .A(n1776), .B(n1775), .C(n1774), .Y(n1172) );
  NAND3XLTS U233 ( .A(n1766), .B(n1765), .C(n1764), .Y(n1173) );
  NAND3XLTS U234 ( .A(n948), .B(n947), .C(n946), .Y(n1290) );
  NAND3XLTS U235 ( .A(n942), .B(n941), .C(n940), .Y(n1291) );
  NAND3XLTS U236 ( .A(n937), .B(n936), .C(n935), .Y(n1292) );
  NAND3XLTS U237 ( .A(n929), .B(n928), .C(n927), .Y(n1293) );
  NAND3XLTS U238 ( .A(n1761), .B(n1760), .C(n1759), .Y(n1182) );
  NAND3XLTS U239 ( .A(n1756), .B(n1755), .C(n1754), .Y(n1183) );
  NAND3XLTS U240 ( .A(n1746), .B(n1745), .C(n1744), .Y(n1184) );
  NAND3XLTS U241 ( .A(n1737), .B(n1736), .C(n1735), .Y(n1185) );
  NAND3XLTS U242 ( .A(n924), .B(n923), .C(n922), .Y(n1294) );
  NAND3XLTS U243 ( .A(n919), .B(n918), .C(n917), .Y(n1295) );
  NAND3XLTS U244 ( .A(n916), .B(n915), .C(n914), .Y(n1296) );
  NAND3XLTS U245 ( .A(n912), .B(n911), .C(n910), .Y(n1297) );
  NAND3XLTS U246 ( .A(n1523), .B(n1522), .C(n1521), .Y(n1232) );
  NAND3XLTS U247 ( .A(n1516), .B(n1515), .C(n1514), .Y(n1233) );
  NAND3XLTS U248 ( .A(n1509), .B(n1508), .C(n1507), .Y(n1234) );
  NAND3XLTS U249 ( .A(n1502), .B(n1501), .C(n1500), .Y(n1235) );
  NAND3XLTS U250 ( .A(n1492), .B(n1491), .C(n1490), .Y(n1236) );
  NAND3XLTS U251 ( .A(n1482), .B(n1481), .C(n1480), .Y(n1237) );
  NAND3XLTS U252 ( .A(n1576), .B(n1575), .C(n1574), .Y(n1226) );
  NAND3XLTS U253 ( .A(n1566), .B(n1565), .C(n1564), .Y(n1227) );
  NAND3XLTS U254 ( .A(n1557), .B(n1556), .C(n1555), .Y(n1228) );
  NAND3XLTS U255 ( .A(n1549), .B(n1548), .C(n1547), .Y(n1229) );
  NAND3XLTS U256 ( .A(n1541), .B(n1540), .C(n1539), .Y(n1230) );
  NAND3XLTS U257 ( .A(n1532), .B(n1531), .C(n1530), .Y(n1231) );
  NAND3XLTS U258 ( .A(n1084), .B(n1083), .C(n1082), .Y(n1268) );
  NAND3XLTS U259 ( .A(n1079), .B(n1078), .C(n1077), .Y(n1269) );
  NAND3XLTS U260 ( .A(n1072), .B(n1071), .C(n1070), .Y(n1270) );
  NAND3XLTS U261 ( .A(n1068), .B(n1067), .C(n1066), .Y(n1271) );
  NAND3XLTS U262 ( .A(n1062), .B(n1061), .C(n1060), .Y(n1272) );
  NAND3XLTS U263 ( .A(n1057), .B(n1056), .C(n1055), .Y(n1273) );
  NAND3XLTS U264 ( .A(n1851), .B(n1850), .C(n1849), .Y(n1146) );
  NAND3XLTS U265 ( .A(n1844), .B(n1843), .C(n1842), .Y(n1147) );
  NAND3XLTS U266 ( .A(n1835), .B(n1834), .C(n1833), .Y(n1148) );
  NAND3XLTS U267 ( .A(n1828), .B(n1827), .C(n1826), .Y(n1149) );
  NAND3XLTS U268 ( .A(n990), .B(n989), .C(n988), .Y(n1282) );
  NAND3XLTS U269 ( .A(n985), .B(n984), .C(n983), .Y(n1283) );
  NAND3XLTS U270 ( .A(n981), .B(n980), .C(n979), .Y(n1284) );
  NAND3XLTS U271 ( .A(n977), .B(n976), .C(n975), .Y(n1285) );
  AOI211XLTS U272 ( .A0(n492), .A1(n527), .B0(n491), .C0(n490), .Y(n493) );
  XOR2XLTS U273 ( .A(n526), .B(n495), .Y(n491) );
  OAI21XLTS U274 ( .A0(n492), .A1(n527), .B0(n489), .Y(n490) );
  NOR2XLTS U275 ( .A(n1642), .B(n1639), .Y(n187) );
  OR2X1TS U276 ( .A(n320), .B(n998), .Y(n358) );
  NAND2X1TS U277 ( .A(n28), .B(n25), .Y(n26) );
  OR2X1TS U278 ( .A(n1603), .B(n230), .Y(n1) );
  OR2X1TS U279 ( .A(n1659), .B(n400), .Y(n2) );
  OR2X1TS U280 ( .A(n1589), .B(n90), .Y(n3) );
  OR2X1TS U281 ( .A(n1614), .B(n279), .Y(n4) );
  OR2X1TS U282 ( .A(n1662), .B(n400), .Y(n5) );
  OR2X1TS U283 ( .A(n1649), .B(n325), .Y(n6) );
  OA21XLTS U284 ( .A0(n19), .A1(n83), .B0(n22), .Y(n7) );
  OR2X1TS U285 ( .A(n21), .B(n508), .Y(n8) );
  OR2X1TS U286 ( .A(n443), .B(n1597), .Y(n9) );
  OR2X1TS U287 ( .A(n443), .B(n1643), .Y(n10) );
  OR2X1TS U288 ( .A(n395), .B(n1030), .Y(n425) );
  NOR2XLTS U289 ( .A(n26), .B(n133), .Y(n129) );
  NOR3XLTS U290 ( .A(n1670), .B(n1663), .C(n399), .Y(n394) );
  NOR3XLTS U291 ( .A(n1585), .B(n1580), .C(n37), .Y(n32) );
  NOR3XLTS U292 ( .A(n1596), .B(n1591), .C(n89), .Y(n84) );
  NOR3XLTS U293 ( .A(n1609), .B(n1604), .C(n229), .Y(n224) );
  NOR3XLTS U294 ( .A(n1621), .B(n1615), .C(n278), .Y(n274) );
  NOR3XLTS U295 ( .A(n1642), .B(n1636), .C(n188), .Y(n184) );
  NOR3XLTS U296 ( .A(n1656), .B(n1650), .C(n323), .Y(n317) );
  OR2X1TS U297 ( .A(n275), .B(n1622), .Y(n11) );
  OR2X1TS U298 ( .A(n443), .B(n1671), .Y(n12) );
  NOR2XLTS U299 ( .A(n845), .B(n520), .Y(n692) );
  NOR2XLTS U300 ( .A(n845), .B(n519), .Y(n545) );
  INVX2TS U301 ( .A(destinationAddressIn_EAST[6]), .Y(n70) );
  INVX2TS U302 ( .A(destinationAddressIn_EAST[4]), .Y(n62) );
  INVX2TS U303 ( .A(destinationAddressIn_EAST[7]), .Y(n65) );
  INVX2TS U304 ( .A(destinationAddressIn_EAST[5]), .Y(n73) );
  INVX2TS U305 ( .A(destinationAddressIn_EAST[11]), .Y(n47) );
  INVX2TS U306 ( .A(destinationAddressIn_EAST[10]), .Y(n51) );
  INVX2TS U307 ( .A(destinationAddressIn_EAST[9]), .Y(n33) );
  INVX2TS U308 ( .A(destinationAddressIn_EAST[8]), .Y(n41) );
  INVX2TS U309 ( .A(writeIn_EAST), .Y(n55) );
  CLKBUFX2TS U310 ( .A(n1955), .Y(n13) );
  INVX2TS U326 ( .A(n1962), .Y(n497) );
  INVX2TS U327 ( .A(n1958), .Y(n448) );
  ADDFHX1TS U328 ( .A(selectBit_SOUTH), .B(selectBit_NORTH), .CI(
        selectBit_EAST), .CO(n466), .S(n461) );
  INVX2TS U329 ( .A(n15), .Y(n78) );
  INVX2TS U330 ( .A(n78), .Y(n122) );
  INVX2TS U331 ( .A(selectBit_WEST), .Y(n456) );
  INVX2TS U332 ( .A(n1583), .Y(n1585) );
  INVX2TS U333 ( .A(n1954), .Y(n460) );
  INVX2TS U334 ( .A(selectBit_SOUTH), .Y(n508) );
  INVX2TS U335 ( .A(n8), .Y(n222) );
  INVX2TS U336 ( .A(n1962), .Y(n83) );
  INVX2TS U337 ( .A(n1962), .Y(n487) );
  NAND2X1TS U338 ( .A(n18), .B(n487), .Y(n22) );
  INVX2TS U339 ( .A(n7), .Y(n80) );
  NAND2X1TS U340 ( .A(selectBit_SOUTH), .B(n21), .Y(n20) );
  OAI21XLTS U341 ( .A0(selectBit_SOUTH), .A1(n21), .B0(n81), .Y(n269) );
  NAND2X1TS U342 ( .A(n314), .B(n269), .Y(n125) );
  INVX2TS U343 ( .A(selectBit_EAST), .Y(n515) );
  INVX2TS U344 ( .A(n515), .Y(n512) );
  INVX2TS U345 ( .A(n22), .Y(n126) );
  INVX2TS U346 ( .A(n1959), .Y(n453) );
  AOI22X1TS U347 ( .A0(n482), .A1(n22), .B0(n126), .B1(n453), .Y(n23) );
  INVX2TS U348 ( .A(n23), .Y(n24) );
  INVX2TS U349 ( .A(n24), .Y(n25) );
  INVX2TS U350 ( .A(n26), .Y(n121) );
  INVX2TS U351 ( .A(n121), .Y(n27) );
  NAND2X1TS U352 ( .A(n454), .B(n126), .Y(n31) );
  INVX2TS U353 ( .A(n25), .Y(n29) );
  INVX2TS U354 ( .A(n508), .Y(n507) );
  INVX2TS U355 ( .A(n456), .Y(n513) );
  INVX2TS U356 ( .A(readReady), .Y(n183) );
  INVX2TS U357 ( .A(n183), .Y(n516) );
  NOR3XLTS U358 ( .A(n513), .B(selectBit_EAST), .C(n516), .Y(n509) );
  NAND2X1TS U359 ( .A(n540), .B(n509), .Y(n525) );
  INVX2TS U360 ( .A(n130), .Y(n452) );
  INVX2TS U361 ( .A(n452), .Y(n85) );
  INVX2TS U362 ( .A(n85), .Y(n30) );
  AOI31XLTS U363 ( .A0(n36), .A1(n31), .A2(n1578), .B0(n30), .Y(n35) );
  INVX2TS U364 ( .A(n1958), .Y(n449) );
  INVX2TS U365 ( .A(n1960), .Y(n273) );
  INVX2TS U366 ( .A(n183), .Y(n514) );
  NAND2X1TS U367 ( .A(n35), .B(n1586), .Y(n37) );
  INVX2TS U368 ( .A(n32), .Y(n887) );
  INVX2TS U369 ( .A(n887), .Y(n1569) );
  CLKBUFX2TS U370 ( .A(n1569), .Y(n46) );
  INVX2TS U371 ( .A(n46), .Y(n69) );
  INVX2TS U372 ( .A(destinationAddressIn_EAST[9]), .Y(n237) );
  INVX2TS U373 ( .A(n34), .Y(n886) );
  INVX2TS U374 ( .A(n886), .Y(n1673) );
  INVX2TS U375 ( .A(n1542), .Y(n52) );
  OR2X1TS U376 ( .A(n1583), .B(n37), .Y(n56) );
  INVX2TS U377 ( .A(n56), .Y(n1680) );
  CLKBUFX2TS U378 ( .A(destinationAddressIn_WEST[9]), .Y(n411) );
  CLKBUFX2TS U379 ( .A(n411), .Y(n732) );
  AOI22X1TS U380 ( .A0(n52), .A1(\destinationAddressbuffer[7][9] ), .B0(n1680), 
        .B1(n732), .Y(n40) );
  INVX2TS U381 ( .A(n43), .Y(n1527) );
  INVX2TS U382 ( .A(n1527), .Y(n1563) );
  INVX2TS U383 ( .A(n151), .Y(n733) );
  OR2X1TS U384 ( .A(n1579), .B(n38), .Y(n59) );
  INVX2TS U385 ( .A(n59), .Y(n1561) );
  INVX2TS U386 ( .A(n1561), .Y(n875) );
  INVX2TS U387 ( .A(n875), .Y(n1572) );
  CLKBUFX2TS U388 ( .A(destinationAddressIn_NORTH[9]), .Y(n735) );
  CLKBUFX2TS U389 ( .A(n735), .Y(n350) );
  AOI22X1TS U390 ( .A0(n1563), .A1(n733), .B0(n1572), .B1(n350), .Y(n39) );
  OAI211XLTS U391 ( .A0(n69), .A1(n237), .B0(n40), .C0(n39), .Y(n1200) );
  INVX2TS U392 ( .A(destinationAddressIn_EAST[8]), .Y(n234) );
  INVX2TS U393 ( .A(n56), .Y(n42) );
  INVX2TS U394 ( .A(n42), .Y(n879) );
  INVX2TS U395 ( .A(n879), .Y(n66) );
  CLKBUFX2TS U396 ( .A(destinationAddressIn_WEST[8]), .Y(n416) );
  CLKBUFX2TS U397 ( .A(n416), .Y(n717) );
  AOI22X1TS U398 ( .A0(n52), .A1(\destinationAddressbuffer[7][8] ), .B0(n66), 
        .B1(n717), .Y(n45) );
  INVX2TS U399 ( .A(n43), .Y(n57) );
  INVX2TS U400 ( .A(n57), .Y(n1698) );
  INVX2TS U401 ( .A(n146), .Y(n718) );
  CLKBUFX2TS U402 ( .A(destinationAddressIn_NORTH[8]), .Y(n719) );
  CLKBUFX2TS U403 ( .A(n719), .Y(n334) );
  AOI22X1TS U404 ( .A0(n1698), .A1(n718), .B0(n1561), .B1(n334), .Y(n44) );
  OAI211XLTS U405 ( .A0(n69), .A1(n234), .B0(n45), .C0(n44), .Y(n1201) );
  INVX2TS U406 ( .A(n46), .Y(n77) );
  INVX2TS U407 ( .A(destinationAddressIn_EAST[11]), .Y(n242) );
  CLKBUFX2TS U408 ( .A(destinationAddressIn_WEST[11]), .Y(n397) );
  CLKBUFX2TS U409 ( .A(n397), .Y(n764) );
  AOI22X1TS U410 ( .A0(n52), .A1(\destinationAddressbuffer[7][11] ), .B0(n66), 
        .B1(n764), .Y(n50) );
  INVX2TS U411 ( .A(n57), .Y(n1538) );
  INVX2TS U412 ( .A(n142), .Y(n767) );
  INVX2TS U413 ( .A(n59), .Y(n48) );
  CLKBUFX2TS U414 ( .A(destinationAddressIn_NORTH[11]), .Y(n768) );
  CLKBUFX2TS U415 ( .A(n768), .Y(n340) );
  AOI22X1TS U416 ( .A0(n1538), .A1(n767), .B0(n48), .B1(n340), .Y(n49) );
  OAI211XLTS U417 ( .A0(n77), .A1(n242), .B0(n50), .C0(n49), .Y(n1198) );
  INVX2TS U418 ( .A(destinationAddressIn_EAST[10]), .Y(n247) );
  INVX2TS U419 ( .A(n56), .Y(n1688) );
  CLKBUFX2TS U420 ( .A(destinationAddressIn_WEST[10]), .Y(n405) );
  CLKBUFX2TS U421 ( .A(n405), .Y(n749) );
  AOI22X1TS U422 ( .A0(n52), .A1(\destinationAddressbuffer[7][10] ), .B0(n1688), .B1(n749), .Y(n54) );
  INVX2TS U423 ( .A(n57), .Y(n888) );
  INVX2TS U424 ( .A(n138), .Y(n752) );
  INVX2TS U425 ( .A(n59), .Y(n1681) );
  CLKBUFX2TS U426 ( .A(destinationAddressIn_NORTH[10]), .Y(n753) );
  CLKBUFX2TS U427 ( .A(n753), .Y(n328) );
  AOI22X1TS U428 ( .A0(n888), .A1(n752), .B0(n1681), .B1(n328), .Y(n53) );
  OAI211XLTS U429 ( .A0(n69), .A1(n247), .B0(n54), .C0(n53), .Y(n1199) );
  INVX2TS U430 ( .A(n1587), .Y(n1694) );
  INVX2TS U431 ( .A(n56), .Y(n1526) );
  AOI22X1TS U432 ( .A0(n1694), .A1(writeOutbuffer[7]), .B0(n1526), .B1(
        writeIn_WEST), .Y(n61) );
  INVX2TS U433 ( .A(n57), .Y(n58) );
  INVX2TS U434 ( .A(writeIn_SOUTH), .Y(n155) );
  INVX2TS U435 ( .A(n155), .Y(n546) );
  INVX2TS U436 ( .A(n59), .Y(n1689) );
  AOI22X1TS U437 ( .A0(n58), .A1(n546), .B0(n1689), .B1(writeIn_NORTH), .Y(n60) );
  OAI211XLTS U438 ( .A0(n77), .A1(n295), .B0(n61), .C0(n60), .Y(n1225) );
  INVX2TS U439 ( .A(destinationAddressIn_EAST[4]), .Y(n262) );
  INVX2TS U440 ( .A(n1542), .Y(n74) );
  CLKBUFX2TS U441 ( .A(destinationAddressIn_WEST[4]), .Y(n158) );
  CLKBUFX2TS U442 ( .A(n158), .Y(n659) );
  AOI22X1TS U443 ( .A0(n74), .A1(\destinationAddressbuffer[7][4] ), .B0(n1688), 
        .B1(n659), .Y(n64) );
  INVX2TS U444 ( .A(destinationAddressIn_SOUTH[4]), .Y(n161) );
  INVX2TS U445 ( .A(n161), .Y(n661) );
  AOI22X1TS U446 ( .A0(n888), .A1(n661), .B0(n1681), .B1(
        destinationAddressIn_NORTH[4]), .Y(n63) );
  OAI211XLTS U447 ( .A0(n77), .A1(n262), .B0(n64), .C0(n63), .Y(n1205) );
  INVX2TS U448 ( .A(destinationAddressIn_EAST[7]), .Y(n266) );
  CLKBUFX2TS U449 ( .A(destinationAddressIn_WEST[7]), .Y(n164) );
  CLKBUFX2TS U450 ( .A(n164), .Y(n706) );
  AOI22X1TS U451 ( .A0(n74), .A1(\destinationAddressbuffer[7][7] ), .B0(n66), 
        .B1(n706), .Y(n68) );
  INVX2TS U452 ( .A(destinationAddressIn_SOUTH[7]), .Y(n167) );
  INVX2TS U453 ( .A(n167), .Y(n707) );
  AOI22X1TS U454 ( .A0(n58), .A1(n707), .B0(n1689), .B1(
        destinationAddressIn_NORTH[7]), .Y(n67) );
  OAI211XLTS U455 ( .A0(n69), .A1(n266), .B0(n68), .C0(n67), .Y(n1202) );
  INVX2TS U456 ( .A(destinationAddressIn_EAST[6]), .Y(n253) );
  CLKBUFX2TS U457 ( .A(destinationAddressIn_WEST[6]), .Y(n170) );
  CLKBUFX2TS U458 ( .A(n170), .Y(n691) );
  AOI22X1TS U459 ( .A0(n74), .A1(\destinationAddressbuffer[7][6] ), .B0(n1526), 
        .B1(n691), .Y(n72) );
  INVX2TS U460 ( .A(destinationAddressIn_SOUTH[6]), .Y(n173) );
  INVX2TS U461 ( .A(n173), .Y(n693) );
  AOI22X1TS U462 ( .A0(n1538), .A1(n693), .B0(n1572), .B1(
        destinationAddressIn_NORTH[6]), .Y(n71) );
  OAI211XLTS U463 ( .A0(n887), .A1(n253), .B0(n72), .C0(n71), .Y(n1203) );
  INVX2TS U464 ( .A(destinationAddressIn_EAST[5]), .Y(n256) );
  CLKBUFX2TS U465 ( .A(destinationAddressIn_WEST[5]), .Y(n175) );
  CLKBUFX2TS U466 ( .A(n175), .Y(n672) );
  AOI22X1TS U467 ( .A0(n74), .A1(\destinationAddressbuffer[7][5] ), .B0(n42), 
        .B1(n672), .Y(n76) );
  INVX2TS U468 ( .A(destinationAddressIn_SOUTH[5]), .Y(n179) );
  INVX2TS U469 ( .A(n179), .Y(n673) );
  AOI22X1TS U470 ( .A0(n1698), .A1(n673), .B0(n48), .B1(
        destinationAddressIn_NORTH[5]), .Y(n75) );
  OAI211XLTS U471 ( .A0(n77), .A1(n256), .B0(n76), .C0(n75), .Y(n1204) );
  INVX2TS U472 ( .A(n79), .Y(n181) );
  NAND2X1TS U473 ( .A(n123), .B(n513), .Y(n268) );
  AOI21X1TS U474 ( .A0(n222), .A1(n80), .B0(n314), .Y(n387) );
  NOR3XLTS U475 ( .A(n387), .B(n270), .C(n269), .Y(n1593) );
  INVX2TS U476 ( .A(n1962), .Y(n458) );
  NOR2XLTS U477 ( .A(n449), .B(n506), .Y(n390) );
  NOR3XLTS U478 ( .A(n25), .B(n81), .C(n271), .Y(n1590) );
  AOI31XLTS U479 ( .A0(n454), .A1(n458), .A2(n390), .B0(n1590), .Y(n82) );
  AOI21X1TS U480 ( .A0(n88), .A1(n82), .B0(n275), .Y(n86) );
  INVX2TS U481 ( .A(n1954), .Y(n393) );
  NAND2X1TS U482 ( .A(n86), .B(n1597), .Y(n89) );
  INVX2TS U483 ( .A(n84), .Y(n1485) );
  INVX2TS U484 ( .A(n1485), .Y(n905) );
  CLKBUFX2TS U485 ( .A(n905), .Y(n97) );
  INVX2TS U486 ( .A(n97), .Y(n113) );
  INVX2TS U487 ( .A(n85), .Y(n443) );
  INVX2TS U488 ( .A(n9), .Y(n895) );
  INVX2TS U489 ( .A(n1493), .Y(n101) );
  OR2X1TS U490 ( .A(n1594), .B(n89), .Y(n105) );
  INVX2TS U491 ( .A(n105), .Y(n87) );
  AOI22X1TS U492 ( .A0(n101), .A1(\destinationAddressbuffer[6][8] ), .B0(n87), 
        .B1(n717), .Y(n93) );
  INVX2TS U493 ( .A(n102), .Y(n110) );
  INVX2TS U494 ( .A(n110), .Y(n1721) );
  CLKBUFX2TS U495 ( .A(n719), .Y(n419) );
  INVX2TS U496 ( .A(n3), .Y(n91) );
  INVX2TS U497 ( .A(n146), .Y(n333) );
  AOI22X1TS U498 ( .A0(n1721), .A1(n419), .B0(n91), .B1(n333), .Y(n92) );
  OAI211XLTS U499 ( .A0(n113), .A1(n234), .B0(n93), .C0(n92), .Y(n1189) );
  AOI22X1TS U500 ( .A0(n101), .A1(\destinationAddressbuffer[6][10] ), .B0(n116), .B1(n749), .Y(n96) );
  INVX2TS U501 ( .A(n110), .Y(n94) );
  CLKBUFX2TS U502 ( .A(n753), .Y(n406) );
  INVX2TS U503 ( .A(n3), .Y(n1711) );
  INVX2TS U504 ( .A(n138), .Y(n327) );
  AOI22X1TS U505 ( .A0(n94), .A1(n406), .B0(n1711), .B1(n327), .Y(n95) );
  OAI211XLTS U506 ( .A0(n113), .A1(n247), .B0(n96), .C0(n95), .Y(n1187) );
  INVX2TS U507 ( .A(n97), .Y(n120) );
  INVX2TS U508 ( .A(n105), .Y(n1496) );
  INVX2TS U509 ( .A(n1496), .Y(n896) );
  INVX2TS U510 ( .A(n896), .Y(n98) );
  AOI22X1TS U511 ( .A0(n101), .A1(\destinationAddressbuffer[6][11] ), .B0(n98), 
        .B1(n764), .Y(n100) );
  CLKBUFX2TS U512 ( .A(n768), .Y(n402) );
  INVX2TS U513 ( .A(n3), .Y(n1729) );
  INVX2TS U514 ( .A(n142), .Y(n339) );
  AOI22X1TS U515 ( .A0(n94), .A1(n402), .B0(n1729), .B1(n339), .Y(n99) );
  OAI211XLTS U516 ( .A0(n120), .A1(n242), .B0(n100), .C0(n99), .Y(n1186) );
  INVX2TS U517 ( .A(n896), .Y(n116) );
  AOI22X1TS U518 ( .A0(n101), .A1(\destinationAddressbuffer[6][9] ), .B0(n116), 
        .B1(n732), .Y(n104) );
  INVX2TS U519 ( .A(n102), .Y(n1487) );
  INVX2TS U520 ( .A(n1487), .Y(n901) );
  CLKBUFX2TS U521 ( .A(n735), .Y(n412) );
  INVX2TS U522 ( .A(n3), .Y(n1498) );
  INVX2TS U523 ( .A(n1498), .Y(n897) );
  INVX2TS U524 ( .A(n151), .Y(n348) );
  AOI22X1TS U525 ( .A0(n901), .A1(n412), .B0(n1703), .B1(n348), .Y(n103) );
  OAI211XLTS U526 ( .A0(n113), .A1(n237), .B0(n104), .C0(n103), .Y(n1188) );
  INVX2TS U527 ( .A(n1598), .Y(n1725) );
  INVX2TS U528 ( .A(n105), .Y(n1709) );
  AOI22X1TS U529 ( .A0(n1725), .A1(writeOutbuffer[6]), .B0(n1709), .B1(
        writeIn_WEST), .Y(n107) );
  INVX2TS U530 ( .A(n110), .Y(n1513) );
  CLKBUFX2TS U531 ( .A(writeIn_NORTH), .Y(n355) );
  CLKBUFX2TS U532 ( .A(n355), .Y(n422) );
  INVX2TS U533 ( .A(n155), .Y(n354) );
  AOI22X1TS U534 ( .A0(n1513), .A1(n422), .B0(n1711), .B1(n354), .Y(n106) );
  OAI211XLTS U535 ( .A0(n120), .A1(n295), .B0(n107), .C0(n106), .Y(n1224) );
  INVX2TS U536 ( .A(n1598), .Y(n117) );
  AOI22X1TS U537 ( .A0(n117), .A1(\destinationAddressbuffer[6][4] ), .B0(n98), 
        .B1(n659), .Y(n109) );
  CLKBUFX2TS U538 ( .A(destinationAddressIn_NORTH[4]), .Y(n381) );
  CLKBUFX2TS U539 ( .A(n381), .Y(n431) );
  INVX2TS U540 ( .A(n161), .Y(n380) );
  AOI22X1TS U541 ( .A0(n1721), .A1(n431), .B0(n1729), .B1(n380), .Y(n108) );
  OAI211XLTS U542 ( .A0(n120), .A1(n262), .B0(n109), .C0(n108), .Y(n1193) );
  AOI22X1TS U543 ( .A0(n117), .A1(\destinationAddressbuffer[6][7] ), .B0(n87), 
        .B1(n706), .Y(n112) );
  INVX2TS U544 ( .A(n110), .Y(n1712) );
  CLKBUFX2TS U545 ( .A(destinationAddressIn_NORTH[7]), .Y(n361) );
  CLKBUFX2TS U546 ( .A(n361), .Y(n435) );
  INVX2TS U547 ( .A(n167), .Y(n360) );
  AOI22X1TS U548 ( .A0(n1712), .A1(n435), .B0(n1498), .B1(n360), .Y(n111) );
  OAI211XLTS U549 ( .A0(n113), .A1(n266), .B0(n112), .C0(n111), .Y(n1190) );
  AOI22X1TS U550 ( .A0(n117), .A1(\destinationAddressbuffer[6][6] ), .B0(n1709), .B1(n691), .Y(n115) );
  CLKBUFX2TS U551 ( .A(destinationAddressIn_NORTH[6]), .Y(n367) );
  CLKBUFX2TS U552 ( .A(n367), .Y(n426) );
  INVX2TS U553 ( .A(n173), .Y(n365) );
  AOI22X1TS U554 ( .A0(n901), .A1(n426), .B0(n91), .B1(n365), .Y(n114) );
  OAI211XLTS U555 ( .A0(n1485), .A1(n253), .B0(n115), .C0(n114), .Y(n1191) );
  AOI22X1TS U556 ( .A0(n117), .A1(\destinationAddressbuffer[6][5] ), .B0(n116), 
        .B1(n672), .Y(n119) );
  CLKBUFX2TS U557 ( .A(destinationAddressIn_NORTH[5]), .Y(n373) );
  CLKBUFX2TS U558 ( .A(n373), .Y(n439) );
  INVX2TS U559 ( .A(n897), .Y(n1720) );
  INVX2TS U560 ( .A(n179), .Y(n372) );
  AOI22X1TS U561 ( .A0(n1712), .A1(n439), .B0(n1720), .B1(n372), .Y(n118) );
  OAI211XLTS U562 ( .A0(n120), .A1(n256), .B0(n119), .C0(n118), .Y(n1192) );
  INVX2TS U563 ( .A(n1959), .Y(n446) );
  NAND2X1TS U564 ( .A(n126), .B(n446), .Y(n127) );
  INVX2TS U565 ( .A(n130), .Y(n275) );
  AOI31XLTS U566 ( .A0(n128), .A1(n27), .A2(n127), .B0(n275), .Y(n132) );
  INVX2TS U567 ( .A(n1959), .Y(n444) );
  INVX2TS U568 ( .A(n129), .Y(n964) );
  INVX2TS U569 ( .A(n964), .Y(n1409) );
  CLKBUFX2TS U570 ( .A(n1409), .Y(n143) );
  INVX2TS U571 ( .A(n143), .Y(n168) );
  INVX2TS U572 ( .A(n130), .Y(n318) );
  INVX2TS U573 ( .A(n131), .Y(n1382) );
  INVX2TS U574 ( .A(n1382), .Y(n956) );
  INVX2TS U575 ( .A(n1632), .Y(n148) );
  NOR3XLTS U576 ( .A(n1630), .B(n1625), .C(n134), .Y(n147) );
  INVX2TS U577 ( .A(n147), .Y(n156) );
  INVX2TS U578 ( .A(n156), .Y(n1383) );
  AOI22X1TS U579 ( .A0(n148), .A1(\destinationAddressbuffer[3][10] ), .B0(
        n1383), .B1(destinationAddressIn_EAST[10]), .Y(n137) );
  OR2X1TS U580 ( .A(n121), .B(n133), .Y(n162) );
  INVX2TS U581 ( .A(n162), .Y(n1805) );
  INVX2TS U582 ( .A(n135), .Y(n152) );
  INVX2TS U583 ( .A(n152), .Y(n1820) );
  CLKBUFX2TS U584 ( .A(n405), .Y(n321) );
  AOI22X1TS U585 ( .A0(n1805), .A1(n328), .B0(n1820), .B1(n321), .Y(n136) );
  OAI211XLTS U586 ( .A0(n168), .A1(n138), .B0(n137), .C0(n136), .Y(n1151) );
  INVX2TS U587 ( .A(n156), .Y(n1802) );
  AOI22X1TS U588 ( .A0(n148), .A1(\destinationAddressbuffer[3][11] ), .B0(
        n1802), .B1(destinationAddressIn_EAST[11]), .Y(n141) );
  INVX2TS U589 ( .A(n162), .Y(n1812) );
  INVX2TS U590 ( .A(n152), .Y(n139) );
  INVX2TS U591 ( .A(n139), .Y(n950) );
  INVX2TS U592 ( .A(n950), .Y(n176) );
  CLKBUFX2TS U593 ( .A(n397), .Y(n338) );
  AOI22X1TS U594 ( .A0(n1812), .A1(n340), .B0(n176), .B1(n338), .Y(n140) );
  OAI211XLTS U595 ( .A0(n964), .A1(n142), .B0(n141), .C0(n140), .Y(n1150) );
  INVX2TS U596 ( .A(n143), .Y(n180) );
  AOI22X1TS U597 ( .A0(n148), .A1(\destinationAddressbuffer[3][8] ), .B0(n1383), .B1(destinationAddressIn_EAST[8]), .Y(n145) );
  INVX2TS U598 ( .A(n162), .Y(n1402) );
  INVX2TS U599 ( .A(n152), .Y(n1804) );
  CLKBUFX2TS U600 ( .A(n416), .Y(n332) );
  AOI22X1TS U601 ( .A0(n1402), .A1(n334), .B0(n1804), .B1(n332), .Y(n144) );
  OAI211XLTS U602 ( .A0(n180), .A1(n146), .B0(n145), .C0(n144), .Y(n1153) );
  INVX2TS U603 ( .A(n147), .Y(n957) );
  INVX2TS U604 ( .A(n957), .Y(n169) );
  AOI22X1TS U605 ( .A0(n148), .A1(\destinationAddressbuffer[3][9] ), .B0(n169), 
        .B1(destinationAddressIn_EAST[9]), .Y(n150) );
  INVX2TS U606 ( .A(n1812), .Y(n1388) );
  INVX2TS U607 ( .A(n1388), .Y(n965) );
  CLKBUFX2TS U608 ( .A(n411), .Y(n345) );
  AOI22X1TS U609 ( .A0(n965), .A1(n350), .B0(n1804), .B1(n345), .Y(n149) );
  OAI211XLTS U610 ( .A0(n168), .A1(n151), .B0(n150), .C0(n149), .Y(n1152) );
  INVX2TS U611 ( .A(n1632), .Y(n1816) );
  INVX2TS U612 ( .A(n156), .Y(n1810) );
  AOI22X1TS U613 ( .A0(n1816), .A1(writeOutbuffer[3]), .B0(n1810), .B1(
        writeIn_EAST), .Y(n154) );
  INVX2TS U614 ( .A(n152), .Y(n1408) );
  CLKBUFX2TS U615 ( .A(writeIn_WEST), .Y(n544) );
  CLKBUFX2TS U616 ( .A(n544), .Y(n353) );
  AOI22X1TS U617 ( .A0(n1805), .A1(n355), .B0(n1408), .B1(n353), .Y(n153) );
  OAI211XLTS U618 ( .A0(n168), .A1(n155), .B0(n154), .C0(n153), .Y(n1221) );
  INVX2TS U619 ( .A(n1392), .Y(n174) );
  INVX2TS U620 ( .A(n156), .Y(n157) );
  AOI22X1TS U621 ( .A0(n174), .A1(\destinationAddressbuffer[3][4] ), .B0(n169), 
        .B1(destinationAddressIn_EAST[4]), .Y(n160) );
  CLKBUFX2TS U622 ( .A(n158), .Y(n377) );
  AOI22X1TS U623 ( .A0(n1812), .A1(n381), .B0(n1820), .B1(n377), .Y(n159) );
  OAI211XLTS U624 ( .A0(n180), .A1(n161), .B0(n160), .C0(n159), .Y(n1157) );
  AOI22X1TS U625 ( .A0(n174), .A1(\destinationAddressbuffer[3][7] ), .B0(n1810), .B1(destinationAddressIn_EAST[7]), .Y(n166) );
  INVX2TS U626 ( .A(n162), .Y(n163) );
  CLKBUFX2TS U627 ( .A(n164), .Y(n359) );
  AOI22X1TS U628 ( .A0(n163), .A1(n361), .B0(n1408), .B1(n359), .Y(n165) );
  OAI211XLTS U629 ( .A0(n168), .A1(n167), .B0(n166), .C0(n165), .Y(n1154) );
  AOI22X1TS U630 ( .A0(n174), .A1(\destinationAddressbuffer[3][6] ), .B0(n169), 
        .B1(destinationAddressIn_EAST[6]), .Y(n172) );
  CLKBUFX2TS U631 ( .A(n170), .Y(n364) );
  AOI22X1TS U632 ( .A0(n965), .A1(n367), .B0(n139), .B1(n364), .Y(n171) );
  OAI211XLTS U633 ( .A0(n180), .A1(n173), .B0(n172), .C0(n171), .Y(n1155) );
  AOI22X1TS U634 ( .A0(n174), .A1(\destinationAddressbuffer[3][5] ), .B0(n1802), .B1(destinationAddressIn_EAST[5]), .Y(n178) );
  CLKBUFX2TS U635 ( .A(n175), .Y(n371) );
  AOI22X1TS U636 ( .A0(n965), .A1(n373), .B0(n176), .B1(n371), .Y(n177) );
  OAI211XLTS U637 ( .A0(n180), .A1(n179), .B0(n178), .C0(n177), .Y(n1156) );
  INVX2TS U638 ( .A(n269), .Y(n315) );
  INVX2TS U639 ( .A(n315), .Y(n385) );
  NOR3XLTS U640 ( .A(n387), .B(n385), .C(n386), .Y(n1639) );
  AOI31XLTS U641 ( .A0(n497), .A1(n390), .A2(n453), .B0(n1635), .Y(n182) );
  AOI21X1TS U642 ( .A0(n187), .A1(n182), .B0(n443), .Y(n185) );
  INVX2TS U643 ( .A(n183), .Y(n511) );
  NAND2X1TS U644 ( .A(n185), .B(n1643), .Y(n188) );
  INVX2TS U645 ( .A(n184), .Y(n1346) );
  INVX2TS U646 ( .A(n1346), .Y(n987) );
  CLKBUFX2TS U647 ( .A(n987), .Y(n197) );
  INVX2TS U648 ( .A(n197), .Y(n214) );
  INVX2TS U649 ( .A(n10), .Y(n978) );
  INVX2TS U650 ( .A(n1357), .Y(n202) );
  OR2X1TS U651 ( .A(n1640), .B(n188), .Y(n201) );
  INVX2TS U652 ( .A(n201), .Y(n186) );
  INVX2TS U653 ( .A(n186), .Y(n986) );
  INVX2TS U654 ( .A(n986), .Y(n208) );
  AOI22X1TS U655 ( .A0(n202), .A1(\destinationAddressbuffer[2][8] ), .B0(n208), 
        .B1(n332), .Y(n192) );
  INVX2TS U656 ( .A(n193), .Y(n211) );
  INVX2TS U657 ( .A(n211), .Y(n1360) );
  INVX2TS U658 ( .A(n190), .Y(n203) );
  INVX2TS U659 ( .A(n190), .Y(n974) );
  INVX2TS U660 ( .A(n974), .Y(n215) );
  AOI22X1TS U661 ( .A0(n1360), .A1(n334), .B0(n215), .B1(n333), .Y(n191) );
  OAI211XLTS U662 ( .A0(n214), .A1(n234), .B0(n192), .C0(n191), .Y(n1141) );
  INVX2TS U663 ( .A(n201), .Y(n1839) );
  AOI22X1TS U664 ( .A0(n202), .A1(\destinationAddressbuffer[2][9] ), .B0(n1839), .B1(n345), .Y(n196) );
  INVX2TS U665 ( .A(n193), .Y(n1353) );
  INVX2TS U666 ( .A(n1353), .Y(n982) );
  INVX2TS U667 ( .A(n203), .Y(n1831) );
  INVX2TS U668 ( .A(n203), .Y(n194) );
  AOI22X1TS U669 ( .A0(n982), .A1(n350), .B0(n194), .B1(n348), .Y(n195) );
  OAI211XLTS U670 ( .A0(n214), .A1(n237), .B0(n196), .C0(n195), .Y(n1140) );
  INVX2TS U671 ( .A(n197), .Y(n221) );
  INVX2TS U672 ( .A(n201), .Y(n1830) );
  AOI22X1TS U673 ( .A0(n202), .A1(\destinationAddressbuffer[2][10] ), .B0(
        n1830), .B1(n321), .Y(n200) );
  INVX2TS U674 ( .A(n211), .Y(n198) );
  AOI22X1TS U675 ( .A0(n198), .A1(n328), .B0(n215), .B1(n327), .Y(n199) );
  OAI211XLTS U676 ( .A0(n221), .A1(n247), .B0(n200), .C0(n199), .Y(n1139) );
  INVX2TS U677 ( .A(n201), .Y(n1370) );
  AOI22X1TS U678 ( .A0(n202), .A1(\destinationAddressbuffer[2][11] ), .B0(
        n1370), .B1(n338), .Y(n205) );
  AOI22X1TS U679 ( .A0(n198), .A1(n340), .B0(n190), .B1(n339), .Y(n204) );
  OAI211XLTS U680 ( .A0(n214), .A1(n242), .B0(n205), .C0(n204), .Y(n1138) );
  INVX2TS U681 ( .A(n1644), .Y(n1845) );
  AOI22X1TS U682 ( .A0(n1845), .A1(writeOutbuffer[2]), .B0(n208), .B1(n353), 
        .Y(n207) );
  INVX2TS U683 ( .A(n211), .Y(n1832) );
  AOI22X1TS U684 ( .A0(n1832), .A1(writeIn_NORTH), .B0(n1378), .B1(n354), .Y(
        n206) );
  OAI211XLTS U685 ( .A0(n221), .A1(n295), .B0(n207), .C0(n206), .Y(n1220) );
  INVX2TS U686 ( .A(n1357), .Y(n218) );
  AOI22X1TS U687 ( .A0(n218), .A1(\destinationAddressbuffer[2][4] ), .B0(n208), 
        .B1(n377), .Y(n210) );
  AOI22X1TS U688 ( .A0(n1360), .A1(destinationAddressIn_NORTH[4]), .B0(n190), 
        .B1(n380), .Y(n209) );
  OAI211XLTS U689 ( .A0(n221), .A1(n262), .B0(n210), .C0(n209), .Y(n1145) );
  AOI22X1TS U690 ( .A0(n218), .A1(\destinationAddressbuffer[2][5] ), .B0(n1830), .B1(n371), .Y(n213) );
  INVX2TS U691 ( .A(n211), .Y(n1841) );
  INVX2TS U692 ( .A(n974), .Y(n1371) );
  AOI22X1TS U693 ( .A0(n1841), .A1(destinationAddressIn_NORTH[5]), .B0(n1371), 
        .B1(n372), .Y(n212) );
  OAI211XLTS U694 ( .A0(n214), .A1(n256), .B0(n213), .C0(n212), .Y(n1144) );
  AOI22X1TS U695 ( .A0(n218), .A1(\destinationAddressbuffer[2][6] ), .B0(n186), 
        .B1(n364), .Y(n217) );
  AOI22X1TS U696 ( .A0(n982), .A1(destinationAddressIn_NORTH[6]), .B0(n215), 
        .B1(n365), .Y(n216) );
  OAI211XLTS U697 ( .A0(n1346), .A1(n253), .B0(n217), .C0(n216), .Y(n1143) );
  AOI22X1TS U698 ( .A0(n218), .A1(\destinationAddressbuffer[2][7] ), .B0(n1370), .B1(n359), .Y(n220) );
  AOI22X1TS U699 ( .A0(n1841), .A1(destinationAddressIn_NORTH[7]), .B0(n1831), 
        .B1(n360), .Y(n219) );
  OAI211XLTS U700 ( .A0(n221), .A1(n266), .B0(n220), .C0(n219), .Y(n1142) );
  CLKINVX1TS U701 ( .A(n1606), .Y(n1604) );
  INVX2TS U702 ( .A(n1957), .Y(n392) );
  AOI31XLTS U703 ( .A0(n228), .A1(n1600), .A2(n223), .B0(n318), .Y(n226) );
  INVX2TS U704 ( .A(n1957), .Y(n389) );
  NAND2X1TS U705 ( .A(n226), .B(n1610), .Y(n229) );
  INVX2TS U706 ( .A(n224), .Y(n1451) );
  INVX2TS U707 ( .A(n1451), .Y(n921) );
  CLKBUFX2TS U708 ( .A(n921), .Y(n238) );
  INVX2TS U709 ( .A(n238), .Y(n257) );
  INVX2TS U710 ( .A(n225), .Y(n1445) );
  INVX2TS U711 ( .A(n1445), .Y(n913) );
  INVX2TS U712 ( .A(n1456), .Y(n244) );
  OR2X1TS U713 ( .A(n1607), .B(n229), .Y(n243) );
  INVX2TS U714 ( .A(n243), .Y(n227) );
  INVX2TS U715 ( .A(n227), .Y(n920) );
  INVX2TS U716 ( .A(n920), .Y(n258) );
  AOI22X1TS U717 ( .A0(n244), .A1(\destinationAddressbuffer[5][8] ), .B0(n258), 
        .B1(n717), .Y(n233) );
  INVX2TS U718 ( .A(n1600), .Y(n1603) );
  INVX2TS U719 ( .A(n1), .Y(n1743) );
  INVX2TS U720 ( .A(n1743), .Y(n1452) );
  INVX2TS U721 ( .A(n1452), .Y(n259) );
  OR2X1TS U722 ( .A(n1600), .B(n230), .Y(n248) );
  INVX2TS U723 ( .A(n248), .Y(n231) );
  INVX2TS U724 ( .A(n231), .Y(n909) );
  INVX2TS U725 ( .A(n909), .Y(n239) );
  AOI22X1TS U726 ( .A0(n259), .A1(n419), .B0(n239), .B1(n333), .Y(n232) );
  OAI211XLTS U727 ( .A0(n257), .A1(n234), .B0(n233), .C0(n232), .Y(n1177) );
  INVX2TS U728 ( .A(n243), .Y(n1457) );
  AOI22X1TS U729 ( .A0(n244), .A1(\destinationAddressbuffer[5][9] ), .B0(n1457), .B1(n732), .Y(n236) );
  INVX2TS U730 ( .A(n248), .Y(n1467) );
  AOI22X1TS U731 ( .A0(n1743), .A1(n412), .B0(n239), .B1(n348), .Y(n235) );
  OAI211XLTS U732 ( .A0(n257), .A1(n237), .B0(n236), .C0(n235), .Y(n1176) );
  INVX2TS U733 ( .A(n238), .Y(n267) );
  INVX2TS U734 ( .A(n243), .Y(n1741) );
  AOI22X1TS U735 ( .A0(n244), .A1(\destinationAddressbuffer[5][11] ), .B0(
        n1741), .B1(n764), .Y(n241) );
  INVX2TS U736 ( .A(n1), .Y(n1458) );
  AOI22X1TS U737 ( .A0(n1458), .A1(n402), .B0(n239), .B1(n339), .Y(n240) );
  OAI211XLTS U738 ( .A0(n267), .A1(n242), .B0(n241), .C0(n240), .Y(n1174) );
  INVX2TS U739 ( .A(n243), .Y(n1462) );
  AOI22X1TS U740 ( .A0(n244), .A1(\destinationAddressbuffer[5][10] ), .B0(
        n1462), .B1(n749), .Y(n246) );
  INVX2TS U741 ( .A(n1), .Y(n1468) );
  INVX2TS U742 ( .A(n248), .Y(n1742) );
  AOI22X1TS U743 ( .A0(n1753), .A1(n406), .B0(n1742), .B1(n327), .Y(n245) );
  OAI211XLTS U744 ( .A0(n257), .A1(n247), .B0(n246), .C0(n245), .Y(n1175) );
  INVX2TS U745 ( .A(n1611), .Y(n1757) );
  AOI22X1TS U746 ( .A0(n1757), .A1(writeOutbuffer[5]), .B0(n258), .B1(n544), 
        .Y(n250) );
  INVX2TS U747 ( .A(n248), .Y(n1463) );
  AOI22X1TS U748 ( .A0(n1743), .A1(n422), .B0(n1463), .B1(n354), .Y(n249) );
  OAI211XLTS U749 ( .A0(n267), .A1(n295), .B0(n250), .C0(n249), .Y(n1223) );
  INVX2TS U750 ( .A(n1611), .Y(n263) );
  AOI22X1TS U751 ( .A0(n263), .A1(\destinationAddressbuffer[5][6] ), .B0(n227), 
        .B1(n691), .Y(n252) );
  AOI22X1TS U752 ( .A0(n1468), .A1(n426), .B0(n1752), .B1(n365), .Y(n251) );
  OAI211XLTS U753 ( .A0(n267), .A1(n253), .B0(n252), .C0(n251), .Y(n1179) );
  AOI22X1TS U754 ( .A0(n263), .A1(\destinationAddressbuffer[5][5] ), .B0(n1462), .B1(n672), .Y(n255) );
  AOI22X1TS U755 ( .A0(n1458), .A1(n439), .B0(n1742), .B1(n372), .Y(n254) );
  OAI211XLTS U756 ( .A0(n257), .A1(n256), .B0(n255), .C0(n254), .Y(n1180) );
  AOI22X1TS U757 ( .A0(n263), .A1(\destinationAddressbuffer[5][4] ), .B0(n258), 
        .B1(n659), .Y(n261) );
  AOI22X1TS U758 ( .A0(n259), .A1(n431), .B0(n239), .B1(n380), .Y(n260) );
  OAI211XLTS U759 ( .A0(n1451), .A1(n262), .B0(n261), .C0(n260), .Y(n1181) );
  AOI22X1TS U760 ( .A0(n263), .A1(\destinationAddressbuffer[5][7] ), .B0(n1741), .B1(n706), .Y(n265) );
  INVX2TS U761 ( .A(n1), .Y(n1446) );
  AOI22X1TS U762 ( .A0(n1446), .A1(n435), .B0(n1463), .B1(n360), .Y(n264) );
  OAI211XLTS U763 ( .A0(n267), .A1(n266), .B0(n265), .C0(n264), .Y(n1178) );
  AOI31XLTS U764 ( .A0(n273), .A1(n390), .A2(n392), .B0(n1614), .Y(n272) );
  AOI21X1TS U765 ( .A0(n277), .A1(n272), .B0(n275), .Y(n276) );
  NAND2X1TS U766 ( .A(n276), .B(n1622), .Y(n278) );
  INVX2TS U767 ( .A(n274), .Y(n1420) );
  INVX2TS U768 ( .A(n1420), .Y(n943) );
  CLKBUFX2TS U769 ( .A(n943), .Y(n287) );
  INVX2TS U770 ( .A(n287), .Y(n305) );
  INVX2TS U771 ( .A(n11), .Y(n930) );
  INVX2TS U772 ( .A(n1425), .Y(n291) );
  OR2X1TS U773 ( .A(n1618), .B(n278), .Y(n290) );
  INVX2TS U774 ( .A(n290), .Y(n1436) );
  AOI22X1TS U775 ( .A0(n291), .A1(\destinationAddressbuffer[4][11] ), .B0(
        n1436), .B1(n338), .Y(n282) );
  INVX2TS U776 ( .A(n292), .Y(n297) );
  INVX2TS U777 ( .A(n297), .Y(n1763) );
  INVX2TS U778 ( .A(n4), .Y(n280) );
  AOI22X1TS U779 ( .A0(n1763), .A1(n767), .B0(n280), .B1(n402), .Y(n281) );
  OAI211XLTS U780 ( .A0(n305), .A1(n47), .B0(n282), .C0(n281), .Y(n1162) );
  INVX2TS U781 ( .A(n290), .Y(n283) );
  AOI22X1TS U782 ( .A0(n291), .A1(\destinationAddressbuffer[4][8] ), .B0(n283), 
        .B1(n332), .Y(n286) );
  INVX2TS U783 ( .A(n297), .Y(n284) );
  AOI22X1TS U784 ( .A0(n1773), .A1(n718), .B0(n310), .B1(n419), .Y(n285) );
  OAI211XLTS U785 ( .A0(n305), .A1(n41), .B0(n286), .C0(n285), .Y(n1165) );
  INVX2TS U786 ( .A(n287), .Y(n313) );
  INVX2TS U787 ( .A(n290), .Y(n1782) );
  INVX2TS U788 ( .A(n1782), .Y(n931) );
  INVX2TS U789 ( .A(n931), .Y(n302) );
  AOI22X1TS U790 ( .A0(n291), .A1(\destinationAddressbuffer[4][9] ), .B0(n302), 
        .B1(n345), .Y(n289) );
  INVX2TS U791 ( .A(n297), .Y(n1784) );
  INVX2TS U792 ( .A(n4), .Y(n1783) );
  INVX2TS U793 ( .A(n1783), .Y(n1421) );
  INVX2TS U794 ( .A(n1421), .Y(n933) );
  AOI22X1TS U795 ( .A0(n1784), .A1(n733), .B0(n933), .B1(n412), .Y(n288) );
  OAI211XLTS U796 ( .A0(n313), .A1(n33), .B0(n289), .C0(n288), .Y(n1164) );
  INVX2TS U797 ( .A(n290), .Y(n1771) );
  AOI22X1TS U798 ( .A0(n291), .A1(\destinationAddressbuffer[4][10] ), .B0(
        n1771), .B1(n321), .Y(n294) );
  INVX2TS U799 ( .A(n292), .Y(n1427) );
  INVX2TS U800 ( .A(n1427), .Y(n306) );
  AOI22X1TS U801 ( .A0(n306), .A1(n752), .B0(n280), .B1(n406), .Y(n293) );
  OAI211XLTS U802 ( .A0(n305), .A1(n51), .B0(n294), .C0(n293), .Y(n1163) );
  INVX2TS U803 ( .A(n1623), .Y(n1788) );
  INVX2TS U804 ( .A(n931), .Y(n296) );
  AOI22X1TS U805 ( .A0(n1788), .A1(writeOutbuffer[4]), .B0(n296), .B1(n353), 
        .Y(n299) );
  INVX2TS U806 ( .A(n297), .Y(n1414) );
  INVX2TS U807 ( .A(n4), .Y(n1772) );
  AOI22X1TS U808 ( .A0(n1414), .A1(n546), .B0(n1772), .B1(n422), .Y(n298) );
  OAI211XLTS U809 ( .A0(n313), .A1(n55), .B0(n299), .C0(n298), .Y(n1222) );
  INVX2TS U810 ( .A(n1623), .Y(n309) );
  AOI22X1TS U811 ( .A0(n309), .A1(\destinationAddressbuffer[4][7] ), .B0(n1436), .B1(n359), .Y(n301) );
  AOI22X1TS U812 ( .A0(n306), .A1(n707), .B0(n1772), .B1(n435), .Y(n300) );
  OAI211XLTS U813 ( .A0(n313), .A1(n65), .B0(n301), .C0(n300), .Y(n1166) );
  AOI22X1TS U814 ( .A0(n309), .A1(\destinationAddressbuffer[4][6] ), .B0(n302), 
        .B1(n364), .Y(n304) );
  AOI22X1TS U815 ( .A0(n306), .A1(n693), .B0(n933), .B1(n426), .Y(n303) );
  OAI211XLTS U816 ( .A0(n305), .A1(n70), .B0(n304), .C0(n303), .Y(n1167) );
  AOI22X1TS U817 ( .A0(n309), .A1(\destinationAddressbuffer[4][4] ), .B0(n283), 
        .B1(n377), .Y(n308) );
  AOI22X1TS U818 ( .A0(n306), .A1(n661), .B0(n933), .B1(n431), .Y(n307) );
  OAI211XLTS U819 ( .A0(n1420), .A1(n62), .B0(n308), .C0(n307), .Y(n1169) );
  AOI22X1TS U820 ( .A0(n309), .A1(\destinationAddressbuffer[4][5] ), .B0(n1771), .B1(n371), .Y(n312) );
  INVX2TS U821 ( .A(n1421), .Y(n310) );
  AOI22X1TS U822 ( .A0(n1414), .A1(n673), .B0(n310), .B1(n439), .Y(n311) );
  OAI211XLTS U823 ( .A0(n313), .A1(n73), .B0(n312), .C0(n311), .Y(n1168) );
  AOI31XLTS U824 ( .A0(n19), .A1(n389), .A2(n453), .B0(n1649), .Y(n316) );
  AOI21X1TS U825 ( .A0(n322), .A1(n316), .B0(n318), .Y(n320) );
  NAND2X1TS U826 ( .A(n320), .B(n1657), .Y(n323) );
  INVX2TS U827 ( .A(n317), .Y(n1087) );
  INVX2TS U828 ( .A(n1087), .Y(n1015) );
  CLKBUFX2TS U829 ( .A(n1015), .Y(n337) );
  INVX2TS U830 ( .A(n337), .Y(n370) );
  INVX2TS U831 ( .A(n319), .Y(n1085) );
  INVX2TS U832 ( .A(n1085), .Y(n998) );
  CLKBUFX2TS U833 ( .A(n358), .Y(n1006) );
  INVX2TS U834 ( .A(n1006), .Y(n346) );
  OR2X1TS U835 ( .A(n1653), .B(n323), .Y(n344) );
  INVX2TS U836 ( .A(n344), .Y(n1863) );
  AOI22X1TS U837 ( .A0(n346), .A1(\destinationAddressbuffer[1][10] ), .B0(
        n1863), .B1(n321), .Y(n330) );
  INVX2TS U838 ( .A(n6), .Y(n324) );
  INVX2TS U839 ( .A(n324), .Y(n1000) );
  INVX2TS U840 ( .A(n1000), .Y(n341) );
  INVX2TS U841 ( .A(n326), .Y(n347) );
  AOI22X1TS U842 ( .A0(n341), .A1(n328), .B0(n366), .B1(n327), .Y(n329) );
  OAI211XLTS U843 ( .A0(n370), .A1(n51), .B0(n330), .C0(n329), .Y(n1127) );
  INVX2TS U844 ( .A(n337), .Y(n376) );
  INVX2TS U845 ( .A(n344), .Y(n331) );
  INVX2TS U846 ( .A(n331), .Y(n1014) );
  INVX2TS U847 ( .A(n1014), .Y(n378) );
  AOI22X1TS U848 ( .A0(n346), .A1(\destinationAddressbuffer[1][8] ), .B0(n378), 
        .B1(n332), .Y(n336) );
  INVX2TS U849 ( .A(n326), .Y(n1017) );
  INVX2TS U850 ( .A(n1017), .Y(n366) );
  AOI22X1TS U851 ( .A0(n341), .A1(n334), .B0(n366), .B1(n333), .Y(n335) );
  OAI211XLTS U852 ( .A0(n376), .A1(n41), .B0(n336), .C0(n335), .Y(n1129) );
  INVX2TS U853 ( .A(n344), .Y(n1111) );
  AOI22X1TS U854 ( .A0(n346), .A1(\destinationAddressbuffer[1][11] ), .B0(
        n1111), .B1(n338), .Y(n343) );
  AOI22X1TS U855 ( .A0(n341), .A1(n340), .B0(n326), .B1(n339), .Y(n342) );
  OAI211XLTS U856 ( .A0(n370), .A1(n47), .B0(n343), .C0(n342), .Y(n1126) );
  INVX2TS U857 ( .A(n344), .Y(n1875) );
  AOI22X1TS U858 ( .A0(n346), .A1(\destinationAddressbuffer[1][9] ), .B0(n1875), .B1(n345), .Y(n352) );
  INVX2TS U859 ( .A(n1000), .Y(n1008) );
  INVX2TS U860 ( .A(n347), .Y(n1101) );
  INVX2TS U861 ( .A(n347), .Y(n349) );
  AOI22X1TS U862 ( .A0(n1008), .A1(n350), .B0(n349), .B1(n348), .Y(n351) );
  OAI211XLTS U863 ( .A0(n370), .A1(n33), .B0(n352), .C0(n351), .Y(n1128) );
  INVX2TS U864 ( .A(n358), .Y(n1882) );
  AOI22X1TS U865 ( .A0(n1882), .A1(writeOutbuffer[1]), .B0(n378), .B1(n353), 
        .Y(n357) );
  AOI22X1TS U866 ( .A0(n1102), .A1(n355), .B0(n1342), .B1(n354), .Y(n356) );
  OAI211XLTS U867 ( .A0(n376), .A1(n55), .B0(n357), .C0(n356), .Y(n1219) );
  INVX2TS U868 ( .A(n358), .Y(n379) );
  AOI22X1TS U869 ( .A0(n379), .A1(\destinationAddressbuffer[1][7] ), .B0(n1111), .B1(n359), .Y(n363) );
  INVX2TS U870 ( .A(n6), .Y(n1866) );
  AOI22X1TS U871 ( .A0(n1866), .A1(n361), .B0(n1101), .B1(n360), .Y(n362) );
  OAI211XLTS U872 ( .A0(n376), .A1(n65), .B0(n363), .C0(n362), .Y(n1130) );
  AOI22X1TS U873 ( .A0(n379), .A1(\destinationAddressbuffer[1][6] ), .B0(n331), 
        .B1(n364), .Y(n369) );
  INVX2TS U874 ( .A(n1000), .Y(n1888) );
  AOI22X1TS U875 ( .A0(n1888), .A1(n367), .B0(n366), .B1(n365), .Y(n368) );
  OAI211XLTS U876 ( .A0(n370), .A1(n70), .B0(n369), .C0(n368), .Y(n1131) );
  AOI22X1TS U877 ( .A0(n379), .A1(\destinationAddressbuffer[1][5] ), .B0(n1863), .B1(n371), .Y(n375) );
  INVX2TS U878 ( .A(n347), .Y(n1877) );
  AOI22X1TS U879 ( .A0(n1866), .A1(n373), .B0(n1877), .B1(n372), .Y(n374) );
  OAI211XLTS U880 ( .A0(n376), .A1(n73), .B0(n375), .C0(n374), .Y(n1132) );
  AOI22X1TS U881 ( .A0(n379), .A1(\destinationAddressbuffer[1][4] ), .B0(n378), 
        .B1(n377), .Y(n383) );
  AOI22X1TS U882 ( .A0(n341), .A1(n381), .B0(n326), .B1(n380), .Y(n382) );
  OAI211XLTS U883 ( .A0(n1087), .A1(n62), .B0(n383), .C0(n382), .Y(n1133) );
  AOI31XLTS U884 ( .A0(n390), .A1(n389), .A2(n444), .B0(n1662), .Y(n391) );
  AOI21X1TS U885 ( .A0(n398), .A1(n391), .B0(n452), .Y(n395) );
  NAND2X1TS U886 ( .A(n395), .B(n1671), .Y(n399) );
  INVX2TS U887 ( .A(n394), .Y(n1052) );
  INVX2TS U888 ( .A(n1052), .Y(n1044) );
  CLKBUFX2TS U889 ( .A(n1044), .Y(n410) );
  INVX2TS U890 ( .A(n410), .Y(n434) );
  INVX2TS U891 ( .A(n12), .Y(n1030) );
  INVX2TS U892 ( .A(n425), .Y(n417) );
  OR2X1TS U893 ( .A(n1667), .B(n399), .Y(n415) );
  INVX2TS U894 ( .A(n415), .Y(n396) );
  INVX2TS U895 ( .A(n396), .Y(n1043) );
  INVX2TS U896 ( .A(n1043), .Y(n430) );
  AOI22X1TS U897 ( .A0(n417), .A1(\destinationAddressbuffer[0][11] ), .B0(n430), .B1(n397), .Y(n404) );
  INVX2TS U898 ( .A(n2), .Y(n1076) );
  INVX2TS U899 ( .A(n5), .Y(n401) );
  INVX2TS U900 ( .A(n401), .Y(n1024) );
  INVX2TS U901 ( .A(n1024), .Y(n407) );
  AOI22X1TS U902 ( .A0(n1076), .A1(n767), .B0(n407), .B1(n402), .Y(n403) );
  OAI211XLTS U903 ( .A0(n434), .A1(n47), .B0(n404), .C0(n403), .Y(n1114) );
  INVX2TS U904 ( .A(n415), .Y(n1074) );
  AOI22X1TS U905 ( .A0(n417), .A1(\destinationAddressbuffer[0][10] ), .B0(
        n1074), .B1(n405), .Y(n409) );
  AOI22X1TS U906 ( .A0(n418), .A1(n752), .B0(n407), .B1(n406), .Y(n408) );
  OAI211XLTS U907 ( .A0(n434), .A1(n51), .B0(n409), .C0(n408), .Y(n1115) );
  INVX2TS U908 ( .A(n410), .Y(n442) );
  INVX2TS U909 ( .A(n415), .Y(n1916) );
  AOI22X1TS U910 ( .A0(n417), .A1(\destinationAddressbuffer[0][9] ), .B0(n396), 
        .B1(n411), .Y(n414) );
  INVX2TS U911 ( .A(n2), .Y(n1930) );
  INVX2TS U912 ( .A(n5), .Y(n1918) );
  AOI22X1TS U913 ( .A0(n1930), .A1(n733), .B0(n1918), .B1(n412), .Y(n413) );
  OAI211XLTS U914 ( .A0(n442), .A1(n33), .B0(n414), .C0(n413), .Y(n1116) );
  INVX2TS U915 ( .A(n415), .Y(n1903) );
  AOI22X1TS U916 ( .A0(n417), .A1(\destinationAddressbuffer[0][8] ), .B0(n1903), .B1(n416), .Y(n421) );
  INVX2TS U917 ( .A(n2), .Y(n418) );
  INVX2TS U918 ( .A(n418), .Y(n1046) );
  INVX2TS U919 ( .A(n1046), .Y(n427) );
  INVX2TS U920 ( .A(n5), .Y(n1075) );
  AOI22X1TS U921 ( .A0(n427), .A1(n718), .B0(n1075), .B1(n419), .Y(n420) );
  OAI211XLTS U922 ( .A0(n434), .A1(n41), .B0(n421), .C0(n420), .Y(n1117) );
  INVX2TS U923 ( .A(n425), .Y(n1923) );
  AOI22X1TS U924 ( .A0(n1923), .A1(writeOutbuffer[0]), .B0(n1074), .B1(
        writeIn_WEST), .Y(n424) );
  INVX2TS U925 ( .A(n2), .Y(n1907) );
  INVX2TS U926 ( .A(n5), .Y(n1054) );
  AOI22X1TS U927 ( .A0(n1907), .A1(n546), .B0(n1054), .B1(n422), .Y(n423) );
  OAI211XLTS U928 ( .A0(n442), .A1(n55), .B0(n424), .C0(n423), .Y(n1218) );
  CLKBUFX2TS U929 ( .A(n425), .Y(n1063) );
  INVX2TS U930 ( .A(n1063), .Y(n438) );
  AOI22X1TS U931 ( .A0(n438), .A1(\destinationAddressbuffer[0][6] ), .B0(n1903), .B1(destinationAddressIn_WEST[6]), .Y(n429) );
  AOI22X1TS U932 ( .A0(n427), .A1(n693), .B0(n401), .B1(n426), .Y(n428) );
  OAI211XLTS U933 ( .A0(n442), .A1(n70), .B0(n429), .C0(n428), .Y(n1119) );
  AOI22X1TS U934 ( .A0(n438), .A1(\destinationAddressbuffer[0][4] ), .B0(n430), 
        .B1(destinationAddressIn_WEST[4]), .Y(n433) );
  AOI22X1TS U935 ( .A0(n418), .A1(n661), .B0(n1075), .B1(n431), .Y(n432) );
  OAI211XLTS U936 ( .A0(n434), .A1(n62), .B0(n433), .C0(n432), .Y(n1121) );
  AOI22X1TS U937 ( .A0(n438), .A1(\destinationAddressbuffer[0][7] ), .B0(n430), 
        .B1(destinationAddressIn_WEST[7]), .Y(n437) );
  AOI22X1TS U938 ( .A0(n418), .A1(n707), .B0(n1054), .B1(n435), .Y(n436) );
  OAI211XLTS U939 ( .A0(n1052), .A1(n65), .B0(n437), .C0(n436), .Y(n1118) );
  AOI22X1TS U940 ( .A0(n438), .A1(\destinationAddressbuffer[0][5] ), .B0(n1916), .B1(destinationAddressIn_WEST[5]), .Y(n441) );
  AOI22X1TS U941 ( .A0(n1907), .A1(n673), .B0(n407), .B1(n439), .Y(n440) );
  OAI211XLTS U942 ( .A0(n442), .A1(n73), .B0(n441), .C0(n440), .Y(n1120) );
  INVX2TS U943 ( .A(n1961), .Y(n529) );
  INVX2TS U944 ( .A(n1961), .Y(n526) );
  INVX2TS U945 ( .A(n1955), .Y(n532) );
  NAND2X1TS U946 ( .A(n526), .B(n532), .Y(n530) );
  OAI21XLTS U947 ( .A0(n529), .A1(n1956), .B0(n530), .Y(n504) );
  INVX2TS U948 ( .A(n1952), .Y(n533) );
  INVX2TS U949 ( .A(n1952), .Y(n528) );
  NOR2XLTS U950 ( .A(n530), .B(n528), .Y(n839) );
  CLKBUFX2TS U951 ( .A(n839), .Y(n797) );
  CLKBUFX2TS U952 ( .A(n797), .Y(n816) );
  AOI21X1TS U953 ( .A0(n530), .A1(n533), .B0(n816), .Y(n501) );
  OAI22X1TS U954 ( .A0(n487), .A1(n504), .B0(n444), .B1(n501), .Y(n445) );
  AOI221XLTS U955 ( .A0(n504), .A1(n458), .B0(n446), .B1(n501), .C0(n445), .Y(
        n450) );
  INVX2TS U956 ( .A(n1949), .Y(n447) );
  NAND2X1TS U957 ( .A(n448), .B(n447), .Y(n463) );
  OAI21XLTS U958 ( .A0(n449), .A1(n1961), .B0(n463), .Y(n467) );
  AOI21X1TS U959 ( .A0(n450), .A1(n467), .B0(n1951), .Y(n451) );
  INVX2TS U960 ( .A(reset), .Y(n494) );
  NAND2X1TS U961 ( .A(n494), .B(n1951), .Y(n505) );
  NOR2XLTS U962 ( .A(reset), .B(n452), .Y(n499) );
  INVX2TS U963 ( .A(n1957), .Y(n464) );
  INVX2TS U964 ( .A(n1960), .Y(n454) );
  INVX2TS U965 ( .A(n1953), .Y(n531) );
  AOI22X1TS U966 ( .A0(n454), .A1(n528), .B0(n531), .B1(n453), .Y(n457) );
  INVX2TS U967 ( .A(n456), .Y(n462) );
  INVX2TS U968 ( .A(n477), .Y(n474) );
  AOI21X1TS U969 ( .A0(n529), .A1(n460), .B0(n459), .Y(n473) );
  ADDHXLTS U970 ( .A(n466), .B(n465), .CO(n477), .S(n479) );
  INVX2TS U971 ( .A(n479), .Y(n468) );
  AOI21X1TS U972 ( .A0(n469), .A1(n468), .B0(n467), .Y(n471) );
  OAI22X1TS U973 ( .A0(n469), .A1(n468), .B0(n475), .B1(n474), .Y(n470) );
  AOI21X1TS U974 ( .A0(n478), .A1(n471), .B0(n470), .Y(n472) );
  AOI211X1TS U975 ( .A0(n475), .A1(n474), .B0(n473), .C0(n472), .Y(n476) );
  INVX2TS U976 ( .A(n476), .Y(n480) );
  NAND2X1TS U977 ( .A(n480), .B(n477), .Y(n484) );
  INVX2TS U978 ( .A(n498), .Y(n492) );
  INVX2TS U979 ( .A(n1953), .Y(n527) );
  ADDHXLTS U980 ( .A(n448), .B(n485), .CO(n488), .S(n495) );
  XNOR2X1TS U981 ( .A(n1956), .B(n496), .Y(n489) );
  OAI2BB2XLTS U982 ( .B0(n1963), .B1(n505), .A0N(n499), .A1N(n493), .Y(N2624)
         );
  NAND2X1TS U983 ( .A(n494), .B(n1950), .Y(n503) );
  AOI22X1TS U984 ( .A0(n1949), .A1(n505), .B0(n503), .B1(n447), .Y(n1336) );
  INVX2TS U985 ( .A(n501), .Y(n502) );
  OAI22X1TS U986 ( .A0(n533), .A1(n505), .B0(n502), .B1(n503), .Y(n1331) );
  OAI22X1TS U987 ( .A0(n13), .A1(n505), .B0(n504), .B1(n503), .Y(n1330) );
  CLKBUFX2TS U988 ( .A(readIn_SOUTH), .Y(n1661) );
  CLKBUFX2TS U989 ( .A(n1661), .Y(n1602) );
  CLKBUFX2TS U990 ( .A(n1950), .Y(n845) );
  CLKBUFX2TS U991 ( .A(n545), .Y(n628) );
  CLKBUFX2TS U992 ( .A(n628), .Y(n854) );
  CLKBUFX2TS U993 ( .A(readIn_WEST), .Y(n1669) );
  CLKBUFX2TS U994 ( .A(n1669), .Y(n1655) );
  INVX2TS U995 ( .A(n1950), .Y(n522) );
  NAND2X1TS U996 ( .A(n540), .B(n522), .Y(n510) );
  NOR4XLTS U997 ( .A(n514), .B(n512), .C(n456), .D(n510), .Y(n613) );
  CLKBUFX2TS U998 ( .A(n613), .Y(n629) );
  CLKBUFX2TS U999 ( .A(n629), .Y(n808) );
  CLKBUFX2TS U1000 ( .A(n808), .Y(n566) );
  AOI22X1TS U1001 ( .A0(n1602), .A1(n854), .B0(n1655), .B1(n566), .Y(n543) );
  CLKBUFX2TS U1002 ( .A(readIn_NORTH), .Y(n1660) );
  CLKBUFX2TS U1003 ( .A(n1660), .Y(n1601) );
  CLKBUFX2TS U1004 ( .A(n692), .Y(n627) );
  CLKBUFX2TS U1005 ( .A(n627), .Y(n565) );
  NOR4XLTS U1006 ( .A(selectBit_WEST), .B(n516), .C(n515), .D(n510), .Y(n647)
         );
  CLKBUFX2TS U1007 ( .A(n647), .Y(n778) );
  CLKBUFX2TS U1008 ( .A(n778), .Y(n670) );
  CLKBUFX2TS U1009 ( .A(n670), .Y(n827) );
  AOI22X1TS U1010 ( .A0(n1601), .A1(n565), .B0(readIn_EAST), .B1(n827), .Y(
        n542) );
  NOR3XLTS U1011 ( .A(n512), .B(n511), .C(n456), .Y(n518) );
  NOR3XLTS U1012 ( .A(selectBit_WEST), .B(n516), .C(n515), .Y(n517) );
  OAI31X1TS U1013 ( .A0(n518), .A1(n539), .A2(n517), .B0(n540), .Y(n521) );
  NAND4XLTS U1014 ( .A(n522), .B(n521), .C(n520), .D(n519), .Y(n675) );
  INVX2TS U1015 ( .A(n675), .Y(n523) );
  INVX2TS U1016 ( .A(n523), .Y(n630) );
  INVX2TS U1017 ( .A(n630), .Y(n524) );
  CLKBUFX2TS U1018 ( .A(n1950), .Y(n601) );
  NOR3XLTS U1019 ( .A(n526), .B(n527), .C(n1955), .Y(n720) );
  CLKBUFX2TS U1020 ( .A(n720), .Y(n631) );
  CLKBUFX2TS U1021 ( .A(n631), .Y(n568) );
  NOR3XLTS U1022 ( .A(n529), .B(n1956), .C(n527), .Y(n694) );
  CLKBUFX2TS U1023 ( .A(n694), .Y(n632) );
  CLKBUFX2TS U1024 ( .A(n632), .Y(n567) );
  AOI22X1TS U1025 ( .A0(readOutbuffer[2]), .A1(n568), .B0(readOutbuffer[0]), 
        .B1(n567), .Y(n537) );
  NOR3XLTS U1026 ( .A(n526), .B(n13), .C(n528), .Y(n721) );
  CLKBUFX2TS U1027 ( .A(n721), .Y(n633) );
  CLKBUFX2TS U1028 ( .A(n633), .Y(n570) );
  NOR3XLTS U1029 ( .A(n529), .B(n532), .C(n533), .Y(n695) );
  CLKBUFX2TS U1030 ( .A(n695), .Y(n634) );
  CLKBUFX2TS U1031 ( .A(n634), .Y(n569) );
  AOI22X1TS U1032 ( .A0(readOutbuffer[6]), .A1(n570), .B0(readOutbuffer[4]), 
        .B1(n569), .Y(n536) );
  NOR2XLTS U1033 ( .A(n531), .B(n530), .Y(n722) );
  CLKBUFX2TS U1034 ( .A(n722), .Y(n635) );
  CLKBUFX2TS U1035 ( .A(n635), .Y(n572) );
  NOR3XLTS U1036 ( .A(n532), .B(n531), .C(n1961), .Y(n696) );
  CLKBUFX2TS U1037 ( .A(n696), .Y(n636) );
  CLKBUFX2TS U1038 ( .A(n636), .Y(n571) );
  AOI22X1TS U1039 ( .A0(readOutbuffer[3]), .A1(n572), .B0(readOutbuffer[1]), 
        .B1(n571), .Y(n535) );
  CLKBUFX2TS U1040 ( .A(n839), .Y(n861) );
  NOR3XLTS U1041 ( .A(n1956), .B(n447), .C(n533), .Y(n862) );
  CLKBUFX2TS U1042 ( .A(n862), .Y(n637) );
  CLKBUFX2TS U1043 ( .A(n637), .Y(n573) );
  AOI22X1TS U1044 ( .A0(readOutbuffer[7]), .A1(n861), .B0(readOutbuffer[5]), 
        .B1(n573), .Y(n534) );
  NAND4XLTS U1045 ( .A(n537), .B(n536), .C(n535), .D(n534), .Y(n538) );
  AOI22X1TS U1046 ( .A0(readOut), .A1(n552), .B0(n601), .B1(n538), .Y(n541) );
  CLKBUFX2TS U1047 ( .A(n670), .Y(n750) );
  AOI22X1TS U1048 ( .A0(writeIn_EAST), .A1(n750), .B0(n544), .B1(n566), .Y(
        n555) );
  CLKBUFX2TS U1049 ( .A(n628), .Y(n766) );
  AOI22X1TS U1050 ( .A0(writeIn_NORTH), .A1(n565), .B0(n546), .B1(n766), .Y(
        n554) );
  AOI22X1TS U1051 ( .A0(writeOutbuffer[2]), .A1(n568), .B0(writeOutbuffer[0]), 
        .B1(n567), .Y(n550) );
  AOI22X1TS U1052 ( .A0(writeOutbuffer[6]), .A1(n570), .B0(writeOutbuffer[4]), 
        .B1(n569), .Y(n549) );
  AOI22X1TS U1053 ( .A0(writeOutbuffer[3]), .A1(n572), .B0(writeOutbuffer[1]), 
        .B1(n571), .Y(n548) );
  AOI22X1TS U1054 ( .A0(writeOutbuffer[7]), .A1(n861), .B0(writeOutbuffer[5]), 
        .B1(n573), .Y(n547) );
  NAND4XLTS U1055 ( .A(n550), .B(n549), .C(n548), .D(n547), .Y(n551) );
  AOI22X1TS U1056 ( .A0(writeOut), .A1(n552), .B0(n601), .B1(n551), .Y(n553)
         );
  CLKBUFX2TS U1057 ( .A(requesterAddressIn_NORTH[0]), .Y(n1025) );
  CLKBUFX2TS U1058 ( .A(n1025), .Y(n993) );
  CLKBUFX2TS U1059 ( .A(requesterAddressIn_EAST[0]), .Y(n1023) );
  CLKBUFX2TS U1060 ( .A(n1023), .Y(n992) );
  CLKBUFX2TS U1061 ( .A(n670), .Y(n590) );
  AOI22X1TS U1062 ( .A0(n993), .A1(n565), .B0(n992), .B1(n590), .Y(n564) );
  CLKBUFX2TS U1063 ( .A(requesterAddressIn_SOUTH[0]), .Y(n1026) );
  CLKBUFX2TS U1064 ( .A(n1026), .Y(n994) );
  CLKBUFX2TS U1065 ( .A(n545), .Y(n660) );
  CLKBUFX2TS U1066 ( .A(requesterAddressIn_WEST[0]), .Y(n925) );
  CLKBUFX2TS U1067 ( .A(n925), .Y(n951) );
  AOI22X1TS U1068 ( .A0(n994), .A1(n660), .B0(n951), .B1(n566), .Y(n563) );
  INVX2TS U1069 ( .A(n675), .Y(n702) );
  CLKBUFX2TS U1070 ( .A(n601), .Y(n596) );
  AOI22X1TS U1071 ( .A0(\requesterAddressbuffer[2][0] ), .A1(n568), .B0(
        \requesterAddressbuffer[0][0] ), .B1(n567), .Y(n559) );
  AOI22X1TS U1072 ( .A0(\requesterAddressbuffer[6][0] ), .A1(n570), .B0(
        \requesterAddressbuffer[4][0] ), .B1(n569), .Y(n558) );
  AOI22X1TS U1073 ( .A0(\requesterAddressbuffer[3][0] ), .A1(n572), .B0(
        \requesterAddressbuffer[1][0] ), .B1(n571), .Y(n557) );
  CLKBUFX2TS U1074 ( .A(n797), .Y(n754) );
  CLKBUFX2TS U1075 ( .A(n754), .Y(n602) );
  AOI22X1TS U1076 ( .A0(\requesterAddressbuffer[7][0] ), .A1(n602), .B0(
        \requesterAddressbuffer[5][0] ), .B1(n573), .Y(n556) );
  NAND4XLTS U1077 ( .A(n559), .B(n558), .C(n557), .D(n556), .Y(n560) );
  AOI22X1TS U1078 ( .A0(requesterAddressOut[0]), .A1(n702), .B0(n596), .B1(
        n560), .Y(n562) );
  INVX2TS U1079 ( .A(readRequesterAddress[0]), .Y(n949) );
  INVX2TS U1080 ( .A(n949), .Y(n991) );
  INVX2TS U1081 ( .A(n561), .Y(n597) );
  NAND2X1TS U1082 ( .A(n991), .B(n597), .Y(n608) );
  CLKBUFX2TS U1083 ( .A(requesterAddressIn_NORTH[1]), .Y(n1032) );
  CLKBUFX2TS U1084 ( .A(n1032), .Y(n1001) );
  CLKBUFX2TS U1085 ( .A(requesterAddressIn_EAST[1]), .Y(n1031) );
  CLKBUFX2TS U1086 ( .A(n1031), .Y(n999) );
  AOI22X1TS U1087 ( .A0(n1001), .A1(n565), .B0(n999), .B1(n590), .Y(n581) );
  CLKBUFX2TS U1088 ( .A(requesterAddressIn_SOUTH[1]), .Y(n1033) );
  CLKBUFX2TS U1089 ( .A(n1033), .Y(n1002) );
  CLKBUFX2TS U1090 ( .A(n628), .Y(n809) );
  CLKBUFX2TS U1091 ( .A(requesterAddressIn_WEST[1]), .Y(n932) );
  CLKBUFX2TS U1092 ( .A(n932), .Y(n958) );
  AOI22X1TS U1093 ( .A0(n1002), .A1(n809), .B0(n958), .B1(n566), .Y(n580) );
  AOI22X1TS U1094 ( .A0(\requesterAddressbuffer[2][1] ), .A1(n568), .B0(
        \requesterAddressbuffer[0][1] ), .B1(n567), .Y(n577) );
  AOI22X1TS U1095 ( .A0(\requesterAddressbuffer[6][1] ), .A1(n570), .B0(
        \requesterAddressbuffer[4][1] ), .B1(n569), .Y(n576) );
  AOI22X1TS U1096 ( .A0(\requesterAddressbuffer[3][1] ), .A1(n572), .B0(
        \requesterAddressbuffer[1][1] ), .B1(n571), .Y(n575) );
  AOI22X1TS U1097 ( .A0(\requesterAddressbuffer[7][1] ), .A1(n602), .B0(
        \requesterAddressbuffer[5][1] ), .B1(n573), .Y(n574) );
  NAND4XLTS U1098 ( .A(n577), .B(n576), .C(n575), .D(n574), .Y(n578) );
  AOI22X1TS U1099 ( .A0(requesterAddressOut[1]), .A1(n524), .B0(n596), .B1(
        n578), .Y(n579) );
  INVX2TS U1100 ( .A(readRequesterAddress[1]), .Y(n955) );
  INVX2TS U1101 ( .A(n955), .Y(n1677) );
  NAND2X1TS U1102 ( .A(n1677), .B(n597), .Y(n623) );
  CLKBUFX2TS U1103 ( .A(requesterAddressIn_NORTH[2]), .Y(n1038) );
  CLKBUFX2TS U1104 ( .A(n1038), .Y(n1009) );
  CLKBUFX2TS U1105 ( .A(n627), .Y(n612) );
  CLKBUFX2TS U1106 ( .A(requesterAddressIn_EAST[2]), .Y(n1037) );
  CLKBUFX2TS U1107 ( .A(n1037), .Y(n1007) );
  AOI22X1TS U1108 ( .A0(n1009), .A1(n612), .B0(n1007), .B1(n590), .Y(n589) );
  CLKBUFX2TS U1109 ( .A(requesterAddressIn_SOUTH[2]), .Y(n1039) );
  CLKBUFX2TS U1110 ( .A(n1039), .Y(n1010) );
  CLKBUFX2TS U1111 ( .A(requesterAddressIn_WEST[2]), .Y(n938) );
  CLKBUFX2TS U1112 ( .A(n938), .Y(n963) );
  AOI22X1TS U1113 ( .A0(n1010), .A1(n660), .B0(n963), .B1(n629), .Y(n588) );
  INVX2TS U1114 ( .A(n675), .Y(n745) );
  CLKBUFX2TS U1115 ( .A(n631), .Y(n614) );
  AOI22X1TS U1116 ( .A0(\requesterAddressbuffer[2][2] ), .A1(n614), .B0(
        \requesterAddressbuffer[0][2] ), .B1(n694), .Y(n585) );
  CLKBUFX2TS U1117 ( .A(n633), .Y(n615) );
  AOI22X1TS U1118 ( .A0(\requesterAddressbuffer[6][2] ), .A1(n615), .B0(
        \requesterAddressbuffer[4][2] ), .B1(n695), .Y(n584) );
  CLKBUFX2TS U1119 ( .A(n635), .Y(n616) );
  AOI22X1TS U1120 ( .A0(\requesterAddressbuffer[3][2] ), .A1(n616), .B0(
        \requesterAddressbuffer[1][2] ), .B1(n696), .Y(n583) );
  CLKBUFX2TS U1121 ( .A(n637), .Y(n617) );
  AOI22X1TS U1122 ( .A0(\requesterAddressbuffer[7][2] ), .A1(n602), .B0(
        \requesterAddressbuffer[5][2] ), .B1(n617), .Y(n582) );
  NAND4XLTS U1123 ( .A(n585), .B(n584), .C(n583), .D(n582), .Y(n586) );
  AOI22X1TS U1124 ( .A0(requesterAddressOut[2]), .A1(n745), .B0(n596), .B1(
        n586), .Y(n587) );
  INVX2TS U1125 ( .A(readRequesterAddress[2]), .Y(n962) );
  INVX2TS U1126 ( .A(n962), .Y(n1686) );
  NAND2X1TS U1127 ( .A(n1686), .B(n597), .Y(n643) );
  CLKBUFX2TS U1128 ( .A(requesterAddressIn_NORTH[3]), .Y(n1047) );
  CLKBUFX2TS U1129 ( .A(n1047), .Y(n1018) );
  CLKBUFX2TS U1130 ( .A(requesterAddressIn_EAST[3]), .Y(n1045) );
  CLKBUFX2TS U1131 ( .A(n1045), .Y(n1016) );
  AOI22X1TS U1132 ( .A0(n1018), .A1(n612), .B0(n1016), .B1(n590), .Y(n600) );
  CLKBUFX2TS U1133 ( .A(requesterAddressIn_SOUTH[3]), .Y(n1048) );
  CLKBUFX2TS U1134 ( .A(n1048), .Y(n1019) );
  CLKBUFX2TS U1135 ( .A(requesterAddressIn_WEST[3]), .Y(n944) );
  CLKBUFX2TS U1136 ( .A(n944), .Y(n970) );
  AOI22X1TS U1137 ( .A0(n1019), .A1(n809), .B0(n970), .B1(n613), .Y(n599) );
  AOI22X1TS U1138 ( .A0(\requesterAddressbuffer[2][3] ), .A1(n614), .B0(
        \requesterAddressbuffer[0][3] ), .B1(n694), .Y(n594) );
  AOI22X1TS U1139 ( .A0(\requesterAddressbuffer[6][3] ), .A1(n615), .B0(
        \requesterAddressbuffer[4][3] ), .B1(n695), .Y(n593) );
  AOI22X1TS U1140 ( .A0(\requesterAddressbuffer[3][3] ), .A1(n616), .B0(
        \requesterAddressbuffer[1][3] ), .B1(n696), .Y(n592) );
  CLKBUFX2TS U1141 ( .A(n754), .Y(n648) );
  AOI22X1TS U1142 ( .A0(\requesterAddressbuffer[7][3] ), .A1(n648), .B0(
        \requesterAddressbuffer[5][3] ), .B1(n617), .Y(n591) );
  NAND4XLTS U1143 ( .A(n594), .B(n593), .C(n592), .D(n591), .Y(n595) );
  AOI22X1TS U1144 ( .A0(requesterAddressOut[3]), .A1(n745), .B0(n596), .B1(
        n595), .Y(n598) );
  INVX2TS U1145 ( .A(readRequesterAddress[3]), .Y(n969) );
  INVX2TS U1146 ( .A(n969), .Y(n1695) );
  NAND2X1TS U1147 ( .A(n1695), .B(n597), .Y(n655) );
  CLKBUFX2TS U1148 ( .A(destinationAddressIn_NORTH[0]), .Y(n1702) );
  CLKBUFX2TS U1149 ( .A(destinationAddressIn_EAST[0]), .Y(n1853) );
  CLKBUFX2TS U1150 ( .A(n1853), .Y(n1734) );
  AOI22X1TS U1151 ( .A0(n1702), .A1(n612), .B0(n1734), .B1(n778), .Y(n611) );
  CLKBUFX2TS U1152 ( .A(destinationAddressIn_WEST[0]), .Y(n1893) );
  CLKBUFX2TS U1153 ( .A(n1893), .Y(n1797) );
  AOI22X1TS U1154 ( .A0(destinationAddressIn_SOUTH[0]), .A1(n660), .B0(n1797), 
        .B1(n613), .Y(n610) );
  CLKBUFX2TS U1155 ( .A(n601), .Y(n654) );
  AOI22X1TS U1156 ( .A0(\destinationAddressbuffer[2][0] ), .A1(n614), .B0(
        \destinationAddressbuffer[0][0] ), .B1(n632), .Y(n606) );
  AOI22X1TS U1157 ( .A0(\destinationAddressbuffer[6][0] ), .A1(n615), .B0(
        \destinationAddressbuffer[4][0] ), .B1(n634), .Y(n605) );
  AOI22X1TS U1158 ( .A0(\destinationAddressbuffer[3][0] ), .A1(n616), .B0(
        \destinationAddressbuffer[1][0] ), .B1(n636), .Y(n604) );
  AOI22X1TS U1159 ( .A0(\destinationAddressbuffer[7][0] ), .A1(n602), .B0(
        \destinationAddressbuffer[5][0] ), .B1(n617), .Y(n603) );
  NAND4XLTS U1160 ( .A(n606), .B(n605), .C(n604), .D(n603), .Y(n607) );
  AOI22X1TS U1161 ( .A0(destinationAddressOut[0]), .A1(n745), .B0(n654), .B1(
        n607), .Y(n609) );
  CLKBUFX2TS U1162 ( .A(destinationAddressIn_NORTH[1]), .Y(n1710) );
  CLKBUFX2TS U1163 ( .A(destinationAddressIn_EAST[1]), .Y(n1862) );
  CLKBUFX2TS U1164 ( .A(n1862), .Y(n1739) );
  AOI22X1TS U1165 ( .A0(n1710), .A1(n612), .B0(n1739), .B1(n647), .Y(n626) );
  CLKBUFX2TS U1166 ( .A(destinationAddressIn_WEST[1]), .Y(n1902) );
  CLKBUFX2TS U1167 ( .A(n1902), .Y(n1803) );
  AOI22X1TS U1168 ( .A0(destinationAddressIn_SOUTH[1]), .A1(n809), .B0(n1803), 
        .B1(n613), .Y(n625) );
  AOI22X1TS U1169 ( .A0(\destinationAddressbuffer[2][1] ), .A1(n614), .B0(
        \destinationAddressbuffer[0][1] ), .B1(n632), .Y(n621) );
  AOI22X1TS U1170 ( .A0(\destinationAddressbuffer[6][1] ), .A1(n615), .B0(
        \destinationAddressbuffer[4][1] ), .B1(n634), .Y(n620) );
  AOI22X1TS U1171 ( .A0(\destinationAddressbuffer[3][1] ), .A1(n616), .B0(
        \destinationAddressbuffer[1][1] ), .B1(n636), .Y(n619) );
  AOI22X1TS U1172 ( .A0(\destinationAddressbuffer[7][1] ), .A1(n648), .B0(
        \destinationAddressbuffer[5][1] ), .B1(n617), .Y(n618) );
  NAND4XLTS U1173 ( .A(n621), .B(n620), .C(n619), .D(n618), .Y(n622) );
  AOI22X1TS U1174 ( .A0(destinationAddressOut[1]), .A1(n702), .B0(n654), .B1(
        n622), .Y(n624) );
  CLKBUFX2TS U1175 ( .A(destinationAddressIn_NORTH[2]), .Y(n1719) );
  CLKBUFX2TS U1176 ( .A(n627), .Y(n674) );
  CLKBUFX2TS U1177 ( .A(destinationAddressIn_EAST[2]), .Y(n1873) );
  CLKBUFX2TS U1178 ( .A(n1873), .Y(n1749) );
  AOI22X1TS U1179 ( .A0(n1719), .A1(n674), .B0(n1749), .B1(n647), .Y(n646) );
  CLKBUFX2TS U1180 ( .A(n628), .Y(n790) );
  CLKBUFX2TS U1181 ( .A(destinationAddressIn_WEST[2]), .Y(n1915) );
  CLKBUFX2TS U1182 ( .A(n1915), .Y(n1811) );
  CLKBUFX2TS U1183 ( .A(n629), .Y(n671) );
  AOI22X1TS U1184 ( .A0(destinationAddressIn_SOUTH[2]), .A1(n790), .B0(n1811), 
        .B1(n671), .Y(n645) );
  INVX2TS U1185 ( .A(n630), .Y(n869) );
  CLKBUFX2TS U1186 ( .A(n631), .Y(n677) );
  CLKBUFX2TS U1187 ( .A(n632), .Y(n676) );
  AOI22X1TS U1188 ( .A0(\destinationAddressbuffer[2][2] ), .A1(n677), .B0(
        \destinationAddressbuffer[0][2] ), .B1(n676), .Y(n641) );
  CLKBUFX2TS U1189 ( .A(n633), .Y(n679) );
  CLKBUFX2TS U1190 ( .A(n634), .Y(n678) );
  AOI22X1TS U1191 ( .A0(\destinationAddressbuffer[6][2] ), .A1(n679), .B0(
        \destinationAddressbuffer[4][2] ), .B1(n678), .Y(n640) );
  CLKBUFX2TS U1192 ( .A(n635), .Y(n681) );
  CLKBUFX2TS U1193 ( .A(n636), .Y(n680) );
  AOI22X1TS U1194 ( .A0(\destinationAddressbuffer[3][2] ), .A1(n681), .B0(
        \destinationAddressbuffer[1][2] ), .B1(n680), .Y(n639) );
  CLKBUFX2TS U1195 ( .A(n637), .Y(n682) );
  AOI22X1TS U1196 ( .A0(\destinationAddressbuffer[7][2] ), .A1(n648), .B0(
        \destinationAddressbuffer[5][2] ), .B1(n682), .Y(n638) );
  NAND4XLTS U1197 ( .A(n641), .B(n640), .C(n639), .D(n638), .Y(n642) );
  AOI22X1TS U1198 ( .A0(destinationAddressOut[2]), .A1(n869), .B0(n654), .B1(
        n642), .Y(n644) );
  CLKBUFX2TS U1199 ( .A(destinationAddressIn_NORTH[3]), .Y(n1728) );
  CLKBUFX2TS U1200 ( .A(destinationAddressIn_EAST[3]), .Y(n1884) );
  CLKBUFX2TS U1201 ( .A(n1884), .Y(n1758) );
  AOI22X1TS U1202 ( .A0(n1728), .A1(n674), .B0(n1758), .B1(n647), .Y(n658) );
  CLKBUFX2TS U1203 ( .A(destinationAddressIn_WEST[3]), .Y(n1927) );
  CLKBUFX2TS U1204 ( .A(n1927), .Y(n1819) );
  AOI22X1TS U1205 ( .A0(destinationAddressIn_SOUTH[3]), .A1(n790), .B0(n1819), 
        .B1(n671), .Y(n657) );
  AOI22X1TS U1206 ( .A0(\destinationAddressbuffer[2][3] ), .A1(n677), .B0(
        \destinationAddressbuffer[0][3] ), .B1(n676), .Y(n652) );
  AOI22X1TS U1207 ( .A0(\destinationAddressbuffer[6][3] ), .A1(n679), .B0(
        \destinationAddressbuffer[4][3] ), .B1(n678), .Y(n651) );
  AOI22X1TS U1208 ( .A0(\destinationAddressbuffer[3][3] ), .A1(n681), .B0(
        \destinationAddressbuffer[1][3] ), .B1(n680), .Y(n650) );
  AOI22X1TS U1209 ( .A0(\destinationAddressbuffer[7][3] ), .A1(n648), .B0(
        \destinationAddressbuffer[5][3] ), .B1(n682), .Y(n649) );
  NAND4XLTS U1210 ( .A(n652), .B(n651), .C(n650), .D(n649), .Y(n653) );
  AOI22X1TS U1211 ( .A0(destinationAddressOut[3]), .A1(n524), .B0(n654), .B1(
        n653), .Y(n656) );
  AOI22X1TS U1212 ( .A0(destinationAddressIn_EAST[4]), .A1(n750), .B0(n659), 
        .B1(n671), .Y(n669) );
  AOI22X1TS U1213 ( .A0(destinationAddressIn_NORTH[4]), .A1(n674), .B0(n661), 
        .B1(n660), .Y(n668) );
  INVX2TS U1214 ( .A(n1951), .Y(n769) );
  CLKBUFX2TS U1215 ( .A(n769), .Y(n868) );
  AOI22X1TS U1216 ( .A0(\destinationAddressbuffer[2][4] ), .A1(n677), .B0(
        \destinationAddressbuffer[0][4] ), .B1(n676), .Y(n665) );
  AOI22X1TS U1217 ( .A0(\destinationAddressbuffer[6][4] ), .A1(n679), .B0(
        \destinationAddressbuffer[4][4] ), .B1(n678), .Y(n664) );
  AOI22X1TS U1218 ( .A0(\destinationAddressbuffer[3][4] ), .A1(n681), .B0(
        \destinationAddressbuffer[1][4] ), .B1(n680), .Y(n663) );
  CLKBUFX2TS U1219 ( .A(n754), .Y(n708) );
  AOI22X1TS U1220 ( .A0(\destinationAddressbuffer[7][4] ), .A1(n708), .B0(
        \destinationAddressbuffer[5][4] ), .B1(n682), .Y(n662) );
  NAND4XLTS U1221 ( .A(n665), .B(n664), .C(n663), .D(n662), .Y(n666) );
  AOI22X1TS U1222 ( .A0(destinationAddressOut[4]), .A1(n702), .B0(n868), .B1(
        n666), .Y(n667) );
  CLKBUFX2TS U1223 ( .A(n670), .Y(n765) );
  AOI22X1TS U1224 ( .A0(destinationAddressIn_EAST[5]), .A1(n765), .B0(n672), 
        .B1(n671), .Y(n690) );
  CLKBUFX2TS U1225 ( .A(n545), .Y(n751) );
  AOI22X1TS U1226 ( .A0(destinationAddressIn_NORTH[5]), .A1(n674), .B0(n673), 
        .B1(n751), .Y(n689) );
  INVX2TS U1227 ( .A(n675), .Y(n834) );
  AOI22X1TS U1228 ( .A0(\destinationAddressbuffer[2][5] ), .A1(n677), .B0(
        \destinationAddressbuffer[0][5] ), .B1(n676), .Y(n686) );
  AOI22X1TS U1229 ( .A0(\destinationAddressbuffer[6][5] ), .A1(n679), .B0(
        \destinationAddressbuffer[4][5] ), .B1(n678), .Y(n685) );
  AOI22X1TS U1230 ( .A0(\destinationAddressbuffer[3][5] ), .A1(n681), .B0(
        \destinationAddressbuffer[1][5] ), .B1(n680), .Y(n684) );
  AOI22X1TS U1231 ( .A0(\destinationAddressbuffer[7][5] ), .A1(n708), .B0(
        \destinationAddressbuffer[5][5] ), .B1(n682), .Y(n683) );
  NAND4XLTS U1232 ( .A(n686), .B(n685), .C(n684), .D(n683), .Y(n687) );
  AOI22X1TS U1233 ( .A0(destinationAddressOut[5]), .A1(n834), .B0(n868), .B1(
        n687), .Y(n688) );
  CLKBUFX2TS U1234 ( .A(n808), .Y(n731) );
  AOI22X1TS U1235 ( .A0(destinationAddressIn_EAST[6]), .A1(n765), .B0(n691), 
        .B1(n731), .Y(n705) );
  CLKBUFX2TS U1236 ( .A(n692), .Y(n734) );
  AOI22X1TS U1237 ( .A0(destinationAddressIn_NORTH[6]), .A1(n734), .B0(n693), 
        .B1(n751), .Y(n704) );
  CLKBUFX2TS U1238 ( .A(n694), .Y(n810) );
  CLKBUFX2TS U1239 ( .A(n810), .Y(n736) );
  AOI22X1TS U1240 ( .A0(\destinationAddressbuffer[2][6] ), .A1(n720), .B0(
        \destinationAddressbuffer[0][6] ), .B1(n736), .Y(n700) );
  CLKBUFX2TS U1241 ( .A(n695), .Y(n812) );
  CLKBUFX2TS U1242 ( .A(n812), .Y(n737) );
  AOI22X1TS U1243 ( .A0(\destinationAddressbuffer[6][6] ), .A1(n721), .B0(
        \destinationAddressbuffer[4][6] ), .B1(n737), .Y(n699) );
  CLKBUFX2TS U1244 ( .A(n696), .Y(n814) );
  CLKBUFX2TS U1245 ( .A(n814), .Y(n738) );
  AOI22X1TS U1246 ( .A0(\destinationAddressbuffer[3][6] ), .A1(n722), .B0(
        \destinationAddressbuffer[1][6] ), .B1(n738), .Y(n698) );
  CLKBUFX2TS U1247 ( .A(n862), .Y(n828) );
  CLKBUFX2TS U1248 ( .A(n828), .Y(n739) );
  AOI22X1TS U1249 ( .A0(\destinationAddressbuffer[7][6] ), .A1(n708), .B0(
        \destinationAddressbuffer[5][6] ), .B1(n739), .Y(n697) );
  NAND4XLTS U1250 ( .A(n700), .B(n699), .C(n698), .D(n697), .Y(n701) );
  AOI22X1TS U1251 ( .A0(destinationAddressOut[6]), .A1(n702), .B0(n868), .B1(
        n701), .Y(n703) );
  AOI22X1TS U1252 ( .A0(destinationAddressIn_EAST[7]), .A1(n827), .B0(n706), 
        .B1(n731), .Y(n716) );
  AOI22X1TS U1253 ( .A0(destinationAddressIn_NORTH[7]), .A1(n734), .B0(n707), 
        .B1(n766), .Y(n715) );
  CLKBUFX2TS U1254 ( .A(n769), .Y(n760) );
  AOI22X1TS U1255 ( .A0(\destinationAddressbuffer[2][7] ), .A1(n720), .B0(
        \destinationAddressbuffer[0][7] ), .B1(n736), .Y(n712) );
  AOI22X1TS U1256 ( .A0(\destinationAddressbuffer[6][7] ), .A1(n721), .B0(
        \destinationAddressbuffer[4][7] ), .B1(n737), .Y(n711) );
  AOI22X1TS U1257 ( .A0(\destinationAddressbuffer[3][7] ), .A1(n722), .B0(
        \destinationAddressbuffer[1][7] ), .B1(n738), .Y(n710) );
  AOI22X1TS U1258 ( .A0(\destinationAddressbuffer[7][7] ), .A1(n708), .B0(
        \destinationAddressbuffer[5][7] ), .B1(n739), .Y(n709) );
  NAND4XLTS U1259 ( .A(n712), .B(n711), .C(n710), .D(n709), .Y(n713) );
  AOI22X1TS U1260 ( .A0(destinationAddressOut[7]), .A1(n523), .B0(n760), .B1(
        n713), .Y(n714) );
  AOI22X1TS U1261 ( .A0(destinationAddressIn_EAST[8]), .A1(n750), .B0(n717), 
        .B1(n731), .Y(n730) );
  AOI22X1TS U1262 ( .A0(n719), .A1(n734), .B0(n718), .B1(n751), .Y(n729) );
  CLKBUFX2TS U1263 ( .A(n720), .Y(n811) );
  AOI22X1TS U1264 ( .A0(\destinationAddressbuffer[2][8] ), .A1(n811), .B0(
        \destinationAddressbuffer[0][8] ), .B1(n736), .Y(n726) );
  CLKBUFX2TS U1265 ( .A(n721), .Y(n813) );
  AOI22X1TS U1266 ( .A0(\destinationAddressbuffer[6][8] ), .A1(n813), .B0(
        \destinationAddressbuffer[4][8] ), .B1(n737), .Y(n725) );
  CLKBUFX2TS U1267 ( .A(n722), .Y(n815) );
  AOI22X1TS U1268 ( .A0(\destinationAddressbuffer[3][8] ), .A1(n815), .B0(
        \destinationAddressbuffer[1][8] ), .B1(n738), .Y(n724) );
  AOI22X1TS U1269 ( .A0(\destinationAddressbuffer[7][8] ), .A1(n816), .B0(
        \destinationAddressbuffer[5][8] ), .B1(n739), .Y(n723) );
  NAND4XLTS U1270 ( .A(n726), .B(n725), .C(n724), .D(n723), .Y(n727) );
  AOI22X1TS U1271 ( .A0(destinationAddressOut[8]), .A1(n869), .B0(n760), .B1(
        n727), .Y(n728) );
  AOI22X1TS U1272 ( .A0(destinationAddressIn_EAST[9]), .A1(n765), .B0(n732), 
        .B1(n731), .Y(n748) );
  AOI22X1TS U1273 ( .A0(n735), .A1(n734), .B0(n733), .B1(n766), .Y(n747) );
  AOI22X1TS U1274 ( .A0(\destinationAddressbuffer[2][9] ), .A1(n811), .B0(
        \destinationAddressbuffer[0][9] ), .B1(n736), .Y(n743) );
  AOI22X1TS U1275 ( .A0(\destinationAddressbuffer[6][9] ), .A1(n813), .B0(
        \destinationAddressbuffer[4][9] ), .B1(n737), .Y(n742) );
  AOI22X1TS U1276 ( .A0(\destinationAddressbuffer[3][9] ), .A1(n815), .B0(
        \destinationAddressbuffer[1][9] ), .B1(n738), .Y(n741) );
  AOI22X1TS U1277 ( .A0(\destinationAddressbuffer[7][9] ), .A1(n816), .B0(
        \destinationAddressbuffer[5][9] ), .B1(n739), .Y(n740) );
  NAND4XLTS U1278 ( .A(n743), .B(n742), .C(n741), .D(n740), .Y(n744) );
  AOI22X1TS U1279 ( .A0(destinationAddressOut[9]), .A1(n745), .B0(n760), .B1(
        n744), .Y(n746) );
  CLKBUFX2TS U1280 ( .A(n808), .Y(n789) );
  AOI22X1TS U1281 ( .A0(destinationAddressIn_EAST[10]), .A1(n750), .B0(n749), 
        .B1(n789), .Y(n763) );
  CLKBUFX2TS U1282 ( .A(n692), .Y(n788) );
  AOI22X1TS U1283 ( .A0(n753), .A1(n788), .B0(n752), .B1(n751), .Y(n762) );
  CLKBUFX2TS U1284 ( .A(n811), .Y(n791) );
  CLKBUFX2TS U1285 ( .A(n810), .Y(n792) );
  AOI22X1TS U1286 ( .A0(\destinationAddressbuffer[2][10] ), .A1(n791), .B0(
        \destinationAddressbuffer[0][10] ), .B1(n792), .Y(n758) );
  CLKBUFX2TS U1287 ( .A(n813), .Y(n793) );
  CLKBUFX2TS U1288 ( .A(n812), .Y(n794) );
  AOI22X1TS U1289 ( .A0(\destinationAddressbuffer[6][10] ), .A1(n793), .B0(
        \destinationAddressbuffer[4][10] ), .B1(n794), .Y(n757) );
  CLKBUFX2TS U1290 ( .A(n815), .Y(n795) );
  CLKBUFX2TS U1291 ( .A(n814), .Y(n796) );
  AOI22X1TS U1292 ( .A0(\destinationAddressbuffer[3][10] ), .A1(n795), .B0(
        \destinationAddressbuffer[1][10] ), .B1(n796), .Y(n756) );
  CLKBUFX2TS U1293 ( .A(n828), .Y(n798) );
  AOI22X1TS U1294 ( .A0(\destinationAddressbuffer[7][10] ), .A1(n754), .B0(
        \destinationAddressbuffer[5][10] ), .B1(n798), .Y(n755) );
  NAND4XLTS U1295 ( .A(n758), .B(n757), .C(n756), .D(n755), .Y(n759) );
  AOI22X1TS U1296 ( .A0(destinationAddressOut[10]), .A1(n869), .B0(n760), .B1(
        n759), .Y(n761) );
  AOI22X1TS U1297 ( .A0(destinationAddressIn_EAST[11]), .A1(n765), .B0(n764), 
        .B1(n789), .Y(n777) );
  AOI22X1TS U1298 ( .A0(n768), .A1(n788), .B0(n767), .B1(n766), .Y(n776) );
  CLKBUFX2TS U1299 ( .A(n769), .Y(n822) );
  AOI22X1TS U1300 ( .A0(\destinationAddressbuffer[2][11] ), .A1(n791), .B0(
        \destinationAddressbuffer[0][11] ), .B1(n792), .Y(n773) );
  AOI22X1TS U1301 ( .A0(\destinationAddressbuffer[6][11] ), .A1(n793), .B0(
        \destinationAddressbuffer[4][11] ), .B1(n794), .Y(n772) );
  AOI22X1TS U1302 ( .A0(\destinationAddressbuffer[3][11] ), .A1(n795), .B0(
        \destinationAddressbuffer[1][11] ), .B1(n796), .Y(n771) );
  AOI22X1TS U1303 ( .A0(\destinationAddressbuffer[7][11] ), .A1(n797), .B0(
        \destinationAddressbuffer[5][11] ), .B1(n798), .Y(n770) );
  NAND4XLTS U1304 ( .A(n773), .B(n772), .C(n771), .D(n770), .Y(n774) );
  AOI22X1TS U1305 ( .A0(destinationAddressOut[11]), .A1(n523), .B0(n822), .B1(
        n774), .Y(n775) );
  CLKBUFX2TS U1306 ( .A(dataIn_NORTH[0]), .Y(n1088) );
  CLKBUFX2TS U1307 ( .A(dataIn_EAST[0]), .Y(n1477) );
  CLKBUFX2TS U1308 ( .A(n1477), .Y(n1347) );
  CLKBUFX2TS U1309 ( .A(n778), .Y(n851) );
  AOI22X1TS U1310 ( .A0(n1088), .A1(n788), .B0(n1347), .B1(n851), .Y(n787) );
  CLKBUFX2TS U1311 ( .A(dataIn_WEST[0]), .Y(n1413) );
  CLKBUFX2TS U1312 ( .A(n1413), .Y(n1053) );
  AOI22X1TS U1313 ( .A0(dataIn_SOUTH[0]), .A1(n790), .B0(n1053), .B1(n789), 
        .Y(n786) );
  AOI22X1TS U1314 ( .A0(\dataoutbuffer[0][0] ), .A1(n792), .B0(
        \dataoutbuffer[2][0] ), .B1(n791), .Y(n782) );
  AOI22X1TS U1315 ( .A0(\dataoutbuffer[4][0] ), .A1(n794), .B0(
        \dataoutbuffer[6][0] ), .B1(n793), .Y(n781) );
  AOI22X1TS U1316 ( .A0(\dataoutbuffer[1][0] ), .A1(n796), .B0(
        \dataoutbuffer[3][0] ), .B1(n795), .Y(n780) );
  AOI22X1TS U1317 ( .A0(\dataoutbuffer[5][0] ), .A1(n798), .B0(
        \dataoutbuffer[7][0] ), .B1(n861), .Y(n779) );
  NAND4XLTS U1318 ( .A(n782), .B(n781), .C(n780), .D(n779), .Y(n783) );
  AOI22X1TS U1319 ( .A0(dataOut[0]), .A1(n524), .B0(n822), .B1(n783), .Y(n785)
         );
  INVX2TS U1320 ( .A(cacheDataOut[0]), .Y(n1086) );
  INVX2TS U1321 ( .A(n561), .Y(n846) );
  NAND2X1TS U1322 ( .A(cacheDataOut[0]), .B(n846), .Y(n784) );
  CLKBUFX2TS U1323 ( .A(dataIn_NORTH[1]), .Y(n1094) );
  CLKBUFX2TS U1324 ( .A(dataIn_EAST[1]), .Y(n1486) );
  CLKBUFX2TS U1325 ( .A(n1486), .Y(n1352) );
  AOI22X1TS U1326 ( .A0(n1094), .A1(n788), .B0(n1352), .B1(n827), .Y(n807) );
  CLKBUFX2TS U1327 ( .A(dataIn_WEST[1]), .Y(n1419) );
  CLKBUFX2TS U1328 ( .A(n1419), .Y(n1059) );
  AOI22X1TS U1329 ( .A0(dataIn_SOUTH[1]), .A1(n790), .B0(n1059), .B1(n789), 
        .Y(n806) );
  AOI22X1TS U1330 ( .A0(\dataoutbuffer[0][1] ), .A1(n792), .B0(
        \dataoutbuffer[2][1] ), .B1(n791), .Y(n802) );
  AOI22X1TS U1331 ( .A0(\dataoutbuffer[4][1] ), .A1(n794), .B0(
        \dataoutbuffer[6][1] ), .B1(n793), .Y(n801) );
  AOI22X1TS U1332 ( .A0(\dataoutbuffer[1][1] ), .A1(n796), .B0(
        \dataoutbuffer[3][1] ), .B1(n795), .Y(n800) );
  AOI22X1TS U1333 ( .A0(\dataoutbuffer[5][1] ), .A1(n798), .B0(
        \dataoutbuffer[7][1] ), .B1(n797), .Y(n799) );
  NAND4XLTS U1334 ( .A(n802), .B(n801), .C(n800), .D(n799), .Y(n803) );
  AOI22X1TS U1335 ( .A0(dataOut[1]), .A1(n834), .B0(n822), .B1(n803), .Y(n805)
         );
  INVX2TS U1336 ( .A(cacheDataOut[1]), .Y(n1092) );
  INVX2TS U1337 ( .A(n561), .Y(n870) );
  NAND2X1TS U1338 ( .A(cacheDataOut[1]), .B(n870), .Y(n804) );
  CLKBUFX2TS U1339 ( .A(dataIn_NORTH[2]), .Y(n1100) );
  CLKBUFX2TS U1340 ( .A(n692), .Y(n852) );
  CLKBUFX2TS U1341 ( .A(dataIn_EAST[2]), .Y(n1495) );
  CLKBUFX2TS U1342 ( .A(n1495), .Y(n1358) );
  AOI22X1TS U1343 ( .A0(n1100), .A1(n852), .B0(n1358), .B1(n851), .Y(n826) );
  CLKBUFX2TS U1344 ( .A(dataIn_WEST[2]), .Y(n1426) );
  CLKBUFX2TS U1345 ( .A(n1426), .Y(n1064) );
  CLKBUFX2TS U1346 ( .A(n808), .Y(n853) );
  AOI22X1TS U1347 ( .A0(dataIn_SOUTH[2]), .A1(n809), .B0(n1064), .B1(n853), 
        .Y(n825) );
  CLKBUFX2TS U1348 ( .A(n810), .Y(n856) );
  CLKBUFX2TS U1349 ( .A(n811), .Y(n855) );
  AOI22X1TS U1350 ( .A0(\dataoutbuffer[0][2] ), .A1(n856), .B0(
        \dataoutbuffer[2][2] ), .B1(n855), .Y(n820) );
  CLKBUFX2TS U1351 ( .A(n812), .Y(n858) );
  CLKBUFX2TS U1352 ( .A(n813), .Y(n857) );
  AOI22X1TS U1353 ( .A0(\dataoutbuffer[4][2] ), .A1(n858), .B0(
        \dataoutbuffer[6][2] ), .B1(n857), .Y(n819) );
  CLKBUFX2TS U1354 ( .A(n814), .Y(n860) );
  CLKBUFX2TS U1355 ( .A(n815), .Y(n859) );
  AOI22X1TS U1356 ( .A0(\dataoutbuffer[1][2] ), .A1(n860), .B0(
        \dataoutbuffer[3][2] ), .B1(n859), .Y(n818) );
  AOI22X1TS U1357 ( .A0(\dataoutbuffer[5][2] ), .A1(n828), .B0(
        \dataoutbuffer[7][2] ), .B1(n816), .Y(n817) );
  NAND4XLTS U1358 ( .A(n820), .B(n819), .C(n818), .D(n817), .Y(n821) );
  AOI22X1TS U1359 ( .A0(dataOut[2]), .A1(n834), .B0(n822), .B1(n821), .Y(n824)
         );
  INVX2TS U1360 ( .A(cacheDataOut[2]), .Y(n1098) );
  NAND2X1TS U1361 ( .A(cacheDataOut[2]), .B(n846), .Y(n823) );
  CLKBUFX2TS U1362 ( .A(dataIn_NORTH[3]), .Y(n1107) );
  CLKBUFX2TS U1363 ( .A(dataIn_EAST[3]), .Y(n1504) );
  CLKBUFX2TS U1364 ( .A(n1504), .Y(n1364) );
  AOI22X1TS U1365 ( .A0(n1107), .A1(n852), .B0(n1364), .B1(n827), .Y(n838) );
  CLKBUFX2TS U1366 ( .A(dataIn_WEST[3]), .Y(n1431) );
  CLKBUFX2TS U1367 ( .A(n1431), .Y(n1069) );
  AOI22X1TS U1368 ( .A0(dataIn_SOUTH[3]), .A1(n854), .B0(n1069), .B1(n853), 
        .Y(n837) );
  AOI22X1TS U1369 ( .A0(\dataoutbuffer[0][3] ), .A1(n856), .B0(
        \dataoutbuffer[2][3] ), .B1(n855), .Y(n832) );
  AOI22X1TS U1370 ( .A0(\dataoutbuffer[4][3] ), .A1(n858), .B0(
        \dataoutbuffer[6][3] ), .B1(n857), .Y(n831) );
  AOI22X1TS U1371 ( .A0(\dataoutbuffer[1][3] ), .A1(n860), .B0(
        \dataoutbuffer[3][3] ), .B1(n859), .Y(n830) );
  AOI22X1TS U1372 ( .A0(\dataoutbuffer[5][3] ), .A1(n828), .B0(
        \dataoutbuffer[7][3] ), .B1(n839), .Y(n829) );
  NAND4XLTS U1373 ( .A(n832), .B(n831), .C(n830), .D(n829), .Y(n833) );
  AOI22X1TS U1374 ( .A0(dataOut[3]), .A1(n834), .B0(n845), .B1(n833), .Y(n836)
         );
  INVX2TS U1375 ( .A(cacheDataOut[3]), .Y(n1106) );
  NAND2X1TS U1376 ( .A(cacheDataOut[3]), .B(n870), .Y(n835) );
  CLKBUFX2TS U1377 ( .A(dataIn_NORTH[4]), .Y(n1112) );
  CLKBUFX2TS U1378 ( .A(dataIn_EAST[4]), .Y(n1510) );
  CLKBUFX2TS U1379 ( .A(n1510), .Y(n1369) );
  AOI22X1TS U1380 ( .A0(n1112), .A1(n852), .B0(n1369), .B1(n851), .Y(n850) );
  CLKBUFX2TS U1381 ( .A(dataIn_WEST[4]), .Y(n1435) );
  CLKBUFX2TS U1382 ( .A(n1435), .Y(n1073) );
  AOI22X1TS U1383 ( .A0(dataIn_SOUTH[4]), .A1(n854), .B0(n1073), .B1(n853), 
        .Y(n849) );
  AOI22X1TS U1384 ( .A0(\dataoutbuffer[0][4] ), .A1(n856), .B0(
        \dataoutbuffer[2][4] ), .B1(n855), .Y(n843) );
  AOI22X1TS U1385 ( .A0(\dataoutbuffer[4][4] ), .A1(n858), .B0(
        \dataoutbuffer[6][4] ), .B1(n857), .Y(n842) );
  AOI22X1TS U1386 ( .A0(\dataoutbuffer[1][4] ), .A1(n860), .B0(
        \dataoutbuffer[3][4] ), .B1(n859), .Y(n841) );
  AOI22X1TS U1387 ( .A0(\dataoutbuffer[5][4] ), .A1(n862), .B0(
        \dataoutbuffer[7][4] ), .B1(n839), .Y(n840) );
  NAND4XLTS U1388 ( .A(n843), .B(n842), .C(n841), .D(n840), .Y(n844) );
  AOI22X1TS U1389 ( .A0(dataOut[4]), .A1(n524), .B0(n845), .B1(n844), .Y(n848)
         );
  INVX2TS U1390 ( .A(cacheDataOut[4]), .Y(n1401) );
  NAND2X1TS U1391 ( .A(cacheDataOut[4]), .B(n846), .Y(n847) );
  CLKBUFX2TS U1392 ( .A(dataIn_NORTH[5]), .Y(n1341) );
  CLKBUFX2TS U1393 ( .A(dataIn_EAST[5]), .Y(n1518) );
  CLKBUFX2TS U1394 ( .A(n1518), .Y(n1377) );
  AOI22X1TS U1395 ( .A0(n1341), .A1(n852), .B0(n1377), .B1(n851), .Y(n874) );
  CLKBUFX2TS U1396 ( .A(dataIn_WEST[5]), .Y(n1441) );
  CLKBUFX2TS U1397 ( .A(n1441), .Y(n1081) );
  AOI22X1TS U1398 ( .A0(dataIn_SOUTH[5]), .A1(n854), .B0(n1081), .B1(n853), 
        .Y(n873) );
  AOI22X1TS U1399 ( .A0(\dataoutbuffer[0][5] ), .A1(n856), .B0(
        \dataoutbuffer[2][5] ), .B1(n855), .Y(n866) );
  AOI22X1TS U1400 ( .A0(\dataoutbuffer[4][5] ), .A1(n858), .B0(
        \dataoutbuffer[6][5] ), .B1(n857), .Y(n865) );
  AOI22X1TS U1401 ( .A0(\dataoutbuffer[1][5] ), .A1(n860), .B0(
        \dataoutbuffer[3][5] ), .B1(n859), .Y(n864) );
  AOI22X1TS U1402 ( .A0(\dataoutbuffer[5][5] ), .A1(n862), .B0(
        \dataoutbuffer[7][5] ), .B1(n861), .Y(n863) );
  NAND4XLTS U1403 ( .A(n866), .B(n865), .C(n864), .D(n863), .Y(n867) );
  AOI22X1TS U1404 ( .A0(dataOut[5]), .A1(n869), .B0(n868), .B1(n867), .Y(n872)
         );
  INVX2TS U1405 ( .A(cacheDataOut[5]), .Y(n1406) );
  NAND2X1TS U1406 ( .A(cacheDataOut[5]), .B(n870), .Y(n871) );
  INVX2TS U1407 ( .A(n949), .Y(n1796) );
  INVX2TS U1408 ( .A(n1587), .Y(n1685) );
  AOI22X1TS U1409 ( .A0(n1796), .A1(n1673), .B0(n1685), .B1(
        \requesterAddressbuffer[7][0] ), .Y(n878) );
  INVX2TS U1410 ( .A(n887), .Y(n1679) );
  AOI22X1TS U1411 ( .A0(n1680), .A1(n951), .B0(n1679), .B1(
        requesterAddressIn_EAST[0]), .Y(n877) );
  CLKBUFX2TS U1412 ( .A(n1026), .Y(n926) );
  INVX2TS U1413 ( .A(n875), .Y(n1697) );
  AOI22X1TS U1414 ( .A0(n1538), .A1(n926), .B0(n1697), .B1(n993), .Y(n876) );
  INVX2TS U1415 ( .A(n886), .Y(n1678) );
  AOI22X1TS U1416 ( .A0(n1678), .A1(n1677), .B0(n1694), .B1(
        \requesterAddressbuffer[7][1] ), .Y(n882) );
  INVX2TS U1417 ( .A(n879), .Y(n1552) );
  AOI22X1TS U1418 ( .A0(n1552), .A1(n958), .B0(n1679), .B1(
        requesterAddressIn_EAST[1]), .Y(n881) );
  CLKBUFX2TS U1419 ( .A(n1033), .Y(n934) );
  AOI22X1TS U1420 ( .A0(n888), .A1(n934), .B0(n48), .B1(n1001), .Y(n880) );
  INVX2TS U1421 ( .A(n1587), .Y(n1533) );
  AOI22X1TS U1422 ( .A0(n34), .A1(n1686), .B0(n1533), .B1(
        \requesterAddressbuffer[7][2] ), .Y(n885) );
  INVX2TS U1423 ( .A(n887), .Y(n1687) );
  AOI22X1TS U1424 ( .A0(n1552), .A1(n963), .B0(n1687), .B1(
        requesterAddressIn_EAST[2]), .Y(n884) );
  CLKBUFX2TS U1425 ( .A(n1039), .Y(n939) );
  AOI22X1TS U1426 ( .A0(n1563), .A1(n939), .B0(n1697), .B1(n1009), .Y(n883) );
  INVX2TS U1427 ( .A(n886), .Y(n1696) );
  AOI22X1TS U1428 ( .A0(n1696), .A1(n1695), .B0(n1533), .B1(
        \requesterAddressbuffer[7][3] ), .Y(n891) );
  AOI22X1TS U1429 ( .A0(n1526), .A1(n970), .B0(n1569), .B1(
        requesterAddressIn_EAST[3]), .Y(n890) );
  CLKBUFX2TS U1430 ( .A(n1048), .Y(n945) );
  AOI22X1TS U1431 ( .A0(n888), .A1(n945), .B0(n1681), .B1(n1018), .Y(n889) );
  INVX2TS U1432 ( .A(n949), .Y(n1852) );
  INVX2TS U1433 ( .A(n1493), .Y(n1716) );
  AOI22X1TS U1434 ( .A0(n1852), .A1(n895), .B0(n1716), .B1(
        \requesterAddressbuffer[6][0] ), .Y(n894) );
  INVX2TS U1435 ( .A(n1485), .Y(n1708) );
  AOI22X1TS U1436 ( .A0(n925), .A1(n1496), .B0(n1023), .B1(n1708), .Y(n893) );
  AOI22X1TS U1437 ( .A0(n926), .A1(n1498), .B0(n993), .B1(n1712), .Y(n892) );
  INVX2TS U1438 ( .A(n955), .Y(n1768) );
  AOI22X1TS U1439 ( .A0(n1768), .A1(n895), .B0(n1725), .B1(
        \requesterAddressbuffer[6][1] ), .Y(n900) );
  INVX2TS U1440 ( .A(n896), .Y(n1727) );
  INVX2TS U1441 ( .A(n1485), .Y(n1718) );
  AOI22X1TS U1442 ( .A0(n932), .A1(n1727), .B0(n1031), .B1(n1718), .Y(n899) );
  INVX2TS U1443 ( .A(n897), .Y(n1703) );
  AOI22X1TS U1444 ( .A0(n934), .A1(n1703), .B0(n1001), .B1(n1730), .Y(n898) );
  INVX2TS U1445 ( .A(n962), .Y(n1779) );
  INVX2TS U1446 ( .A(n9), .Y(n1707) );
  INVX2TS U1447 ( .A(n1598), .Y(n1483) );
  AOI22X1TS U1448 ( .A0(n1779), .A1(n1707), .B0(n1483), .B1(
        \requesterAddressbuffer[6][2] ), .Y(n904) );
  AOI22X1TS U1449 ( .A0(n938), .A1(n116), .B0(n1037), .B1(n905), .Y(n903) );
  AOI22X1TS U1450 ( .A0(n939), .A1(n1711), .B0(n1009), .B1(n901), .Y(n902) );
  INVX2TS U1451 ( .A(n969), .Y(n1790) );
  INVX2TS U1452 ( .A(n9), .Y(n1717) );
  AOI22X1TS U1453 ( .A0(n1790), .A1(n1717), .B0(n1483), .B1(
        \requesterAddressbuffer[6][3] ), .Y(n908) );
  AOI22X1TS U1454 ( .A0(n944), .A1(n98), .B0(n1045), .B1(n905), .Y(n907) );
  AOI22X1TS U1455 ( .A0(n945), .A1(n1720), .B0(n1018), .B1(n1513), .Y(n906) );
  INVX2TS U1456 ( .A(n1456), .Y(n1747) );
  AOI22X1TS U1457 ( .A0(n991), .A1(n913), .B0(n1747), .B1(
        \requesterAddressbuffer[5][0] ), .Y(n912) );
  INVX2TS U1458 ( .A(n1451), .Y(n1740) );
  AOI22X1TS U1459 ( .A0(n925), .A1(n1457), .B0(n1023), .B1(n1740), .Y(n911) );
  INVX2TS U1460 ( .A(n909), .Y(n1752) );
  AOI22X1TS U1461 ( .A0(n926), .A1(n1752), .B0(requesterAddressIn_NORTH[0]), 
        .B1(n1446), .Y(n910) );
  AOI22X1TS U1462 ( .A0(n1677), .A1(n913), .B0(n1757), .B1(
        \requesterAddressbuffer[5][1] ), .Y(n916) );
  INVX2TS U1463 ( .A(n1451), .Y(n1750) );
  AOI22X1TS U1464 ( .A0(n932), .A1(n1751), .B0(n1031), .B1(n1750), .Y(n915) );
  AOI22X1TS U1465 ( .A0(n934), .A1(n1467), .B0(requesterAddressIn_NORTH[1]), 
        .B1(n1468), .Y(n914) );
  INVX2TS U1466 ( .A(n1445), .Y(n1738) );
  INVX2TS U1467 ( .A(n1611), .Y(n1450) );
  AOI22X1TS U1468 ( .A0(n1686), .A1(n1738), .B0(n1450), .B1(
        \requesterAddressbuffer[5][2] ), .Y(n919) );
  AOI22X1TS U1469 ( .A0(n938), .A1(n1462), .B0(n1037), .B1(n921), .Y(n918) );
  AOI22X1TS U1470 ( .A0(n939), .A1(n1463), .B0(requesterAddressIn_NORTH[2]), 
        .B1(n1468), .Y(n917) );
  INVX2TS U1471 ( .A(n1445), .Y(n1748) );
  AOI22X1TS U1472 ( .A0(n1695), .A1(n1748), .B0(n1450), .B1(
        \requesterAddressbuffer[5][3] ), .Y(n924) );
  INVX2TS U1473 ( .A(n920), .Y(n1751) );
  AOI22X1TS U1474 ( .A0(n944), .A1(n1751), .B0(n1045), .B1(n921), .Y(n923) );
  AOI22X1TS U1475 ( .A0(n945), .A1(n231), .B0(requesterAddressIn_NORTH[3]), 
        .B1(n1458), .Y(n922) );
  INVX2TS U1476 ( .A(n1425), .Y(n1777) );
  AOI22X1TS U1477 ( .A0(n991), .A1(n930), .B0(n1777), .B1(
        \requesterAddressbuffer[4][0] ), .Y(n929) );
  INVX2TS U1478 ( .A(n1420), .Y(n1769) );
  AOI22X1TS U1479 ( .A0(n925), .A1(n1782), .B0(requesterAddressIn_EAST[0]), 
        .B1(n1769), .Y(n928) );
  AOI22X1TS U1480 ( .A0(n926), .A1(n1763), .B0(requesterAddressIn_NORTH[0]), 
        .B1(n310), .Y(n927) );
  INVX2TS U1481 ( .A(n955), .Y(n1901) );
  AOI22X1TS U1482 ( .A0(n1901), .A1(n930), .B0(n1788), .B1(
        \requesterAddressbuffer[4][1] ), .Y(n937) );
  INVX2TS U1483 ( .A(n1420), .Y(n1780) );
  AOI22X1TS U1484 ( .A0(n932), .A1(n302), .B0(requesterAddressIn_EAST[1]), 
        .B1(n1780), .Y(n936) );
  AOI22X1TS U1485 ( .A0(n934), .A1(n1414), .B0(requesterAddressIn_NORTH[1]), 
        .B1(n933), .Y(n935) );
  INVX2TS U1486 ( .A(n962), .Y(n1913) );
  INVX2TS U1487 ( .A(n11), .Y(n1767) );
  INVX2TS U1488 ( .A(n1623), .Y(n1418) );
  AOI22X1TS U1489 ( .A0(n1913), .A1(n1767), .B0(n1418), .B1(
        \requesterAddressbuffer[4][2] ), .Y(n942) );
  AOI22X1TS U1490 ( .A0(n938), .A1(n1771), .B0(requesterAddressIn_EAST[2]), 
        .B1(n943), .Y(n941) );
  AOI22X1TS U1491 ( .A0(n939), .A1(n1784), .B0(requesterAddressIn_NORTH[2]), 
        .B1(n1783), .Y(n940) );
  INVX2TS U1492 ( .A(n969), .Y(n1925) );
  INVX2TS U1493 ( .A(n11), .Y(n1778) );
  AOI22X1TS U1494 ( .A0(n1925), .A1(n1778), .B0(n1418), .B1(
        \requesterAddressbuffer[4][3] ), .Y(n948) );
  AOI22X1TS U1495 ( .A0(n944), .A1(n296), .B0(requesterAddressIn_EAST[3]), 
        .B1(n943), .Y(n947) );
  AOI22X1TS U1496 ( .A0(n945), .A1(n284), .B0(requesterAddressIn_NORTH[3]), 
        .B1(n1772), .Y(n946) );
  INVX2TS U1497 ( .A(n949), .Y(n1892) );
  INVX2TS U1498 ( .A(n1392), .Y(n1809) );
  AOI22X1TS U1499 ( .A0(n1892), .A1(n956), .B0(n1809), .B1(
        \requesterAddressbuffer[3][0] ), .Y(n954) );
  INVX2TS U1500 ( .A(n950), .Y(n1393) );
  AOI22X1TS U1501 ( .A0(n951), .A1(n1393), .B0(n992), .B1(n157), .Y(n953) );
  INVX2TS U1502 ( .A(n964), .Y(n1397) );
  AOI22X1TS U1503 ( .A0(n994), .A1(n1397), .B0(n1025), .B1(n1805), .Y(n952) );
  INVX2TS U1504 ( .A(n955), .Y(n1861) );
  AOI22X1TS U1505 ( .A0(n1861), .A1(n956), .B0(n1816), .B1(
        \requesterAddressbuffer[3][1] ), .Y(n961) );
  INVX2TS U1506 ( .A(n957), .Y(n1818) );
  AOI22X1TS U1507 ( .A0(n958), .A1(n135), .B0(n999), .B1(n1818), .Y(n960) );
  AOI22X1TS U1508 ( .A0(n1002), .A1(n129), .B0(n1032), .B1(n163), .Y(n959) );
  INVX2TS U1509 ( .A(n962), .Y(n1872) );
  INVX2TS U1510 ( .A(n1382), .Y(n1801) );
  INVX2TS U1511 ( .A(n1632), .Y(n1387) );
  AOI22X1TS U1512 ( .A0(n1872), .A1(n1801), .B0(n1387), .B1(
        \requesterAddressbuffer[3][2] ), .Y(n968) );
  AOI22X1TS U1513 ( .A0(n963), .A1(n1820), .B0(n1007), .B1(n1383), .Y(n967) );
  INVX2TS U1514 ( .A(n964), .Y(n1821) );
  AOI22X1TS U1515 ( .A0(n1010), .A1(n1821), .B0(n1038), .B1(n965), .Y(n966) );
  INVX2TS U1516 ( .A(n969), .Y(n1883) );
  AOI22X1TS U1517 ( .A0(n1883), .A1(n131), .B0(n1387), .B1(
        \requesterAddressbuffer[3][3] ), .Y(n973) );
  AOI22X1TS U1518 ( .A0(n970), .A1(n1393), .B0(n1016), .B1(n1810), .Y(n972) );
  AOI22X1TS U1519 ( .A0(n1019), .A1(n1397), .B0(n1047), .B1(n1402), .Y(n971)
         );
  INVX2TS U1520 ( .A(n1644), .Y(n1836) );
  AOI22X1TS U1521 ( .A0(n1796), .A1(n978), .B0(n1836), .B1(
        \requesterAddressbuffer[2][0] ), .Y(n977) );
  INVX2TS U1522 ( .A(n1346), .Y(n1838) );
  AOI22X1TS U1523 ( .A0(requesterAddressIn_WEST[0]), .A1(n1839), .B0(n992), 
        .B1(n1838), .Y(n976) );
  INVX2TS U1524 ( .A(n974), .Y(n1378) );
  AOI22X1TS U1525 ( .A0(n994), .A1(n1378), .B0(n1025), .B1(n1841), .Y(n975) );
  AOI22X1TS U1526 ( .A0(n1901), .A1(n978), .B0(n1845), .B1(
        \requesterAddressbuffer[2][1] ), .Y(n981) );
  INVX2TS U1527 ( .A(n1346), .Y(n1847) );
  AOI22X1TS U1528 ( .A0(requesterAddressIn_WEST[1]), .A1(n1359), .B0(n999), 
        .B1(n1847), .Y(n980) );
  INVX2TS U1529 ( .A(n203), .Y(n1840) );
  AOI22X1TS U1530 ( .A0(n1002), .A1(n1840), .B0(n1032), .B1(n1848), .Y(n979)
         );
  INVX2TS U1531 ( .A(n10), .Y(n1829) );
  INVX2TS U1532 ( .A(n1644), .Y(n1351) );
  AOI22X1TS U1533 ( .A0(n1913), .A1(n1829), .B0(n1351), .B1(
        \requesterAddressbuffer[2][2] ), .Y(n985) );
  AOI22X1TS U1534 ( .A0(requesterAddressIn_WEST[2]), .A1(n1830), .B0(n1007), 
        .B1(n987), .Y(n984) );
  AOI22X1TS U1535 ( .A0(n1010), .A1(n1831), .B0(n1038), .B1(n982), .Y(n983) );
  INVX2TS U1536 ( .A(n10), .Y(n1837) );
  AOI22X1TS U1537 ( .A0(n1925), .A1(n1837), .B0(n1351), .B1(
        \requesterAddressbuffer[2][3] ), .Y(n990) );
  INVX2TS U1538 ( .A(n986), .Y(n1359) );
  AOI22X1TS U1539 ( .A0(requesterAddressIn_WEST[3]), .A1(n1359), .B0(n1016), 
        .B1(n987), .Y(n989) );
  AOI22X1TS U1540 ( .A0(n1019), .A1(n194), .B0(n1047), .B1(n1832), .Y(n988) );
  INVX2TS U1541 ( .A(n1006), .Y(n1870) );
  AOI22X1TS U1542 ( .A0(n991), .A1(n998), .B0(n1870), .B1(
        \requesterAddressbuffer[1][0] ), .Y(n997) );
  INVX2TS U1543 ( .A(n1087), .Y(n1874) );
  AOI22X1TS U1544 ( .A0(requesterAddressIn_WEST[0]), .A1(n1875), .B0(n992), 
        .B1(n1874), .Y(n996) );
  AOI22X1TS U1545 ( .A0(n994), .A1(n1101), .B0(n993), .B1(n1866), .Y(n995) );
  AOI22X1TS U1546 ( .A0(n1768), .A1(n998), .B0(n1882), .B1(
        \requesterAddressbuffer[1][1] ), .Y(n1005) );
  INVX2TS U1547 ( .A(n1087), .Y(n1885) );
  AOI22X1TS U1548 ( .A0(requesterAddressIn_WEST[1]), .A1(n1099), .B0(n999), 
        .B1(n1885), .Y(n1004) );
  INVX2TS U1549 ( .A(n1017), .Y(n1855) );
  INVX2TS U1550 ( .A(n1000), .Y(n1102) );
  AOI22X1TS U1551 ( .A0(n1002), .A1(n1855), .B0(n1001), .B1(n1102), .Y(n1003)
         );
  INVX2TS U1552 ( .A(n1085), .Y(n1860) );
  INVX2TS U1553 ( .A(n1006), .Y(n1093) );
  AOI22X1TS U1554 ( .A0(n1779), .A1(n1860), .B0(n1093), .B1(
        \requesterAddressbuffer[1][2] ), .Y(n1013) );
  AOI22X1TS U1555 ( .A0(requesterAddressIn_WEST[2]), .A1(n1863), .B0(n1007), 
        .B1(n1015), .Y(n1012) );
  AOI22X1TS U1556 ( .A0(n1010), .A1(n349), .B0(n1009), .B1(n1008), .Y(n1011)
         );
  INVX2TS U1557 ( .A(n1085), .Y(n1871) );
  AOI22X1TS U1558 ( .A0(n1790), .A1(n1871), .B0(n1093), .B1(
        \requesterAddressbuffer[1][3] ), .Y(n1022) );
  INVX2TS U1559 ( .A(n1014), .Y(n1099) );
  AOI22X1TS U1560 ( .A0(requesterAddressIn_WEST[3]), .A1(n1099), .B0(n1016), 
        .B1(n1015), .Y(n1021) );
  INVX2TS U1561 ( .A(n1017), .Y(n1342) );
  AOI22X1TS U1562 ( .A0(n1019), .A1(n1342), .B0(n1018), .B1(n324), .Y(n1020)
         );
  INVX2TS U1563 ( .A(n1063), .Y(n1911) );
  AOI22X1TS U1564 ( .A0(readRequesterAddress[0]), .A1(n1030), .B0(n1911), .B1(
        \requesterAddressbuffer[0][0] ), .Y(n1029) );
  INVX2TS U1565 ( .A(n1052), .Y(n1914) );
  AOI22X1TS U1566 ( .A0(requesterAddressIn_WEST[0]), .A1(n1916), .B0(n1023), 
        .B1(n1914), .Y(n1028) );
  INVX2TS U1567 ( .A(n1024), .Y(n1905) );
  AOI22X1TS U1568 ( .A0(n1026), .A1(n1076), .B0(n1025), .B1(n1905), .Y(n1027)
         );
  AOI22X1TS U1569 ( .A0(n1861), .A1(n1030), .B0(n1923), .B1(
        \requesterAddressbuffer[0][1] ), .Y(n1036) );
  INVX2TS U1570 ( .A(n1052), .Y(n1926) );
  AOI22X1TS U1571 ( .A0(requesterAddressIn_WEST[1]), .A1(n1065), .B0(n1031), 
        .B1(n1926), .Y(n1035) );
  AOI22X1TS U1572 ( .A0(n1033), .A1(n1907), .B0(n1032), .B1(n1905), .Y(n1034)
         );
  INVX2TS U1573 ( .A(n12), .Y(n1900) );
  INVX2TS U1574 ( .A(n1063), .Y(n1058) );
  AOI22X1TS U1575 ( .A0(n1872), .A1(n1900), .B0(n1058), .B1(
        \requesterAddressbuffer[0][2] ), .Y(n1042) );
  AOI22X1TS U1576 ( .A0(requesterAddressIn_WEST[2]), .A1(n1903), .B0(n1037), 
        .B1(n1044), .Y(n1041) );
  AOI22X1TS U1577 ( .A0(n1039), .A1(n1930), .B0(n1038), .B1(n1918), .Y(n1040)
         );
  INVX2TS U1578 ( .A(n12), .Y(n1912) );
  AOI22X1TS U1579 ( .A0(n1883), .A1(n1912), .B0(n1058), .B1(
        \requesterAddressbuffer[0][3] ), .Y(n1051) );
  INVX2TS U1580 ( .A(n1043), .Y(n1065) );
  AOI22X1TS U1581 ( .A0(requesterAddressIn_WEST[3]), .A1(n1065), .B0(n1045), 
        .B1(n1044), .Y(n1050) );
  INVX2TS U1582 ( .A(n1046), .Y(n1896) );
  AOI22X1TS U1583 ( .A0(n1048), .A1(n1896), .B0(n1047), .B1(n1054), .Y(n1049)
         );
  INVX2TS U1584 ( .A(n12), .Y(n1924) );
  INVX2TS U1585 ( .A(n1086), .Y(n1476) );
  AOI22X1TS U1586 ( .A0(n1924), .A1(n1476), .B0(n1058), .B1(
        \dataoutbuffer[0][0] ), .Y(n1057) );
  AOI22X1TS U1587 ( .A0(n1065), .A1(n1053), .B0(n1044), .B1(n1347), .Y(n1056)
         );
  CLKBUFX2TS U1588 ( .A(n1088), .Y(n1479) );
  AOI22X1TS U1589 ( .A0(n1930), .A1(dataIn_SOUTH[0]), .B0(n1054), .B1(n1479), 
        .Y(n1055) );
  INVX2TS U1590 ( .A(n1092), .Y(n1484) );
  AOI22X1TS U1591 ( .A0(n1900), .A1(n1484), .B0(n1058), .B1(
        \dataoutbuffer[0][1] ), .Y(n1062) );
  AOI22X1TS U1592 ( .A0(n396), .A1(n1059), .B0(n1914), .B1(n1352), .Y(n1061)
         );
  CLKBUFX2TS U1593 ( .A(n1094), .Y(n1489) );
  AOI22X1TS U1594 ( .A0(n1896), .A1(dataIn_SOUTH[1]), .B0(n401), .B1(n1489), 
        .Y(n1060) );
  INVX2TS U1595 ( .A(n1098), .Y(n1494) );
  INVX2TS U1596 ( .A(n1063), .Y(n1080) );
  AOI22X1TS U1597 ( .A0(n1912), .A1(n1494), .B0(n1080), .B1(
        \dataoutbuffer[0][2] ), .Y(n1068) );
  AOI22X1TS U1598 ( .A0(n1065), .A1(n1064), .B0(n1926), .B1(n1358), .Y(n1067)
         );
  CLKBUFX2TS U1599 ( .A(n1100), .Y(n1499) );
  AOI22X1TS U1600 ( .A0(n1076), .A1(dataIn_SOUTH[2]), .B0(n1905), .B1(n1499), 
        .Y(n1066) );
  INVX2TS U1601 ( .A(n1106), .Y(n1503) );
  AOI22X1TS U1602 ( .A0(n1924), .A1(n1503), .B0(n1080), .B1(
        \dataoutbuffer[0][3] ), .Y(n1072) );
  AOI22X1TS U1603 ( .A0(n1074), .A1(n1069), .B0(n394), .B1(n1364), .Y(n1071)
         );
  CLKBUFX2TS U1604 ( .A(n1107), .Y(n1506) );
  AOI22X1TS U1605 ( .A0(n1896), .A1(dataIn_SOUTH[3]), .B0(n1075), .B1(n1506), 
        .Y(n1070) );
  INVX2TS U1606 ( .A(n1401), .Y(n1368) );
  AOI22X1TS U1607 ( .A0(n1900), .A1(n1368), .B0(n1080), .B1(
        \dataoutbuffer[0][4] ), .Y(n1079) );
  AOI22X1TS U1608 ( .A0(n1074), .A1(n1073), .B0(n394), .B1(n1369), .Y(n1078)
         );
  CLKBUFX2TS U1609 ( .A(n1112), .Y(n1512) );
  AOI22X1TS U1610 ( .A0(n1076), .A1(dataIn_SOUTH[4]), .B0(n1075), .B1(n1512), 
        .Y(n1077) );
  INVX2TS U1611 ( .A(n1406), .Y(n1376) );
  AOI22X1TS U1612 ( .A0(n1912), .A1(n1376), .B0(n1080), .B1(
        \dataoutbuffer[0][5] ), .Y(n1084) );
  AOI22X1TS U1613 ( .A0(n396), .A1(n1081), .B0(n1914), .B1(n1377), .Y(n1083)
         );
  CLKBUFX2TS U1614 ( .A(n1341), .Y(n1520) );
  AOI22X1TS U1615 ( .A0(n427), .A1(dataIn_SOUTH[5]), .B0(n401), .B1(n1520), 
        .Y(n1082) );
  INVX2TS U1616 ( .A(n1086), .Y(n1524) );
  AOI22X1TS U1617 ( .A0(n319), .A1(n1524), .B0(n1093), .B1(
        \dataoutbuffer[1][0] ), .Y(n1091) );
  AOI22X1TS U1618 ( .A0(n1099), .A1(dataIn_WEST[0]), .B0(n317), .B1(n1347), 
        .Y(n1090) );
  CLKBUFX2TS U1619 ( .A(n1088), .Y(n1528) );
  CLKBUFX2TS U1620 ( .A(dataIn_SOUTH[0]), .Y(n1529) );
  CLKBUFX2TS U1621 ( .A(n1529), .Y(n1478) );
  AOI22X1TS U1622 ( .A0(n1102), .A1(n1528), .B0(n349), .B1(n1478), .Y(n1089)
         );
  INVX2TS U1623 ( .A(n1092), .Y(n1534) );
  AOI22X1TS U1624 ( .A0(n1860), .A1(n1534), .B0(n1093), .B1(
        \dataoutbuffer[1][1] ), .Y(n1097) );
  AOI22X1TS U1625 ( .A0(n331), .A1(dataIn_WEST[1]), .B0(n1874), .B1(n1352), 
        .Y(n1096) );
  CLKBUFX2TS U1626 ( .A(n1094), .Y(n1536) );
  CLKBUFX2TS U1627 ( .A(dataIn_SOUTH[1]), .Y(n1537) );
  CLKBUFX2TS U1628 ( .A(n1537), .Y(n1488) );
  AOI22X1TS U1629 ( .A0(n1888), .A1(n1536), .B0(n1855), .B1(n1488), .Y(n1095)
         );
  INVX2TS U1630 ( .A(n1098), .Y(n1543) );
  INVX2TS U1631 ( .A(n1006), .Y(n1340) );
  AOI22X1TS U1632 ( .A0(n1871), .A1(n1543), .B0(n1340), .B1(
        \dataoutbuffer[1][2] ), .Y(n1105) );
  AOI22X1TS U1633 ( .A0(n1099), .A1(dataIn_WEST[2]), .B0(n1885), .B1(n1358), 
        .Y(n1104) );
  CLKBUFX2TS U1634 ( .A(n1100), .Y(n1545) );
  CLKBUFX2TS U1635 ( .A(dataIn_SOUTH[2]), .Y(n1546) );
  CLKBUFX2TS U1636 ( .A(n1546), .Y(n1497) );
  AOI22X1TS U1637 ( .A0(n1102), .A1(n1545), .B0(n1101), .B1(n1497), .Y(n1103)
         );
  INVX2TS U1638 ( .A(n1106), .Y(n1550) );
  AOI22X1TS U1639 ( .A0(n998), .A1(n1550), .B0(n1340), .B1(
        \dataoutbuffer[1][3] ), .Y(n1110) );
  AOI22X1TS U1640 ( .A0(n1111), .A1(dataIn_WEST[3]), .B0(n317), .B1(n1364), 
        .Y(n1109) );
  CLKBUFX2TS U1641 ( .A(n1107), .Y(n1553) );
  CLKBUFX2TS U1642 ( .A(dataIn_SOUTH[3]), .Y(n1554) );
  CLKBUFX2TS U1643 ( .A(n1554), .Y(n1505) );
  AOI22X1TS U1644 ( .A0(n324), .A1(n1553), .B0(n1342), .B1(n1505), .Y(n1108)
         );
  AOI22X1TS U1645 ( .A0(n1860), .A1(n1368), .B0(n1340), .B1(
        \dataoutbuffer[1][4] ), .Y(n1339) );
  AOI22X1TS U1646 ( .A0(n1111), .A1(dataIn_WEST[4]), .B0(n317), .B1(n1369), 
        .Y(n1338) );
  CLKBUFX2TS U1647 ( .A(n1112), .Y(n1560) );
  CLKBUFX2TS U1648 ( .A(dataIn_SOUTH[4]), .Y(n1562) );
  CLKBUFX2TS U1649 ( .A(n1562), .Y(n1511) );
  AOI22X1TS U1650 ( .A0(n324), .A1(n1560), .B0(n1877), .B1(n1511), .Y(n1337)
         );
  AOI22X1TS U1651 ( .A0(n1871), .A1(n1376), .B0(n1340), .B1(
        \dataoutbuffer[1][5] ), .Y(n1345) );
  AOI22X1TS U1652 ( .A0(n331), .A1(dataIn_WEST[5]), .B0(n1874), .B1(n1377), 
        .Y(n1344) );
  CLKBUFX2TS U1653 ( .A(n1341), .Y(n1571) );
  CLKBUFX2TS U1654 ( .A(dataIn_SOUTH[5]), .Y(n1573) );
  CLKBUFX2TS U1655 ( .A(n1573), .Y(n1519) );
  AOI22X1TS U1656 ( .A0(n1888), .A1(n1571), .B0(n1342), .B1(n1519), .Y(n1343)
         );
  INVX2TS U1657 ( .A(n10), .Y(n1846) );
  AOI22X1TS U1658 ( .A0(n1846), .A1(n1476), .B0(n1351), .B1(
        \dataoutbuffer[2][0] ), .Y(n1350) );
  AOI22X1TS U1659 ( .A0(n1359), .A1(n1413), .B0(n184), .B1(n1347), .Y(n1349)
         );
  AOI22X1TS U1660 ( .A0(n1360), .A1(n1528), .B0(n1840), .B1(dataIn_SOUTH[0]), 
        .Y(n1348) );
  AOI22X1TS U1661 ( .A0(n1829), .A1(n1484), .B0(n1351), .B1(
        \dataoutbuffer[2][1] ), .Y(n1356) );
  AOI22X1TS U1662 ( .A0(n186), .A1(n1419), .B0(n1838), .B1(n1352), .Y(n1355)
         );
  INVX2TS U1663 ( .A(n1353), .Y(n1848) );
  AOI22X1TS U1664 ( .A0(n1848), .A1(n1536), .B0(n1371), .B1(dataIn_SOUTH[1]), 
        .Y(n1354) );
  INVX2TS U1665 ( .A(n1357), .Y(n1375) );
  AOI22X1TS U1666 ( .A0(n1837), .A1(n1494), .B0(n1375), .B1(
        \dataoutbuffer[2][2] ), .Y(n1363) );
  AOI22X1TS U1667 ( .A0(n1359), .A1(n1426), .B0(n1847), .B1(n1358), .Y(n1362)
         );
  AOI22X1TS U1668 ( .A0(n1360), .A1(n1545), .B0(n215), .B1(dataIn_SOUTH[2]), 
        .Y(n1361) );
  AOI22X1TS U1669 ( .A0(n1846), .A1(n1503), .B0(n1375), .B1(
        \dataoutbuffer[2][3] ), .Y(n1367) );
  AOI22X1TS U1670 ( .A0(n1370), .A1(n1431), .B0(n184), .B1(n1364), .Y(n1366)
         );
  AOI22X1TS U1671 ( .A0(n982), .A1(n1553), .B0(n1378), .B1(dataIn_SOUTH[3]), 
        .Y(n1365) );
  AOI22X1TS U1672 ( .A0(n1829), .A1(n1368), .B0(n1375), .B1(
        \dataoutbuffer[2][4] ), .Y(n1374) );
  AOI22X1TS U1673 ( .A0(n1370), .A1(n1435), .B0(n184), .B1(n1369), .Y(n1373)
         );
  AOI22X1TS U1674 ( .A0(n1832), .A1(n1560), .B0(n1371), .B1(dataIn_SOUTH[4]), 
        .Y(n1372) );
  AOI22X1TS U1675 ( .A0(n1837), .A1(n1376), .B0(n1375), .B1(
        \dataoutbuffer[2][5] ), .Y(n1381) );
  AOI22X1TS U1676 ( .A0(n186), .A1(n1441), .B0(n1838), .B1(n1377), .Y(n1380)
         );
  AOI22X1TS U1677 ( .A0(n1848), .A1(n1571), .B0(n1378), .B1(dataIn_SOUTH[5]), 
        .Y(n1379) );
  INVX2TS U1678 ( .A(n1382), .Y(n1817) );
  AOI22X1TS U1679 ( .A0(n1817), .A1(n1476), .B0(n1387), .B1(
        \dataoutbuffer[3][0] ), .Y(n1386) );
  AOI22X1TS U1680 ( .A0(n176), .A1(n1413), .B0(n1383), .B1(dataIn_EAST[0]), 
        .Y(n1385) );
  AOI22X1TS U1681 ( .A0(n163), .A1(n1479), .B0(n1397), .B1(n1478), .Y(n1384)
         );
  AOI22X1TS U1682 ( .A0(n1801), .A1(n1484), .B0(n1387), .B1(
        \dataoutbuffer[3][1] ), .Y(n1391) );
  AOI22X1TS U1683 ( .A0(n1393), .A1(n1419), .B0(n1818), .B1(dataIn_EAST[1]), 
        .Y(n1390) );
  INVX2TS U1684 ( .A(n1388), .Y(n1822) );
  AOI22X1TS U1685 ( .A0(n1822), .A1(n1489), .B0(n143), .B1(n1488), .Y(n1389)
         );
  INVX2TS U1686 ( .A(n1392), .Y(n1407) );
  AOI22X1TS U1687 ( .A0(n131), .A1(n1494), .B0(n1407), .B1(
        \dataoutbuffer[3][2] ), .Y(n1396) );
  AOI22X1TS U1688 ( .A0(n1393), .A1(n1426), .B0(n157), .B1(dataIn_EAST[2]), 
        .Y(n1395) );
  AOI22X1TS U1689 ( .A0(n163), .A1(n1499), .B0(n1821), .B1(n1497), .Y(n1394)
         );
  AOI22X1TS U1690 ( .A0(n1817), .A1(n1503), .B0(n1407), .B1(
        \dataoutbuffer[3][3] ), .Y(n1400) );
  AOI22X1TS U1691 ( .A0(n139), .A1(n1431), .B0(n169), .B1(dataIn_EAST[3]), .Y(
        n1399) );
  AOI22X1TS U1692 ( .A0(n1402), .A1(n1506), .B0(n1397), .B1(n1505), .Y(n1398)
         );
  INVX2TS U1693 ( .A(n1401), .Y(n1558) );
  AOI22X1TS U1694 ( .A0(n1801), .A1(n1558), .B0(n1407), .B1(
        \dataoutbuffer[3][4] ), .Y(n1405) );
  AOI22X1TS U1695 ( .A0(n1408), .A1(n1435), .B0(n157), .B1(dataIn_EAST[4]), 
        .Y(n1404) );
  AOI22X1TS U1696 ( .A0(n1402), .A1(n1512), .B0(n1409), .B1(n1511), .Y(n1403)
         );
  INVX2TS U1697 ( .A(n1406), .Y(n1568) );
  AOI22X1TS U1698 ( .A0(n956), .A1(n1568), .B0(n1407), .B1(
        \dataoutbuffer[3][5] ), .Y(n1412) );
  AOI22X1TS U1699 ( .A0(n1408), .A1(n1441), .B0(n1818), .B1(dataIn_EAST[5]), 
        .Y(n1411) );
  AOI22X1TS U1700 ( .A0(n1822), .A1(n1520), .B0(n1409), .B1(n1519), .Y(n1410)
         );
  INVX2TS U1701 ( .A(n11), .Y(n1789) );
  AOI22X1TS U1702 ( .A0(n1789), .A1(n1524), .B0(n1418), .B1(
        \dataoutbuffer[4][0] ), .Y(n1417) );
  CLKBUFX2TS U1703 ( .A(n1413), .Y(n1525) );
  AOI22X1TS U1704 ( .A0(n283), .A1(n1525), .B0(n1780), .B1(dataIn_EAST[0]), 
        .Y(n1416) );
  AOI22X1TS U1705 ( .A0(n1414), .A1(n1529), .B0(n280), .B1(n1528), .Y(n1415)
         );
  AOI22X1TS U1706 ( .A0(n1767), .A1(n1534), .B0(n1418), .B1(
        \dataoutbuffer[4][1] ), .Y(n1424) );
  CLKBUFX2TS U1707 ( .A(n1419), .Y(n1535) );
  AOI22X1TS U1708 ( .A0(n296), .A1(n1535), .B0(n943), .B1(dataIn_EAST[1]), .Y(
        n1423) );
  INVX2TS U1709 ( .A(n1421), .Y(n1792) );
  AOI22X1TS U1710 ( .A0(n1784), .A1(n1537), .B0(n1792), .B1(n1536), .Y(n1422)
         );
  INVX2TS U1711 ( .A(n1425), .Y(n1440) );
  AOI22X1TS U1712 ( .A0(n1778), .A1(n1543), .B0(n1440), .B1(
        \dataoutbuffer[4][2] ), .Y(n1430) );
  CLKBUFX2TS U1713 ( .A(n1426), .Y(n1544) );
  AOI22X1TS U1714 ( .A0(n283), .A1(n1544), .B0(n1769), .B1(dataIn_EAST[2]), 
        .Y(n1429) );
  INVX2TS U1715 ( .A(n1427), .Y(n1773) );
  AOI22X1TS U1716 ( .A0(n1773), .A1(n1546), .B0(n280), .B1(n1545), .Y(n1428)
         );
  AOI22X1TS U1717 ( .A0(n1789), .A1(n1550), .B0(n1440), .B1(
        \dataoutbuffer[4][3] ), .Y(n1434) );
  CLKBUFX2TS U1718 ( .A(n1431), .Y(n1551) );
  AOI22X1TS U1719 ( .A0(n1436), .A1(n1551), .B0(n1780), .B1(dataIn_EAST[3]), 
        .Y(n1433) );
  AOI22X1TS U1720 ( .A0(n284), .A1(n1554), .B0(n1792), .B1(n1553), .Y(n1432)
         );
  AOI22X1TS U1721 ( .A0(n1767), .A1(n1558), .B0(n1440), .B1(
        \dataoutbuffer[4][4] ), .Y(n1439) );
  CLKBUFX2TS U1722 ( .A(n1435), .Y(n1559) );
  AOI22X1TS U1723 ( .A0(n1436), .A1(n1559), .B0(n274), .B1(dataIn_EAST[4]), 
        .Y(n1438) );
  AOI22X1TS U1724 ( .A0(n1763), .A1(n1562), .B0(n310), .B1(n1560), .Y(n1437)
         );
  AOI22X1TS U1725 ( .A0(n1778), .A1(n1568), .B0(n1440), .B1(
        \dataoutbuffer[4][5] ), .Y(n1444) );
  CLKBUFX2TS U1726 ( .A(n1441), .Y(n1570) );
  AOI22X1TS U1727 ( .A0(n302), .A1(n1570), .B0(n1769), .B1(dataIn_EAST[5]), 
        .Y(n1443) );
  AOI22X1TS U1728 ( .A0(n1773), .A1(n1573), .B0(n1792), .B1(n1571), .Y(n1442)
         );
  AOI22X1TS U1729 ( .A0(n225), .A1(n1524), .B0(n1450), .B1(
        \dataoutbuffer[5][0] ), .Y(n1449) );
  AOI22X1TS U1730 ( .A0(n1457), .A1(n1525), .B0(n1750), .B1(n1477), .Y(n1448)
         );
  AOI22X1TS U1731 ( .A0(n1446), .A1(n1479), .B0(n1467), .B1(n1478), .Y(n1447)
         );
  AOI22X1TS U1732 ( .A0(n1738), .A1(n1534), .B0(n1450), .B1(
        \dataoutbuffer[5][1] ), .Y(n1455) );
  AOI22X1TS U1733 ( .A0(n258), .A1(n1535), .B0(n921), .B1(n1486), .Y(n1454) );
  INVX2TS U1734 ( .A(n1452), .Y(n1753) );
  AOI22X1TS U1735 ( .A0(n1753), .A1(n1489), .B0(n231), .B1(n1488), .Y(n1453)
         );
  INVX2TS U1736 ( .A(n1456), .Y(n1472) );
  AOI22X1TS U1737 ( .A0(n1748), .A1(n1543), .B0(n1472), .B1(
        \dataoutbuffer[5][2] ), .Y(n1461) );
  AOI22X1TS U1738 ( .A0(n1457), .A1(n1544), .B0(n1740), .B1(n1495), .Y(n1460)
         );
  AOI22X1TS U1739 ( .A0(n1458), .A1(n1499), .B0(n1752), .B1(n1497), .Y(n1459)
         );
  AOI22X1TS U1740 ( .A0(n913), .A1(n1550), .B0(n1472), .B1(
        \dataoutbuffer[5][3] ), .Y(n1466) );
  AOI22X1TS U1741 ( .A0(n1462), .A1(n1551), .B0(n1750), .B1(n1504), .Y(n1465)
         );
  AOI22X1TS U1742 ( .A0(n259), .A1(n1506), .B0(n1463), .B1(n1505), .Y(n1464)
         );
  AOI22X1TS U1743 ( .A0(n1738), .A1(n1558), .B0(n1472), .B1(
        \dataoutbuffer[5][4] ), .Y(n1471) );
  AOI22X1TS U1744 ( .A0(n1741), .A1(n1559), .B0(n224), .B1(n1510), .Y(n1470)
         );
  AOI22X1TS U1745 ( .A0(n1468), .A1(n1512), .B0(n1467), .B1(n1511), .Y(n1469)
         );
  AOI22X1TS U1746 ( .A0(n1748), .A1(n1568), .B0(n1472), .B1(
        \dataoutbuffer[5][5] ), .Y(n1475) );
  AOI22X1TS U1747 ( .A0(n227), .A1(n1570), .B0(n1740), .B1(n1518), .Y(n1474)
         );
  AOI22X1TS U1748 ( .A0(n259), .A1(n1520), .B0(n231), .B1(n1519), .Y(n1473) );
  INVX2TS U1749 ( .A(n9), .Y(n1726) );
  AOI22X1TS U1750 ( .A0(n1726), .A1(n1476), .B0(n1483), .B1(
        \dataoutbuffer[6][0] ), .Y(n1482) );
  AOI22X1TS U1751 ( .A0(n1496), .A1(n1525), .B0(n1718), .B1(n1477), .Y(n1481)
         );
  AOI22X1TS U1752 ( .A0(n901), .A1(n1479), .B0(n1729), .B1(n1478), .Y(n1480)
         );
  AOI22X1TS U1753 ( .A0(n1707), .A1(n1484), .B0(n1483), .B1(
        \dataoutbuffer[6][1] ), .Y(n1492) );
  AOI22X1TS U1754 ( .A0(n1727), .A1(n1535), .B0(n905), .B1(n1486), .Y(n1491)
         );
  INVX2TS U1755 ( .A(n1487), .Y(n1730) );
  AOI22X1TS U1756 ( .A0(n1730), .A1(n1489), .B0(n1703), .B1(n1488), .Y(n1490)
         );
  INVX2TS U1757 ( .A(n1493), .Y(n1517) );
  AOI22X1TS U1758 ( .A0(n1717), .A1(n1494), .B0(n1517), .B1(
        \dataoutbuffer[6][2] ), .Y(n1502) );
  AOI22X1TS U1759 ( .A0(n1496), .A1(n1544), .B0(n1708), .B1(n1495), .Y(n1501)
         );
  AOI22X1TS U1760 ( .A0(n94), .A1(n1499), .B0(n1498), .B1(n1497), .Y(n1500) );
  AOI22X1TS U1761 ( .A0(n1726), .A1(n1503), .B0(n1517), .B1(
        \dataoutbuffer[6][3] ), .Y(n1509) );
  AOI22X1TS U1762 ( .A0(n98), .A1(n1551), .B0(n1718), .B1(n1504), .Y(n1508) );
  AOI22X1TS U1763 ( .A0(n1513), .A1(n1506), .B0(n91), .B1(n1505), .Y(n1507) );
  AOI22X1TS U1764 ( .A0(n1707), .A1(n1368), .B0(n1517), .B1(
        \dataoutbuffer[6][4] ), .Y(n1516) );
  AOI22X1TS U1765 ( .A0(n1709), .A1(n1559), .B0(n84), .B1(n1510), .Y(n1515) );
  AOI22X1TS U1766 ( .A0(n1513), .A1(n1512), .B0(n1720), .B1(n1511), .Y(n1514)
         );
  AOI22X1TS U1767 ( .A0(n1717), .A1(n1376), .B0(n1517), .B1(
        \dataoutbuffer[6][5] ), .Y(n1523) );
  AOI22X1TS U1768 ( .A0(n1727), .A1(n1570), .B0(n1708), .B1(n1518), .Y(n1522)
         );
  AOI22X1TS U1769 ( .A0(n1730), .A1(n1520), .B0(n91), .B1(n1519), .Y(n1521) );
  AOI22X1TS U1770 ( .A0(n1678), .A1(n1524), .B0(n1533), .B1(
        \dataoutbuffer[7][0] ), .Y(n1532) );
  AOI22X1TS U1771 ( .A0(n1526), .A1(n1525), .B0(n1687), .B1(dataIn_EAST[0]), 
        .Y(n1531) );
  INVX2TS U1772 ( .A(n1527), .Y(n1690) );
  AOI22X1TS U1773 ( .A0(n1690), .A1(n1529), .B0(n1561), .B1(n1528), .Y(n1530)
         );
  AOI22X1TS U1774 ( .A0(n34), .A1(n1534), .B0(n1533), .B1(
        \dataoutbuffer[7][1] ), .Y(n1541) );
  AOI22X1TS U1775 ( .A0(n66), .A1(n1535), .B0(n32), .B1(dataIn_EAST[1]), .Y(
        n1540) );
  AOI22X1TS U1776 ( .A0(n1538), .A1(n1537), .B0(n1697), .B1(n1536), .Y(n1539)
         );
  INVX2TS U1777 ( .A(n1542), .Y(n1567) );
  AOI22X1TS U1778 ( .A0(n1696), .A1(n1543), .B0(n1567), .B1(
        \dataoutbuffer[7][2] ), .Y(n1549) );
  AOI22X1TS U1779 ( .A0(n1552), .A1(n1544), .B0(n1679), .B1(dataIn_EAST[2]), 
        .Y(n1548) );
  AOI22X1TS U1780 ( .A0(n1690), .A1(n1546), .B0(n48), .B1(n1545), .Y(n1547) );
  AOI22X1TS U1781 ( .A0(n1678), .A1(n1550), .B0(n1567), .B1(
        \dataoutbuffer[7][3] ), .Y(n1557) );
  AOI22X1TS U1782 ( .A0(n1552), .A1(n1551), .B0(n1687), .B1(dataIn_EAST[3]), 
        .Y(n1556) );
  AOI22X1TS U1783 ( .A0(n1690), .A1(n1554), .B0(n1572), .B1(n1553), .Y(n1555)
         );
  AOI22X1TS U1784 ( .A0(n34), .A1(n1558), .B0(n1567), .B1(
        \dataoutbuffer[7][4] ), .Y(n1566) );
  AOI22X1TS U1785 ( .A0(n1680), .A1(n1559), .B0(n1569), .B1(dataIn_EAST[4]), 
        .Y(n1565) );
  AOI22X1TS U1786 ( .A0(n1563), .A1(n1562), .B0(n1561), .B1(n1560), .Y(n1564)
         );
  AOI22X1TS U1787 ( .A0(n1696), .A1(n1568), .B0(n1567), .B1(
        \dataoutbuffer[7][5] ), .Y(n1576) );
  AOI22X1TS U1788 ( .A0(n42), .A1(n1570), .B0(n1569), .B1(dataIn_EAST[5]), .Y(
        n1575) );
  AOI22X1TS U1789 ( .A0(n1563), .A1(n1573), .B0(n1572), .B1(n1571), .Y(n1574)
         );
  CLKBUFX2TS U1790 ( .A(n1669), .Y(n1620) );
  INVX2TS U1791 ( .A(n1577), .Y(n1665) );
  AOI22X1TS U1792 ( .A0(n1579), .A1(n1602), .B0(n1601), .B1(n1578), .Y(n1581)
         );
  AOI22X1TS U1793 ( .A0(n1582), .A1(n1665), .B0(n1581), .B1(n1580), .Y(n1584)
         );
  AOI22X1TS U1794 ( .A0(n1585), .A1(n1620), .B0(n1584), .B1(n1583), .Y(n1588)
         );
  AOI32X1TS U1795 ( .A0(n1588), .A1(n1587), .A2(n1586), .B0(n1694), .B1(n1964), 
        .Y(n1217) );
  INVX2TS U1796 ( .A(n1577), .Y(n1638) );
  AOI22X1TS U1797 ( .A0(n1590), .A1(n1602), .B0(n1601), .B1(n1589), .Y(n1592)
         );
  AOI22X1TS U1798 ( .A0(n1593), .A1(n1638), .B0(n1592), .B1(n1591), .Y(n1595)
         );
  AOI22X1TS U1799 ( .A0(n1596), .A1(n1620), .B0(n1595), .B1(n1594), .Y(n1599)
         );
  AOI32X1TS U1800 ( .A0(n1599), .A1(n1598), .A2(n1597), .B0(n1725), .B1(n1965), 
        .Y(n1216) );
  AOI22X1TS U1801 ( .A0(n1603), .A1(n1602), .B0(n1601), .B1(n1600), .Y(n1605)
         );
  AOI22X1TS U1802 ( .A0(n1606), .A1(n1638), .B0(n1605), .B1(n1604), .Y(n1608)
         );
  AOI22X1TS U1803 ( .A0(n1609), .A1(n1620), .B0(n1608), .B1(n1607), .Y(n1612)
         );
  AOI32X1TS U1804 ( .A0(n1612), .A1(n1611), .A2(n1610), .B0(n1757), .B1(n1966), 
        .Y(n1215) );
  CLKBUFX2TS U1805 ( .A(n1661), .Y(n1648) );
  CLKBUFX2TS U1806 ( .A(n1660), .Y(n1647) );
  AOI22X1TS U1807 ( .A0(n1614), .A1(n1648), .B0(n1647), .B1(n1613), .Y(n1616)
         );
  AOI22X1TS U1808 ( .A0(n1617), .A1(n1665), .B0(n1616), .B1(n1615), .Y(n1619)
         );
  AOI22X1TS U1809 ( .A0(n1621), .A1(n1620), .B0(n1619), .B1(n1618), .Y(n1624)
         );
  AOI32X1TS U1810 ( .A0(n1624), .A1(n1623), .A2(n1622), .B0(n1788), .B1(n1967), 
        .Y(n1214) );
  AOI22X1TS U1811 ( .A0(n121), .A1(n1648), .B0(n1647), .B1(n26), .Y(n1626) );
  AOI22X1TS U1812 ( .A0(n1627), .A1(n1638), .B0(n1626), .B1(n1625), .Y(n1629)
         );
  AOI22X1TS U1813 ( .A0(n1630), .A1(n1669), .B0(n1629), .B1(n1628), .Y(n1633)
         );
  AOI32X1TS U1814 ( .A0(n1633), .A1(n1632), .A2(n1631), .B0(n1816), .B1(n1968), 
        .Y(n1213) );
  AOI22X1TS U1815 ( .A0(n1635), .A1(n1648), .B0(n1647), .B1(n1634), .Y(n1637)
         );
  AOI22X1TS U1816 ( .A0(n1639), .A1(n1638), .B0(n1637), .B1(n1636), .Y(n1641)
         );
  AOI22X1TS U1817 ( .A0(n1642), .A1(n1655), .B0(n1641), .B1(n1640), .Y(n1645)
         );
  AOI32X1TS U1818 ( .A0(n1645), .A1(n1644), .A2(n1643), .B0(n1845), .B1(n1969), 
        .Y(n1212) );
  AOI22X1TS U1819 ( .A0(n1649), .A1(n1648), .B0(n1647), .B1(n1646), .Y(n1651)
         );
  AOI22X1TS U1820 ( .A0(n1652), .A1(n1665), .B0(n1651), .B1(n1650), .Y(n1654)
         );
  AOI22X1TS U1821 ( .A0(n1656), .A1(n1655), .B0(n1654), .B1(n1653), .Y(n1658)
         );
  AOI32X1TS U1822 ( .A0(n1658), .A1(n358), .A2(n1657), .B0(n1882), .B1(n1970), 
        .Y(n1211) );
  AOI22X1TS U1823 ( .A0(n1662), .A1(n1661), .B0(n1660), .B1(n1659), .Y(n1664)
         );
  AOI22X1TS U1824 ( .A0(n1666), .A1(n1665), .B0(n1664), .B1(n1663), .Y(n1668)
         );
  AOI22X1TS U1825 ( .A0(n1670), .A1(n1669), .B0(n1668), .B1(n1667), .Y(n1672)
         );
  AOI32X1TS U1826 ( .A0(n1672), .A1(n425), .A2(n1671), .B0(n1923), .B1(n1971), 
        .Y(n1210) );
  AOI22X1TS U1827 ( .A0(n1852), .A1(n1673), .B0(n1685), .B1(
        \destinationAddressbuffer[7][0] ), .Y(n1676) );
  CLKBUFX2TS U1828 ( .A(n1893), .Y(n1762) );
  AOI22X1TS U1829 ( .A0(n1688), .A1(n1762), .B0(n32), .B1(n1734), .Y(n1675) );
  CLKBUFX2TS U1830 ( .A(n1702), .Y(n1856) );
  AOI22X1TS U1831 ( .A0(n58), .A1(destinationAddressIn_SOUTH[0]), .B0(n1689), 
        .B1(n1856), .Y(n1674) );
  AOI22X1TS U1832 ( .A0(n1678), .A1(n1677), .B0(n1685), .B1(
        \destinationAddressbuffer[7][1] ), .Y(n1684) );
  CLKBUFX2TS U1833 ( .A(n1902), .Y(n1770) );
  AOI22X1TS U1834 ( .A0(n1680), .A1(n1770), .B0(n1679), .B1(n1739), .Y(n1683)
         );
  CLKBUFX2TS U1835 ( .A(n1710), .Y(n1865) );
  AOI22X1TS U1836 ( .A0(n1698), .A1(destinationAddressIn_SOUTH[1]), .B0(n1681), 
        .B1(n1865), .Y(n1682) );
  AOI22X1TS U1837 ( .A0(n1673), .A1(n1686), .B0(n1685), .B1(
        \destinationAddressbuffer[7][2] ), .Y(n1693) );
  CLKBUFX2TS U1838 ( .A(n1915), .Y(n1781) );
  AOI22X1TS U1839 ( .A0(n1688), .A1(n1781), .B0(n1687), .B1(n1749), .Y(n1692)
         );
  CLKBUFX2TS U1840 ( .A(n1719), .Y(n1878) );
  AOI22X1TS U1841 ( .A0(n1690), .A1(destinationAddressIn_SOUTH[2]), .B0(n1689), 
        .B1(n1878), .Y(n1691) );
  AOI22X1TS U1842 ( .A0(n1696), .A1(n1695), .B0(n1694), .B1(
        \destinationAddressbuffer[7][3] ), .Y(n1701) );
  CLKBUFX2TS U1843 ( .A(n1927), .Y(n1791) );
  AOI22X1TS U1844 ( .A0(n42), .A1(n1791), .B0(n32), .B1(n1758), .Y(n1700) );
  CLKBUFX2TS U1845 ( .A(n1728), .Y(n1887) );
  AOI22X1TS U1846 ( .A0(n1698), .A1(destinationAddressIn_SOUTH[3]), .B0(n1697), 
        .B1(n1887), .Y(n1699) );
  AOI22X1TS U1847 ( .A0(n1892), .A1(n1726), .B0(n1716), .B1(
        \destinationAddressbuffer[6][0] ), .Y(n1706) );
  AOI22X1TS U1848 ( .A0(n87), .A1(n1762), .B0(n84), .B1(n1734), .Y(n1705) );
  CLKBUFX2TS U1849 ( .A(n1702), .Y(n1894) );
  CLKBUFX2TS U1850 ( .A(destinationAddressIn_SOUTH[0]), .Y(n1895) );
  CLKBUFX2TS U1851 ( .A(n1895), .Y(n1854) );
  AOI22X1TS U1852 ( .A0(n1721), .A1(n1894), .B0(n1703), .B1(n1854), .Y(n1704)
         );
  AOI22X1TS U1853 ( .A0(n1768), .A1(n1707), .B0(n1716), .B1(
        \destinationAddressbuffer[6][1] ), .Y(n1715) );
  AOI22X1TS U1854 ( .A0(n1709), .A1(n1770), .B0(n1708), .B1(n1739), .Y(n1714)
         );
  CLKBUFX2TS U1855 ( .A(n1710), .Y(n1904) );
  CLKBUFX2TS U1856 ( .A(destinationAddressIn_SOUTH[1]), .Y(n1906) );
  CLKBUFX2TS U1857 ( .A(n1906), .Y(n1864) );
  AOI22X1TS U1858 ( .A0(n1712), .A1(n1904), .B0(n1711), .B1(n1864), .Y(n1713)
         );
  AOI22X1TS U1859 ( .A0(n1779), .A1(n1717), .B0(n1716), .B1(
        \destinationAddressbuffer[6][2] ), .Y(n1724) );
  AOI22X1TS U1860 ( .A0(n87), .A1(n1781), .B0(n1718), .B1(n1749), .Y(n1723) );
  CLKBUFX2TS U1861 ( .A(n1719), .Y(n1917) );
  CLKBUFX2TS U1862 ( .A(destinationAddressIn_SOUTH[2]), .Y(n1919) );
  CLKBUFX2TS U1863 ( .A(n1919), .Y(n1876) );
  AOI22X1TS U1864 ( .A0(n1721), .A1(n1917), .B0(n1720), .B1(n1876), .Y(n1722)
         );
  AOI22X1TS U1865 ( .A0(n1790), .A1(n1726), .B0(n1725), .B1(
        \destinationAddressbuffer[6][3] ), .Y(n1733) );
  AOI22X1TS U1866 ( .A0(n1727), .A1(n1791), .B0(n84), .B1(n1758), .Y(n1732) );
  CLKBUFX2TS U1867 ( .A(n1728), .Y(n1928) );
  CLKBUFX2TS U1868 ( .A(destinationAddressIn_SOUTH[3]), .Y(n1929) );
  CLKBUFX2TS U1869 ( .A(n1929), .Y(n1886) );
  AOI22X1TS U1870 ( .A0(n1730), .A1(n1928), .B0(n1729), .B1(n1886), .Y(n1731)
         );
  AOI22X1TS U1871 ( .A0(n1892), .A1(n225), .B0(n1747), .B1(
        \destinationAddressbuffer[5][0] ), .Y(n1737) );
  AOI22X1TS U1872 ( .A0(n1751), .A1(n1762), .B0(n224), .B1(n1734), .Y(n1736)
         );
  AOI22X1TS U1873 ( .A0(n1753), .A1(n1894), .B0(n1742), .B1(
        destinationAddressIn_SOUTH[0]), .Y(n1735) );
  AOI22X1TS U1874 ( .A0(readRequesterAddress[1]), .A1(n1738), .B0(n1747), .B1(
        \destinationAddressbuffer[5][1] ), .Y(n1746) );
  AOI22X1TS U1875 ( .A0(n1741), .A1(n1770), .B0(n1740), .B1(n1739), .Y(n1745)
         );
  AOI22X1TS U1876 ( .A0(n1743), .A1(n1904), .B0(n1742), .B1(
        destinationAddressIn_SOUTH[1]), .Y(n1744) );
  AOI22X1TS U1877 ( .A0(readRequesterAddress[2]), .A1(n1748), .B0(n1747), .B1(
        \destinationAddressbuffer[5][2] ), .Y(n1756) );
  AOI22X1TS U1878 ( .A0(n1751), .A1(n1781), .B0(n1750), .B1(n1749), .Y(n1755)
         );
  AOI22X1TS U1879 ( .A0(n1753), .A1(n1917), .B0(n1752), .B1(
        destinationAddressIn_SOUTH[2]), .Y(n1754) );
  AOI22X1TS U1880 ( .A0(readRequesterAddress[3]), .A1(n225), .B0(n1757), .B1(
        \destinationAddressbuffer[5][3] ), .Y(n1761) );
  AOI22X1TS U1881 ( .A0(n227), .A1(n1791), .B0(n224), .B1(n1758), .Y(n1760) );
  AOI22X1TS U1882 ( .A0(n1446), .A1(n1928), .B0(n1467), .B1(
        destinationAddressIn_SOUTH[3]), .Y(n1759) );
  AOI22X1TS U1883 ( .A0(n1796), .A1(n1789), .B0(n1777), .B1(
        \destinationAddressbuffer[4][0] ), .Y(n1766) );
  AOI22X1TS U1884 ( .A0(n1782), .A1(n1762), .B0(n274), .B1(
        destinationAddressIn_EAST[0]), .Y(n1765) );
  AOI22X1TS U1885 ( .A0(n1763), .A1(n1895), .B0(n1783), .B1(n1894), .Y(n1764)
         );
  AOI22X1TS U1886 ( .A0(n1768), .A1(n1767), .B0(n1777), .B1(
        \destinationAddressbuffer[4][1] ), .Y(n1776) );
  AOI22X1TS U1887 ( .A0(n1771), .A1(n1770), .B0(n1769), .B1(
        destinationAddressIn_EAST[1]), .Y(n1775) );
  AOI22X1TS U1888 ( .A0(n1773), .A1(n1906), .B0(n1772), .B1(n1904), .Y(n1774)
         );
  AOI22X1TS U1889 ( .A0(n1779), .A1(n1778), .B0(n1777), .B1(
        \destinationAddressbuffer[4][2] ), .Y(n1787) );
  AOI22X1TS U1890 ( .A0(n1782), .A1(n1781), .B0(n1780), .B1(
        destinationAddressIn_EAST[2]), .Y(n1786) );
  AOI22X1TS U1891 ( .A0(n1784), .A1(n1919), .B0(n1783), .B1(n1917), .Y(n1785)
         );
  AOI22X1TS U1892 ( .A0(n1790), .A1(n1789), .B0(n1788), .B1(
        \destinationAddressbuffer[4][3] ), .Y(n1795) );
  AOI22X1TS U1893 ( .A0(n296), .A1(n1791), .B0(n274), .B1(
        destinationAddressIn_EAST[3]), .Y(n1794) );
  AOI22X1TS U1894 ( .A0(n284), .A1(n1929), .B0(n1792), .B1(n1928), .Y(n1793)
         );
  AOI22X1TS U1895 ( .A0(n1796), .A1(n1817), .B0(n1809), .B1(
        \destinationAddressbuffer[3][0] ), .Y(n1800) );
  AOI22X1TS U1896 ( .A0(n1804), .A1(n1797), .B0(n1802), .B1(
        destinationAddressIn_EAST[0]), .Y(n1799) );
  AOI22X1TS U1897 ( .A0(n1822), .A1(n1856), .B0(n1409), .B1(n1854), .Y(n1798)
         );
  AOI22X1TS U1898 ( .A0(n1861), .A1(n1801), .B0(n1809), .B1(
        \destinationAddressbuffer[3][1] ), .Y(n1808) );
  AOI22X1TS U1899 ( .A0(n1804), .A1(n1803), .B0(n1802), .B1(
        destinationAddressIn_EAST[1]), .Y(n1807) );
  AOI22X1TS U1900 ( .A0(n1805), .A1(n1865), .B0(n1821), .B1(n1864), .Y(n1806)
         );
  AOI22X1TS U1901 ( .A0(n1872), .A1(n131), .B0(n1809), .B1(
        \destinationAddressbuffer[3][2] ), .Y(n1815) );
  AOI22X1TS U1902 ( .A0(n139), .A1(n1811), .B0(n1810), .B1(
        destinationAddressIn_EAST[2]), .Y(n1814) );
  AOI22X1TS U1903 ( .A0(n1812), .A1(n1878), .B0(n129), .B1(n1876), .Y(n1813)
         );
  AOI22X1TS U1904 ( .A0(n1883), .A1(n1817), .B0(n1816), .B1(
        \destinationAddressbuffer[3][3] ), .Y(n1825) );
  AOI22X1TS U1905 ( .A0(n1820), .A1(n1819), .B0(n1818), .B1(
        destinationAddressIn_EAST[3]), .Y(n1824) );
  AOI22X1TS U1906 ( .A0(n1822), .A1(n1887), .B0(n1821), .B1(n1886), .Y(n1823)
         );
  AOI22X1TS U1907 ( .A0(n1852), .A1(n1846), .B0(n1836), .B1(
        \destinationAddressbuffer[2][0] ), .Y(n1828) );
  AOI22X1TS U1908 ( .A0(n1839), .A1(destinationAddressIn_WEST[0]), .B0(n1847), 
        .B1(n1853), .Y(n1827) );
  AOI22X1TS U1909 ( .A0(n198), .A1(n1856), .B0(n1840), .B1(n1854), .Y(n1826)
         );
  AOI22X1TS U1910 ( .A0(n1901), .A1(n1829), .B0(n1836), .B1(
        \destinationAddressbuffer[2][1] ), .Y(n1835) );
  AOI22X1TS U1911 ( .A0(n1830), .A1(destinationAddressIn_WEST[1]), .B0(n987), 
        .B1(n1862), .Y(n1834) );
  AOI22X1TS U1912 ( .A0(n1832), .A1(n1865), .B0(n1831), .B1(n1864), .Y(n1833)
         );
  AOI22X1TS U1913 ( .A0(n1913), .A1(n1837), .B0(n1836), .B1(
        \destinationAddressbuffer[2][2] ), .Y(n1844) );
  AOI22X1TS U1914 ( .A0(n1839), .A1(destinationAddressIn_WEST[2]), .B0(n1838), 
        .B1(n1873), .Y(n1843) );
  AOI22X1TS U1915 ( .A0(n1841), .A1(n1878), .B0(n1840), .B1(n1876), .Y(n1842)
         );
  AOI22X1TS U1916 ( .A0(n1925), .A1(n1846), .B0(n1845), .B1(
        \destinationAddressbuffer[2][3] ), .Y(n1851) );
  AOI22X1TS U1917 ( .A0(n208), .A1(destinationAddressIn_WEST[3]), .B0(n1847), 
        .B1(n1884), .Y(n1850) );
  AOI22X1TS U1918 ( .A0(n1848), .A1(n1887), .B0(n194), .B1(n1886), .Y(n1849)
         );
  AOI22X1TS U1919 ( .A0(n1852), .A1(n319), .B0(n1870), .B1(
        \destinationAddressbuffer[1][0] ), .Y(n1859) );
  AOI22X1TS U1920 ( .A0(n1875), .A1(n1893), .B0(n1885), .B1(n1853), .Y(n1858)
         );
  AOI22X1TS U1921 ( .A0(n1008), .A1(n1856), .B0(n1855), .B1(n1854), .Y(n1857)
         );
  AOI22X1TS U1922 ( .A0(n1861), .A1(n1860), .B0(n1870), .B1(
        \destinationAddressbuffer[1][1] ), .Y(n1869) );
  AOI22X1TS U1923 ( .A0(n1863), .A1(n1902), .B0(n1015), .B1(n1862), .Y(n1868)
         );
  AOI22X1TS U1924 ( .A0(n1866), .A1(n1865), .B0(n349), .B1(n1864), .Y(n1867)
         );
  AOI22X1TS U1925 ( .A0(n1872), .A1(n1871), .B0(n1870), .B1(
        \destinationAddressbuffer[1][2] ), .Y(n1881) );
  AOI22X1TS U1926 ( .A0(n1875), .A1(n1915), .B0(n1874), .B1(n1873), .Y(n1880)
         );
  AOI22X1TS U1927 ( .A0(n1008), .A1(n1878), .B0(n1877), .B1(n1876), .Y(n1879)
         );
  AOI22X1TS U1928 ( .A0(n1883), .A1(n319), .B0(n1882), .B1(
        \destinationAddressbuffer[1][3] ), .Y(n1891) );
  AOI22X1TS U1929 ( .A0(n378), .A1(n1927), .B0(n1885), .B1(n1884), .Y(n1890)
         );
  AOI22X1TS U1930 ( .A0(n1888), .A1(n1887), .B0(n366), .B1(n1886), .Y(n1889)
         );
  AOI22X1TS U1931 ( .A0(n1892), .A1(n1924), .B0(n1911), .B1(
        \destinationAddressbuffer[0][0] ), .Y(n1899) );
  AOI22X1TS U1932 ( .A0(n1916), .A1(n1893), .B0(n1926), .B1(
        destinationAddressIn_EAST[0]), .Y(n1898) );
  AOI22X1TS U1933 ( .A0(n1896), .A1(n1895), .B0(n1918), .B1(n1894), .Y(n1897)
         );
  AOI22X1TS U1934 ( .A0(n1901), .A1(n1900), .B0(n1911), .B1(
        \destinationAddressbuffer[0][1] ), .Y(n1910) );
  AOI22X1TS U1935 ( .A0(n1903), .A1(n1902), .B0(n410), .B1(
        destinationAddressIn_EAST[1]), .Y(n1909) );
  AOI22X1TS U1936 ( .A0(n1907), .A1(n1906), .B0(n1905), .B1(n1904), .Y(n1908)
         );
  AOI22X1TS U1937 ( .A0(n1913), .A1(n1912), .B0(n1911), .B1(
        \destinationAddressbuffer[0][2] ), .Y(n1922) );
  AOI22X1TS U1938 ( .A0(n1916), .A1(n1915), .B0(n1914), .B1(
        destinationAddressIn_EAST[2]), .Y(n1921) );
  AOI22X1TS U1939 ( .A0(n427), .A1(n1919), .B0(n1918), .B1(n1917), .Y(n1920)
         );
  AOI22X1TS U1940 ( .A0(n1925), .A1(n1924), .B0(n1923), .B1(
        \destinationAddressbuffer[0][3] ), .Y(n1933) );
  AOI22X1TS U1941 ( .A0(n430), .A1(n1927), .B0(n1926), .B1(
        destinationAddressIn_EAST[3]), .Y(n1932) );
  AOI22X1TS U1942 ( .A0(n1930), .A1(n1929), .B0(n407), .B1(n1928), .Y(n1931)
         );
endmodule


module outputPortArbiter_1 ( clk, reset, selectBit_NORTH, 
        destinationAddressIn_NORTH, requesterAddressIn_NORTH, readIn_NORTH, 
        writeIn_NORTH, dataIn_NORTH, selectBit_SOUTH, 
        destinationAddressIn_SOUTH, requesterAddressIn_SOUTH, readIn_SOUTH, 
        writeIn_SOUTH, dataIn_SOUTH, selectBit_EAST, destinationAddressIn_EAST, 
        requesterAddressIn_EAST, readIn_EAST, writeIn_EAST, dataIn_EAST, 
        selectBit_WEST, destinationAddressIn_WEST, requesterAddressIn_WEST, 
        readIn_WEST, writeIn_WEST, dataIn_WEST, readReady, 
        readRequesterAddress, cacheDataOut, destinationAddressOut, 
        requesterAddressOut, readOut, writeOut, dataOut );
  input [11:0] destinationAddressIn_NORTH;
  input [3:0] requesterAddressIn_NORTH;
  input [5:0] dataIn_NORTH;
  input [11:0] destinationAddressIn_SOUTH;
  input [3:0] requesterAddressIn_SOUTH;
  input [5:0] dataIn_SOUTH;
  input [11:0] destinationAddressIn_EAST;
  input [3:0] requesterAddressIn_EAST;
  input [5:0] dataIn_EAST;
  input [11:0] destinationAddressIn_WEST;
  input [3:0] requesterAddressIn_WEST;
  input [5:0] dataIn_WEST;
  input [3:0] readRequesterAddress;
  input [5:0] cacheDataOut;
  output [11:0] destinationAddressOut;
  output [3:0] requesterAddressOut;
  output [5:0] dataOut;
  input clk, reset, selectBit_NORTH, readIn_NORTH, writeIn_NORTH,
         selectBit_SOUTH, readIn_SOUTH, writeIn_SOUTH, selectBit_EAST,
         readIn_EAST, writeIn_EAST, selectBit_WEST, readIn_WEST, writeIn_WEST,
         readReady;
  output readOut, writeOut;
  wire   \requesterAddressbuffer[0][3] , \requesterAddressbuffer[0][2] ,
         \requesterAddressbuffer[0][1] , \requesterAddressbuffer[0][0] ,
         \requesterAddressbuffer[1][3] , \requesterAddressbuffer[1][2] ,
         \requesterAddressbuffer[1][1] , \requesterAddressbuffer[1][0] ,
         \requesterAddressbuffer[2][3] , \requesterAddressbuffer[2][2] ,
         \requesterAddressbuffer[2][1] , \requesterAddressbuffer[2][0] ,
         \requesterAddressbuffer[3][3] , \requesterAddressbuffer[3][2] ,
         \requesterAddressbuffer[3][1] , \requesterAddressbuffer[3][0] ,
         \requesterAddressbuffer[4][3] , \requesterAddressbuffer[4][2] ,
         \requesterAddressbuffer[4][1] , \requesterAddressbuffer[4][0] ,
         \requesterAddressbuffer[5][3] , \requesterAddressbuffer[5][2] ,
         \requesterAddressbuffer[5][1] , \requesterAddressbuffer[5][0] ,
         \requesterAddressbuffer[6][3] , \requesterAddressbuffer[6][2] ,
         \requesterAddressbuffer[6][1] , \requesterAddressbuffer[6][0] ,
         \requesterAddressbuffer[7][3] , \requesterAddressbuffer[7][2] ,
         \requesterAddressbuffer[7][1] , \requesterAddressbuffer[7][0] ,
         \destinationAddressbuffer[0][11] , \destinationAddressbuffer[0][10] ,
         \destinationAddressbuffer[0][9] , \destinationAddressbuffer[0][8] ,
         \destinationAddressbuffer[0][7] , \destinationAddressbuffer[0][6] ,
         \destinationAddressbuffer[0][5] , \destinationAddressbuffer[0][4] ,
         \destinationAddressbuffer[0][3] , \destinationAddressbuffer[0][2] ,
         \destinationAddressbuffer[0][1] , \destinationAddressbuffer[0][0] ,
         \destinationAddressbuffer[1][11] , \destinationAddressbuffer[1][10] ,
         \destinationAddressbuffer[1][9] , \destinationAddressbuffer[1][8] ,
         \destinationAddressbuffer[1][7] , \destinationAddressbuffer[1][6] ,
         \destinationAddressbuffer[1][5] , \destinationAddressbuffer[1][4] ,
         \destinationAddressbuffer[1][3] , \destinationAddressbuffer[1][2] ,
         \destinationAddressbuffer[1][1] , \destinationAddressbuffer[1][0] ,
         \destinationAddressbuffer[2][11] , \destinationAddressbuffer[2][10] ,
         \destinationAddressbuffer[2][9] , \destinationAddressbuffer[2][8] ,
         \destinationAddressbuffer[2][7] , \destinationAddressbuffer[2][6] ,
         \destinationAddressbuffer[2][5] , \destinationAddressbuffer[2][4] ,
         \destinationAddressbuffer[2][3] , \destinationAddressbuffer[2][2] ,
         \destinationAddressbuffer[2][1] , \destinationAddressbuffer[2][0] ,
         \destinationAddressbuffer[3][11] , \destinationAddressbuffer[3][10] ,
         \destinationAddressbuffer[3][9] , \destinationAddressbuffer[3][8] ,
         \destinationAddressbuffer[3][7] , \destinationAddressbuffer[3][6] ,
         \destinationAddressbuffer[3][5] , \destinationAddressbuffer[3][4] ,
         \destinationAddressbuffer[3][3] , \destinationAddressbuffer[3][2] ,
         \destinationAddressbuffer[3][1] , \destinationAddressbuffer[3][0] ,
         \destinationAddressbuffer[4][11] , \destinationAddressbuffer[4][10] ,
         \destinationAddressbuffer[4][9] , \destinationAddressbuffer[4][8] ,
         \destinationAddressbuffer[4][7] , \destinationAddressbuffer[4][6] ,
         \destinationAddressbuffer[4][5] , \destinationAddressbuffer[4][4] ,
         \destinationAddressbuffer[4][3] , \destinationAddressbuffer[4][2] ,
         \destinationAddressbuffer[4][1] , \destinationAddressbuffer[4][0] ,
         \destinationAddressbuffer[5][11] , \destinationAddressbuffer[5][10] ,
         \destinationAddressbuffer[5][9] , \destinationAddressbuffer[5][8] ,
         \destinationAddressbuffer[5][7] , \destinationAddressbuffer[5][6] ,
         \destinationAddressbuffer[5][5] , \destinationAddressbuffer[5][4] ,
         \destinationAddressbuffer[5][3] , \destinationAddressbuffer[5][2] ,
         \destinationAddressbuffer[5][1] , \destinationAddressbuffer[5][0] ,
         \destinationAddressbuffer[6][11] , \destinationAddressbuffer[6][10] ,
         \destinationAddressbuffer[6][9] , \destinationAddressbuffer[6][8] ,
         \destinationAddressbuffer[6][7] , \destinationAddressbuffer[6][6] ,
         \destinationAddressbuffer[6][5] , \destinationAddressbuffer[6][4] ,
         \destinationAddressbuffer[6][3] , \destinationAddressbuffer[6][2] ,
         \destinationAddressbuffer[6][1] , \destinationAddressbuffer[6][0] ,
         \destinationAddressbuffer[7][11] , \destinationAddressbuffer[7][10] ,
         \destinationAddressbuffer[7][9] , \destinationAddressbuffer[7][8] ,
         \destinationAddressbuffer[7][7] , \destinationAddressbuffer[7][6] ,
         \destinationAddressbuffer[7][5] , \destinationAddressbuffer[7][4] ,
         \destinationAddressbuffer[7][3] , \destinationAddressbuffer[7][2] ,
         \destinationAddressbuffer[7][1] , \destinationAddressbuffer[7][0] ,
         \dataoutbuffer[7][5] , \dataoutbuffer[7][4] , \dataoutbuffer[7][3] ,
         \dataoutbuffer[7][2] , \dataoutbuffer[7][1] , \dataoutbuffer[7][0] ,
         \dataoutbuffer[6][5] , \dataoutbuffer[6][4] , \dataoutbuffer[6][3] ,
         \dataoutbuffer[6][2] , \dataoutbuffer[6][1] , \dataoutbuffer[6][0] ,
         \dataoutbuffer[5][5] , \dataoutbuffer[5][4] , \dataoutbuffer[5][3] ,
         \dataoutbuffer[5][2] , \dataoutbuffer[5][1] , \dataoutbuffer[5][0] ,
         \dataoutbuffer[4][5] , \dataoutbuffer[4][4] , \dataoutbuffer[4][3] ,
         \dataoutbuffer[4][2] , \dataoutbuffer[4][1] , \dataoutbuffer[4][0] ,
         \dataoutbuffer[3][5] , \dataoutbuffer[3][4] , \dataoutbuffer[3][3] ,
         \dataoutbuffer[3][2] , \dataoutbuffer[3][1] , \dataoutbuffer[3][0] ,
         \dataoutbuffer[2][5] , \dataoutbuffer[2][4] , \dataoutbuffer[2][3] ,
         \dataoutbuffer[2][2] , \dataoutbuffer[2][1] , \dataoutbuffer[2][0] ,
         \dataoutbuffer[1][5] , \dataoutbuffer[1][4] , \dataoutbuffer[1][3] ,
         \dataoutbuffer[1][2] , \dataoutbuffer[1][1] , \dataoutbuffer[1][0] ,
         \dataoutbuffer[0][5] , \dataoutbuffer[0][4] , \dataoutbuffer[0][3] ,
         \dataoutbuffer[0][2] , \dataoutbuffer[0][1] , \dataoutbuffer[0][0] ,
         N2624, n1, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
         n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
         n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
         n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
         n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
         n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
         n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188;
  wire   [0:7] writeOutbuffer;
  wire   [0:7] readOutbuffer;

  DFFNSRX1TS full_reg_reg ( .D(N2624), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(
        n1957) );
  DFFNSRX1TS \requesterAddressbuffer_reg[2][0]  ( .D(n2017), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[2][1]  ( .D(n2018), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[2][2]  ( .D(n2019), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[2][3]  ( .D(n2020), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][0]  ( .D(n2153), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][1]  ( .D(n2154), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][2]  ( .D(n2155), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][3]  ( .D(n2156), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][0]  ( .D(n2029), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][1]  ( .D(n2030), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][2]  ( .D(n2031), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][3]  ( .D(n2032), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][4]  ( .D(n2033), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][5]  ( .D(n2034), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][5] ) );
  DFFNSRX1TS \writeOutbuffer_reg[7]  ( .D(n2077), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[7]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][4]  ( .D(n2097), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][5]  ( .D(n2098), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][6]  ( .D(n2099), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][7]  ( .D(n2100), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][8]  ( .D(n2101), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][9]  ( .D(n2102), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][11]  ( .D(n2104), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[6]  ( .D(n2078), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[6]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][4]  ( .D(n2109), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][5]  ( .D(n2110), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][6]  ( .D(n2111), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][7]  ( .D(n2112), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][8]  ( .D(n2113), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][9]  ( .D(n2114), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][10]  ( .D(n2115), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][11]  ( .D(n2116), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[3]  ( .D(n2081), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[3]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][4]  ( .D(n2145), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][5]  ( .D(n2146), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][6]  ( .D(n2147), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][7]  ( .D(n2148), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][8]  ( .D(n2149), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][9]  ( .D(n2150), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][10]  ( .D(n2151), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][11]  ( .D(n2152), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[2]  ( .D(n2082), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[2]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][4]  ( .D(n2157), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][5]  ( .D(n2158), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][6]  ( .D(n2159), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][7]  ( .D(n2160), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][8]  ( .D(n2161), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][9]  ( .D(n2162), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][10]  ( .D(n2163), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][11]  ( .D(n2164), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][11] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][0]  ( .D(n2071), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][1]  ( .D(n2072), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][2]  ( .D(n2073), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][3]  ( .D(n2074), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][4]  ( .D(n2075), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][5]  ( .D(n2076), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][0]  ( .D(n2065), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][1]  ( .D(n2066), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][2]  ( .D(n2067), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][3]  ( .D(n2068), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][4]  ( .D(n2069), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][5]  ( .D(n2070), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][5] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[5][0]  ( .D(n2005), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[5][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[5][1]  ( .D(n2006), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[5][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[5][2]  ( .D(n2007), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[5][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[5][3]  ( .D(n2008), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[5][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][0]  ( .D(n2117), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][1]  ( .D(n2118), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][2]  ( .D(n2119), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][3]  ( .D(n2120), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[4][0]  ( .D(n2009), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[4][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[4][1]  ( .D(n2010), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[4][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[4][2]  ( .D(n2011), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[4][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[4][3]  ( .D(n2012), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[4][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][0]  ( .D(n2129), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][1]  ( .D(n2130), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][2]  ( .D(n2131), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][3]  ( .D(n2132), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][0]  ( .D(n2047), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][1]  ( .D(n2048), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][2]  ( .D(n2049), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][3]  ( .D(n2050), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][4]  ( .D(n2051), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][5]  ( .D(n2052), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][0]  ( .D(n2041), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][1]  ( .D(n2042), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][2]  ( .D(n2043), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][3]  ( .D(n2044), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][4]  ( .D(n2045), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][5]  ( .D(n2046), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][5] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[1][0]  ( .D(n2021), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[1][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[1][1]  ( .D(n2022), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[1][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[1][2]  ( .D(n2023), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[1][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[1][3]  ( .D(n2024), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[1][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][0]  ( .D(n2165), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][1]  ( .D(n2166), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][2]  ( .D(n2167), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][3]  ( .D(n2168), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[0][0]  ( .D(n2025), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[0][1]  ( .D(n2026), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[0][2]  ( .D(n2027), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[0][3]  ( .D(n2028), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][0]  ( .D(n2177), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][1]  ( .D(n2178), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][2]  ( .D(n2179), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][3]  ( .D(n2180), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[7][0]  ( .D(n1997), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[7][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[7][1]  ( .D(n1998), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[7][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[7][2]  ( .D(n1999), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[7][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[7][3]  ( .D(n2000), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[7][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][0]  ( .D(n2093), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][1]  ( .D(n2094), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][2]  ( .D(n2095), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][3]  ( .D(n2096), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[6][0]  ( .D(n2001), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[6][1]  ( .D(n2002), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[6][2]  ( .D(n2003), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[6][3]  ( .D(n2004), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][0]  ( .D(n2105), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][1]  ( .D(n2106), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][2]  ( .D(n2107), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][3]  ( .D(n2108), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][0]  ( .D(n2059), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][1]  ( .D(n2060), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][2]  ( .D(n2061), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][3]  ( .D(n2062), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][4]  ( .D(n2063), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][5]  ( .D(n2064), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][0]  ( .D(n2053), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][1]  ( .D(n2054), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][2]  ( .D(n2055), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][3]  ( .D(n2056), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][4]  ( .D(n2057), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][5]  ( .D(n2058), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][5] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[3][0]  ( .D(n2013), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[3][1]  ( .D(n2014), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[3][2]  ( .D(n2015), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[3][3]  ( .D(n2016), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][0]  ( .D(n2141), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][1]  ( .D(n2142), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][2]  ( .D(n2143), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][3]  ( .D(n2144), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][0]  ( .D(n2035), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][1]  ( .D(n2036), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][2]  ( .D(n2037), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][3]  ( .D(n2038), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][4]  ( .D(n2039), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][5]  ( .D(n2040), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][5] ) );
  DFFNSRX1TS \writeOutbuffer_reg[5]  ( .D(n2079), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[5]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][4]  ( .D(n2121), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][5]  ( .D(n2122), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][6]  ( .D(n2123), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][7]  ( .D(n2124), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][8]  ( .D(n2125), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][9]  ( .D(n2126), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][10]  ( .D(n2127), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][11]  ( .D(n2128), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[4]  ( .D(n2080), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[4]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][4]  ( .D(n2133), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][5]  ( .D(n2134), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][6]  ( .D(n2135), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][7]  ( .D(n2136), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][8]  ( .D(n2137), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][9]  ( .D(n2138), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][10]  ( .D(n2139), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][11]  ( .D(n2140), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[1]  ( .D(n2083), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[1]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][4]  ( .D(n2169), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][5]  ( .D(n2170), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][6]  ( .D(n2171), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][7]  ( .D(n2172), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][8]  ( .D(n2173), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][9]  ( .D(n2174), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][10]  ( .D(n2175), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][11]  ( .D(n2176), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[0]  ( .D(n2084), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[0]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][4]  ( .D(n2181), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][5]  ( .D(n2182), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][6]  ( .D(n2183), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][7]  ( .D(n2184), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][8]  ( .D(n2185), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][9]  ( .D(n2186), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][10]  ( .D(n2187), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][11]  ( .D(n2188), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][11] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][10]  ( .D(n2103), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][10] ) );
  DFFNSRX1TS writeOut_reg ( .D(n1974), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        writeOut) );
  DFFNSRX1TS \destinationAddressOut_reg[4]  ( .D(n1983), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[4]) );
  DFFNSRX1TS \destinationAddressOut_reg[5]  ( .D(n1984), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[5]) );
  DFFNSRX1TS \destinationAddressOut_reg[6]  ( .D(n1985), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[6]) );
  DFFNSRX1TS \destinationAddressOut_reg[7]  ( .D(n1986), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[7]) );
  DFFNSRX1TS \destinationAddressOut_reg[8]  ( .D(n1987), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[8]) );
  DFFNSRX1TS \destinationAddressOut_reg[9]  ( .D(n1988), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[9]) );
  DFFNSRX1TS \destinationAddressOut_reg[10]  ( .D(n1989), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[10]) );
  DFFNSRX1TS \destinationAddressOut_reg[11]  ( .D(n1990), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[11]) );
  DFFNSRX1TS readOut_reg ( .D(n1973), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        readOut) );
  DFFNSRX1TS \requesterAddressOut_reg[0]  ( .D(n1975), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[0]) );
  DFFNSRX1TS \requesterAddressOut_reg[1]  ( .D(n1976), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[1]) );
  DFFNSRX1TS \requesterAddressOut_reg[2]  ( .D(n1977), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[2]) );
  DFFNSRX1TS \requesterAddressOut_reg[3]  ( .D(n1978), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[3]) );
  DFFNSRX1TS \destinationAddressOut_reg[0]  ( .D(n1979), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[0]) );
  DFFNSRX1TS \destinationAddressOut_reg[1]  ( .D(n1980), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[1]) );
  DFFNSRX1TS \destinationAddressOut_reg[2]  ( .D(n1981), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[2]) );
  DFFNSRX1TS \destinationAddressOut_reg[3]  ( .D(n1982), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[3]) );
  DFFNSRX1TS \dataOut_reg[0]  ( .D(n1991), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[0]) );
  DFFNSRX1TS \dataOut_reg[1]  ( .D(n1992), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[1]) );
  DFFNSRX1TS \dataOut_reg[2]  ( .D(n1993), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[2]) );
  DFFNSRX1TS \dataOut_reg[3]  ( .D(n1994), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[3]) );
  DFFNSRX1TS \dataOut_reg[4]  ( .D(n1995), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[4]) );
  DFFNSRX1TS \dataOut_reg[5]  ( .D(n1996), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[5]) );
  DFFNSRX1TS \read_reg_reg[1]  ( .D(n1972), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1950), .QN(n1949) );
  DFFNSRX1TS \write_reg_reg[0]  ( .D(n1967), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1948), .QN(n1952) );
  DFFNSRX1TS \write_reg_reg[2]  ( .D(n1969), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1953), .QN(n1954) );
  DFFNSRX1TS \read_reg_reg[0]  ( .D(n1966), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1943), .QN(n1955) );
  DFFNSRX1TS \read_reg_reg[2]  ( .D(n1971), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1946), .QN(n1947) );
  DFFNSRX1TS empty_reg_reg ( .D(n1970), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        n1945), .QN(n1944) );
  DFFNSRX1TS \readOutbuffer_reg[7]  ( .D(n2085), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[7]), .QN(n1958) );
  DFFNSRX1TS \readOutbuffer_reg[4]  ( .D(n2088), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[4]), .QN(n1961) );
  DFFNSRX1TS \readOutbuffer_reg[6]  ( .D(n2086), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[6]), .QN(n1959) );
  DFFNSRX1TS \readOutbuffer_reg[5]  ( .D(n2087), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[5]), .QN(n1960) );
  DFFNSRX1TS \readOutbuffer_reg[1]  ( .D(n2091), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[1]), .QN(n1964) );
  DFFNSRX1TS \readOutbuffer_reg[2]  ( .D(n2090), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[2]), .QN(n1963) );
  DFFNSRX1TS \readOutbuffer_reg[0]  ( .D(n2092), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[0]), .QN(n1965) );
  DFFNSRX1TS \readOutbuffer_reg[3]  ( .D(n2089), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[3]), .QN(n1962) );
  DFFNSRX1TS \write_reg_reg[1]  ( .D(n1968), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1951), .QN(n1956) );
  CLKBUFX2TS U3 ( .A(n16), .Y(n218) );
  CMPR32X2TS U4 ( .A(n470), .B(n501), .C(n18), .CO(n19), .S(n16) );
  CMPR32X2TS U5 ( .A(n536), .B(n468), .C(n467), .CO(n459), .S(n473) );
  ADDFX1TS U6 ( .A(selectBit_SOUTH), .B(selectBit_NORTH), .CI(selectBit_EAST), 
        .CO(n470), .S(n465) );
  CLKBUFX2TS U7 ( .A(n20), .Y(n21) );
  CLKBUFX2TS U8 ( .A(n22), .Y(n82) );
  NOR3XLTS U9 ( .A(n518), .B(selectBit_EAST), .C(n520), .Y(n513) );
  NOR2XLTS U10 ( .A(n1608), .B(n280), .Y(n293) );
  NOR2XLTS U11 ( .A(n1573), .B(n40), .Y(n45) );
  NOR2XLTS U12 ( .A(n126), .B(n390), .Y(n1622) );
  ADDHXLTS U13 ( .A(n452), .B(n465), .CO(n18), .S(n17) );
  INVX2TS U14 ( .A(n1612), .Y(n1610) );
  INVX2TS U15 ( .A(n1601), .Y(n1599) );
  INVX2TS U16 ( .A(n1588), .Y(n1586) );
  INVX2TS U17 ( .A(n1577), .Y(n1575) );
  INVX2TS U18 ( .A(n1651), .Y(n1648) );
  INVX2TS U19 ( .A(n1591), .Y(n1589) );
  NOR2XLTS U20 ( .A(selectBit_NORTH), .B(n511), .Y(n544) );
  NOR2XLTS U21 ( .A(n1641), .B(n325), .Y(n326) );
  NOR2XLTS U22 ( .A(n1623), .B(n135), .Y(n136) );
  NOR2XLTS U23 ( .A(n319), .B(n1652), .Y(n320) );
  NOR2XLTS U24 ( .A(n319), .B(n1626), .Y(n132) );
  NOR2XLTS U25 ( .A(n275), .B(n1617), .Y(n276) );
  NOR3XLTS U26 ( .A(n1604), .B(n1599), .C(n226), .Y(n222) );
  NOR2XLTS U27 ( .A(n447), .B(n1592), .Y(n87) );
  NOR2XLTS U28 ( .A(n1581), .B(n32), .Y(n36) );
  NOR2XLTS U29 ( .A(n1629), .B(n185), .Y(n186) );
  NOR2XLTS U30 ( .A(n28), .B(n134), .Y(n131) );
  OAI21XLTS U31 ( .A0(n496), .A1(n531), .B0(n493), .Y(n494) );
  AOI211XLTS U32 ( .A0(n496), .A1(n531), .B0(n495), .C0(n494), .Y(n497) );
  NOR3XLTS U33 ( .A(n1637), .B(n1631), .C(n183), .Y(n1) );
  NOR2X1TS U34 ( .A(n1598), .B(n227), .Y(n237) );
  NOR2X1TS U35 ( .A(n1644), .B(n325), .Y(n332) );
  NOR2X1TS U36 ( .A(n1630), .B(n185), .Y(n194) );
  NAND2BXLTS U37 ( .AN(n91), .B(n90), .Y(n93) );
  NAND2BXLTS U38 ( .AN(n403), .B(n402), .Y(n404) );
  NAND2BXLTS U39 ( .AN(n279), .B(n278), .Y(n280) );
  NAND2BXLTS U40 ( .AN(n183), .B(n182), .Y(n185) );
  NAND2BXLTS U41 ( .AN(n324), .B(n323), .Y(n325) );
  NOR2X1TS U42 ( .A(n126), .B(n270), .Y(n1577) );
  XOR2XLTS U43 ( .A(n530), .B(n499), .Y(n495) );
  ADDFX1TS U44 ( .A(n492), .B(n491), .CI(n490), .CO(n485), .S(n500) );
  OAI21X1TS U45 ( .A0(selectBit_SOUTH), .A1(n23), .B0(n82), .Y(n269) );
  NAND3X1TS U46 ( .A(n84), .B(n31), .C(n219), .Y(n1573) );
  INVX1TS U47 ( .A(n1637), .Y(n1635) );
  NAND3X1TS U48 ( .A(n26), .B(n219), .C(n271), .Y(n1595) );
  NOR2X1TS U49 ( .A(n219), .B(n81), .Y(n315) );
  INVX1TS U50 ( .A(n1665), .Y(n1662) );
  INVX1TS U51 ( .A(n1616), .Y(n1613) );
  AND2X2TS U52 ( .A(n529), .B(n1957), .Y(n220) );
  NAND2BX1TS U53 ( .AN(n124), .B(n466), .Y(n388) );
  NOR2X1TS U54 ( .A(n464), .B(n510), .Y(n20) );
  ADDFX1TS U55 ( .A(n466), .B(n520), .CI(n465), .CO(n469), .S(n482) );
  CLKBUFX2TS U56 ( .A(n58), .Y(n296) );
  CLKBUFX2TS U57 ( .A(readIn_EAST), .Y(n1572) );
  INVX1TS U58 ( .A(n1954), .Y(n486) );
  OR3X1TS U59 ( .A(n1651), .B(n1645), .C(n324), .Y(n4) );
  INVX2TS U60 ( .A(n4), .Y(n318) );
  NOR2X1TS U61 ( .A(n11), .B(n81), .Y(n30) );
  OAI21X1TS U62 ( .A0(n30), .A1(n27), .B0(n29), .Y(n125) );
  NAND2BX1TS U63 ( .AN(n125), .B(selectBit_EAST), .Y(n390) );
  NOR3X1TS U64 ( .A(n316), .B(n315), .C(n270), .Y(n1601) );
  NOR3BX1TS U65 ( .AN(n391), .B(n270), .C(n269), .Y(n1612) );
  NOR2XLTS U66 ( .A(n1604), .B(n1601), .Y(n225) );
  NOR3BXLTS U67 ( .AN(readReady), .B(n518), .C(n517), .Y(n543) );
  NAND2BXLTS U68 ( .AN(n135), .B(n130), .Y(n134) );
  NAND2X1TS U69 ( .A(n133), .B(n1626), .Y(n135) );
  OR2X1TS U70 ( .A(n277), .B(n937), .Y(n1422) );
  OR2X1TS U71 ( .A(n223), .B(n919), .Y(n1453) );
  OR2X1TS U72 ( .A(n181), .B(n992), .Y(n1358) );
  OR2X1TS U73 ( .A(n133), .B(n967), .Y(n1391) );
  OR2X1TS U74 ( .A(n88), .B(n900), .Y(n1487) );
  OR2X1TS U75 ( .A(n37), .B(n1668), .Y(n1537) );
  CLKAND2X2TS U76 ( .A(n484), .B(n483), .Y(n490) );
  NAND4XLTS U77 ( .A(n462), .B(n452), .C(n515), .D(n448), .Y(n1626) );
  INVX2TS U78 ( .A(n1625), .Y(n1623) );
  CLKBUFX2TS U79 ( .A(n1391), .Y(n1627) );
  NOR3XLTS U80 ( .A(n16), .B(n123), .C(n388), .Y(n1665) );
  INVX2TS U81 ( .A(n1661), .Y(n1658) );
  NOR3XLTS U82 ( .A(n17), .B(n179), .C(n388), .Y(n1637) );
  INVX2TS U83 ( .A(n1634), .Y(n1631) );
  CLKBUFX2TS U84 ( .A(n1358), .Y(n1639) );
  NAND4XLTS U85 ( .A(n453), .B(n515), .C(n450), .D(n396), .Y(n1652) );
  NOR3XLTS U86 ( .A(n16), .B(n80), .C(n388), .Y(n1651) );
  INVX2TS U87 ( .A(n1647), .Y(n1645) );
  NOR3X1TS U88 ( .A(n218), .B(n80), .C(n268), .Y(n1604) );
  CLKBUFX2TS U89 ( .A(n1453), .Y(n1606) );
  NAND4XLTS U90 ( .A(n84), .B(n458), .C(n516), .D(n397), .Y(n1592) );
  NOR3XLTS U91 ( .A(n17), .B(n179), .C(n268), .Y(n1591) );
  CLKBUFX2TS U92 ( .A(n1487), .Y(n1593) );
  NAND4XLTS U93 ( .A(n273), .B(n515), .C(n397), .D(n393), .Y(n1617) );
  NOR3XLTS U94 ( .A(n218), .B(n17), .C(n268), .Y(n1616) );
  CLKBUFX2TS U95 ( .A(n1422), .Y(n1618) );
  NAND4XLTS U96 ( .A(n1948), .B(n501), .C(n486), .D(n520), .Y(n1581) );
  CLKBUFX2TS U97 ( .A(n1537), .Y(n1582) );
  NAND3XLTS U98 ( .A(n544), .B(n1945), .C(n543), .Y(n565) );
  CLKAND2X2TS U99 ( .A(n529), .B(n527), .Y(n556) );
  INVX2TS U100 ( .A(selectBit_NORTH), .Y(n510) );
  NOR2XLTS U101 ( .A(n1616), .B(n1612), .Y(n278) );
  NOR2XLTS U102 ( .A(n1591), .B(n1588), .Y(n90) );
  NOR2XLTS U103 ( .A(n1580), .B(n1577), .Y(n38) );
  NOR2XLTS U104 ( .A(n1665), .B(n1661), .Y(n402) );
  AO21X1TS U105 ( .A0(n464), .A1(n510), .B0(n21), .Y(n23) );
  NAND3XLTS U106 ( .A(selectBit_NORTH), .B(n513), .C(n512), .Y(n524) );
  NAND3XLTS U107 ( .A(n511), .B(n513), .C(n510), .Y(n523) );
  NOR2XLTS U108 ( .A(n1651), .B(n1647), .Y(n323) );
  NOR2XLTS U109 ( .A(n1625), .B(n1622), .Y(n130) );
  NAND2BXLTS U110 ( .AN(n226), .B(n225), .Y(n227) );
  NAND3XLTS U111 ( .A(n21), .B(n458), .C(n396), .Y(n221) );
  NOR2XLTS U112 ( .A(n1637), .B(n1634), .Y(n182) );
  NAND2BXLTS U113 ( .AN(n39), .B(n38), .Y(n40) );
  XOR2XLTS U114 ( .A(n459), .B(n461), .Y(n479) );
  OAI21XLTS U115 ( .A0(n462), .A1(n1949), .B0(n461), .Y(n463) );
  INVX2TS U116 ( .A(n271), .Y(n392) );
  XOR2X1TS U117 ( .A(n486), .B(n19), .Y(n124) );
  NOR2XLTS U118 ( .A(n86), .B(reset), .Y(n504) );
  NOR3X1TS U119 ( .A(n179), .B(n80), .C(n388), .Y(n1625) );
  INVX2TS U120 ( .A(n1622), .Y(n1620) );
  NAND4XLTS U121 ( .A(n516), .B(n397), .C(n396), .D(n448), .Y(n1666) );
  NOR3XLTS U122 ( .A(n31), .B(n392), .C(n82), .Y(n1657) );
  INVX2TS U123 ( .A(n1657), .Y(n1654) );
  NOR3BXLTS U124 ( .AN(n391), .B(n390), .C(n389), .Y(n1661) );
  NAND4XLTS U125 ( .A(n491), .B(n516), .C(n397), .D(n450), .Y(n1638) );
  NOR3XLTS U126 ( .A(n31), .B(n82), .C(n271), .Y(n1630) );
  INVX2TS U127 ( .A(n1630), .Y(n1629) );
  NOR3XLTS U128 ( .A(n31), .B(n392), .C(n11), .Y(n1644) );
  INVX2TS U129 ( .A(n1644), .Y(n1641) );
  NOR3XLTS U130 ( .A(n316), .B(n315), .C(n390), .Y(n1647) );
  NAND4XLTS U131 ( .A(n453), .B(n458), .C(readReady), .D(n393), .Y(n1605) );
  INVX2TS U132 ( .A(n1595), .Y(n1598) );
  INVX2TS U133 ( .A(n1604), .Y(n1602) );
  INVX2TS U134 ( .A(n1585), .Y(n1584) );
  NOR3XLTS U135 ( .A(n392), .B(n22), .C(n25), .Y(n1609) );
  INVX2TS U136 ( .A(n1609), .Y(n1608) );
  NAND4XLTS U137 ( .A(n218), .B(n123), .C(n124), .D(n466), .Y(n1578) );
  INVX2TS U138 ( .A(n1573), .Y(n1574) );
  INVX2TS U139 ( .A(destinationAddressIn_SOUTH[11]), .Y(n152) );
  INVX2TS U140 ( .A(destinationAddressIn_SOUTH[10]), .Y(n139) );
  INVX2TS U141 ( .A(destinationAddressIn_SOUTH[9]), .Y(n147) );
  INVX2TS U142 ( .A(destinationAddressIn_SOUTH[8]), .Y(n142) );
  CLKAND2X2TS U143 ( .A(n484), .B(n482), .Y(n489) );
  AO22XLTS U144 ( .A0(n1953), .A1(n504), .B0(n503), .B1(n502), .Y(n1969) );
  AO22XLTS U145 ( .A0(n1948), .A1(n504), .B0(n503), .B1(n499), .Y(n1967) );
  AO22XLTS U146 ( .A0(n501), .A1(n504), .B0(n503), .B1(n500), .Y(n1968) );
  OAI21XLTS U147 ( .A0(n86), .A1(n455), .B0(n498), .Y(n1970) );
  NAND4XLTS U148 ( .A(n878), .B(n877), .C(n876), .D(n875), .Y(n1996) );
  NAND4XLTS U149 ( .A(n854), .B(n853), .C(n852), .D(n851), .Y(n1995) );
  NAND4XLTS U150 ( .A(n842), .B(n841), .C(n840), .D(n839), .Y(n1994) );
  NAND4XLTS U151 ( .A(n830), .B(n829), .C(n828), .D(n827), .Y(n1993) );
  NAND4XLTS U152 ( .A(n811), .B(n810), .C(n809), .D(n808), .Y(n1992) );
  NAND4XLTS U153 ( .A(n791), .B(n790), .C(n789), .D(n788), .Y(n1991) );
  NAND4XLTS U154 ( .A(n662), .B(n661), .C(n660), .D(n659), .Y(n1982) );
  NAND4XLTS U155 ( .A(n650), .B(n649), .C(n648), .D(n647), .Y(n1981) );
  NAND4XLTS U156 ( .A(n630), .B(n629), .C(n628), .D(n627), .Y(n1980) );
  NAND4XLTS U157 ( .A(n615), .B(n614), .C(n613), .D(n612), .Y(n1979) );
  NAND4XLTS U158 ( .A(n604), .B(n603), .C(n602), .D(n659), .Y(n1978) );
  NAND4XLTS U159 ( .A(n593), .B(n592), .C(n591), .D(n647), .Y(n1977) );
  NAND4XLTS U160 ( .A(n585), .B(n584), .C(n583), .D(n627), .Y(n1976) );
  NAND4XLTS U161 ( .A(n568), .B(n567), .C(n566), .D(n612), .Y(n1975) );
  NAND4XLTS U162 ( .A(n547), .B(n546), .C(n545), .D(n565), .Y(n1973) );
  NAND3XLTS U163 ( .A(n781), .B(n780), .C(n779), .Y(n1990) );
  NAND3XLTS U164 ( .A(n767), .B(n766), .C(n765), .Y(n1989) );
  NAND3XLTS U165 ( .A(n752), .B(n751), .C(n750), .Y(n1988) );
  NAND3XLTS U166 ( .A(n734), .B(n733), .C(n732), .Y(n1987) );
  NAND3XLTS U167 ( .A(n720), .B(n719), .C(n718), .Y(n1986) );
  NAND3XLTS U168 ( .A(n709), .B(n708), .C(n707), .Y(n1985) );
  NAND3XLTS U169 ( .A(n694), .B(n693), .C(n692), .Y(n1984) );
  NAND3XLTS U170 ( .A(n673), .B(n672), .C(n671), .Y(n1983) );
  NAND3XLTS U171 ( .A(n559), .B(n558), .C(n557), .Y(n1974) );
  NAND3XLTS U172 ( .A(n1347), .B(n1346), .C(n1345), .Y(n2040) );
  NAND3XLTS U173 ( .A(n1341), .B(n1340), .C(n1339), .Y(n2039) );
  NAND3XLTS U174 ( .A(n1112), .B(n1111), .C(n1110), .Y(n2038) );
  NAND3XLTS U175 ( .A(n1106), .B(n1105), .C(n1104), .Y(n2037) );
  NAND3XLTS U176 ( .A(n1098), .B(n1097), .C(n1096), .Y(n2036) );
  NAND3XLTS U177 ( .A(n1092), .B(n1091), .C(n1090), .Y(n2035) );
  NAND3XLTS U178 ( .A(n1818), .B(n1817), .C(n1816), .Y(n2144) );
  NAND3XLTS U179 ( .A(n1809), .B(n1808), .C(n1807), .Y(n2143) );
  NAND3XLTS U180 ( .A(n1803), .B(n1802), .C(n1801), .Y(n2142) );
  NAND3XLTS U181 ( .A(n1795), .B(n1794), .C(n1793), .Y(n2141) );
  NAND3XLTS U182 ( .A(n988), .B(n987), .C(n986), .Y(n2016) );
  NAND3XLTS U183 ( .A(n982), .B(n981), .C(n980), .Y(n2015) );
  NAND3XLTS U184 ( .A(n974), .B(n973), .C(n972), .Y(n2014) );
  NAND3XLTS U185 ( .A(n965), .B(n964), .C(n963), .Y(n2013) );
  NAND3XLTS U186 ( .A(n1441), .B(n1440), .C(n1439), .Y(n2058) );
  NAND3XLTS U187 ( .A(n1435), .B(n1434), .C(n1433), .Y(n2057) );
  NAND3XLTS U188 ( .A(n1431), .B(n1430), .C(n1429), .Y(n2056) );
  NAND3XLTS U189 ( .A(n1427), .B(n1426), .C(n1425), .Y(n2055) );
  NAND3XLTS U190 ( .A(n1420), .B(n1419), .C(n1418), .Y(n2054) );
  NAND3XLTS U191 ( .A(n1413), .B(n1412), .C(n1411), .Y(n2053) );
  NAND3XLTS U192 ( .A(n1469), .B(n1468), .C(n1467), .Y(n2064) );
  NAND3XLTS U193 ( .A(n1465), .B(n1464), .C(n1463), .Y(n2063) );
  NAND3XLTS U194 ( .A(n1461), .B(n1460), .C(n1459), .Y(n2062) );
  NAND3XLTS U195 ( .A(n1457), .B(n1456), .C(n1455), .Y(n2061) );
  NAND3XLTS U196 ( .A(n1452), .B(n1451), .C(n1450), .Y(n2060) );
  NAND3XLTS U197 ( .A(n1447), .B(n1446), .C(n1445), .Y(n2059) );
  NAND3XLTS U198 ( .A(n1726), .B(n1725), .C(n1724), .Y(n2108) );
  NAND3XLTS U199 ( .A(n1718), .B(n1717), .C(n1716), .Y(n2107) );
  NAND3XLTS U200 ( .A(n1710), .B(n1709), .C(n1708), .Y(n2106) );
  NAND3XLTS U201 ( .A(n1701), .B(n1700), .C(n1699), .Y(n2105) );
  NAND3XLTS U202 ( .A(n914), .B(n913), .C(n912), .Y(n2004) );
  NAND3XLTS U203 ( .A(n910), .B(n909), .C(n908), .Y(n2003) );
  NAND3XLTS U204 ( .A(n906), .B(n905), .C(n904), .Y(n2002) );
  NAND3XLTS U205 ( .A(n899), .B(n898), .C(n897), .Y(n2001) );
  NAND3XLTS U206 ( .A(n1696), .B(n1695), .C(n1694), .Y(n2096) );
  NAND3XLTS U207 ( .A(n1688), .B(n1687), .C(n1686), .Y(n2095) );
  NAND3XLTS U208 ( .A(n1680), .B(n1679), .C(n1678), .Y(n2094) );
  NAND3XLTS U209 ( .A(n1673), .B(n1672), .C(n1671), .Y(n2093) );
  NAND3XLTS U210 ( .A(n896), .B(n895), .C(n894), .Y(n2000) );
  NAND3XLTS U211 ( .A(n891), .B(n890), .C(n889), .Y(n1999) );
  NAND3XLTS U212 ( .A(n887), .B(n886), .C(n885), .Y(n1998) );
  NAND3XLTS U213 ( .A(n884), .B(n883), .C(n882), .Y(n1997) );
  NAND3XLTS U214 ( .A(n1927), .B(n1926), .C(n1925), .Y(n2180) );
  NAND3XLTS U215 ( .A(n1918), .B(n1917), .C(n1916), .Y(n2179) );
  NAND3XLTS U216 ( .A(n1906), .B(n1905), .C(n1904), .Y(n2178) );
  NAND3XLTS U217 ( .A(n1896), .B(n1895), .C(n1894), .Y(n2177) );
  NAND3XLTS U218 ( .A(n1061), .B(n1060), .C(n1059), .Y(n2028) );
  NAND3XLTS U219 ( .A(n1054), .B(n1053), .C(n1052), .Y(n2027) );
  NAND3XLTS U220 ( .A(n1049), .B(n1048), .C(n1047), .Y(n2026) );
  NAND3XLTS U221 ( .A(n1043), .B(n1042), .C(n1041), .Y(n2025) );
  NAND3XLTS U222 ( .A(n1888), .B(n1887), .C(n1886), .Y(n2168) );
  NAND3XLTS U223 ( .A(n1878), .B(n1877), .C(n1876), .Y(n2167) );
  NAND3XLTS U224 ( .A(n1865), .B(n1864), .C(n1863), .Y(n2166) );
  NAND3XLTS U225 ( .A(n1854), .B(n1853), .C(n1852), .Y(n2165) );
  NAND3XLTS U226 ( .A(n1036), .B(n1035), .C(n1034), .Y(n2024) );
  NAND3XLTS U227 ( .A(n1027), .B(n1026), .C(n1025), .Y(n2023) );
  NAND3XLTS U228 ( .A(n1019), .B(n1018), .C(n1017), .Y(n2022) );
  NAND3XLTS U229 ( .A(n1012), .B(n1011), .C(n1010), .Y(n2021) );
  NAND3XLTS U230 ( .A(n1380), .B(n1379), .C(n1378), .Y(n2046) );
  NAND3XLTS U231 ( .A(n1375), .B(n1374), .C(n1373), .Y(n2045) );
  NAND3XLTS U232 ( .A(n1371), .B(n1370), .C(n1369), .Y(n2044) );
  NAND3XLTS U233 ( .A(n1366), .B(n1365), .C(n1364), .Y(n2043) );
  NAND3XLTS U234 ( .A(n1357), .B(n1356), .C(n1355), .Y(n2042) );
  NAND3XLTS U235 ( .A(n1351), .B(n1350), .C(n1349), .Y(n2041) );
  NAND3XLTS U236 ( .A(n1408), .B(n1407), .C(n1406), .Y(n2052) );
  NAND3XLTS U237 ( .A(n1403), .B(n1402), .C(n1401), .Y(n2051) );
  NAND3XLTS U238 ( .A(n1397), .B(n1396), .C(n1395), .Y(n2050) );
  NAND3XLTS U239 ( .A(n1394), .B(n1393), .C(n1392), .Y(n2049) );
  NAND3XLTS U240 ( .A(n1389), .B(n1388), .C(n1387), .Y(n2048) );
  NAND3XLTS U241 ( .A(n1384), .B(n1383), .C(n1382), .Y(n2047) );
  NAND3XLTS U242 ( .A(n1789), .B(n1788), .C(n1787), .Y(n2132) );
  NAND3XLTS U243 ( .A(n1782), .B(n1781), .C(n1780), .Y(n2131) );
  NAND3XLTS U244 ( .A(n1774), .B(n1773), .C(n1772), .Y(n2130) );
  NAND3XLTS U245 ( .A(n1765), .B(n1764), .C(n1763), .Y(n2129) );
  NAND3XLTS U246 ( .A(n958), .B(n957), .C(n956), .Y(n2012) );
  NAND3XLTS U247 ( .A(n951), .B(n950), .C(n949), .Y(n2011) );
  NAND3XLTS U248 ( .A(n945), .B(n944), .C(n943), .Y(n2010) );
  NAND3XLTS U249 ( .A(n936), .B(n935), .C(n934), .Y(n2009) );
  NAND3XLTS U250 ( .A(n1760), .B(n1759), .C(n1758), .Y(n2120) );
  NAND3XLTS U251 ( .A(n1753), .B(n1752), .C(n1751), .Y(n2119) );
  NAND3XLTS U252 ( .A(n1742), .B(n1741), .C(n1740), .Y(n2118) );
  NAND3XLTS U253 ( .A(n1732), .B(n1731), .C(n1730), .Y(n2117) );
  NAND3XLTS U254 ( .A(n930), .B(n929), .C(n928), .Y(n2008) );
  NAND3XLTS U255 ( .A(n925), .B(n924), .C(n923), .Y(n2007) );
  NAND3XLTS U256 ( .A(n922), .B(n921), .C(n920), .Y(n2006) );
  NAND3XLTS U257 ( .A(n918), .B(n917), .C(n916), .Y(n2005) );
  NAND3XLTS U258 ( .A(n1519), .B(n1518), .C(n1517), .Y(n2070) );
  NAND3XLTS U259 ( .A(n1510), .B(n1509), .C(n1508), .Y(n2069) );
  NAND3XLTS U260 ( .A(n1503), .B(n1502), .C(n1501), .Y(n2068) );
  NAND3XLTS U261 ( .A(n1495), .B(n1494), .C(n1493), .Y(n2067) );
  NAND3XLTS U262 ( .A(n1485), .B(n1484), .C(n1483), .Y(n2066) );
  NAND3XLTS U263 ( .A(n1477), .B(n1476), .C(n1475), .Y(n2065) );
  NAND3XLTS U264 ( .A(n1571), .B(n1570), .C(n1569), .Y(n2076) );
  NAND3XLTS U265 ( .A(n1562), .B(n1561), .C(n1560), .Y(n2075) );
  NAND3XLTS U266 ( .A(n1552), .B(n1551), .C(n1550), .Y(n2074) );
  NAND3XLTS U267 ( .A(n1544), .B(n1543), .C(n1542), .Y(n2073) );
  NAND3XLTS U268 ( .A(n1536), .B(n1535), .C(n1534), .Y(n2072) );
  NAND3XLTS U269 ( .A(n1528), .B(n1527), .C(n1526), .Y(n2071) );
  NAND3XLTS U270 ( .A(n1087), .B(n1086), .C(n1085), .Y(n2034) );
  NAND3XLTS U271 ( .A(n1083), .B(n1082), .C(n1081), .Y(n2033) );
  NAND3XLTS U272 ( .A(n1079), .B(n1078), .C(n1077), .Y(n2032) );
  NAND3XLTS U273 ( .A(n1076), .B(n1075), .C(n1074), .Y(n2031) );
  NAND3XLTS U274 ( .A(n1070), .B(n1069), .C(n1068), .Y(n2030) );
  NAND3XLTS U275 ( .A(n1065), .B(n1064), .C(n1063), .Y(n2029) );
  NAND3XLTS U276 ( .A(n1845), .B(n1844), .C(n1843), .Y(n2156) );
  NAND3XLTS U277 ( .A(n1838), .B(n1837), .C(n1836), .Y(n2155) );
  NAND3XLTS U278 ( .A(n1829), .B(n1828), .C(n1827), .Y(n2154) );
  NAND3XLTS U279 ( .A(n1822), .B(n1821), .C(n1820), .Y(n2153) );
  NAND3XLTS U280 ( .A(n1005), .B(n1004), .C(n1003), .Y(n2020) );
  NAND3XLTS U281 ( .A(n1000), .B(n999), .C(n998), .Y(n2019) );
  NAND3XLTS U282 ( .A(n995), .B(n994), .C(n993), .Y(n2018) );
  NAND3XLTS U283 ( .A(n991), .B(n990), .C(n989), .Y(n2017) );
  OR2X1TS U284 ( .A(n321), .B(n1013), .Y(n359) );
  NAND2X1TS U285 ( .A(n30), .B(n27), .Y(n28) );
  OR2X1TS U286 ( .A(n1654), .B(n404), .Y(n5) );
  OR2X1TS U287 ( .A(n1584), .B(n93), .Y(n6) );
  OR2X1TS U288 ( .A(n1657), .B(n404), .Y(n7) );
  OR2X1TS U289 ( .A(n1609), .B(n280), .Y(n8) );
  OR2X1TS U290 ( .A(n1585), .B(n93), .Y(n9) );
  OA21XLTS U291 ( .A0(n21), .A1(n84), .B0(n24), .Y(n10) );
  OR2X1TS U292 ( .A(n23), .B(n512), .Y(n11) );
  OR2X1TS U293 ( .A(n447), .B(n1638), .Y(n12) );
  OR2X1TS U294 ( .A(n399), .B(n1044), .Y(n429) );
  NOR3XLTS U295 ( .A(n1665), .B(n1658), .C(n403), .Y(n398) );
  NOR3XLTS U296 ( .A(n1580), .B(n1575), .C(n39), .Y(n34) );
  NOR3XLTS U297 ( .A(n1591), .B(n1586), .C(n91), .Y(n85) );
  NOR3XLTS U298 ( .A(n1616), .B(n1610), .C(n279), .Y(n274) );
  OR2X1TS U299 ( .A(n456), .B(n1605), .Y(n13) );
  OR2X1TS U300 ( .A(n447), .B(n1666), .Y(n14) );
  NOR2XLTS U301 ( .A(n849), .B(n524), .Y(n696) );
  NOR2XLTS U302 ( .A(n849), .B(n523), .Y(n549) );
  INVX2TS U303 ( .A(destinationAddressIn_EAST[11]), .Y(n43) );
  INVX2TS U304 ( .A(destinationAddressIn_EAST[10]), .Y(n53) );
  INVX2TS U305 ( .A(destinationAddressIn_EAST[9]), .Y(n35) );
  INVX2TS U306 ( .A(destinationAddressIn_EAST[8]), .Y(n50) );
  INVX2TS U307 ( .A(writeIn_EAST), .Y(n58) );
  INVX2TS U308 ( .A(destinationAddressIn_EAST[7]), .Y(n72) );
  INVX2TS U309 ( .A(destinationAddressIn_EAST[6]), .Y(n64) );
  INVX2TS U310 ( .A(destinationAddressIn_EAST[5]), .Y(n67) );
  INVX2TS U311 ( .A(destinationAddressIn_EAST[4]), .Y(n75) );
  CLKBUFX2TS U312 ( .A(n1949), .Y(n15) );
  INVX2TS U328 ( .A(n1956), .Y(n501) );
  INVX2TS U329 ( .A(n1952), .Y(n452) );
  INVX2TS U330 ( .A(n17), .Y(n80) );
  INVX2TS U331 ( .A(n80), .Y(n123) );
  INVX2TS U332 ( .A(selectBit_WEST), .Y(n460) );
  INVX2TS U333 ( .A(n1578), .Y(n1580) );
  INVX2TS U334 ( .A(n1948), .Y(n464) );
  INVX2TS U335 ( .A(selectBit_SOUTH), .Y(n512) );
  INVX2TS U336 ( .A(n11), .Y(n219) );
  INVX2TS U337 ( .A(n1956), .Y(n84) );
  INVX2TS U338 ( .A(n1956), .Y(n491) );
  NAND2X1TS U339 ( .A(n20), .B(n491), .Y(n24) );
  INVX2TS U340 ( .A(n10), .Y(n81) );
  NAND2X1TS U341 ( .A(selectBit_SOUTH), .B(n23), .Y(n22) );
  NAND2X1TS U342 ( .A(n315), .B(n269), .Y(n126) );
  INVX2TS U343 ( .A(selectBit_EAST), .Y(n519) );
  INVX2TS U344 ( .A(n519), .Y(n517) );
  INVX2TS U345 ( .A(n1954), .Y(n273) );
  INVX2TS U346 ( .A(n24), .Y(n127) );
  INVX2TS U347 ( .A(n1953), .Y(n457) );
  AOI22X1TS U348 ( .A0(n273), .A1(n24), .B0(n127), .B1(n457), .Y(n25) );
  INVX2TS U349 ( .A(n25), .Y(n26) );
  INVX2TS U350 ( .A(n26), .Y(n27) );
  INVX2TS U351 ( .A(n28), .Y(n122) );
  INVX2TS U352 ( .A(n122), .Y(n29) );
  NAND2X1TS U353 ( .A(n517), .B(n125), .Y(n270) );
  NAND2X1TS U354 ( .A(n273), .B(n127), .Y(n33) );
  INVX2TS U355 ( .A(n27), .Y(n31) );
  INVX2TS U356 ( .A(n512), .Y(n511) );
  INVX2TS U357 ( .A(n460), .Y(n518) );
  INVX2TS U358 ( .A(readReady), .Y(n129) );
  INVX2TS U359 ( .A(n129), .Y(n520) );
  NAND2X1TS U360 ( .A(n544), .B(n513), .Y(n529) );
  INVX2TS U361 ( .A(n220), .Y(n319) );
  INVX2TS U362 ( .A(n319), .Y(n86) );
  INVX2TS U363 ( .A(n86), .Y(n32) );
  AOI31XLTS U364 ( .A0(n38), .A1(n33), .A2(n1573), .B0(n32), .Y(n37) );
  NAND2X1TS U365 ( .A(n37), .B(n1581), .Y(n39) );
  INVX2TS U366 ( .A(n34), .Y(n893) );
  INVX2TS U367 ( .A(n893), .Y(n1683) );
  CLKBUFX2TS U368 ( .A(n1683), .Y(n49) );
  INVX2TS U369 ( .A(n49), .Y(n71) );
  INVX2TS U370 ( .A(destinationAddressIn_EAST[9]), .Y(n240) );
  INVX2TS U371 ( .A(n36), .Y(n892) );
  INVX2TS U372 ( .A(n892), .Y(n1668) );
  INVX2TS U373 ( .A(n1537), .Y(n55) );
  OR2X1TS U374 ( .A(n1578), .B(n39), .Y(n54) );
  INVX2TS U375 ( .A(n54), .Y(n1684) );
  CLKBUFX2TS U376 ( .A(destinationAddressIn_WEST[9]), .Y(n415) );
  CLKBUFX2TS U377 ( .A(n415), .Y(n736) );
  AOI22X1TS U378 ( .A0(n55), .A1(\destinationAddressbuffer[7][9] ), .B0(n44), 
        .B1(n736), .Y(n42) );
  INVX2TS U379 ( .A(n45), .Y(n880) );
  INVX2TS U380 ( .A(n880), .Y(n1677) );
  INVX2TS U381 ( .A(n147), .Y(n737) );
  OR2X1TS U382 ( .A(n1574), .B(n40), .Y(n61) );
  INVX2TS U383 ( .A(n61), .Y(n1524) );
  INVX2TS U384 ( .A(n1524), .Y(n881) );
  INVX2TS U385 ( .A(n881), .Y(n888) );
  CLKBUFX2TS U386 ( .A(destinationAddressIn_NORTH[9]), .Y(n739) );
  CLKBUFX2TS U387 ( .A(n739), .Y(n328) );
  AOI22X1TS U388 ( .A0(n1677), .A1(n737), .B0(n888), .B1(n328), .Y(n41) );
  OAI211XLTS U389 ( .A0(n71), .A1(n240), .B0(n42), .C0(n41), .Y(n2102) );
  INVX2TS U390 ( .A(destinationAddressIn_EAST[11]), .Y(n245) );
  INVX2TS U391 ( .A(n54), .Y(n44) );
  INVX2TS U392 ( .A(n44), .Y(n879) );
  INVX2TS U393 ( .A(n879), .Y(n68) );
  CLKBUFX2TS U394 ( .A(destinationAddressIn_WEST[11]), .Y(n401) );
  CLKBUFX2TS U395 ( .A(n401), .Y(n768) );
  AOI22X1TS U396 ( .A0(n55), .A1(\destinationAddressbuffer[7][11] ), .B0(n68), 
        .B1(n768), .Y(n48) );
  INVX2TS U397 ( .A(n45), .Y(n59) );
  INVX2TS U398 ( .A(n59), .Y(n1559) );
  INVX2TS U399 ( .A(n152), .Y(n771) );
  INVX2TS U400 ( .A(n61), .Y(n46) );
  CLKBUFX2TS U401 ( .A(destinationAddressIn_NORTH[11]), .Y(n772) );
  CLKBUFX2TS U402 ( .A(n772), .Y(n351) );
  AOI22X1TS U403 ( .A0(n1559), .A1(n771), .B0(n46), .B1(n351), .Y(n47) );
  OAI211XLTS U404 ( .A0(n71), .A1(n245), .B0(n48), .C0(n47), .Y(n2104) );
  INVX2TS U405 ( .A(n49), .Y(n79) );
  INVX2TS U406 ( .A(destinationAddressIn_EAST[8]), .Y(n231) );
  INVX2TS U407 ( .A(n54), .Y(n1670) );
  CLKBUFX2TS U408 ( .A(destinationAddressIn_WEST[8]), .Y(n421) );
  CLKBUFX2TS U409 ( .A(n421), .Y(n721) );
  AOI22X1TS U410 ( .A0(n55), .A1(\destinationAddressbuffer[7][8] ), .B0(n1670), 
        .B1(n721), .Y(n52) );
  INVX2TS U411 ( .A(n59), .Y(n1693) );
  INVX2TS U412 ( .A(n142), .Y(n722) );
  CLKBUFX2TS U413 ( .A(destinationAddressIn_NORTH[8]), .Y(n723) );
  CLKBUFX2TS U414 ( .A(n723), .Y(n343) );
  AOI22X1TS U415 ( .A0(n1693), .A1(n722), .B0(n1524), .B1(n343), .Y(n51) );
  OAI211XLTS U416 ( .A0(n79), .A1(n231), .B0(n52), .C0(n51), .Y(n2101) );
  INVX2TS U417 ( .A(destinationAddressIn_EAST[10]), .Y(n235) );
  INVX2TS U418 ( .A(n54), .Y(n1522) );
  CLKBUFX2TS U419 ( .A(destinationAddressIn_WEST[10]), .Y(n409) );
  CLKBUFX2TS U420 ( .A(n409), .Y(n753) );
  AOI22X1TS U421 ( .A0(n55), .A1(\destinationAddressbuffer[7][10] ), .B0(n1522), .B1(n753), .Y(n57) );
  INVX2TS U422 ( .A(n59), .Y(n1685) );
  INVX2TS U423 ( .A(n139), .Y(n756) );
  INVX2TS U424 ( .A(n61), .Y(n1557) );
  CLKBUFX2TS U425 ( .A(destinationAddressIn_NORTH[10]), .Y(n757) );
  CLKBUFX2TS U426 ( .A(n757), .Y(n336) );
  AOI22X1TS U427 ( .A0(n1685), .A1(n756), .B0(n1557), .B1(n336), .Y(n56) );
  OAI211XLTS U428 ( .A0(n71), .A1(n235), .B0(n57), .C0(n56), .Y(n2103) );
  INVX2TS U429 ( .A(n1582), .Y(n1689) );
  AOI22X1TS U430 ( .A0(n1689), .A1(writeOutbuffer[7]), .B0(n1522), .B1(
        writeIn_WEST), .Y(n63) );
  INVX2TS U431 ( .A(n59), .Y(n60) );
  INVX2TS U432 ( .A(writeIn_SOUTH), .Y(n156) );
  INVX2TS U433 ( .A(n156), .Y(n550) );
  INVX2TS U434 ( .A(n61), .Y(n1676) );
  AOI22X1TS U435 ( .A0(n60), .A1(n550), .B0(n1676), .B1(writeIn_NORTH), .Y(n62) );
  OAI211XLTS U436 ( .A0(n79), .A1(n296), .B0(n63), .C0(n62), .Y(n2077) );
  INVX2TS U437 ( .A(destinationAddressIn_EAST[6]), .Y(n259) );
  INVX2TS U438 ( .A(n1537), .Y(n76) );
  AOI22X1TS U439 ( .A0(n76), .A1(\destinationAddressbuffer[7][6] ), .B0(n1684), 
        .B1(destinationAddressIn_WEST[6]), .Y(n66) );
  INVX2TS U440 ( .A(destinationAddressIn_SOUTH[6]), .Y(n162) );
  INVX2TS U441 ( .A(n162), .Y(n697) );
  AOI22X1TS U442 ( .A0(n1685), .A1(n697), .B0(n888), .B1(
        destinationAddressIn_NORTH[6]), .Y(n65) );
  OAI211XLTS U443 ( .A0(n79), .A1(n259), .B0(n66), .C0(n65), .Y(n2099) );
  INVX2TS U444 ( .A(destinationAddressIn_EAST[5]), .Y(n251) );
  AOI22X1TS U445 ( .A0(n76), .A1(\destinationAddressbuffer[7][5] ), .B0(n68), 
        .B1(destinationAddressIn_WEST[5]), .Y(n70) );
  INVX2TS U446 ( .A(destinationAddressIn_SOUTH[5]), .Y(n166) );
  INVX2TS U447 ( .A(n166), .Y(n677) );
  AOI22X1TS U448 ( .A0(n1693), .A1(n677), .B0(n46), .B1(
        destinationAddressIn_NORTH[5]), .Y(n69) );
  OAI211XLTS U449 ( .A0(n71), .A1(n251), .B0(n70), .C0(n69), .Y(n2098) );
  INVX2TS U450 ( .A(destinationAddressIn_EAST[7]), .Y(n254) );
  AOI22X1TS U451 ( .A0(n76), .A1(\destinationAddressbuffer[7][7] ), .B0(n1670), 
        .B1(destinationAddressIn_WEST[7]), .Y(n74) );
  INVX2TS U452 ( .A(destinationAddressIn_SOUTH[7]), .Y(n177) );
  INVX2TS U453 ( .A(n177), .Y(n711) );
  AOI22X1TS U454 ( .A0(n60), .A1(n711), .B0(n1676), .B1(
        destinationAddressIn_NORTH[7]), .Y(n73) );
  OAI211XLTS U455 ( .A0(n893), .A1(n254), .B0(n74), .C0(n73), .Y(n2100) );
  INVX2TS U456 ( .A(destinationAddressIn_EAST[4]), .Y(n266) );
  AOI22X1TS U457 ( .A0(n76), .A1(\destinationAddressbuffer[7][4] ), .B0(n68), 
        .B1(destinationAddressIn_WEST[4]), .Y(n78) );
  INVX2TS U458 ( .A(destinationAddressIn_SOUTH[4]), .Y(n172) );
  INVX2TS U459 ( .A(n172), .Y(n665) );
  AOI22X1TS U460 ( .A0(n1559), .A1(n665), .B0(n1557), .B1(
        destinationAddressIn_NORTH[4]), .Y(n77) );
  OAI211XLTS U461 ( .A0(n79), .A1(n266), .B0(n78), .C0(n77), .Y(n2097) );
  INVX2TS U462 ( .A(n218), .Y(n179) );
  NAND2X1TS U463 ( .A(n124), .B(n518), .Y(n268) );
  AOI21X1TS U464 ( .A0(n219), .A1(n81), .B0(n315), .Y(n391) );
  NOR3XLTS U465 ( .A(n391), .B(n270), .C(n269), .Y(n1588) );
  INVX2TS U466 ( .A(n1956), .Y(n462) );
  INVX2TS U467 ( .A(n1952), .Y(n453) );
  NOR2XLTS U468 ( .A(n453), .B(n510), .Y(n394) );
  INVX2TS U469 ( .A(n10), .Y(n271) );
  NOR3XLTS U470 ( .A(n27), .B(n82), .C(n271), .Y(n1585) );
  AOI31XLTS U471 ( .A0(n273), .A1(n462), .A2(n394), .B0(n1585), .Y(n83) );
  AOI21X1TS U472 ( .A0(n90), .A1(n83), .B0(n275), .Y(n88) );
  INVX2TS U473 ( .A(n129), .Y(n516) );
  INVX2TS U474 ( .A(n1948), .Y(n397) );
  NAND2X1TS U475 ( .A(n88), .B(n1592), .Y(n91) );
  INVX2TS U476 ( .A(n85), .Y(n1471) );
  INVX2TS U477 ( .A(n1471), .Y(n911) );
  CLKBUFX2TS U478 ( .A(n911), .Y(n99) );
  INVX2TS U479 ( .A(n99), .Y(n115) );
  INVX2TS U480 ( .A(n86), .Y(n447) );
  INVX2TS U481 ( .A(n87), .Y(n1486) );
  INVX2TS U482 ( .A(n1486), .Y(n900) );
  INVX2TS U483 ( .A(n1487), .Y(n103) );
  OR2X1TS U484 ( .A(n1589), .B(n91), .Y(n102) );
  INVX2TS U485 ( .A(n102), .Y(n89) );
  AOI22X1TS U486 ( .A0(n103), .A1(\destinationAddressbuffer[6][11] ), .B0(n89), 
        .B1(n768), .Y(n96) );
  INVX2TS U487 ( .A(n9), .Y(n92) );
  INVX2TS U488 ( .A(n92), .Y(n903) );
  INVX2TS U489 ( .A(n903), .Y(n104) );
  CLKBUFX2TS U490 ( .A(n772), .Y(n406) );
  INVX2TS U491 ( .A(n6), .Y(n94) );
  INVX2TS U492 ( .A(n152), .Y(n350) );
  AOI22X1TS U493 ( .A0(n104), .A1(n406), .B0(n94), .B1(n350), .Y(n95) );
  OAI211XLTS U494 ( .A0(n115), .A1(n245), .B0(n96), .C0(n95), .Y(n2116) );
  INVX2TS U495 ( .A(n102), .Y(n1490) );
  INVX2TS U496 ( .A(n1490), .Y(n901) );
  INVX2TS U497 ( .A(n901), .Y(n112) );
  AOI22X1TS U498 ( .A0(n103), .A1(\destinationAddressbuffer[6][9] ), .B0(n112), 
        .B1(n736), .Y(n98) );
  INVX2TS U499 ( .A(n903), .Y(n907) );
  CLKBUFX2TS U500 ( .A(n739), .Y(n417) );
  INVX2TS U501 ( .A(n6), .Y(n1706) );
  INVX2TS U502 ( .A(n147), .Y(n327) );
  AOI22X1TS U503 ( .A0(n907), .A1(n417), .B0(n1706), .B1(n327), .Y(n97) );
  OAI211XLTS U504 ( .A0(n115), .A1(n240), .B0(n98), .C0(n97), .Y(n2114) );
  INVX2TS U505 ( .A(n99), .Y(n121) );
  AOI22X1TS U506 ( .A0(n103), .A1(\destinationAddressbuffer[6][8] ), .B0(n109), 
        .B1(n721), .Y(n101) );
  INVX2TS U507 ( .A(n9), .Y(n1698) );
  CLKBUFX2TS U508 ( .A(n723), .Y(n423) );
  INVX2TS U509 ( .A(n6), .Y(n1515) );
  INVX2TS U510 ( .A(n142), .Y(n342) );
  AOI22X1TS U511 ( .A0(n1698), .A1(n423), .B0(n1515), .B1(n342), .Y(n100) );
  OAI211XLTS U512 ( .A0(n121), .A1(n231), .B0(n101), .C0(n100), .Y(n2113) );
  INVX2TS U513 ( .A(n102), .Y(n1704) );
  AOI22X1TS U514 ( .A0(n103), .A1(\destinationAddressbuffer[6][10] ), .B0(
        n1704), .B1(n753), .Y(n106) );
  CLKBUFX2TS U515 ( .A(n757), .Y(n410) );
  INVX2TS U516 ( .A(n6), .Y(n1723) );
  INVX2TS U517 ( .A(n1723), .Y(n902) );
  INVX2TS U518 ( .A(n139), .Y(n334) );
  AOI22X1TS U519 ( .A0(n104), .A1(n410), .B0(n1714), .B1(n334), .Y(n105) );
  OAI211XLTS U520 ( .A0(n115), .A1(n235), .B0(n106), .C0(n105), .Y(n2115) );
  INVX2TS U521 ( .A(n1593), .Y(n1719) );
  AOI22X1TS U522 ( .A0(n1719), .A1(writeOutbuffer[6]), .B0(n1704), .B1(
        writeIn_WEST), .Y(n108) );
  INVX2TS U523 ( .A(n9), .Y(n1715) );
  CLKBUFX2TS U524 ( .A(writeIn_NORTH), .Y(n356) );
  CLKBUFX2TS U525 ( .A(n356), .Y(n426) );
  INVX2TS U526 ( .A(n156), .Y(n355) );
  AOI22X1TS U527 ( .A0(n1715), .A1(n426), .B0(n1515), .B1(n355), .Y(n107) );
  OAI211XLTS U528 ( .A0(n121), .A1(n296), .B0(n108), .C0(n107), .Y(n2078) );
  INVX2TS U529 ( .A(n1593), .Y(n118) );
  INVX2TS U530 ( .A(n901), .Y(n109) );
  AOI22X1TS U531 ( .A0(n118), .A1(\destinationAddressbuffer[6][4] ), .B0(n109), 
        .B1(destinationAddressIn_WEST[4]), .Y(n111) );
  CLKBUFX2TS U532 ( .A(destinationAddressIn_NORTH[4]), .Y(n363) );
  CLKBUFX2TS U533 ( .A(n363), .Y(n443) );
  INVX2TS U534 ( .A(n172), .Y(n362) );
  AOI22X1TS U535 ( .A0(n1698), .A1(n443), .B0(n1706), .B1(n362), .Y(n110) );
  OAI211XLTS U536 ( .A0(n121), .A1(n266), .B0(n111), .C0(n110), .Y(n2109) );
  AOI22X1TS U537 ( .A0(n118), .A1(\destinationAddressbuffer[6][6] ), .B0(n112), 
        .B1(destinationAddressIn_WEST[6]), .Y(n114) );
  CLKBUFX2TS U538 ( .A(destinationAddressIn_NORTH[6]), .Y(n370) );
  CLKBUFX2TS U539 ( .A(n370), .Y(n433) );
  INVX2TS U540 ( .A(n162), .Y(n368) );
  AOI22X1TS U541 ( .A0(n907), .A1(n433), .B0(n94), .B1(n368), .Y(n113) );
  OAI211XLTS U542 ( .A0(n115), .A1(n259), .B0(n114), .C0(n113), .Y(n2111) );
  AOI22X1TS U543 ( .A0(n118), .A1(\destinationAddressbuffer[6][7] ), .B0(n112), 
        .B1(destinationAddressIn_WEST[7]), .Y(n117) );
  INVX2TS U544 ( .A(n9), .Y(n1707) );
  CLKBUFX2TS U545 ( .A(destinationAddressIn_NORTH[7]), .Y(n377) );
  CLKBUFX2TS U546 ( .A(n377), .Y(n430) );
  INVX2TS U547 ( .A(n177), .Y(n376) );
  AOI22X1TS U548 ( .A0(n1707), .A1(n430), .B0(n1723), .B1(n376), .Y(n116) );
  OAI211XLTS U549 ( .A0(n1471), .A1(n254), .B0(n117), .C0(n116), .Y(n2112) );
  AOI22X1TS U550 ( .A0(n118), .A1(\destinationAddressbuffer[6][5] ), .B0(n89), 
        .B1(destinationAddressIn_WEST[5]), .Y(n120) );
  CLKBUFX2TS U551 ( .A(destinationAddressIn_NORTH[5]), .Y(n384) );
  CLKBUFX2TS U552 ( .A(n384), .Y(n438) );
  INVX2TS U553 ( .A(n902), .Y(n1499) );
  INVX2TS U554 ( .A(n166), .Y(n383) );
  AOI22X1TS U555 ( .A0(n1707), .A1(n438), .B0(n1499), .B1(n383), .Y(n119) );
  OAI211XLTS U556 ( .A0(n121), .A1(n251), .B0(n120), .C0(n119), .Y(n2110) );
  INVX2TS U557 ( .A(n1953), .Y(n450) );
  NAND2X1TS U558 ( .A(n127), .B(n450), .Y(n128) );
  INVX2TS U559 ( .A(n220), .Y(n456) );
  AOI31XLTS U560 ( .A0(n130), .A1(n29), .A2(n128), .B0(n456), .Y(n133) );
  INVX2TS U561 ( .A(n129), .Y(n515) );
  INVX2TS U562 ( .A(n1953), .Y(n448) );
  INVX2TS U563 ( .A(n131), .Y(n977) );
  INVX2TS U564 ( .A(n977), .Y(n1386) );
  CLKBUFX2TS U565 ( .A(n1386), .Y(n143) );
  INVX2TS U566 ( .A(n143), .Y(n167) );
  INVX2TS U567 ( .A(n132), .Y(n1390) );
  INVX2TS U568 ( .A(n1390), .Y(n967) );
  INVX2TS U569 ( .A(n1627), .Y(n148) );
  NOR3XLTS U570 ( .A(n1625), .B(n1620), .C(n135), .Y(n144) );
  INVX2TS U571 ( .A(n144), .Y(n168) );
  INVX2TS U572 ( .A(n168), .Y(n1381) );
  AOI22X1TS U573 ( .A0(n148), .A1(\destinationAddressbuffer[3][10] ), .B0(
        n1381), .B1(destinationAddressIn_EAST[10]), .Y(n138) );
  OR2X1TS U574 ( .A(n122), .B(n134), .Y(n158) );
  INVX2TS U575 ( .A(n158), .Y(n1800) );
  INVX2TS U576 ( .A(n136), .Y(n153) );
  INVX2TS U577 ( .A(n153), .Y(n1792) );
  CLKBUFX2TS U578 ( .A(n409), .Y(n331) );
  AOI22X1TS U579 ( .A0(n1800), .A1(n336), .B0(n1792), .B1(n331), .Y(n137) );
  OAI211XLTS U580 ( .A0(n167), .A1(n139), .B0(n138), .C0(n137), .Y(n2151) );
  AOI22X1TS U581 ( .A0(n148), .A1(\destinationAddressbuffer[3][8] ), .B0(n1381), .B1(destinationAddressIn_EAST[8]), .Y(n141) );
  INVX2TS U582 ( .A(n158), .Y(n1806) );
  INVX2TS U583 ( .A(n153), .Y(n1399) );
  CLKBUFX2TS U584 ( .A(n421), .Y(n341) );
  AOI22X1TS U585 ( .A0(n1806), .A1(n343), .B0(n1399), .B1(n341), .Y(n140) );
  OAI211XLTS U586 ( .A0(n977), .A1(n142), .B0(n141), .C0(n140), .Y(n2149) );
  INVX2TS U587 ( .A(n143), .Y(n178) );
  INVX2TS U588 ( .A(n144), .Y(n968) );
  INVX2TS U589 ( .A(n968), .Y(n157) );
  AOI22X1TS U590 ( .A0(n148), .A1(\destinationAddressbuffer[3][9] ), .B0(n157), 
        .B1(destinationAddressIn_EAST[9]), .Y(n146) );
  INVX2TS U591 ( .A(n158), .Y(n1400) );
  INVX2TS U592 ( .A(n970), .Y(n978) );
  CLKBUFX2TS U593 ( .A(n415), .Y(n322) );
  AOI22X1TS U594 ( .A0(n978), .A1(n328), .B0(n1399), .B1(n322), .Y(n145) );
  OAI211XLTS U595 ( .A0(n178), .A1(n147), .B0(n146), .C0(n145), .Y(n2150) );
  INVX2TS U596 ( .A(n168), .Y(n1797) );
  AOI22X1TS U597 ( .A0(n148), .A1(\destinationAddressbuffer[3][11] ), .B0(
        n1797), .B1(destinationAddressIn_EAST[11]), .Y(n151) );
  INVX2TS U598 ( .A(n153), .Y(n149) );
  INVX2TS U599 ( .A(n149), .Y(n960) );
  INVX2TS U600 ( .A(n960), .Y(n163) );
  CLKBUFX2TS U601 ( .A(n401), .Y(n347) );
  AOI22X1TS U602 ( .A0(n1400), .A1(n351), .B0(n163), .B1(n347), .Y(n150) );
  OAI211XLTS U603 ( .A0(n167), .A1(n152), .B0(n151), .C0(n150), .Y(n2152) );
  INVX2TS U604 ( .A(n1627), .Y(n1810) );
  INVX2TS U605 ( .A(n168), .Y(n1398) );
  AOI22X1TS U606 ( .A0(n1810), .A1(writeOutbuffer[3]), .B0(n1398), .B1(
        writeIn_EAST), .Y(n155) );
  INVX2TS U607 ( .A(n153), .Y(n1814) );
  CLKBUFX2TS U608 ( .A(writeIn_WEST), .Y(n548) );
  CLKBUFX2TS U609 ( .A(n548), .Y(n354) );
  AOI22X1TS U610 ( .A0(n1800), .A1(n356), .B0(n1814), .B1(n354), .Y(n154) );
  OAI211XLTS U611 ( .A0(n167), .A1(n156), .B0(n155), .C0(n154), .Y(n2081) );
  INVX2TS U612 ( .A(n1391), .Y(n173) );
  AOI22X1TS U613 ( .A0(n173), .A1(\destinationAddressbuffer[3][6] ), .B0(n157), 
        .B1(destinationAddressIn_EAST[6]), .Y(n161) );
  INVX2TS U614 ( .A(n158), .Y(n159) );
  INVX2TS U615 ( .A(n159), .Y(n970) );
  INVX2TS U616 ( .A(n970), .Y(n174) );
  CLKBUFX2TS U617 ( .A(destinationAddressIn_WEST[6]), .Y(n695) );
  CLKBUFX2TS U618 ( .A(n695), .Y(n366) );
  AOI22X1TS U619 ( .A0(n174), .A1(n370), .B0(n1792), .B1(n366), .Y(n160) );
  OAI211XLTS U620 ( .A0(n178), .A1(n162), .B0(n161), .C0(n160), .Y(n2147) );
  AOI22X1TS U621 ( .A0(n173), .A1(\destinationAddressbuffer[3][5] ), .B0(n1797), .B1(destinationAddressIn_EAST[5]), .Y(n165) );
  CLKBUFX2TS U622 ( .A(destinationAddressIn_WEST[5]), .Y(n676) );
  CLKBUFX2TS U623 ( .A(n676), .Y(n381) );
  AOI22X1TS U624 ( .A0(n978), .A1(n384), .B0(n163), .B1(n381), .Y(n164) );
  OAI211XLTS U625 ( .A0(n167), .A1(n166), .B0(n165), .C0(n164), .Y(n2146) );
  INVX2TS U626 ( .A(n168), .Y(n169) );
  AOI22X1TS U627 ( .A0(n173), .A1(\destinationAddressbuffer[3][4] ), .B0(n157), 
        .B1(destinationAddressIn_EAST[4]), .Y(n171) );
  CLKBUFX2TS U628 ( .A(destinationAddressIn_WEST[4]), .Y(n663) );
  CLKBUFX2TS U629 ( .A(n663), .Y(n360) );
  AOI22X1TS U630 ( .A0(n1400), .A1(n363), .B0(n149), .B1(n360), .Y(n170) );
  OAI211XLTS U631 ( .A0(n178), .A1(n172), .B0(n171), .C0(n170), .Y(n2145) );
  AOI22X1TS U632 ( .A0(n173), .A1(\destinationAddressbuffer[3][7] ), .B0(n1398), .B1(destinationAddressIn_EAST[7]), .Y(n176) );
  CLKBUFX2TS U633 ( .A(destinationAddressIn_WEST[7]), .Y(n710) );
  CLKBUFX2TS U634 ( .A(n710), .Y(n374) );
  AOI22X1TS U635 ( .A0(n174), .A1(n377), .B0(n1814), .B1(n374), .Y(n175) );
  OAI211XLTS U636 ( .A0(n178), .A1(n177), .B0(n176), .C0(n175), .Y(n2148) );
  INVX2TS U637 ( .A(n269), .Y(n316) );
  INVX2TS U638 ( .A(n316), .Y(n389) );
  NOR3XLTS U639 ( .A(n391), .B(n389), .C(n390), .Y(n1634) );
  AOI31XLTS U640 ( .A0(n501), .A1(n394), .A2(n457), .B0(n1630), .Y(n180) );
  AOI21X1TS U641 ( .A0(n182), .A1(n180), .B0(n447), .Y(n181) );
  NAND2X1TS U642 ( .A(n181), .B(n1638), .Y(n183) );
  INVX2TS U643 ( .A(n1), .Y(n1359) );
  INVX2TS U644 ( .A(n1359), .Y(n1002) );
  CLKBUFX2TS U645 ( .A(n1002), .Y(n193) );
  INVX2TS U646 ( .A(n193), .Y(n209) );
  INVX2TS U647 ( .A(n12), .Y(n992) );
  INVX2TS U648 ( .A(n1358), .Y(n198) );
  OR2X1TS U649 ( .A(n1635), .B(n183), .Y(n197) );
  INVX2TS U650 ( .A(n197), .Y(n1825) );
  AOI22X1TS U651 ( .A0(n198), .A1(\destinationAddressbuffer[2][10] ), .B0(
        n1825), .B1(n331), .Y(n189) );
  INVX2TS U652 ( .A(n194), .Y(n204) );
  INVX2TS U653 ( .A(n204), .Y(n184) );
  INVX2TS U654 ( .A(n186), .Y(n199) );
  INVX2TS U655 ( .A(n199), .Y(n1841) );
  INVX2TS U656 ( .A(n199), .Y(n187) );
  AOI22X1TS U657 ( .A0(n184), .A1(n336), .B0(n187), .B1(n334), .Y(n188) );
  OAI211XLTS U658 ( .A0(n209), .A1(n235), .B0(n189), .C0(n188), .Y(n2163) );
  INVX2TS U659 ( .A(n197), .Y(n190) );
  INVX2TS U660 ( .A(n190), .Y(n1001) );
  INVX2TS U661 ( .A(n1001), .Y(n213) );
  AOI22X1TS U662 ( .A0(n198), .A1(\destinationAddressbuffer[2][8] ), .B0(n213), 
        .B1(n341), .Y(n192) );
  INVX2TS U663 ( .A(n204), .Y(n1363) );
  AOI22X1TS U664 ( .A0(n1363), .A1(n343), .B0(n186), .B1(n342), .Y(n191) );
  OAI211XLTS U665 ( .A0(n209), .A1(n231), .B0(n192), .C0(n191), .Y(n2161) );
  INVX2TS U666 ( .A(n193), .Y(n217) );
  INVX2TS U667 ( .A(n197), .Y(n1819) );
  AOI22X1TS U668 ( .A0(n198), .A1(\destinationAddressbuffer[2][9] ), .B0(n1819), .B1(n322), .Y(n196) );
  INVX2TS U669 ( .A(n194), .Y(n1354) );
  INVX2TS U670 ( .A(n1354), .Y(n997) );
  AOI22X1TS U671 ( .A0(n997), .A1(n328), .B0(n210), .B1(n327), .Y(n195) );
  OAI211XLTS U672 ( .A0(n217), .A1(n240), .B0(n196), .C0(n195), .Y(n2162) );
  INVX2TS U673 ( .A(n197), .Y(n1833) );
  AOI22X1TS U674 ( .A0(n198), .A1(\destinationAddressbuffer[2][11] ), .B0(
        n1833), .B1(n347), .Y(n201) );
  INVX2TS U675 ( .A(n186), .Y(n996) );
  INVX2TS U676 ( .A(n996), .Y(n210) );
  AOI22X1TS U677 ( .A0(n184), .A1(n351), .B0(n210), .B1(n350), .Y(n200) );
  OAI211XLTS U678 ( .A0(n209), .A1(n245), .B0(n201), .C0(n200), .Y(n2164) );
  INVX2TS U679 ( .A(n1639), .Y(n1839) );
  AOI22X1TS U680 ( .A0(n1839), .A1(writeOutbuffer[2]), .B0(n213), .B1(n354), 
        .Y(n203) );
  INVX2TS U681 ( .A(n204), .Y(n1826) );
  AOI22X1TS U682 ( .A0(n1826), .A1(writeIn_NORTH), .B0(n186), .B1(n355), .Y(
        n202) );
  OAI211XLTS U683 ( .A0(n217), .A1(n296), .B0(n203), .C0(n202), .Y(n2082) );
  INVX2TS U684 ( .A(n1358), .Y(n214) );
  AOI22X1TS U685 ( .A0(n214), .A1(\destinationAddressbuffer[2][7] ), .B0(n1833), .B1(n374), .Y(n206) );
  INVX2TS U686 ( .A(n204), .Y(n1835) );
  AOI22X1TS U687 ( .A0(n1835), .A1(destinationAddressIn_NORTH[7]), .B0(n1841), 
        .B1(n376), .Y(n205) );
  OAI211XLTS U688 ( .A0(n217), .A1(n254), .B0(n206), .C0(n205), .Y(n2160) );
  AOI22X1TS U689 ( .A0(n214), .A1(\destinationAddressbuffer[2][5] ), .B0(n1825), .B1(n381), .Y(n208) );
  INVX2TS U690 ( .A(n996), .Y(n1368) );
  AOI22X1TS U691 ( .A0(n1835), .A1(destinationAddressIn_NORTH[5]), .B0(n1368), 
        .B1(n383), .Y(n207) );
  OAI211XLTS U692 ( .A0(n209), .A1(n251), .B0(n208), .C0(n207), .Y(n2158) );
  AOI22X1TS U693 ( .A0(n214), .A1(\destinationAddressbuffer[2][6] ), .B0(n190), 
        .B1(n366), .Y(n212) );
  AOI22X1TS U694 ( .A0(n997), .A1(destinationAddressIn_NORTH[6]), .B0(n210), 
        .B1(n368), .Y(n211) );
  OAI211XLTS U695 ( .A0(n1359), .A1(n259), .B0(n212), .C0(n211), .Y(n2159) );
  AOI22X1TS U696 ( .A0(n214), .A1(\destinationAddressbuffer[2][4] ), .B0(n213), 
        .B1(n360), .Y(n216) );
  AOI22X1TS U697 ( .A0(n1363), .A1(destinationAddressIn_NORTH[4]), .B0(n1362), 
        .B1(n362), .Y(n215) );
  OAI211XLTS U698 ( .A0(n217), .A1(n266), .B0(n216), .C0(n215), .Y(n2157) );
  INVX2TS U699 ( .A(n1951), .Y(n396) );
  INVX2TS U700 ( .A(n220), .Y(n275) );
  AOI31XLTS U701 ( .A0(n225), .A1(n1595), .A2(n221), .B0(n275), .Y(n223) );
  INVX2TS U702 ( .A(n1951), .Y(n393) );
  NAND2X1TS U703 ( .A(n223), .B(n1605), .Y(n226) );
  INVX2TS U704 ( .A(n222), .Y(n1442) );
  INVX2TS U705 ( .A(n1442), .Y(n927) );
  CLKBUFX2TS U706 ( .A(n927), .Y(n236) );
  INVX2TS U707 ( .A(n236), .Y(n255) );
  INVX2TS U708 ( .A(n13), .Y(n919) );
  INVX2TS U709 ( .A(n1453), .Y(n242) );
  OR2X1TS U710 ( .A(n1602), .B(n226), .Y(n241) );
  INVX2TS U711 ( .A(n241), .Y(n224) );
  INVX2TS U712 ( .A(n224), .Y(n926) );
  INVX2TS U713 ( .A(n926), .Y(n260) );
  AOI22X1TS U714 ( .A0(n242), .A1(\destinationAddressbuffer[5][8] ), .B0(n260), 
        .B1(n721), .Y(n230) );
  INVX2TS U715 ( .A(n237), .Y(n262) );
  INVX2TS U716 ( .A(n262), .Y(n1449) );
  OR2X1TS U717 ( .A(n1595), .B(n227), .Y(n248) );
  INVX2TS U718 ( .A(n248), .Y(n228) );
  INVX2TS U719 ( .A(n228), .Y(n915) );
  INVX2TS U720 ( .A(n915), .Y(n263) );
  AOI22X1TS U721 ( .A0(n1449), .A1(n423), .B0(n263), .B1(n342), .Y(n229) );
  OAI211XLTS U722 ( .A0(n255), .A1(n231), .B0(n230), .C0(n229), .Y(n2125) );
  INVX2TS U723 ( .A(n241), .Y(n1458) );
  AOI22X1TS U724 ( .A0(n242), .A1(\destinationAddressbuffer[5][10] ), .B0(
        n1458), .B1(n753), .Y(n234) );
  INVX2TS U725 ( .A(n262), .Y(n232) );
  INVX2TS U726 ( .A(n248), .Y(n1462) );
  AOI22X1TS U727 ( .A0(n232), .A1(n410), .B0(n1462), .B1(n334), .Y(n233) );
  OAI211XLTS U728 ( .A0(n255), .A1(n235), .B0(n234), .C0(n233), .Y(n2127) );
  INVX2TS U729 ( .A(n236), .Y(n267) );
  INVX2TS U730 ( .A(n241), .Y(n1454) );
  AOI22X1TS U731 ( .A0(n242), .A1(\destinationAddressbuffer[5][9] ), .B0(n1454), .B1(n736), .Y(n239) );
  INVX2TS U732 ( .A(n237), .Y(n1443) );
  INVX2TS U733 ( .A(n1443), .Y(n256) );
  INVX2TS U734 ( .A(n248), .Y(n1749) );
  AOI22X1TS U735 ( .A0(n256), .A1(n417), .B0(n1749), .B1(n327), .Y(n238) );
  OAI211XLTS U736 ( .A0(n267), .A1(n240), .B0(n239), .C0(n238), .Y(n2126) );
  INVX2TS U737 ( .A(n241), .Y(n1737) );
  AOI22X1TS U738 ( .A0(n242), .A1(\destinationAddressbuffer[5][11] ), .B0(
        n1737), .B1(n768), .Y(n244) );
  AOI22X1TS U739 ( .A0(n1449), .A1(n406), .B0(n1462), .B1(n350), .Y(n243) );
  OAI211XLTS U740 ( .A0(n255), .A1(n245), .B0(n244), .C0(n243), .Y(n2128) );
  INVX2TS U741 ( .A(n1606), .Y(n1754) );
  AOI22X1TS U742 ( .A0(n1754), .A1(writeOutbuffer[5]), .B0(n260), .B1(n548), 
        .Y(n247) );
  AOI22X1TS U743 ( .A0(n256), .A1(n426), .B0(n263), .B1(n355), .Y(n246) );
  OAI211XLTS U744 ( .A0(n267), .A1(n296), .B0(n247), .C0(n246), .Y(n2079) );
  INVX2TS U745 ( .A(n1606), .Y(n261) );
  AOI22X1TS U746 ( .A0(n261), .A1(\destinationAddressbuffer[5][5] ), .B0(n1458), .B1(n676), .Y(n250) );
  INVX2TS U747 ( .A(n248), .Y(n1444) );
  AOI22X1TS U748 ( .A0(n232), .A1(n438), .B0(n1444), .B1(n383), .Y(n249) );
  OAI211XLTS U749 ( .A0(n267), .A1(n251), .B0(n250), .C0(n249), .Y(n2122) );
  AOI22X1TS U750 ( .A0(n261), .A1(\destinationAddressbuffer[5][7] ), .B0(n1737), .B1(n710), .Y(n253) );
  INVX2TS U751 ( .A(n262), .Y(n1729) );
  AOI22X1TS U752 ( .A0(n1729), .A1(n430), .B0(n1444), .B1(n376), .Y(n252) );
  OAI211XLTS U753 ( .A0(n255), .A1(n254), .B0(n253), .C0(n252), .Y(n2124) );
  AOI22X1TS U754 ( .A0(n261), .A1(\destinationAddressbuffer[5][6] ), .B0(n224), 
        .B1(n695), .Y(n258) );
  AOI22X1TS U755 ( .A0(n256), .A1(n433), .B0(n228), .B1(n368), .Y(n257) );
  OAI211XLTS U756 ( .A0(n1442), .A1(n259), .B0(n258), .C0(n257), .Y(n2123) );
  AOI22X1TS U757 ( .A0(n261), .A1(\destinationAddressbuffer[5][4] ), .B0(n260), 
        .B1(n663), .Y(n265) );
  INVX2TS U758 ( .A(n262), .Y(n1750) );
  AOI22X1TS U759 ( .A0(n1750), .A1(n443), .B0(n263), .B1(n362), .Y(n264) );
  OAI211XLTS U760 ( .A0(n267), .A1(n266), .B0(n265), .C0(n264), .Y(n2121) );
  AOI31XLTS U761 ( .A0(n486), .A1(n394), .A2(n396), .B0(n1609), .Y(n272) );
  AOI21X1TS U762 ( .A0(n278), .A1(n272), .B0(n275), .Y(n277) );
  NAND2X1TS U763 ( .A(n277), .B(n1617), .Y(n279) );
  INVX2TS U764 ( .A(n274), .Y(n1409) );
  INVX2TS U765 ( .A(n1409), .Y(n952) );
  CLKBUFX2TS U766 ( .A(n952), .Y(n287) );
  INVX2TS U767 ( .A(n287), .Y(n307) );
  INVX2TS U768 ( .A(n276), .Y(n1421) );
  INVX2TS U769 ( .A(n1421), .Y(n937) );
  INVX2TS U770 ( .A(n1422), .Y(n292) );
  OR2X1TS U771 ( .A(n1613), .B(n279), .Y(n291) );
  INVX2TS U772 ( .A(n291), .Y(n1779) );
  AOI22X1TS U773 ( .A0(n292), .A1(\destinationAddressbuffer[4][11] ), .B0(
        n1779), .B1(n347), .Y(n283) );
  INVX2TS U774 ( .A(n293), .Y(n304) );
  INVX2TS U775 ( .A(n304), .Y(n1424) );
  INVX2TS U776 ( .A(n8), .Y(n281) );
  AOI22X1TS U777 ( .A0(n1424), .A1(n771), .B0(n281), .B1(n406), .Y(n282) );
  OAI211XLTS U778 ( .A0(n307), .A1(n43), .B0(n283), .C0(n282), .Y(n2140) );
  INVX2TS U779 ( .A(n291), .Y(n1761) );
  INVX2TS U780 ( .A(n1761), .Y(n938) );
  INVX2TS U781 ( .A(n938), .Y(n303) );
  AOI22X1TS U782 ( .A0(n292), .A1(\destinationAddressbuffer[4][9] ), .B0(n303), 
        .B1(n322), .Y(n286) );
  INVX2TS U783 ( .A(n304), .Y(n284) );
  INVX2TS U784 ( .A(n8), .Y(n1762) );
  INVX2TS U785 ( .A(n1762), .Y(n1417) );
  INVX2TS U786 ( .A(n1417), .Y(n941) );
  AOI22X1TS U787 ( .A0(n1771), .A1(n737), .B0(n941), .B1(n417), .Y(n285) );
  OAI211XLTS U788 ( .A0(n307), .A1(n35), .B0(n286), .C0(n285), .Y(n2138) );
  INVX2TS U789 ( .A(n287), .Y(n314) );
  INVX2TS U790 ( .A(n291), .Y(n288) );
  AOI22X1TS U791 ( .A0(n292), .A1(\destinationAddressbuffer[4][8] ), .B0(n288), 
        .B1(n341), .Y(n290) );
  INVX2TS U792 ( .A(n304), .Y(n1786) );
  AOI22X1TS U793 ( .A0(n1786), .A1(n722), .B0(n300), .B1(n423), .Y(n289) );
  OAI211XLTS U794 ( .A0(n314), .A1(n50), .B0(n290), .C0(n289), .Y(n2137) );
  INVX2TS U795 ( .A(n291), .Y(n1769) );
  AOI22X1TS U796 ( .A0(n292), .A1(\destinationAddressbuffer[4][10] ), .B0(
        n1769), .B1(n331), .Y(n295) );
  INVX2TS U797 ( .A(n293), .Y(n1416) );
  INVX2TS U798 ( .A(n1416), .Y(n311) );
  AOI22X1TS U799 ( .A0(n311), .A1(n756), .B0(n281), .B1(n410), .Y(n294) );
  OAI211XLTS U800 ( .A0(n307), .A1(n53), .B0(n295), .C0(n294), .Y(n2139) );
  INVX2TS U801 ( .A(n1618), .Y(n1783) );
  INVX2TS U802 ( .A(n938), .Y(n297) );
  AOI22X1TS U803 ( .A0(n1783), .A1(writeOutbuffer[4]), .B0(n297), .B1(n354), 
        .Y(n299) );
  INVX2TS U804 ( .A(n8), .Y(n1770) );
  AOI22X1TS U805 ( .A0(n1786), .A1(n550), .B0(n1770), .B1(n426), .Y(n298) );
  OAI211XLTS U806 ( .A0(n314), .A1(n58), .B0(n299), .C0(n298), .Y(n2080) );
  INVX2TS U807 ( .A(n1618), .Y(n310) );
  AOI22X1TS U808 ( .A0(n310), .A1(\destinationAddressbuffer[4][5] ), .B0(n1769), .B1(n381), .Y(n302) );
  INVX2TS U809 ( .A(n1417), .Y(n300) );
  AOI22X1TS U810 ( .A0(n311), .A1(n677), .B0(n300), .B1(n438), .Y(n301) );
  OAI211XLTS U811 ( .A0(n314), .A1(n67), .B0(n302), .C0(n301), .Y(n2134) );
  AOI22X1TS U812 ( .A0(n310), .A1(\destinationAddressbuffer[4][6] ), .B0(n303), 
        .B1(n366), .Y(n306) );
  INVX2TS U813 ( .A(n304), .Y(n1438) );
  AOI22X1TS U814 ( .A0(n1438), .A1(n697), .B0(n941), .B1(n433), .Y(n305) );
  OAI211XLTS U815 ( .A0(n307), .A1(n64), .B0(n306), .C0(n305), .Y(n2135) );
  AOI22X1TS U816 ( .A0(n310), .A1(\destinationAddressbuffer[4][7] ), .B0(n1779), .B1(n374), .Y(n309) );
  AOI22X1TS U817 ( .A0(n311), .A1(n711), .B0(n1770), .B1(n430), .Y(n308) );
  OAI211XLTS U818 ( .A0(n1409), .A1(n72), .B0(n309), .C0(n308), .Y(n2136) );
  AOI22X1TS U819 ( .A0(n310), .A1(\destinationAddressbuffer[4][4] ), .B0(n288), 
        .B1(n360), .Y(n313) );
  AOI22X1TS U820 ( .A0(n311), .A1(n665), .B0(n941), .B1(n443), .Y(n312) );
  OAI211XLTS U821 ( .A0(n314), .A1(n75), .B0(n313), .C0(n312), .Y(n2133) );
  AOI31XLTS U822 ( .A0(n21), .A1(n393), .A2(n457), .B0(n1644), .Y(n317) );
  AOI21X1TS U823 ( .A0(n323), .A1(n317), .B0(n319), .Y(n321) );
  NAND2X1TS U824 ( .A(n321), .B(n1652), .Y(n324) );
  INVX2TS U825 ( .A(n4), .Y(n1029) );
  CLKBUFX2TS U826 ( .A(n1029), .Y(n339) );
  INVX2TS U827 ( .A(n339), .Y(n373) );
  INVX2TS U828 ( .A(n320), .Y(n1099) );
  INVX2TS U829 ( .A(n1099), .Y(n1013) );
  CLKBUFX2TS U830 ( .A(n359), .Y(n1020) );
  INVX2TS U831 ( .A(n1020), .Y(n348) );
  OR2X1TS U832 ( .A(n1648), .B(n324), .Y(n346) );
  INVX2TS U833 ( .A(n346), .Y(n1848) );
  AOI22X1TS U834 ( .A0(n348), .A1(\destinationAddressbuffer[1][9] ), .B0(n1848), .B1(n322), .Y(n330) );
  INVX2TS U835 ( .A(n332), .Y(n367) );
  INVX2TS U836 ( .A(n367), .Y(n1022) );
  INVX2TS U837 ( .A(n326), .Y(n349) );
  AOI22X1TS U838 ( .A0(n1022), .A1(n328), .B0(n369), .B1(n327), .Y(n329) );
  OAI211XLTS U839 ( .A0(n373), .A1(n35), .B0(n330), .C0(n329), .Y(n2174) );
  INVX2TS U840 ( .A(n339), .Y(n380) );
  INVX2TS U841 ( .A(n346), .Y(n1859) );
  AOI22X1TS U842 ( .A0(n348), .A1(\destinationAddressbuffer[1][10] ), .B0(
        n1859), .B1(n331), .Y(n338) );
  INVX2TS U843 ( .A(n332), .Y(n375) );
  INVX2TS U844 ( .A(n375), .Y(n333) );
  INVX2TS U845 ( .A(n349), .Y(n1883) );
  INVX2TS U846 ( .A(n349), .Y(n335) );
  AOI22X1TS U847 ( .A0(n333), .A1(n336), .B0(n335), .B1(n334), .Y(n337) );
  OAI211XLTS U848 ( .A0(n380), .A1(n53), .B0(n338), .C0(n337), .Y(n2175) );
  INVX2TS U849 ( .A(n339), .Y(n387) );
  INVX2TS U850 ( .A(n346), .Y(n340) );
  INVX2TS U851 ( .A(n340), .Y(n1028) );
  INVX2TS U852 ( .A(n1028), .Y(n361) );
  AOI22X1TS U853 ( .A0(n348), .A1(\destinationAddressbuffer[1][8] ), .B0(n361), 
        .B1(n341), .Y(n345) );
  INVX2TS U854 ( .A(n375), .Y(n1851) );
  AOI22X1TS U855 ( .A0(n1851), .A1(n343), .B0(n326), .B1(n342), .Y(n344) );
  OAI211XLTS U856 ( .A0(n387), .A1(n50), .B0(n345), .C0(n344), .Y(n2173) );
  INVX2TS U857 ( .A(n346), .Y(n1871) );
  AOI22X1TS U858 ( .A0(n348), .A1(\destinationAddressbuffer[1][11] ), .B0(
        n1871), .B1(n347), .Y(n353) );
  INVX2TS U859 ( .A(n326), .Y(n1031) );
  INVX2TS U860 ( .A(n1031), .Y(n369) );
  AOI22X1TS U861 ( .A0(n333), .A1(n351), .B0(n369), .B1(n350), .Y(n352) );
  OAI211XLTS U862 ( .A0(n373), .A1(n43), .B0(n353), .C0(n352), .Y(n2176) );
  INVX2TS U863 ( .A(n359), .Y(n1879) );
  AOI22X1TS U864 ( .A0(n1879), .A1(writeOutbuffer[1]), .B0(n361), .B1(n354), 
        .Y(n358) );
  INVX2TS U865 ( .A(n375), .Y(n1875) );
  AOI22X1TS U866 ( .A0(n1875), .A1(n356), .B0(n326), .B1(n355), .Y(n357) );
  OAI211XLTS U867 ( .A0(n380), .A1(n58), .B0(n358), .C0(n357), .Y(n2083) );
  INVX2TS U868 ( .A(n359), .Y(n382) );
  AOI22X1TS U869 ( .A0(n382), .A1(\destinationAddressbuffer[1][4] ), .B0(n361), 
        .B1(n360), .Y(n365) );
  AOI22X1TS U870 ( .A0(n1851), .A1(n363), .B0(n1103), .B1(n362), .Y(n364) );
  OAI211XLTS U871 ( .A0(n387), .A1(n75), .B0(n365), .C0(n364), .Y(n2169) );
  AOI22X1TS U872 ( .A0(n382), .A1(\destinationAddressbuffer[1][6] ), .B0(n340), 
        .B1(n366), .Y(n372) );
  INVX2TS U873 ( .A(n367), .Y(n1885) );
  AOI22X1TS U874 ( .A0(n1885), .A1(n370), .B0(n369), .B1(n368), .Y(n371) );
  OAI211XLTS U875 ( .A0(n373), .A1(n64), .B0(n372), .C0(n371), .Y(n2171) );
  AOI22X1TS U876 ( .A0(n382), .A1(\destinationAddressbuffer[1][7] ), .B0(n1871), .B1(n374), .Y(n379) );
  INVX2TS U877 ( .A(n375), .Y(n1862) );
  AOI22X1TS U878 ( .A0(n1862), .A1(n377), .B0(n1883), .B1(n376), .Y(n378) );
  OAI211XLTS U879 ( .A0(n380), .A1(n72), .B0(n379), .C0(n378), .Y(n2172) );
  AOI22X1TS U880 ( .A0(n382), .A1(\destinationAddressbuffer[1][5] ), .B0(n1859), .B1(n381), .Y(n386) );
  INVX2TS U881 ( .A(n349), .Y(n1109) );
  AOI22X1TS U882 ( .A0(n1862), .A1(n384), .B0(n1109), .B1(n383), .Y(n385) );
  OAI211XLTS U883 ( .A0(n387), .A1(n67), .B0(n386), .C0(n385), .Y(n2170) );
  AOI31XLTS U884 ( .A0(n394), .A1(n393), .A2(n448), .B0(n1657), .Y(n395) );
  AOI21X1TS U885 ( .A0(n402), .A1(n395), .B0(n456), .Y(n399) );
  NAND2X1TS U886 ( .A(n399), .B(n1666), .Y(n403) );
  INVX2TS U887 ( .A(n398), .Y(n1072) );
  INVX2TS U888 ( .A(n1072), .Y(n1056) );
  CLKBUFX2TS U889 ( .A(n1056), .Y(n414) );
  INVX2TS U890 ( .A(n414), .Y(n436) );
  INVX2TS U891 ( .A(n14), .Y(n1044) );
  INVX2TS U892 ( .A(n429), .Y(n422) );
  OR2X1TS U893 ( .A(n1662), .B(n403), .Y(n420) );
  INVX2TS U894 ( .A(n420), .Y(n400) );
  INVX2TS U895 ( .A(n400), .Y(n1055) );
  INVX2TS U896 ( .A(n1055), .Y(n437) );
  AOI22X1TS U897 ( .A0(n422), .A1(\destinationAddressbuffer[0][11] ), .B0(n437), .B1(n401), .Y(n408) );
  INVX2TS U898 ( .A(n5), .Y(n1915) );
  INVX2TS U899 ( .A(n7), .Y(n405) );
  INVX2TS U900 ( .A(n405), .Y(n1039) );
  INVX2TS U901 ( .A(n1039), .Y(n411) );
  AOI22X1TS U902 ( .A0(n1915), .A1(n771), .B0(n411), .B1(n406), .Y(n407) );
  OAI211XLTS U903 ( .A0(n436), .A1(n43), .B0(n408), .C0(n407), .Y(n2188) );
  INVX2TS U904 ( .A(n420), .Y(n1911) );
  AOI22X1TS U905 ( .A0(n422), .A1(\destinationAddressbuffer[0][10] ), .B0(
        n1911), .B1(n409), .Y(n413) );
  AOI22X1TS U906 ( .A0(n416), .A1(n756), .B0(n411), .B1(n410), .Y(n412) );
  OAI211XLTS U907 ( .A0(n436), .A1(n53), .B0(n413), .C0(n412), .Y(n2187) );
  INVX2TS U908 ( .A(n414), .Y(n446) );
  INVX2TS U909 ( .A(n420), .Y(n1890) );
  AOI22X1TS U910 ( .A0(n422), .A1(\destinationAddressbuffer[0][9] ), .B0(n400), 
        .B1(n415), .Y(n419) );
  INVX2TS U911 ( .A(n5), .Y(n416) );
  INVX2TS U912 ( .A(n416), .Y(n1038) );
  INVX2TS U913 ( .A(n1038), .Y(n439) );
  INVX2TS U914 ( .A(n7), .Y(n1902) );
  AOI22X1TS U915 ( .A0(n439), .A1(n737), .B0(n1902), .B1(n417), .Y(n418) );
  OAI211XLTS U916 ( .A0(n446), .A1(n35), .B0(n419), .C0(n418), .Y(n2186) );
  INVX2TS U917 ( .A(n420), .Y(n1900) );
  AOI22X1TS U918 ( .A0(n422), .A1(\destinationAddressbuffer[0][8] ), .B0(n1900), .B1(n421), .Y(n425) );
  INVX2TS U919 ( .A(n5), .Y(n1067) );
  INVX2TS U920 ( .A(n7), .Y(n1913) );
  AOI22X1TS U921 ( .A0(n1067), .A1(n722), .B0(n1913), .B1(n423), .Y(n424) );
  OAI211XLTS U922 ( .A0(n436), .A1(n50), .B0(n425), .C0(n424), .Y(n2185) );
  INVX2TS U923 ( .A(n429), .Y(n1919) );
  AOI22X1TS U924 ( .A0(n1919), .A1(writeOutbuffer[0]), .B0(n1911), .B1(
        writeIn_WEST), .Y(n428) );
  INVX2TS U925 ( .A(n7), .Y(n1062) );
  AOI22X1TS U926 ( .A0(n1067), .A1(n550), .B0(n1062), .B1(n426), .Y(n427) );
  OAI211XLTS U927 ( .A0(n446), .A1(n58), .B0(n428), .C0(n427), .Y(n2084) );
  CLKBUFX2TS U928 ( .A(n429), .Y(n1071) );
  INVX2TS U929 ( .A(n1071), .Y(n442) );
  AOI22X1TS U930 ( .A0(n442), .A1(\destinationAddressbuffer[0][7] ), .B0(n1900), .B1(destinationAddressIn_WEST[7]), .Y(n432) );
  AOI22X1TS U931 ( .A0(n416), .A1(n711), .B0(n1062), .B1(n430), .Y(n431) );
  OAI211XLTS U932 ( .A0(n446), .A1(n72), .B0(n432), .C0(n431), .Y(n2184) );
  AOI22X1TS U933 ( .A0(n442), .A1(\destinationAddressbuffer[0][6] ), .B0(n1890), .B1(destinationAddressIn_WEST[6]), .Y(n435) );
  INVX2TS U934 ( .A(n5), .Y(n1893) );
  AOI22X1TS U935 ( .A0(n1893), .A1(n697), .B0(n405), .B1(n433), .Y(n434) );
  OAI211XLTS U936 ( .A0(n436), .A1(n64), .B0(n435), .C0(n434), .Y(n2183) );
  AOI22X1TS U937 ( .A0(n442), .A1(\destinationAddressbuffer[0][5] ), .B0(n437), 
        .B1(destinationAddressIn_WEST[5]), .Y(n441) );
  AOI22X1TS U938 ( .A0(n439), .A1(n677), .B0(n411), .B1(n438), .Y(n440) );
  OAI211XLTS U939 ( .A0(n1072), .A1(n67), .B0(n441), .C0(n440), .Y(n2182) );
  AOI22X1TS U940 ( .A0(n442), .A1(\destinationAddressbuffer[0][4] ), .B0(n437), 
        .B1(destinationAddressIn_WEST[4]), .Y(n445) );
  AOI22X1TS U941 ( .A0(n416), .A1(n665), .B0(n1913), .B1(n443), .Y(n444) );
  OAI211XLTS U942 ( .A0(n446), .A1(n75), .B0(n445), .C0(n444), .Y(n2181) );
  INVX2TS U943 ( .A(n1955), .Y(n533) );
  INVX2TS U944 ( .A(n1955), .Y(n530) );
  INVX2TS U945 ( .A(n1949), .Y(n536) );
  NAND2X1TS U946 ( .A(n530), .B(n536), .Y(n534) );
  OAI21XLTS U947 ( .A0(n533), .A1(n1950), .B0(n534), .Y(n508) );
  INVX2TS U948 ( .A(n1946), .Y(n537) );
  INVX2TS U949 ( .A(n1946), .Y(n532) );
  NOR2XLTS U950 ( .A(n534), .B(n532), .Y(n843) );
  CLKBUFX2TS U951 ( .A(n843), .Y(n801) );
  CLKBUFX2TS U952 ( .A(n801), .Y(n820) );
  AOI21X1TS U953 ( .A0(n534), .A1(n537), .B0(n820), .Y(n505) );
  OAI22X1TS U954 ( .A0(n491), .A1(n508), .B0(n448), .B1(n505), .Y(n449) );
  AOI221XLTS U955 ( .A0(n508), .A1(n462), .B0(n450), .B1(n505), .C0(n449), .Y(
        n454) );
  INVX2TS U956 ( .A(n1943), .Y(n451) );
  NAND2X1TS U957 ( .A(n452), .B(n451), .Y(n467) );
  OAI21XLTS U958 ( .A0(n453), .A1(n1955), .B0(n467), .Y(n471) );
  AOI21X1TS U959 ( .A0(n454), .A1(n471), .B0(n1945), .Y(n455) );
  INVX2TS U960 ( .A(reset), .Y(n498) );
  NAND2X1TS U961 ( .A(n498), .B(n1945), .Y(n509) );
  NOR2XLTS U962 ( .A(reset), .B(n456), .Y(n503) );
  INVX2TS U963 ( .A(n1951), .Y(n468) );
  INVX2TS U964 ( .A(n1954), .Y(n458) );
  INVX2TS U965 ( .A(n1947), .Y(n535) );
  AOI22X1TS U966 ( .A0(n458), .A1(n532), .B0(n535), .B1(n457), .Y(n461) );
  INVX2TS U967 ( .A(n460), .Y(n466) );
  INVX2TS U968 ( .A(n481), .Y(n478) );
  AOI21X1TS U969 ( .A0(n533), .A1(n464), .B0(n463), .Y(n477) );
  ADDHXLTS U970 ( .A(n470), .B(n469), .CO(n481), .S(n483) );
  INVX2TS U971 ( .A(n483), .Y(n472) );
  AOI21X1TS U972 ( .A0(n473), .A1(n472), .B0(n471), .Y(n475) );
  OAI22X1TS U973 ( .A0(n473), .A1(n472), .B0(n479), .B1(n478), .Y(n474) );
  AOI21X1TS U974 ( .A0(n482), .A1(n475), .B0(n474), .Y(n476) );
  AOI211X1TS U975 ( .A0(n479), .A1(n478), .B0(n477), .C0(n476), .Y(n480) );
  INVX2TS U976 ( .A(n480), .Y(n484) );
  NAND2X1TS U977 ( .A(n484), .B(n481), .Y(n488) );
  XNOR2X1TS U978 ( .A(n486), .B(n485), .Y(n487) );
  XOR2X1TS U979 ( .A(n488), .B(n487), .Y(n502) );
  INVX2TS U980 ( .A(n502), .Y(n496) );
  INVX2TS U981 ( .A(n1947), .Y(n531) );
  ADDHXLTS U982 ( .A(n452), .B(n489), .CO(n492), .S(n499) );
  XNOR2X1TS U983 ( .A(n1950), .B(n500), .Y(n493) );
  OAI2BB2XLTS U984 ( .B0(n1957), .B1(n509), .A0N(n503), .A1N(n497), .Y(N2624)
         );
  NAND2X1TS U985 ( .A(n498), .B(n1944), .Y(n507) );
  AOI22X1TS U986 ( .A0(n1943), .A1(n509), .B0(n507), .B1(n451), .Y(n1966) );
  INVX2TS U987 ( .A(n505), .Y(n506) );
  OAI22X1TS U988 ( .A0(n537), .A1(n509), .B0(n506), .B1(n507), .Y(n1971) );
  OAI22X1TS U989 ( .A0(n15), .A1(n509), .B0(n508), .B1(n507), .Y(n1972) );
  CLKBUFX2TS U990 ( .A(readIn_SOUTH), .Y(n1656) );
  CLKBUFX2TS U991 ( .A(n1656), .Y(n1597) );
  CLKBUFX2TS U992 ( .A(n1944), .Y(n849) );
  CLKBUFX2TS U993 ( .A(n549), .Y(n632) );
  CLKBUFX2TS U994 ( .A(n632), .Y(n858) );
  CLKBUFX2TS U995 ( .A(readIn_WEST), .Y(n1664) );
  CLKBUFX2TS U996 ( .A(n1664), .Y(n1650) );
  INVX2TS U997 ( .A(n1944), .Y(n526) );
  NAND2X1TS U998 ( .A(n544), .B(n526), .Y(n514) );
  NOR4XLTS U999 ( .A(readReady), .B(n517), .C(n460), .D(n514), .Y(n617) );
  CLKBUFX2TS U1000 ( .A(n617), .Y(n633) );
  CLKBUFX2TS U1001 ( .A(n633), .Y(n812) );
  CLKBUFX2TS U1002 ( .A(n812), .Y(n570) );
  AOI22X1TS U1003 ( .A0(n1597), .A1(n858), .B0(n1650), .B1(n570), .Y(n547) );
  CLKBUFX2TS U1004 ( .A(readIn_NORTH), .Y(n1655) );
  CLKBUFX2TS U1005 ( .A(n1655), .Y(n1596) );
  CLKBUFX2TS U1006 ( .A(n696), .Y(n631) );
  CLKBUFX2TS U1007 ( .A(n631), .Y(n569) );
  NOR4XLTS U1008 ( .A(selectBit_WEST), .B(n515), .C(n519), .D(n514), .Y(n651)
         );
  CLKBUFX2TS U1009 ( .A(n651), .Y(n782) );
  CLKBUFX2TS U1010 ( .A(n782), .Y(n674) );
  CLKBUFX2TS U1011 ( .A(n674), .Y(n831) );
  AOI22X1TS U1012 ( .A0(n1596), .A1(n569), .B0(readIn_EAST), .B1(n831), .Y(
        n546) );
  NOR3XLTS U1013 ( .A(n517), .B(n516), .C(n460), .Y(n522) );
  NOR3XLTS U1014 ( .A(selectBit_WEST), .B(n520), .C(n519), .Y(n521) );
  OAI31X1TS U1015 ( .A0(n522), .A1(n543), .A2(n521), .B0(n544), .Y(n525) );
  NAND4XLTS U1016 ( .A(n526), .B(n525), .C(n524), .D(n523), .Y(n679) );
  INVX2TS U1017 ( .A(n679), .Y(n527) );
  INVX2TS U1018 ( .A(n527), .Y(n634) );
  INVX2TS U1019 ( .A(n634), .Y(n528) );
  CLKBUFX2TS U1020 ( .A(n1944), .Y(n605) );
  NOR3XLTS U1021 ( .A(n530), .B(n531), .C(n1949), .Y(n724) );
  CLKBUFX2TS U1022 ( .A(n724), .Y(n635) );
  CLKBUFX2TS U1023 ( .A(n635), .Y(n572) );
  NOR3XLTS U1024 ( .A(n533), .B(n1950), .C(n531), .Y(n698) );
  CLKBUFX2TS U1025 ( .A(n698), .Y(n636) );
  CLKBUFX2TS U1026 ( .A(n636), .Y(n571) );
  AOI22X1TS U1027 ( .A0(readOutbuffer[2]), .A1(n572), .B0(readOutbuffer[0]), 
        .B1(n571), .Y(n541) );
  NOR3XLTS U1028 ( .A(n530), .B(n15), .C(n532), .Y(n725) );
  CLKBUFX2TS U1029 ( .A(n725), .Y(n637) );
  CLKBUFX2TS U1030 ( .A(n637), .Y(n574) );
  NOR3XLTS U1031 ( .A(n533), .B(n536), .C(n537), .Y(n699) );
  CLKBUFX2TS U1032 ( .A(n699), .Y(n638) );
  CLKBUFX2TS U1033 ( .A(n638), .Y(n573) );
  AOI22X1TS U1034 ( .A0(readOutbuffer[6]), .A1(n574), .B0(readOutbuffer[4]), 
        .B1(n573), .Y(n540) );
  NOR2XLTS U1035 ( .A(n535), .B(n534), .Y(n726) );
  CLKBUFX2TS U1036 ( .A(n726), .Y(n639) );
  CLKBUFX2TS U1037 ( .A(n639), .Y(n576) );
  NOR3XLTS U1038 ( .A(n536), .B(n535), .C(n1955), .Y(n700) );
  CLKBUFX2TS U1039 ( .A(n700), .Y(n640) );
  CLKBUFX2TS U1040 ( .A(n640), .Y(n575) );
  AOI22X1TS U1041 ( .A0(readOutbuffer[3]), .A1(n576), .B0(readOutbuffer[1]), 
        .B1(n575), .Y(n539) );
  CLKBUFX2TS U1042 ( .A(n843), .Y(n865) );
  NOR3XLTS U1043 ( .A(n1950), .B(n451), .C(n537), .Y(n866) );
  CLKBUFX2TS U1044 ( .A(n866), .Y(n641) );
  CLKBUFX2TS U1045 ( .A(n641), .Y(n577) );
  AOI22X1TS U1046 ( .A0(readOutbuffer[7]), .A1(n865), .B0(readOutbuffer[5]), 
        .B1(n577), .Y(n538) );
  NAND4XLTS U1047 ( .A(n541), .B(n540), .C(n539), .D(n538), .Y(n542) );
  AOI22X1TS U1048 ( .A0(readOut), .A1(n556), .B0(n605), .B1(n542), .Y(n545) );
  CLKBUFX2TS U1049 ( .A(n674), .Y(n754) );
  AOI22X1TS U1050 ( .A0(writeIn_EAST), .A1(n754), .B0(n548), .B1(n570), .Y(
        n559) );
  CLKBUFX2TS U1051 ( .A(n632), .Y(n770) );
  AOI22X1TS U1052 ( .A0(writeIn_NORTH), .A1(n569), .B0(n550), .B1(n770), .Y(
        n558) );
  AOI22X1TS U1053 ( .A0(writeOutbuffer[2]), .A1(n572), .B0(writeOutbuffer[0]), 
        .B1(n571), .Y(n554) );
  AOI22X1TS U1054 ( .A0(writeOutbuffer[6]), .A1(n574), .B0(writeOutbuffer[4]), 
        .B1(n573), .Y(n553) );
  AOI22X1TS U1055 ( .A0(writeOutbuffer[3]), .A1(n576), .B0(writeOutbuffer[1]), 
        .B1(n575), .Y(n552) );
  AOI22X1TS U1056 ( .A0(writeOutbuffer[7]), .A1(n865), .B0(writeOutbuffer[5]), 
        .B1(n577), .Y(n551) );
  NAND4XLTS U1057 ( .A(n554), .B(n553), .C(n552), .D(n551), .Y(n555) );
  AOI22X1TS U1058 ( .A0(writeOut), .A1(n556), .B0(n605), .B1(n555), .Y(n557)
         );
  CLKBUFX2TS U1059 ( .A(requesterAddressIn_NORTH[0]), .Y(n1008) );
  CLKBUFX2TS U1060 ( .A(requesterAddressIn_EAST[0]), .Y(n1037) );
  CLKBUFX2TS U1061 ( .A(n1037), .Y(n1007) );
  CLKBUFX2TS U1062 ( .A(n674), .Y(n594) );
  AOI22X1TS U1063 ( .A0(n1008), .A1(n569), .B0(n1007), .B1(n594), .Y(n568) );
  CLKBUFX2TS U1064 ( .A(requesterAddressIn_SOUTH[0]), .Y(n1040) );
  CLKBUFX2TS U1065 ( .A(n1040), .Y(n1009) );
  CLKBUFX2TS U1066 ( .A(n549), .Y(n664) );
  CLKBUFX2TS U1067 ( .A(requesterAddressIn_WEST[0]), .Y(n932) );
  CLKBUFX2TS U1068 ( .A(n932), .Y(n961) );
  AOI22X1TS U1069 ( .A0(n1009), .A1(n664), .B0(n961), .B1(n570), .Y(n567) );
  INVX2TS U1070 ( .A(n679), .Y(n706) );
  CLKBUFX2TS U1071 ( .A(n605), .Y(n600) );
  AOI22X1TS U1072 ( .A0(\requesterAddressbuffer[2][0] ), .A1(n572), .B0(
        \requesterAddressbuffer[0][0] ), .B1(n571), .Y(n563) );
  AOI22X1TS U1073 ( .A0(\requesterAddressbuffer[6][0] ), .A1(n574), .B0(
        \requesterAddressbuffer[4][0] ), .B1(n573), .Y(n562) );
  AOI22X1TS U1074 ( .A0(\requesterAddressbuffer[3][0] ), .A1(n576), .B0(
        \requesterAddressbuffer[1][0] ), .B1(n575), .Y(n561) );
  CLKBUFX2TS U1075 ( .A(n801), .Y(n758) );
  CLKBUFX2TS U1076 ( .A(n758), .Y(n606) );
  AOI22X1TS U1077 ( .A0(\requesterAddressbuffer[7][0] ), .A1(n606), .B0(
        \requesterAddressbuffer[5][0] ), .B1(n577), .Y(n560) );
  NAND4XLTS U1078 ( .A(n563), .B(n562), .C(n561), .D(n560), .Y(n564) );
  AOI22X1TS U1079 ( .A0(requesterAddressOut[0]), .A1(n706), .B0(n600), .B1(
        n564), .Y(n566) );
  INVX2TS U1080 ( .A(readRequesterAddress[0]), .Y(n959) );
  INVX2TS U1081 ( .A(n959), .Y(n1006) );
  INVX2TS U1082 ( .A(n565), .Y(n601) );
  NAND2X1TS U1083 ( .A(n1006), .B(n601), .Y(n612) );
  CLKBUFX2TS U1084 ( .A(requesterAddressIn_NORTH[1]), .Y(n1015) );
  CLKBUFX2TS U1085 ( .A(requesterAddressIn_EAST[1]), .Y(n1045) );
  CLKBUFX2TS U1086 ( .A(n1045), .Y(n1014) );
  AOI22X1TS U1087 ( .A0(n1015), .A1(n569), .B0(n1014), .B1(n594), .Y(n585) );
  CLKBUFX2TS U1088 ( .A(requesterAddressIn_SOUTH[1]), .Y(n1046) );
  CLKBUFX2TS U1089 ( .A(n1046), .Y(n1016) );
  CLKBUFX2TS U1090 ( .A(n632), .Y(n813) );
  CLKBUFX2TS U1091 ( .A(requesterAddressIn_WEST[1]), .Y(n940) );
  CLKBUFX2TS U1092 ( .A(n940), .Y(n969) );
  AOI22X1TS U1093 ( .A0(n1016), .A1(n813), .B0(n969), .B1(n570), .Y(n584) );
  AOI22X1TS U1094 ( .A0(\requesterAddressbuffer[2][1] ), .A1(n572), .B0(
        \requesterAddressbuffer[0][1] ), .B1(n571), .Y(n581) );
  AOI22X1TS U1095 ( .A0(\requesterAddressbuffer[6][1] ), .A1(n574), .B0(
        \requesterAddressbuffer[4][1] ), .B1(n573), .Y(n580) );
  AOI22X1TS U1096 ( .A0(\requesterAddressbuffer[3][1] ), .A1(n576), .B0(
        \requesterAddressbuffer[1][1] ), .B1(n575), .Y(n579) );
  AOI22X1TS U1097 ( .A0(\requesterAddressbuffer[7][1] ), .A1(n606), .B0(
        \requesterAddressbuffer[5][1] ), .B1(n577), .Y(n578) );
  NAND4XLTS U1098 ( .A(n581), .B(n580), .C(n579), .D(n578), .Y(n582) );
  AOI22X1TS U1099 ( .A0(requesterAddressOut[1]), .A1(n528), .B0(n600), .B1(
        n582), .Y(n583) );
  INVX2TS U1100 ( .A(readRequesterAddress[1]), .Y(n966) );
  INVX2TS U1101 ( .A(n966), .Y(n1674) );
  NAND2X1TS U1102 ( .A(n1674), .B(n601), .Y(n627) );
  CLKBUFX2TS U1103 ( .A(requesterAddressIn_NORTH[2]), .Y(n1023) );
  CLKBUFX2TS U1104 ( .A(n631), .Y(n616) );
  CLKBUFX2TS U1105 ( .A(requesterAddressIn_EAST[2]), .Y(n1050) );
  CLKBUFX2TS U1106 ( .A(n1050), .Y(n1021) );
  AOI22X1TS U1107 ( .A0(n1023), .A1(n616), .B0(n1021), .B1(n594), .Y(n593) );
  CLKBUFX2TS U1108 ( .A(requesterAddressIn_SOUTH[2]), .Y(n1051) );
  CLKBUFX2TS U1109 ( .A(n1051), .Y(n1024) );
  CLKBUFX2TS U1110 ( .A(requesterAddressIn_WEST[2]), .Y(n947) );
  CLKBUFX2TS U1111 ( .A(n947), .Y(n976) );
  AOI22X1TS U1112 ( .A0(n1024), .A1(n664), .B0(n976), .B1(n633), .Y(n592) );
  INVX2TS U1113 ( .A(n679), .Y(n749) );
  CLKBUFX2TS U1114 ( .A(n635), .Y(n618) );
  AOI22X1TS U1115 ( .A0(\requesterAddressbuffer[2][2] ), .A1(n618), .B0(
        \requesterAddressbuffer[0][2] ), .B1(n698), .Y(n589) );
  CLKBUFX2TS U1116 ( .A(n637), .Y(n619) );
  AOI22X1TS U1117 ( .A0(\requesterAddressbuffer[6][2] ), .A1(n619), .B0(
        \requesterAddressbuffer[4][2] ), .B1(n699), .Y(n588) );
  CLKBUFX2TS U1118 ( .A(n639), .Y(n620) );
  AOI22X1TS U1119 ( .A0(\requesterAddressbuffer[3][2] ), .A1(n620), .B0(
        \requesterAddressbuffer[1][2] ), .B1(n700), .Y(n587) );
  CLKBUFX2TS U1120 ( .A(n641), .Y(n621) );
  AOI22X1TS U1121 ( .A0(\requesterAddressbuffer[7][2] ), .A1(n606), .B0(
        \requesterAddressbuffer[5][2] ), .B1(n621), .Y(n586) );
  NAND4XLTS U1122 ( .A(n589), .B(n588), .C(n587), .D(n586), .Y(n590) );
  AOI22X1TS U1123 ( .A0(requesterAddressOut[2]), .A1(n749), .B0(n600), .B1(
        n590), .Y(n591) );
  INVX2TS U1124 ( .A(readRequesterAddress[2]), .Y(n975) );
  INVX2TS U1125 ( .A(n975), .Y(n1682) );
  NAND2X1TS U1126 ( .A(n1682), .B(n601), .Y(n647) );
  CLKBUFX2TS U1127 ( .A(requesterAddressIn_NORTH[3]), .Y(n1032) );
  CLKBUFX2TS U1128 ( .A(requesterAddressIn_EAST[3]), .Y(n1057) );
  CLKBUFX2TS U1129 ( .A(n1057), .Y(n1030) );
  AOI22X1TS U1130 ( .A0(n1032), .A1(n616), .B0(n1030), .B1(n594), .Y(n604) );
  CLKBUFX2TS U1131 ( .A(requesterAddressIn_SOUTH[3]), .Y(n1058) );
  CLKBUFX2TS U1132 ( .A(n1058), .Y(n1033) );
  CLKBUFX2TS U1133 ( .A(requesterAddressIn_WEST[3]), .Y(n954) );
  CLKBUFX2TS U1134 ( .A(n954), .Y(n984) );
  AOI22X1TS U1135 ( .A0(n1033), .A1(n813), .B0(n984), .B1(n617), .Y(n603) );
  AOI22X1TS U1136 ( .A0(\requesterAddressbuffer[2][3] ), .A1(n618), .B0(
        \requesterAddressbuffer[0][3] ), .B1(n698), .Y(n598) );
  AOI22X1TS U1137 ( .A0(\requesterAddressbuffer[6][3] ), .A1(n619), .B0(
        \requesterAddressbuffer[4][3] ), .B1(n699), .Y(n597) );
  AOI22X1TS U1138 ( .A0(\requesterAddressbuffer[3][3] ), .A1(n620), .B0(
        \requesterAddressbuffer[1][3] ), .B1(n700), .Y(n596) );
  CLKBUFX2TS U1139 ( .A(n758), .Y(n652) );
  AOI22X1TS U1140 ( .A0(\requesterAddressbuffer[7][3] ), .A1(n652), .B0(
        \requesterAddressbuffer[5][3] ), .B1(n621), .Y(n595) );
  NAND4XLTS U1141 ( .A(n598), .B(n597), .C(n596), .D(n595), .Y(n599) );
  AOI22X1TS U1142 ( .A0(requesterAddressOut[3]), .A1(n749), .B0(n600), .B1(
        n599), .Y(n602) );
  INVX2TS U1143 ( .A(readRequesterAddress[3]), .Y(n983) );
  INVX2TS U1144 ( .A(n983), .Y(n1690) );
  NAND2X1TS U1145 ( .A(n1690), .B(n601), .Y(n659) );
  CLKBUFX2TS U1146 ( .A(destinationAddressIn_NORTH[0]), .Y(n1697) );
  CLKBUFX2TS U1147 ( .A(destinationAddressIn_EAST[0]), .Y(n1847) );
  CLKBUFX2TS U1148 ( .A(n1847), .Y(n1727) );
  AOI22X1TS U1149 ( .A0(n1697), .A1(n616), .B0(n1727), .B1(n782), .Y(n615) );
  CLKBUFX2TS U1150 ( .A(destinationAddressIn_WEST[0]), .Y(n1728) );
  CLKBUFX2TS U1151 ( .A(n1728), .Y(n1791) );
  AOI22X1TS U1152 ( .A0(destinationAddressIn_SOUTH[0]), .A1(n664), .B0(n1791), 
        .B1(n617), .Y(n614) );
  CLKBUFX2TS U1153 ( .A(n605), .Y(n658) );
  AOI22X1TS U1154 ( .A0(\destinationAddressbuffer[2][0] ), .A1(n618), .B0(
        \destinationAddressbuffer[0][0] ), .B1(n636), .Y(n610) );
  AOI22X1TS U1155 ( .A0(\destinationAddressbuffer[6][0] ), .A1(n619), .B0(
        \destinationAddressbuffer[4][0] ), .B1(n638), .Y(n609) );
  AOI22X1TS U1156 ( .A0(\destinationAddressbuffer[3][0] ), .A1(n620), .B0(
        \destinationAddressbuffer[1][0] ), .B1(n640), .Y(n608) );
  AOI22X1TS U1157 ( .A0(\destinationAddressbuffer[7][0] ), .A1(n606), .B0(
        \destinationAddressbuffer[5][0] ), .B1(n621), .Y(n607) );
  NAND4XLTS U1158 ( .A(n610), .B(n609), .C(n608), .D(n607), .Y(n611) );
  AOI22X1TS U1159 ( .A0(destinationAddressOut[0]), .A1(n749), .B0(n658), .B1(
        n611), .Y(n613) );
  CLKBUFX2TS U1160 ( .A(destinationAddressIn_NORTH[1]), .Y(n1705) );
  CLKBUFX2TS U1161 ( .A(destinationAddressIn_EAST[1]), .Y(n1857) );
  CLKBUFX2TS U1162 ( .A(n1857), .Y(n1734) );
  AOI22X1TS U1163 ( .A0(n1705), .A1(n616), .B0(n1734), .B1(n651), .Y(n630) );
  CLKBUFX2TS U1164 ( .A(destinationAddressIn_WEST[1]), .Y(n1736) );
  CLKBUFX2TS U1165 ( .A(n1736), .Y(n1798) );
  AOI22X1TS U1166 ( .A0(destinationAddressIn_SOUTH[1]), .A1(n813), .B0(n1798), 
        .B1(n617), .Y(n629) );
  AOI22X1TS U1167 ( .A0(\destinationAddressbuffer[2][1] ), .A1(n618), .B0(
        \destinationAddressbuffer[0][1] ), .B1(n636), .Y(n625) );
  AOI22X1TS U1168 ( .A0(\destinationAddressbuffer[6][1] ), .A1(n619), .B0(
        \destinationAddressbuffer[4][1] ), .B1(n638), .Y(n624) );
  AOI22X1TS U1169 ( .A0(\destinationAddressbuffer[3][1] ), .A1(n620), .B0(
        \destinationAddressbuffer[1][1] ), .B1(n640), .Y(n623) );
  AOI22X1TS U1170 ( .A0(\destinationAddressbuffer[7][1] ), .A1(n652), .B0(
        \destinationAddressbuffer[5][1] ), .B1(n621), .Y(n622) );
  NAND4XLTS U1171 ( .A(n625), .B(n624), .C(n623), .D(n622), .Y(n626) );
  AOI22X1TS U1172 ( .A0(destinationAddressOut[1]), .A1(n706), .B0(n658), .B1(
        n626), .Y(n628) );
  CLKBUFX2TS U1173 ( .A(destinationAddressIn_NORTH[2]), .Y(n1713) );
  CLKBUFX2TS U1174 ( .A(n631), .Y(n678) );
  CLKBUFX2TS U1175 ( .A(destinationAddressIn_EAST[2]), .Y(n1869) );
  CLKBUFX2TS U1176 ( .A(n1869), .Y(n1745) );
  AOI22X1TS U1177 ( .A0(n1713), .A1(n678), .B0(n1745), .B1(n651), .Y(n650) );
  CLKBUFX2TS U1178 ( .A(n632), .Y(n794) );
  CLKBUFX2TS U1179 ( .A(destinationAddressIn_WEST[2]), .Y(n1747) );
  CLKBUFX2TS U1180 ( .A(n1747), .Y(n1805) );
  CLKBUFX2TS U1181 ( .A(n633), .Y(n675) );
  AOI22X1TS U1182 ( .A0(destinationAddressIn_SOUTH[2]), .A1(n794), .B0(n1805), 
        .B1(n675), .Y(n649) );
  INVX2TS U1183 ( .A(n634), .Y(n873) );
  CLKBUFX2TS U1184 ( .A(n635), .Y(n681) );
  CLKBUFX2TS U1185 ( .A(n636), .Y(n680) );
  AOI22X1TS U1186 ( .A0(\destinationAddressbuffer[2][2] ), .A1(n681), .B0(
        \destinationAddressbuffer[0][2] ), .B1(n680), .Y(n645) );
  CLKBUFX2TS U1187 ( .A(n637), .Y(n683) );
  CLKBUFX2TS U1188 ( .A(n638), .Y(n682) );
  AOI22X1TS U1189 ( .A0(\destinationAddressbuffer[6][2] ), .A1(n683), .B0(
        \destinationAddressbuffer[4][2] ), .B1(n682), .Y(n644) );
  CLKBUFX2TS U1190 ( .A(n639), .Y(n685) );
  CLKBUFX2TS U1191 ( .A(n640), .Y(n684) );
  AOI22X1TS U1192 ( .A0(\destinationAddressbuffer[3][2] ), .A1(n685), .B0(
        \destinationAddressbuffer[1][2] ), .B1(n684), .Y(n643) );
  CLKBUFX2TS U1193 ( .A(n641), .Y(n686) );
  AOI22X1TS U1194 ( .A0(\destinationAddressbuffer[7][2] ), .A1(n652), .B0(
        \destinationAddressbuffer[5][2] ), .B1(n686), .Y(n642) );
  NAND4XLTS U1195 ( .A(n645), .B(n644), .C(n643), .D(n642), .Y(n646) );
  AOI22X1TS U1196 ( .A0(destinationAddressOut[2]), .A1(n873), .B0(n658), .B1(
        n646), .Y(n648) );
  CLKBUFX2TS U1197 ( .A(destinationAddressIn_NORTH[3]), .Y(n1722) );
  CLKBUFX2TS U1198 ( .A(destinationAddressIn_EAST[3]), .Y(n1881) );
  CLKBUFX2TS U1199 ( .A(n1881), .Y(n1756) );
  AOI22X1TS U1200 ( .A0(n1722), .A1(n678), .B0(n1756), .B1(n651), .Y(n662) );
  CLKBUFX2TS U1201 ( .A(destinationAddressIn_WEST[3]), .Y(n1757) );
  CLKBUFX2TS U1202 ( .A(n1757), .Y(n1813) );
  AOI22X1TS U1203 ( .A0(destinationAddressIn_SOUTH[3]), .A1(n794), .B0(n1813), 
        .B1(n675), .Y(n661) );
  AOI22X1TS U1204 ( .A0(\destinationAddressbuffer[2][3] ), .A1(n681), .B0(
        \destinationAddressbuffer[0][3] ), .B1(n680), .Y(n656) );
  AOI22X1TS U1205 ( .A0(\destinationAddressbuffer[6][3] ), .A1(n683), .B0(
        \destinationAddressbuffer[4][3] ), .B1(n682), .Y(n655) );
  AOI22X1TS U1206 ( .A0(\destinationAddressbuffer[3][3] ), .A1(n685), .B0(
        \destinationAddressbuffer[1][3] ), .B1(n684), .Y(n654) );
  AOI22X1TS U1207 ( .A0(\destinationAddressbuffer[7][3] ), .A1(n652), .B0(
        \destinationAddressbuffer[5][3] ), .B1(n686), .Y(n653) );
  NAND4XLTS U1208 ( .A(n656), .B(n655), .C(n654), .D(n653), .Y(n657) );
  AOI22X1TS U1209 ( .A0(destinationAddressOut[3]), .A1(n528), .B0(n658), .B1(
        n657), .Y(n660) );
  AOI22X1TS U1210 ( .A0(destinationAddressIn_EAST[4]), .A1(n754), .B0(n663), 
        .B1(n675), .Y(n673) );
  AOI22X1TS U1211 ( .A0(destinationAddressIn_NORTH[4]), .A1(n678), .B0(n665), 
        .B1(n664), .Y(n672) );
  INVX2TS U1212 ( .A(n1945), .Y(n773) );
  CLKBUFX2TS U1213 ( .A(n773), .Y(n872) );
  AOI22X1TS U1214 ( .A0(\destinationAddressbuffer[2][4] ), .A1(n681), .B0(
        \destinationAddressbuffer[0][4] ), .B1(n680), .Y(n669) );
  AOI22X1TS U1215 ( .A0(\destinationAddressbuffer[6][4] ), .A1(n683), .B0(
        \destinationAddressbuffer[4][4] ), .B1(n682), .Y(n668) );
  AOI22X1TS U1216 ( .A0(\destinationAddressbuffer[3][4] ), .A1(n685), .B0(
        \destinationAddressbuffer[1][4] ), .B1(n684), .Y(n667) );
  CLKBUFX2TS U1217 ( .A(n758), .Y(n712) );
  AOI22X1TS U1218 ( .A0(\destinationAddressbuffer[7][4] ), .A1(n712), .B0(
        \destinationAddressbuffer[5][4] ), .B1(n686), .Y(n666) );
  NAND4XLTS U1219 ( .A(n669), .B(n668), .C(n667), .D(n666), .Y(n670) );
  AOI22X1TS U1220 ( .A0(destinationAddressOut[4]), .A1(n706), .B0(n872), .B1(
        n670), .Y(n671) );
  CLKBUFX2TS U1221 ( .A(n674), .Y(n769) );
  AOI22X1TS U1222 ( .A0(destinationAddressIn_EAST[5]), .A1(n769), .B0(n676), 
        .B1(n675), .Y(n694) );
  CLKBUFX2TS U1223 ( .A(n549), .Y(n755) );
  AOI22X1TS U1224 ( .A0(destinationAddressIn_NORTH[5]), .A1(n678), .B0(n677), 
        .B1(n755), .Y(n693) );
  INVX2TS U1225 ( .A(n679), .Y(n838) );
  AOI22X1TS U1226 ( .A0(\destinationAddressbuffer[2][5] ), .A1(n681), .B0(
        \destinationAddressbuffer[0][5] ), .B1(n680), .Y(n690) );
  AOI22X1TS U1227 ( .A0(\destinationAddressbuffer[6][5] ), .A1(n683), .B0(
        \destinationAddressbuffer[4][5] ), .B1(n682), .Y(n689) );
  AOI22X1TS U1228 ( .A0(\destinationAddressbuffer[3][5] ), .A1(n685), .B0(
        \destinationAddressbuffer[1][5] ), .B1(n684), .Y(n688) );
  AOI22X1TS U1229 ( .A0(\destinationAddressbuffer[7][5] ), .A1(n712), .B0(
        \destinationAddressbuffer[5][5] ), .B1(n686), .Y(n687) );
  NAND4XLTS U1230 ( .A(n690), .B(n689), .C(n688), .D(n687), .Y(n691) );
  AOI22X1TS U1231 ( .A0(destinationAddressOut[5]), .A1(n838), .B0(n872), .B1(
        n691), .Y(n692) );
  CLKBUFX2TS U1232 ( .A(n812), .Y(n735) );
  AOI22X1TS U1233 ( .A0(destinationAddressIn_EAST[6]), .A1(n769), .B0(n695), 
        .B1(n735), .Y(n709) );
  CLKBUFX2TS U1234 ( .A(n696), .Y(n738) );
  AOI22X1TS U1235 ( .A0(destinationAddressIn_NORTH[6]), .A1(n738), .B0(n697), 
        .B1(n755), .Y(n708) );
  CLKBUFX2TS U1236 ( .A(n698), .Y(n814) );
  CLKBUFX2TS U1237 ( .A(n814), .Y(n740) );
  AOI22X1TS U1238 ( .A0(\destinationAddressbuffer[2][6] ), .A1(n724), .B0(
        \destinationAddressbuffer[0][6] ), .B1(n740), .Y(n704) );
  CLKBUFX2TS U1239 ( .A(n699), .Y(n816) );
  CLKBUFX2TS U1240 ( .A(n816), .Y(n741) );
  AOI22X1TS U1241 ( .A0(\destinationAddressbuffer[6][6] ), .A1(n725), .B0(
        \destinationAddressbuffer[4][6] ), .B1(n741), .Y(n703) );
  CLKBUFX2TS U1242 ( .A(n700), .Y(n818) );
  CLKBUFX2TS U1243 ( .A(n818), .Y(n742) );
  AOI22X1TS U1244 ( .A0(\destinationAddressbuffer[3][6] ), .A1(n726), .B0(
        \destinationAddressbuffer[1][6] ), .B1(n742), .Y(n702) );
  CLKBUFX2TS U1245 ( .A(n866), .Y(n832) );
  CLKBUFX2TS U1246 ( .A(n832), .Y(n743) );
  AOI22X1TS U1247 ( .A0(\destinationAddressbuffer[7][6] ), .A1(n712), .B0(
        \destinationAddressbuffer[5][6] ), .B1(n743), .Y(n701) );
  NAND4XLTS U1248 ( .A(n704), .B(n703), .C(n702), .D(n701), .Y(n705) );
  AOI22X1TS U1249 ( .A0(destinationAddressOut[6]), .A1(n706), .B0(n872), .B1(
        n705), .Y(n707) );
  AOI22X1TS U1250 ( .A0(destinationAddressIn_EAST[7]), .A1(n831), .B0(n710), 
        .B1(n735), .Y(n720) );
  AOI22X1TS U1251 ( .A0(destinationAddressIn_NORTH[7]), .A1(n738), .B0(n711), 
        .B1(n770), .Y(n719) );
  CLKBUFX2TS U1252 ( .A(n773), .Y(n764) );
  AOI22X1TS U1253 ( .A0(\destinationAddressbuffer[2][7] ), .A1(n724), .B0(
        \destinationAddressbuffer[0][7] ), .B1(n740), .Y(n716) );
  AOI22X1TS U1254 ( .A0(\destinationAddressbuffer[6][7] ), .A1(n725), .B0(
        \destinationAddressbuffer[4][7] ), .B1(n741), .Y(n715) );
  AOI22X1TS U1255 ( .A0(\destinationAddressbuffer[3][7] ), .A1(n726), .B0(
        \destinationAddressbuffer[1][7] ), .B1(n742), .Y(n714) );
  AOI22X1TS U1256 ( .A0(\destinationAddressbuffer[7][7] ), .A1(n712), .B0(
        \destinationAddressbuffer[5][7] ), .B1(n743), .Y(n713) );
  NAND4XLTS U1257 ( .A(n716), .B(n715), .C(n714), .D(n713), .Y(n717) );
  AOI22X1TS U1258 ( .A0(destinationAddressOut[7]), .A1(n527), .B0(n764), .B1(
        n717), .Y(n718) );
  AOI22X1TS U1259 ( .A0(destinationAddressIn_EAST[8]), .A1(n754), .B0(n721), 
        .B1(n735), .Y(n734) );
  AOI22X1TS U1260 ( .A0(n723), .A1(n738), .B0(n722), .B1(n755), .Y(n733) );
  CLKBUFX2TS U1261 ( .A(n724), .Y(n815) );
  AOI22X1TS U1262 ( .A0(\destinationAddressbuffer[2][8] ), .A1(n815), .B0(
        \destinationAddressbuffer[0][8] ), .B1(n740), .Y(n730) );
  CLKBUFX2TS U1263 ( .A(n725), .Y(n817) );
  AOI22X1TS U1264 ( .A0(\destinationAddressbuffer[6][8] ), .A1(n817), .B0(
        \destinationAddressbuffer[4][8] ), .B1(n741), .Y(n729) );
  CLKBUFX2TS U1265 ( .A(n726), .Y(n819) );
  AOI22X1TS U1266 ( .A0(\destinationAddressbuffer[3][8] ), .A1(n819), .B0(
        \destinationAddressbuffer[1][8] ), .B1(n742), .Y(n728) );
  AOI22X1TS U1267 ( .A0(\destinationAddressbuffer[7][8] ), .A1(n820), .B0(
        \destinationAddressbuffer[5][8] ), .B1(n743), .Y(n727) );
  NAND4XLTS U1268 ( .A(n730), .B(n729), .C(n728), .D(n727), .Y(n731) );
  AOI22X1TS U1269 ( .A0(destinationAddressOut[8]), .A1(n873), .B0(n764), .B1(
        n731), .Y(n732) );
  AOI22X1TS U1270 ( .A0(destinationAddressIn_EAST[9]), .A1(n769), .B0(n736), 
        .B1(n735), .Y(n752) );
  AOI22X1TS U1271 ( .A0(n739), .A1(n738), .B0(n737), .B1(n770), .Y(n751) );
  AOI22X1TS U1272 ( .A0(\destinationAddressbuffer[2][9] ), .A1(n815), .B0(
        \destinationAddressbuffer[0][9] ), .B1(n740), .Y(n747) );
  AOI22X1TS U1273 ( .A0(\destinationAddressbuffer[6][9] ), .A1(n817), .B0(
        \destinationAddressbuffer[4][9] ), .B1(n741), .Y(n746) );
  AOI22X1TS U1274 ( .A0(\destinationAddressbuffer[3][9] ), .A1(n819), .B0(
        \destinationAddressbuffer[1][9] ), .B1(n742), .Y(n745) );
  AOI22X1TS U1275 ( .A0(\destinationAddressbuffer[7][9] ), .A1(n820), .B0(
        \destinationAddressbuffer[5][9] ), .B1(n743), .Y(n744) );
  NAND4XLTS U1276 ( .A(n747), .B(n746), .C(n745), .D(n744), .Y(n748) );
  AOI22X1TS U1277 ( .A0(destinationAddressOut[9]), .A1(n749), .B0(n764), .B1(
        n748), .Y(n750) );
  CLKBUFX2TS U1278 ( .A(n812), .Y(n793) );
  AOI22X1TS U1279 ( .A0(destinationAddressIn_EAST[10]), .A1(n754), .B0(n753), 
        .B1(n793), .Y(n767) );
  CLKBUFX2TS U1280 ( .A(n696), .Y(n792) );
  AOI22X1TS U1281 ( .A0(n757), .A1(n792), .B0(n756), .B1(n755), .Y(n766) );
  CLKBUFX2TS U1282 ( .A(n815), .Y(n795) );
  CLKBUFX2TS U1283 ( .A(n814), .Y(n796) );
  AOI22X1TS U1284 ( .A0(\destinationAddressbuffer[2][10] ), .A1(n795), .B0(
        \destinationAddressbuffer[0][10] ), .B1(n796), .Y(n762) );
  CLKBUFX2TS U1285 ( .A(n817), .Y(n797) );
  CLKBUFX2TS U1286 ( .A(n816), .Y(n798) );
  AOI22X1TS U1287 ( .A0(\destinationAddressbuffer[6][10] ), .A1(n797), .B0(
        \destinationAddressbuffer[4][10] ), .B1(n798), .Y(n761) );
  CLKBUFX2TS U1288 ( .A(n819), .Y(n799) );
  CLKBUFX2TS U1289 ( .A(n818), .Y(n800) );
  AOI22X1TS U1290 ( .A0(\destinationAddressbuffer[3][10] ), .A1(n799), .B0(
        \destinationAddressbuffer[1][10] ), .B1(n800), .Y(n760) );
  CLKBUFX2TS U1291 ( .A(n832), .Y(n802) );
  AOI22X1TS U1292 ( .A0(\destinationAddressbuffer[7][10] ), .A1(n758), .B0(
        \destinationAddressbuffer[5][10] ), .B1(n802), .Y(n759) );
  NAND4XLTS U1293 ( .A(n762), .B(n761), .C(n760), .D(n759), .Y(n763) );
  AOI22X1TS U1294 ( .A0(destinationAddressOut[10]), .A1(n873), .B0(n764), .B1(
        n763), .Y(n765) );
  AOI22X1TS U1295 ( .A0(destinationAddressIn_EAST[11]), .A1(n769), .B0(n768), 
        .B1(n793), .Y(n781) );
  AOI22X1TS U1296 ( .A0(n772), .A1(n792), .B0(n771), .B1(n770), .Y(n780) );
  CLKBUFX2TS U1297 ( .A(n773), .Y(n826) );
  AOI22X1TS U1298 ( .A0(\destinationAddressbuffer[2][11] ), .A1(n795), .B0(
        \destinationAddressbuffer[0][11] ), .B1(n796), .Y(n777) );
  AOI22X1TS U1299 ( .A0(\destinationAddressbuffer[6][11] ), .A1(n797), .B0(
        \destinationAddressbuffer[4][11] ), .B1(n798), .Y(n776) );
  AOI22X1TS U1300 ( .A0(\destinationAddressbuffer[3][11] ), .A1(n799), .B0(
        \destinationAddressbuffer[1][11] ), .B1(n800), .Y(n775) );
  AOI22X1TS U1301 ( .A0(\destinationAddressbuffer[7][11] ), .A1(n801), .B0(
        \destinationAddressbuffer[5][11] ), .B1(n802), .Y(n774) );
  NAND4XLTS U1302 ( .A(n777), .B(n776), .C(n775), .D(n774), .Y(n778) );
  AOI22X1TS U1303 ( .A0(destinationAddressOut[11]), .A1(n527), .B0(n826), .B1(
        n778), .Y(n779) );
  CLKBUFX2TS U1304 ( .A(dataIn_NORTH[0]), .Y(n1089) );
  CLKBUFX2TS U1305 ( .A(dataIn_EAST[0]), .Y(n1472) );
  CLKBUFX2TS U1306 ( .A(n1472), .Y(n1348) );
  CLKBUFX2TS U1307 ( .A(n782), .Y(n855) );
  AOI22X1TS U1308 ( .A0(n1089), .A1(n792), .B0(n1348), .B1(n855), .Y(n791) );
  CLKBUFX2TS U1309 ( .A(dataIn_WEST[0]), .Y(n1521) );
  CLKBUFX2TS U1310 ( .A(n1521), .Y(n1410) );
  AOI22X1TS U1311 ( .A0(dataIn_SOUTH[0]), .A1(n794), .B0(n1410), .B1(n793), 
        .Y(n790) );
  AOI22X1TS U1312 ( .A0(\dataoutbuffer[0][0] ), .A1(n796), .B0(
        \dataoutbuffer[2][0] ), .B1(n795), .Y(n786) );
  AOI22X1TS U1313 ( .A0(\dataoutbuffer[4][0] ), .A1(n798), .B0(
        \dataoutbuffer[6][0] ), .B1(n797), .Y(n785) );
  AOI22X1TS U1314 ( .A0(\dataoutbuffer[1][0] ), .A1(n800), .B0(
        \dataoutbuffer[3][0] ), .B1(n799), .Y(n784) );
  AOI22X1TS U1315 ( .A0(\dataoutbuffer[5][0] ), .A1(n802), .B0(
        \dataoutbuffer[7][0] ), .B1(n865), .Y(n783) );
  NAND4XLTS U1316 ( .A(n786), .B(n785), .C(n784), .D(n783), .Y(n787) );
  AOI22X1TS U1317 ( .A0(dataOut[0]), .A1(n528), .B0(n826), .B1(n787), .Y(n789)
         );
  INVX2TS U1318 ( .A(cacheDataOut[0]), .Y(n1088) );
  INVX2TS U1319 ( .A(n565), .Y(n850) );
  NAND2X1TS U1320 ( .A(cacheDataOut[0]), .B(n850), .Y(n788) );
  CLKBUFX2TS U1321 ( .A(dataIn_NORTH[1]), .Y(n1095) );
  CLKBUFX2TS U1322 ( .A(dataIn_EAST[1]), .Y(n1480) );
  CLKBUFX2TS U1323 ( .A(n1480), .Y(n1353) );
  AOI22X1TS U1324 ( .A0(n1095), .A1(n792), .B0(n1353), .B1(n831), .Y(n811) );
  CLKBUFX2TS U1325 ( .A(dataIn_WEST[1]), .Y(n1531) );
  CLKBUFX2TS U1326 ( .A(n1531), .Y(n1415) );
  AOI22X1TS U1327 ( .A0(dataIn_SOUTH[1]), .A1(n794), .B0(n1415), .B1(n793), 
        .Y(n810) );
  AOI22X1TS U1328 ( .A0(\dataoutbuffer[0][1] ), .A1(n796), .B0(
        \dataoutbuffer[2][1] ), .B1(n795), .Y(n806) );
  AOI22X1TS U1329 ( .A0(\dataoutbuffer[4][1] ), .A1(n798), .B0(
        \dataoutbuffer[6][1] ), .B1(n797), .Y(n805) );
  AOI22X1TS U1330 ( .A0(\dataoutbuffer[1][1] ), .A1(n800), .B0(
        \dataoutbuffer[3][1] ), .B1(n799), .Y(n804) );
  AOI22X1TS U1331 ( .A0(\dataoutbuffer[5][1] ), .A1(n802), .B0(
        \dataoutbuffer[7][1] ), .B1(n801), .Y(n803) );
  NAND4XLTS U1332 ( .A(n806), .B(n805), .C(n804), .D(n803), .Y(n807) );
  AOI22X1TS U1333 ( .A0(dataOut[1]), .A1(n838), .B0(n826), .B1(n807), .Y(n809)
         );
  INVX2TS U1334 ( .A(cacheDataOut[1]), .Y(n1093) );
  INVX2TS U1335 ( .A(n565), .Y(n874) );
  NAND2X1TS U1336 ( .A(cacheDataOut[1]), .B(n874), .Y(n808) );
  CLKBUFX2TS U1337 ( .A(dataIn_NORTH[2]), .Y(n1102) );
  CLKBUFX2TS U1338 ( .A(n696), .Y(n856) );
  CLKBUFX2TS U1339 ( .A(dataIn_EAST[2]), .Y(n1489) );
  CLKBUFX2TS U1340 ( .A(n1489), .Y(n1360) );
  AOI22X1TS U1341 ( .A0(n1102), .A1(n856), .B0(n1360), .B1(n855), .Y(n830) );
  CLKBUFX2TS U1342 ( .A(dataIn_WEST[2]), .Y(n1539) );
  CLKBUFX2TS U1343 ( .A(n1539), .Y(n1423) );
  CLKBUFX2TS U1344 ( .A(n812), .Y(n857) );
  AOI22X1TS U1345 ( .A0(dataIn_SOUTH[2]), .A1(n813), .B0(n1423), .B1(n857), 
        .Y(n829) );
  CLKBUFX2TS U1346 ( .A(n814), .Y(n860) );
  CLKBUFX2TS U1347 ( .A(n815), .Y(n859) );
  AOI22X1TS U1348 ( .A0(\dataoutbuffer[0][2] ), .A1(n860), .B0(
        \dataoutbuffer[2][2] ), .B1(n859), .Y(n824) );
  CLKBUFX2TS U1349 ( .A(n816), .Y(n862) );
  CLKBUFX2TS U1350 ( .A(n817), .Y(n861) );
  AOI22X1TS U1351 ( .A0(\dataoutbuffer[4][2] ), .A1(n862), .B0(
        \dataoutbuffer[6][2] ), .B1(n861), .Y(n823) );
  CLKBUFX2TS U1352 ( .A(n818), .Y(n864) );
  CLKBUFX2TS U1353 ( .A(n819), .Y(n863) );
  AOI22X1TS U1354 ( .A0(\dataoutbuffer[1][2] ), .A1(n864), .B0(
        \dataoutbuffer[3][2] ), .B1(n863), .Y(n822) );
  AOI22X1TS U1355 ( .A0(\dataoutbuffer[5][2] ), .A1(n832), .B0(
        \dataoutbuffer[7][2] ), .B1(n820), .Y(n821) );
  NAND4XLTS U1356 ( .A(n824), .B(n823), .C(n822), .D(n821), .Y(n825) );
  AOI22X1TS U1357 ( .A0(dataOut[2]), .A1(n838), .B0(n826), .B1(n825), .Y(n828)
         );
  INVX2TS U1358 ( .A(cacheDataOut[2]), .Y(n1100) );
  NAND2X1TS U1359 ( .A(cacheDataOut[2]), .B(n850), .Y(n827) );
  CLKBUFX2TS U1360 ( .A(dataIn_NORTH[3]), .Y(n1108) );
  CLKBUFX2TS U1361 ( .A(dataIn_EAST[3]), .Y(n1497) );
  CLKBUFX2TS U1362 ( .A(n1497), .Y(n1367) );
  AOI22X1TS U1363 ( .A0(n1108), .A1(n856), .B0(n1367), .B1(n831), .Y(n842) );
  CLKBUFX2TS U1364 ( .A(dataIn_WEST[3]), .Y(n1546) );
  CLKBUFX2TS U1365 ( .A(n1546), .Y(n1428) );
  AOI22X1TS U1366 ( .A0(dataIn_SOUTH[3]), .A1(n858), .B0(n1428), .B1(n857), 
        .Y(n841) );
  AOI22X1TS U1367 ( .A0(\dataoutbuffer[0][3] ), .A1(n860), .B0(
        \dataoutbuffer[2][3] ), .B1(n859), .Y(n836) );
  AOI22X1TS U1368 ( .A0(\dataoutbuffer[4][3] ), .A1(n862), .B0(
        \dataoutbuffer[6][3] ), .B1(n861), .Y(n835) );
  AOI22X1TS U1369 ( .A0(\dataoutbuffer[1][3] ), .A1(n864), .B0(
        \dataoutbuffer[3][3] ), .B1(n863), .Y(n834) );
  AOI22X1TS U1370 ( .A0(\dataoutbuffer[5][3] ), .A1(n832), .B0(
        \dataoutbuffer[7][3] ), .B1(n843), .Y(n833) );
  NAND4XLTS U1371 ( .A(n836), .B(n835), .C(n834), .D(n833), .Y(n837) );
  AOI22X1TS U1372 ( .A0(dataOut[3]), .A1(n838), .B0(n849), .B1(n837), .Y(n840)
         );
  INVX2TS U1373 ( .A(cacheDataOut[3]), .Y(n1107) );
  NAND2X1TS U1374 ( .A(cacheDataOut[3]), .B(n874), .Y(n839) );
  CLKBUFX2TS U1375 ( .A(dataIn_NORTH[4]), .Y(n1338) );
  CLKBUFX2TS U1376 ( .A(dataIn_EAST[4]), .Y(n1505) );
  CLKBUFX2TS U1377 ( .A(n1505), .Y(n1372) );
  AOI22X1TS U1378 ( .A0(n1338), .A1(n856), .B0(n1372), .B1(n855), .Y(n854) );
  CLKBUFX2TS U1379 ( .A(dataIn_WEST[4]), .Y(n1555) );
  CLKBUFX2TS U1380 ( .A(n1555), .Y(n1432) );
  AOI22X1TS U1381 ( .A0(dataIn_SOUTH[4]), .A1(n858), .B0(n1432), .B1(n857), 
        .Y(n853) );
  AOI22X1TS U1382 ( .A0(\dataoutbuffer[0][4] ), .A1(n860), .B0(
        \dataoutbuffer[2][4] ), .B1(n859), .Y(n847) );
  AOI22X1TS U1383 ( .A0(\dataoutbuffer[4][4] ), .A1(n862), .B0(
        \dataoutbuffer[6][4] ), .B1(n861), .Y(n846) );
  AOI22X1TS U1384 ( .A0(\dataoutbuffer[1][4] ), .A1(n864), .B0(
        \dataoutbuffer[3][4] ), .B1(n863), .Y(n845) );
  AOI22X1TS U1385 ( .A0(\dataoutbuffer[5][4] ), .A1(n866), .B0(
        \dataoutbuffer[7][4] ), .B1(n843), .Y(n844) );
  NAND4XLTS U1386 ( .A(n847), .B(n846), .C(n845), .D(n844), .Y(n848) );
  AOI22X1TS U1387 ( .A0(dataOut[4]), .A1(n528), .B0(n849), .B1(n848), .Y(n852)
         );
  INVX2TS U1388 ( .A(cacheDataOut[4]), .Y(n1337) );
  NAND2X1TS U1389 ( .A(cacheDataOut[4]), .B(n850), .Y(n851) );
  CLKBUFX2TS U1390 ( .A(dataIn_NORTH[5]), .Y(n1344) );
  CLKBUFX2TS U1391 ( .A(dataIn_EAST[5]), .Y(n1513) );
  CLKBUFX2TS U1392 ( .A(n1513), .Y(n1377) );
  AOI22X1TS U1393 ( .A0(n1344), .A1(n856), .B0(n1377), .B1(n855), .Y(n878) );
  CLKBUFX2TS U1394 ( .A(dataIn_WEST[5]), .Y(n1565) );
  CLKBUFX2TS U1395 ( .A(n1565), .Y(n1437) );
  AOI22X1TS U1396 ( .A0(dataIn_SOUTH[5]), .A1(n858), .B0(n1437), .B1(n857), 
        .Y(n877) );
  AOI22X1TS U1397 ( .A0(\dataoutbuffer[0][5] ), .A1(n860), .B0(
        \dataoutbuffer[2][5] ), .B1(n859), .Y(n870) );
  AOI22X1TS U1398 ( .A0(\dataoutbuffer[4][5] ), .A1(n862), .B0(
        \dataoutbuffer[6][5] ), .B1(n861), .Y(n869) );
  AOI22X1TS U1399 ( .A0(\dataoutbuffer[1][5] ), .A1(n864), .B0(
        \dataoutbuffer[3][5] ), .B1(n863), .Y(n868) );
  AOI22X1TS U1400 ( .A0(\dataoutbuffer[5][5] ), .A1(n866), .B0(
        \dataoutbuffer[7][5] ), .B1(n865), .Y(n867) );
  NAND4XLTS U1401 ( .A(n870), .B(n869), .C(n868), .D(n867), .Y(n871) );
  AOI22X1TS U1402 ( .A0(dataOut[5]), .A1(n873), .B0(n872), .B1(n871), .Y(n876)
         );
  INVX2TS U1403 ( .A(cacheDataOut[5]), .Y(n1342) );
  NAND2X1TS U1404 ( .A(cacheDataOut[5]), .B(n874), .Y(n875) );
  INVX2TS U1405 ( .A(n959), .Y(n1790) );
  INVX2TS U1406 ( .A(n1582), .Y(n1681) );
  AOI22X1TS U1407 ( .A0(n1790), .A1(n1668), .B0(n1681), .B1(
        \requesterAddressbuffer[7][0] ), .Y(n884) );
  INVX2TS U1408 ( .A(n879), .Y(n1547) );
  INVX2TS U1409 ( .A(n893), .Y(n1554) );
  CLKBUFX2TS U1410 ( .A(n1037), .Y(n931) );
  AOI22X1TS U1411 ( .A0(n1547), .A1(n961), .B0(n1554), .B1(n931), .Y(n883) );
  INVX2TS U1412 ( .A(n880), .Y(n1568) );
  CLKBUFX2TS U1413 ( .A(n1040), .Y(n933) );
  INVX2TS U1414 ( .A(n881), .Y(n1692) );
  CLKBUFX2TS U1415 ( .A(n1008), .Y(n962) );
  AOI22X1TS U1416 ( .A0(n1568), .A1(n933), .B0(n1692), .B1(n962), .Y(n882) );
  INVX2TS U1417 ( .A(n892), .Y(n1675) );
  AOI22X1TS U1418 ( .A0(n1675), .A1(n1674), .B0(n1689), .B1(
        \requesterAddressbuffer[7][1] ), .Y(n887) );
  INVX2TS U1419 ( .A(n893), .Y(n1669) );
  CLKBUFX2TS U1420 ( .A(n1045), .Y(n939) );
  AOI22X1TS U1421 ( .A0(n1547), .A1(n969), .B0(n1669), .B1(n939), .Y(n886) );
  CLKBUFX2TS U1422 ( .A(n1046), .Y(n942) );
  CLKBUFX2TS U1423 ( .A(n1015), .Y(n971) );
  AOI22X1TS U1424 ( .A0(n1677), .A1(n942), .B0(n1524), .B1(n971), .Y(n885) );
  INVX2TS U1425 ( .A(n1582), .Y(n1529) );
  AOI22X1TS U1426 ( .A0(n36), .A1(n1682), .B0(n1529), .B1(
        \requesterAddressbuffer[7][2] ), .Y(n891) );
  CLKBUFX2TS U1427 ( .A(n1050), .Y(n946) );
  AOI22X1TS U1428 ( .A0(n44), .A1(n976), .B0(n1554), .B1(n946), .Y(n890) );
  CLKBUFX2TS U1429 ( .A(n1051), .Y(n948) );
  CLKBUFX2TS U1430 ( .A(n1023), .Y(n979) );
  AOI22X1TS U1431 ( .A0(n1568), .A1(n948), .B0(n888), .B1(n979), .Y(n889) );
  INVX2TS U1432 ( .A(n892), .Y(n1691) );
  AOI22X1TS U1433 ( .A0(n1691), .A1(n1690), .B0(n1529), .B1(
        \requesterAddressbuffer[7][3] ), .Y(n896) );
  CLKBUFX2TS U1434 ( .A(n1057), .Y(n953) );
  AOI22X1TS U1435 ( .A0(n1522), .A1(n984), .B0(n34), .B1(n953), .Y(n895) );
  CLKBUFX2TS U1436 ( .A(n1058), .Y(n955) );
  CLKBUFX2TS U1437 ( .A(n1032), .Y(n985) );
  AOI22X1TS U1438 ( .A0(n1685), .A1(n955), .B0(n1557), .B1(n985), .Y(n894) );
  INVX2TS U1439 ( .A(n959), .Y(n1846) );
  INVX2TS U1440 ( .A(n1487), .Y(n1711) );
  AOI22X1TS U1441 ( .A0(n1846), .A1(n900), .B0(n1711), .B1(
        \requesterAddressbuffer[6][0] ), .Y(n899) );
  INVX2TS U1442 ( .A(n1471), .Y(n1703) );
  AOI22X1TS U1443 ( .A0(n932), .A1(n1490), .B0(n931), .B1(n1703), .Y(n898) );
  AOI22X1TS U1444 ( .A0(n933), .A1(n1723), .B0(n962), .B1(n1707), .Y(n897) );
  INVX2TS U1445 ( .A(n966), .Y(n1767) );
  AOI22X1TS U1446 ( .A0(n1767), .A1(n900), .B0(n1719), .B1(
        \requesterAddressbuffer[6][1] ), .Y(n906) );
  INVX2TS U1447 ( .A(n901), .Y(n1721) );
  INVX2TS U1448 ( .A(n1471), .Y(n1712) );
  AOI22X1TS U1449 ( .A0(n940), .A1(n1721), .B0(n939), .B1(n1712), .Y(n905) );
  INVX2TS U1450 ( .A(n902), .Y(n1714) );
  AOI22X1TS U1451 ( .A0(n942), .A1(n1714), .B0(n971), .B1(n907), .Y(n904) );
  INVX2TS U1452 ( .A(n975), .Y(n1777) );
  INVX2TS U1453 ( .A(n1486), .Y(n1702) );
  INVX2TS U1454 ( .A(n1593), .Y(n1478) );
  AOI22X1TS U1455 ( .A0(n1777), .A1(n1702), .B0(n1478), .B1(
        \requesterAddressbuffer[6][2] ), .Y(n910) );
  AOI22X1TS U1456 ( .A0(n947), .A1(n112), .B0(n946), .B1(n911), .Y(n909) );
  AOI22X1TS U1457 ( .A0(n948), .A1(n1706), .B0(n979), .B1(n907), .Y(n908) );
  INVX2TS U1458 ( .A(n983), .Y(n1784) );
  AOI22X1TS U1459 ( .A0(n1784), .A1(n87), .B0(n1478), .B1(
        \requesterAddressbuffer[6][3] ), .Y(n914) );
  AOI22X1TS U1460 ( .A0(n954), .A1(n109), .B0(n953), .B1(n911), .Y(n913) );
  AOI22X1TS U1461 ( .A0(n955), .A1(n1499), .B0(n985), .B1(n1715), .Y(n912) );
  INVX2TS U1462 ( .A(n1453), .Y(n1743) );
  AOI22X1TS U1463 ( .A0(n1006), .A1(n919), .B0(n1743), .B1(
        \requesterAddressbuffer[5][0] ), .Y(n918) );
  INVX2TS U1464 ( .A(n1442), .Y(n1735) );
  AOI22X1TS U1465 ( .A0(n932), .A1(n1454), .B0(n931), .B1(n1735), .Y(n917) );
  INVX2TS U1466 ( .A(n915), .Y(n1738) );
  AOI22X1TS U1467 ( .A0(n933), .A1(n1738), .B0(requesterAddressIn_NORTH[0]), 
        .B1(n1449), .Y(n916) );
  AOI22X1TS U1468 ( .A0(n1674), .A1(n919), .B0(n1754), .B1(
        \requesterAddressbuffer[5][1] ), .Y(n922) );
  INVX2TS U1469 ( .A(n1442), .Y(n1746) );
  AOI22X1TS U1470 ( .A0(n940), .A1(n1748), .B0(n939), .B1(n1746), .Y(n921) );
  AOI22X1TS U1471 ( .A0(n942), .A1(n1749), .B0(requesterAddressIn_NORTH[1]), 
        .B1(n1750), .Y(n920) );
  INVX2TS U1472 ( .A(n13), .Y(n1733) );
  INVX2TS U1473 ( .A(n1606), .Y(n1448) );
  AOI22X1TS U1474 ( .A0(n1682), .A1(n1733), .B0(n1448), .B1(
        \requesterAddressbuffer[5][2] ), .Y(n925) );
  AOI22X1TS U1475 ( .A0(n947), .A1(n1458), .B0(n946), .B1(n927), .Y(n924) );
  AOI22X1TS U1476 ( .A0(n948), .A1(n1444), .B0(requesterAddressIn_NORTH[2]), 
        .B1(n1729), .Y(n923) );
  INVX2TS U1477 ( .A(n13), .Y(n1744) );
  AOI22X1TS U1478 ( .A0(n1690), .A1(n1744), .B0(n1448), .B1(
        \requesterAddressbuffer[5][3] ), .Y(n930) );
  INVX2TS U1479 ( .A(n926), .Y(n1748) );
  AOI22X1TS U1480 ( .A0(n954), .A1(n1748), .B0(n953), .B1(n927), .Y(n929) );
  AOI22X1TS U1481 ( .A0(n955), .A1(n228), .B0(requesterAddressIn_NORTH[3]), 
        .B1(n1739), .Y(n928) );
  INVX2TS U1482 ( .A(n1422), .Y(n1775) );
  AOI22X1TS U1483 ( .A0(n1006), .A1(n937), .B0(n1775), .B1(
        \requesterAddressbuffer[4][0] ), .Y(n936) );
  INVX2TS U1484 ( .A(n1409), .Y(n1768) );
  AOI22X1TS U1485 ( .A0(n932), .A1(n1761), .B0(n931), .B1(n1768), .Y(n935) );
  AOI22X1TS U1486 ( .A0(n933), .A1(n284), .B0(requesterAddressIn_NORTH[0]), 
        .B1(n300), .Y(n934) );
  INVX2TS U1487 ( .A(n966), .Y(n1898) );
  AOI22X1TS U1488 ( .A0(n1898), .A1(n937), .B0(n1783), .B1(
        \requesterAddressbuffer[4][1] ), .Y(n945) );
  INVX2TS U1489 ( .A(n1409), .Y(n1778) );
  AOI22X1TS U1490 ( .A0(n940), .A1(n303), .B0(n939), .B1(n1778), .Y(n944) );
  AOI22X1TS U1491 ( .A0(n942), .A1(n1786), .B0(requesterAddressIn_NORTH[1]), 
        .B1(n941), .Y(n943) );
  INVX2TS U1492 ( .A(n975), .Y(n1909) );
  INVX2TS U1493 ( .A(n1421), .Y(n1766) );
  INVX2TS U1494 ( .A(n1618), .Y(n1414) );
  AOI22X1TS U1495 ( .A0(n1909), .A1(n1766), .B0(n1414), .B1(
        \requesterAddressbuffer[4][2] ), .Y(n951) );
  AOI22X1TS U1496 ( .A0(n947), .A1(n1769), .B0(n946), .B1(n952), .Y(n950) );
  AOI22X1TS U1497 ( .A0(n948), .A1(n1438), .B0(requesterAddressIn_NORTH[2]), 
        .B1(n1762), .Y(n949) );
  INVX2TS U1498 ( .A(n983), .Y(n1921) );
  INVX2TS U1499 ( .A(n1421), .Y(n1776) );
  AOI22X1TS U1500 ( .A0(n1921), .A1(n1776), .B0(n1414), .B1(
        \requesterAddressbuffer[4][3] ), .Y(n958) );
  AOI22X1TS U1501 ( .A0(n954), .A1(n297), .B0(n953), .B1(n952), .Y(n957) );
  AOI22X1TS U1502 ( .A0(n955), .A1(n1424), .B0(requesterAddressIn_NORTH[3]), 
        .B1(n1770), .Y(n956) );
  INVX2TS U1503 ( .A(n959), .Y(n1889) );
  INVX2TS U1504 ( .A(n1391), .Y(n1804) );
  AOI22X1TS U1505 ( .A0(n1889), .A1(n967), .B0(n1804), .B1(
        \requesterAddressbuffer[3][0] ), .Y(n965) );
  INVX2TS U1506 ( .A(n960), .Y(n1799) );
  AOI22X1TS U1507 ( .A0(n961), .A1(n1799), .B0(n1007), .B1(n169), .Y(n964) );
  INVX2TS U1508 ( .A(n977), .Y(n1405) );
  AOI22X1TS U1509 ( .A0(n1009), .A1(n1405), .B0(n962), .B1(n1800), .Y(n963) );
  INVX2TS U1510 ( .A(n966), .Y(n1856) );
  AOI22X1TS U1511 ( .A0(n1856), .A1(n967), .B0(n1810), .B1(
        \requesterAddressbuffer[3][1] ), .Y(n974) );
  INVX2TS U1512 ( .A(n968), .Y(n1812) );
  AOI22X1TS U1513 ( .A0(n969), .A1(n136), .B0(n1014), .B1(n1812), .Y(n973) );
  AOI22X1TS U1514 ( .A0(n1016), .A1(n131), .B0(n971), .B1(n978), .Y(n972) );
  INVX2TS U1515 ( .A(n975), .Y(n1868) );
  INVX2TS U1516 ( .A(n1390), .Y(n1796) );
  INVX2TS U1517 ( .A(n1627), .Y(n1385) );
  AOI22X1TS U1518 ( .A0(n1868), .A1(n1796), .B0(n1385), .B1(
        \requesterAddressbuffer[3][2] ), .Y(n982) );
  AOI22X1TS U1519 ( .A0(n976), .A1(n1792), .B0(n1021), .B1(n1381), .Y(n981) );
  INVX2TS U1520 ( .A(n977), .Y(n1815) );
  AOI22X1TS U1521 ( .A0(n1024), .A1(n1815), .B0(n979), .B1(n978), .Y(n980) );
  INVX2TS U1522 ( .A(n983), .Y(n1880) );
  AOI22X1TS U1523 ( .A0(n1880), .A1(n132), .B0(n1385), .B1(
        \requesterAddressbuffer[3][3] ), .Y(n988) );
  AOI22X1TS U1524 ( .A0(n984), .A1(n1799), .B0(n1030), .B1(n1398), .Y(n987) );
  AOI22X1TS U1525 ( .A0(n1033), .A1(n1405), .B0(n985), .B1(n1806), .Y(n986) );
  INVX2TS U1526 ( .A(n1639), .Y(n1830) );
  AOI22X1TS U1527 ( .A0(n1790), .A1(n992), .B0(n1830), .B1(
        \requesterAddressbuffer[2][0] ), .Y(n991) );
  INVX2TS U1528 ( .A(n1359), .Y(n1824) );
  AOI22X1TS U1529 ( .A0(requesterAddressIn_WEST[0]), .A1(n1819), .B0(n1007), 
        .B1(n1824), .Y(n990) );
  AOI22X1TS U1530 ( .A0(n1009), .A1(n1841), .B0(n1008), .B1(n1835), .Y(n989)
         );
  AOI22X1TS U1531 ( .A0(n1898), .A1(n992), .B0(n1839), .B1(
        \requesterAddressbuffer[2][1] ), .Y(n995) );
  INVX2TS U1532 ( .A(n1359), .Y(n1832) );
  AOI22X1TS U1533 ( .A0(requesterAddressIn_WEST[1]), .A1(n1361), .B0(n1014), 
        .B1(n1832), .Y(n994) );
  INVX2TS U1534 ( .A(n199), .Y(n1834) );
  AOI22X1TS U1535 ( .A0(n1016), .A1(n1834), .B0(n1015), .B1(n1842), .Y(n993)
         );
  INVX2TS U1536 ( .A(n12), .Y(n1823) );
  INVX2TS U1537 ( .A(n1639), .Y(n1352) );
  AOI22X1TS U1538 ( .A0(n1909), .A1(n1823), .B0(n1352), .B1(
        \requesterAddressbuffer[2][2] ), .Y(n1000) );
  AOI22X1TS U1539 ( .A0(requesterAddressIn_WEST[2]), .A1(n1825), .B0(n1021), 
        .B1(n1002), .Y(n999) );
  INVX2TS U1540 ( .A(n996), .Y(n1362) );
  AOI22X1TS U1541 ( .A0(n1024), .A1(n1362), .B0(n1023), .B1(n997), .Y(n998) );
  INVX2TS U1542 ( .A(n12), .Y(n1831) );
  AOI22X1TS U1543 ( .A0(n1921), .A1(n1831), .B0(n1352), .B1(
        \requesterAddressbuffer[2][3] ), .Y(n1005) );
  INVX2TS U1544 ( .A(n1001), .Y(n1361) );
  AOI22X1TS U1545 ( .A0(requesterAddressIn_WEST[3]), .A1(n1361), .B0(n1030), 
        .B1(n1002), .Y(n1004) );
  AOI22X1TS U1546 ( .A0(n1033), .A1(n187), .B0(n1032), .B1(n1826), .Y(n1003)
         );
  INVX2TS U1547 ( .A(n1020), .Y(n1866) );
  AOI22X1TS U1548 ( .A0(n1006), .A1(n1013), .B0(n1866), .B1(
        \requesterAddressbuffer[1][0] ), .Y(n1012) );
  INVX2TS U1549 ( .A(n4), .Y(n1858) );
  AOI22X1TS U1550 ( .A0(requesterAddressIn_WEST[0]), .A1(n1848), .B0(n1007), 
        .B1(n1858), .Y(n1011) );
  AOI22X1TS U1551 ( .A0(n1009), .A1(n1883), .B0(n1008), .B1(n1862), .Y(n1010)
         );
  AOI22X1TS U1552 ( .A0(n1767), .A1(n1013), .B0(n1879), .B1(
        \requesterAddressbuffer[1][1] ), .Y(n1019) );
  INVX2TS U1553 ( .A(n4), .Y(n1870) );
  AOI22X1TS U1554 ( .A0(requesterAddressIn_WEST[1]), .A1(n1101), .B0(n1014), 
        .B1(n1870), .Y(n1018) );
  INVX2TS U1555 ( .A(n1031), .Y(n1873) );
  AOI22X1TS U1556 ( .A0(n1016), .A1(n1873), .B0(n1015), .B1(n1022), .Y(n1017)
         );
  INVX2TS U1557 ( .A(n1099), .Y(n1855) );
  INVX2TS U1558 ( .A(n1020), .Y(n1094) );
  AOI22X1TS U1559 ( .A0(n1777), .A1(n1855), .B0(n1094), .B1(
        \requesterAddressbuffer[1][2] ), .Y(n1027) );
  AOI22X1TS U1560 ( .A0(requesterAddressIn_WEST[2]), .A1(n1859), .B0(n1021), 
        .B1(n1029), .Y(n1026) );
  AOI22X1TS U1561 ( .A0(n1024), .A1(n335), .B0(n1023), .B1(n1022), .Y(n1025)
         );
  INVX2TS U1562 ( .A(n1099), .Y(n1867) );
  AOI22X1TS U1563 ( .A0(n1784), .A1(n1867), .B0(n1094), .B1(
        \requesterAddressbuffer[1][3] ), .Y(n1036) );
  INVX2TS U1564 ( .A(n1028), .Y(n1101) );
  AOI22X1TS U1565 ( .A0(requesterAddressIn_WEST[3]), .A1(n1101), .B0(n1030), 
        .B1(n1029), .Y(n1035) );
  INVX2TS U1566 ( .A(n1031), .Y(n1103) );
  AOI22X1TS U1567 ( .A0(n1033), .A1(n1103), .B0(n1032), .B1(n1875), .Y(n1034)
         );
  INVX2TS U1568 ( .A(n1071), .Y(n1907) );
  AOI22X1TS U1569 ( .A0(readRequesterAddress[0]), .A1(n1044), .B0(n1907), .B1(
        \requesterAddressbuffer[0][0] ), .Y(n1043) );
  INVX2TS U1570 ( .A(n1072), .Y(n1899) );
  AOI22X1TS U1571 ( .A0(requesterAddressIn_WEST[0]), .A1(n1890), .B0(n1037), 
        .B1(n1899), .Y(n1042) );
  INVX2TS U1572 ( .A(n1038), .Y(n1924) );
  INVX2TS U1573 ( .A(n1039), .Y(n1080) );
  AOI22X1TS U1574 ( .A0(n1040), .A1(n1924), .B0(requesterAddressIn_NORTH[0]), 
        .B1(n1080), .Y(n1041) );
  AOI22X1TS U1575 ( .A0(n1856), .A1(n1044), .B0(n1919), .B1(
        \requesterAddressbuffer[0][1] ), .Y(n1049) );
  INVX2TS U1576 ( .A(n1072), .Y(n1910) );
  AOI22X1TS U1577 ( .A0(requesterAddressIn_WEST[1]), .A1(n1073), .B0(n1045), 
        .B1(n1910), .Y(n1048) );
  AOI22X1TS U1578 ( .A0(n1046), .A1(n1067), .B0(requesterAddressIn_NORTH[1]), 
        .B1(n1080), .Y(n1047) );
  INVX2TS U1579 ( .A(n14), .Y(n1897) );
  INVX2TS U1580 ( .A(n1071), .Y(n1066) );
  AOI22X1TS U1581 ( .A0(n1868), .A1(n1897), .B0(n1066), .B1(
        \requesterAddressbuffer[0][2] ), .Y(n1054) );
  AOI22X1TS U1582 ( .A0(requesterAddressIn_WEST[2]), .A1(n1900), .B0(n1050), 
        .B1(n1056), .Y(n1053) );
  AOI22X1TS U1583 ( .A0(n1051), .A1(n1893), .B0(requesterAddressIn_NORTH[2]), 
        .B1(n1902), .Y(n1052) );
  INVX2TS U1584 ( .A(n14), .Y(n1908) );
  AOI22X1TS U1585 ( .A0(n1880), .A1(n1908), .B0(n1066), .B1(
        \requesterAddressbuffer[0][3] ), .Y(n1061) );
  INVX2TS U1586 ( .A(n1055), .Y(n1073) );
  AOI22X1TS U1587 ( .A0(requesterAddressIn_WEST[3]), .A1(n1073), .B0(n1057), 
        .B1(n1056), .Y(n1060) );
  AOI22X1TS U1588 ( .A0(n1058), .A1(n1915), .B0(requesterAddressIn_NORTH[3]), 
        .B1(n1062), .Y(n1059) );
  INVX2TS U1589 ( .A(n1088), .Y(n1470) );
  AOI22X1TS U1590 ( .A0(n1897), .A1(n1470), .B0(n1066), .B1(
        \dataoutbuffer[0][0] ), .Y(n1065) );
  AOI22X1TS U1591 ( .A0(n1073), .A1(n1410), .B0(n1899), .B1(n1348), .Y(n1064)
         );
  CLKBUFX2TS U1592 ( .A(n1089), .Y(n1474) );
  AOI22X1TS U1593 ( .A0(n1924), .A1(dataIn_SOUTH[0]), .B0(n1062), .B1(n1474), 
        .Y(n1063) );
  INVX2TS U1594 ( .A(n1093), .Y(n1479) );
  AOI22X1TS U1595 ( .A0(n1908), .A1(n1479), .B0(n1066), .B1(
        \dataoutbuffer[0][1] ), .Y(n1070) );
  AOI22X1TS U1596 ( .A0(n400), .A1(n1415), .B0(n1910), .B1(n1353), .Y(n1069)
         );
  CLKBUFX2TS U1597 ( .A(n1095), .Y(n1482) );
  AOI22X1TS U1598 ( .A0(n1067), .A1(dataIn_SOUTH[1]), .B0(n405), .B1(n1482), 
        .Y(n1068) );
  INVX2TS U1599 ( .A(n14), .Y(n1920) );
  INVX2TS U1600 ( .A(n1100), .Y(n1488) );
  INVX2TS U1601 ( .A(n1071), .Y(n1084) );
  AOI22X1TS U1602 ( .A0(n1920), .A1(n1488), .B0(n1084), .B1(
        \dataoutbuffer[0][2] ), .Y(n1076) );
  AOI22X1TS U1603 ( .A0(n1073), .A1(n1423), .B0(n398), .B1(n1360), .Y(n1075)
         );
  CLKBUFX2TS U1604 ( .A(n1102), .Y(n1492) );
  AOI22X1TS U1605 ( .A0(n1924), .A1(dataIn_SOUTH[2]), .B0(n1080), .B1(n1492), 
        .Y(n1074) );
  INVX2TS U1606 ( .A(n1107), .Y(n1496) );
  AOI22X1TS U1607 ( .A0(n1897), .A1(n1496), .B0(n1084), .B1(
        \dataoutbuffer[0][3] ), .Y(n1079) );
  AOI22X1TS U1608 ( .A0(n1911), .A1(n1428), .B0(n1899), .B1(n1367), .Y(n1078)
         );
  CLKBUFX2TS U1609 ( .A(n1108), .Y(n1500) );
  AOI22X1TS U1610 ( .A0(n439), .A1(dataIn_SOUTH[3]), .B0(n1913), .B1(n1500), 
        .Y(n1077) );
  INVX2TS U1611 ( .A(n1337), .Y(n1504) );
  AOI22X1TS U1612 ( .A0(n1908), .A1(n1504), .B0(n1084), .B1(
        \dataoutbuffer[0][4] ), .Y(n1083) );
  AOI22X1TS U1613 ( .A0(n1890), .A1(n1432), .B0(n1910), .B1(n1372), .Y(n1082)
         );
  CLKBUFX2TS U1614 ( .A(n1338), .Y(n1507) );
  AOI22X1TS U1615 ( .A0(n1915), .A1(dataIn_SOUTH[4]), .B0(n1080), .B1(n1507), 
        .Y(n1081) );
  INVX2TS U1616 ( .A(n1342), .Y(n1512) );
  AOI22X1TS U1617 ( .A0(n1920), .A1(n1512), .B0(n1084), .B1(
        \dataoutbuffer[0][5] ), .Y(n1087) );
  AOI22X1TS U1618 ( .A0(n400), .A1(n1437), .B0(n398), .B1(n1377), .Y(n1086) );
  CLKBUFX2TS U1619 ( .A(n1344), .Y(n1516) );
  AOI22X1TS U1620 ( .A0(n1893), .A1(dataIn_SOUTH[5]), .B0(n405), .B1(n1516), 
        .Y(n1085) );
  INVX2TS U1621 ( .A(n1088), .Y(n1520) );
  AOI22X1TS U1622 ( .A0(n1855), .A1(n1520), .B0(n1094), .B1(
        \dataoutbuffer[1][0] ), .Y(n1092) );
  AOI22X1TS U1623 ( .A0(n1101), .A1(dataIn_WEST[0]), .B0(n1858), .B1(n1348), 
        .Y(n1091) );
  CLKBUFX2TS U1624 ( .A(n1089), .Y(n1523) );
  CLKBUFX2TS U1625 ( .A(dataIn_SOUTH[0]), .Y(n1525) );
  CLKBUFX2TS U1626 ( .A(n1525), .Y(n1473) );
  AOI22X1TS U1627 ( .A0(n1022), .A1(n1523), .B0(n1109), .B1(n1473), .Y(n1090)
         );
  INVX2TS U1628 ( .A(n1093), .Y(n1530) );
  AOI22X1TS U1629 ( .A0(n1867), .A1(n1530), .B0(n1094), .B1(
        \dataoutbuffer[1][1] ), .Y(n1098) );
  AOI22X1TS U1630 ( .A0(n340), .A1(dataIn_WEST[1]), .B0(n1870), .B1(n1353), 
        .Y(n1097) );
  CLKBUFX2TS U1631 ( .A(n1095), .Y(n1532) );
  CLKBUFX2TS U1632 ( .A(dataIn_SOUTH[1]), .Y(n1533) );
  CLKBUFX2TS U1633 ( .A(n1533), .Y(n1481) );
  AOI22X1TS U1634 ( .A0(n1885), .A1(n1532), .B0(n1103), .B1(n1481), .Y(n1096)
         );
  INVX2TS U1635 ( .A(n1100), .Y(n1538) );
  INVX2TS U1636 ( .A(n1020), .Y(n1343) );
  AOI22X1TS U1637 ( .A0(n320), .A1(n1538), .B0(n1343), .B1(
        \dataoutbuffer[1][2] ), .Y(n1106) );
  AOI22X1TS U1638 ( .A0(n1101), .A1(dataIn_WEST[2]), .B0(n318), .B1(n1360), 
        .Y(n1105) );
  CLKBUFX2TS U1639 ( .A(n1102), .Y(n1540) );
  CLKBUFX2TS U1640 ( .A(dataIn_SOUTH[2]), .Y(n1541) );
  CLKBUFX2TS U1641 ( .A(n1541), .Y(n1491) );
  AOI22X1TS U1642 ( .A0(n333), .A1(n1540), .B0(n1103), .B1(n1491), .Y(n1104)
         );
  INVX2TS U1643 ( .A(n1107), .Y(n1545) );
  AOI22X1TS U1644 ( .A0(n1855), .A1(n1545), .B0(n1343), .B1(
        \dataoutbuffer[1][3] ), .Y(n1112) );
  AOI22X1TS U1645 ( .A0(n1871), .A1(dataIn_WEST[3]), .B0(n1858), .B1(n1367), 
        .Y(n1111) );
  CLKBUFX2TS U1646 ( .A(n1108), .Y(n1548) );
  CLKBUFX2TS U1647 ( .A(dataIn_SOUTH[3]), .Y(n1549) );
  CLKBUFX2TS U1648 ( .A(n1549), .Y(n1498) );
  AOI22X1TS U1649 ( .A0(n1875), .A1(n1548), .B0(n1109), .B1(n1498), .Y(n1110)
         );
  INVX2TS U1650 ( .A(n1337), .Y(n1553) );
  AOI22X1TS U1651 ( .A0(n1867), .A1(n1553), .B0(n1343), .B1(
        \dataoutbuffer[1][4] ), .Y(n1341) );
  AOI22X1TS U1652 ( .A0(n1848), .A1(dataIn_WEST[4]), .B0(n1870), .B1(n1372), 
        .Y(n1340) );
  CLKBUFX2TS U1653 ( .A(n1338), .Y(n1556) );
  CLKBUFX2TS U1654 ( .A(dataIn_SOUTH[4]), .Y(n1558) );
  CLKBUFX2TS U1655 ( .A(n1558), .Y(n1506) );
  AOI22X1TS U1656 ( .A0(n1851), .A1(n1556), .B0(n335), .B1(n1506), .Y(n1339)
         );
  INVX2TS U1657 ( .A(n1342), .Y(n1564) );
  AOI22X1TS U1658 ( .A0(n1013), .A1(n1564), .B0(n1343), .B1(
        \dataoutbuffer[1][5] ), .Y(n1347) );
  AOI22X1TS U1659 ( .A0(n340), .A1(dataIn_WEST[5]), .B0(n318), .B1(n1377), .Y(
        n1346) );
  CLKBUFX2TS U1660 ( .A(n1344), .Y(n1566) );
  CLKBUFX2TS U1661 ( .A(dataIn_SOUTH[5]), .Y(n1567) );
  CLKBUFX2TS U1662 ( .A(n1567), .Y(n1514) );
  AOI22X1TS U1663 ( .A0(n1885), .A1(n1566), .B0(n369), .B1(n1514), .Y(n1345)
         );
  AOI22X1TS U1664 ( .A0(n1823), .A1(n1470), .B0(n1352), .B1(
        \dataoutbuffer[2][0] ), .Y(n1351) );
  AOI22X1TS U1665 ( .A0(n1361), .A1(dataIn_WEST[0]), .B0(n1824), .B1(n1348), 
        .Y(n1350) );
  AOI22X1TS U1666 ( .A0(n1363), .A1(n1523), .B0(n1368), .B1(dataIn_SOUTH[0]), 
        .Y(n1349) );
  AOI22X1TS U1667 ( .A0(n1831), .A1(n1479), .B0(n1352), .B1(
        \dataoutbuffer[2][1] ), .Y(n1357) );
  AOI22X1TS U1668 ( .A0(n190), .A1(dataIn_WEST[1]), .B0(n1832), .B1(n1353), 
        .Y(n1356) );
  INVX2TS U1669 ( .A(n1354), .Y(n1842) );
  AOI22X1TS U1670 ( .A0(n1842), .A1(n1532), .B0(n1362), .B1(dataIn_SOUTH[1]), 
        .Y(n1355) );
  INVX2TS U1671 ( .A(n12), .Y(n1840) );
  INVX2TS U1672 ( .A(n1358), .Y(n1376) );
  AOI22X1TS U1673 ( .A0(n1840), .A1(n1488), .B0(n1376), .B1(
        \dataoutbuffer[2][2] ), .Y(n1366) );
  AOI22X1TS U1674 ( .A0(n1361), .A1(dataIn_WEST[2]), .B0(n1), .B1(n1360), .Y(
        n1365) );
  AOI22X1TS U1675 ( .A0(n1363), .A1(n1540), .B0(n1362), .B1(dataIn_SOUTH[2]), 
        .Y(n1364) );
  AOI22X1TS U1676 ( .A0(n1823), .A1(n1496), .B0(n1376), .B1(
        \dataoutbuffer[2][3] ), .Y(n1371) );
  AOI22X1TS U1677 ( .A0(n1833), .A1(dataIn_WEST[3]), .B0(n1824), .B1(n1367), 
        .Y(n1370) );
  AOI22X1TS U1678 ( .A0(n997), .A1(n1548), .B0(n1368), .B1(dataIn_SOUTH[3]), 
        .Y(n1369) );
  AOI22X1TS U1679 ( .A0(n1831), .A1(n1504), .B0(n1376), .B1(
        \dataoutbuffer[2][4] ), .Y(n1375) );
  AOI22X1TS U1680 ( .A0(n1819), .A1(dataIn_WEST[4]), .B0(n1832), .B1(n1372), 
        .Y(n1374) );
  AOI22X1TS U1681 ( .A0(n1826), .A1(n1556), .B0(n1834), .B1(dataIn_SOUTH[4]), 
        .Y(n1373) );
  AOI22X1TS U1682 ( .A0(n1840), .A1(n1512), .B0(n1376), .B1(
        \dataoutbuffer[2][5] ), .Y(n1380) );
  AOI22X1TS U1683 ( .A0(n190), .A1(dataIn_WEST[5]), .B0(n1), .B1(n1377), .Y(
        n1379) );
  AOI22X1TS U1684 ( .A0(n1842), .A1(n1566), .B0(n210), .B1(dataIn_SOUTH[5]), 
        .Y(n1378) );
  AOI22X1TS U1685 ( .A0(n1796), .A1(n1470), .B0(n1385), .B1(
        \dataoutbuffer[3][0] ), .Y(n1384) );
  AOI22X1TS U1686 ( .A0(n1399), .A1(dataIn_WEST[0]), .B0(n1381), .B1(
        dataIn_EAST[0]), .Y(n1383) );
  AOI22X1TS U1687 ( .A0(n159), .A1(n1474), .B0(n1386), .B1(n1473), .Y(n1382)
         );
  AOI22X1TS U1688 ( .A0(n132), .A1(n1479), .B0(n1385), .B1(
        \dataoutbuffer[3][1] ), .Y(n1389) );
  AOI22X1TS U1689 ( .A0(n1814), .A1(dataIn_WEST[1]), .B0(n1812), .B1(
        dataIn_EAST[1]), .Y(n1388) );
  AOI22X1TS U1690 ( .A0(n1400), .A1(n1482), .B0(n1386), .B1(n1481), .Y(n1387)
         );
  INVX2TS U1691 ( .A(n1390), .Y(n1811) );
  INVX2TS U1692 ( .A(n1391), .Y(n1404) );
  AOI22X1TS U1693 ( .A0(n1811), .A1(n1488), .B0(n1404), .B1(
        \dataoutbuffer[3][2] ), .Y(n1394) );
  AOI22X1TS U1694 ( .A0(n163), .A1(dataIn_WEST[2]), .B0(n169), .B1(
        dataIn_EAST[2]), .Y(n1393) );
  AOI22X1TS U1695 ( .A0(n159), .A1(n1492), .B0(n1405), .B1(n1491), .Y(n1392)
         );
  AOI22X1TS U1696 ( .A0(n1796), .A1(n1496), .B0(n1404), .B1(
        \dataoutbuffer[3][3] ), .Y(n1397) );
  AOI22X1TS U1697 ( .A0(n1799), .A1(dataIn_WEST[3]), .B0(n157), .B1(
        dataIn_EAST[3]), .Y(n1396) );
  AOI22X1TS U1698 ( .A0(n1806), .A1(n1500), .B0(n143), .B1(n1498), .Y(n1395)
         );
  AOI22X1TS U1699 ( .A0(n967), .A1(n1504), .B0(n1404), .B1(
        \dataoutbuffer[3][4] ), .Y(n1403) );
  AOI22X1TS U1700 ( .A0(n1399), .A1(dataIn_WEST[4]), .B0(n1398), .B1(
        dataIn_EAST[4]), .Y(n1402) );
  AOI22X1TS U1701 ( .A0(n1400), .A1(n1507), .B0(n1815), .B1(n1506), .Y(n1401)
         );
  AOI22X1TS U1702 ( .A0(n1811), .A1(n1512), .B0(n1404), .B1(
        \dataoutbuffer[3][5] ), .Y(n1408) );
  AOI22X1TS U1703 ( .A0(n149), .A1(dataIn_WEST[5]), .B0(n1812), .B1(
        dataIn_EAST[5]), .Y(n1407) );
  AOI22X1TS U1704 ( .A0(n159), .A1(n1516), .B0(n1405), .B1(n1514), .Y(n1406)
         );
  AOI22X1TS U1705 ( .A0(n1766), .A1(n1520), .B0(n1414), .B1(
        \dataoutbuffer[4][0] ), .Y(n1413) );
  AOI22X1TS U1706 ( .A0(n288), .A1(n1410), .B0(n952), .B1(dataIn_EAST[0]), .Y(
        n1412) );
  AOI22X1TS U1707 ( .A0(n1424), .A1(n1525), .B0(n281), .B1(n1523), .Y(n1411)
         );
  AOI22X1TS U1708 ( .A0(n1776), .A1(n1530), .B0(n1414), .B1(
        \dataoutbuffer[4][1] ), .Y(n1420) );
  AOI22X1TS U1709 ( .A0(n297), .A1(n1415), .B0(n1768), .B1(dataIn_EAST[1]), 
        .Y(n1419) );
  INVX2TS U1710 ( .A(n1416), .Y(n1771) );
  INVX2TS U1711 ( .A(n1417), .Y(n1785) );
  AOI22X1TS U1712 ( .A0(n1771), .A1(n1533), .B0(n1785), .B1(n1532), .Y(n1418)
         );
  INVX2TS U1713 ( .A(n1422), .Y(n1436) );
  AOI22X1TS U1714 ( .A0(n276), .A1(n1538), .B0(n1436), .B1(
        \dataoutbuffer[4][2] ), .Y(n1427) );
  AOI22X1TS U1715 ( .A0(n288), .A1(n1423), .B0(n1778), .B1(dataIn_EAST[2]), 
        .Y(n1426) );
  AOI22X1TS U1716 ( .A0(n1424), .A1(n1541), .B0(n281), .B1(n1540), .Y(n1425)
         );
  AOI22X1TS U1717 ( .A0(n1766), .A1(n1545), .B0(n1436), .B1(
        \dataoutbuffer[4][3] ), .Y(n1431) );
  AOI22X1TS U1718 ( .A0(n1779), .A1(n1428), .B0(n274), .B1(dataIn_EAST[3]), 
        .Y(n1430) );
  AOI22X1TS U1719 ( .A0(n1438), .A1(n1549), .B0(n1785), .B1(n1548), .Y(n1429)
         );
  AOI22X1TS U1720 ( .A0(n1776), .A1(n1553), .B0(n1436), .B1(
        \dataoutbuffer[4][4] ), .Y(n1435) );
  AOI22X1TS U1721 ( .A0(n1761), .A1(n1432), .B0(n1768), .B1(dataIn_EAST[4]), 
        .Y(n1434) );
  AOI22X1TS U1722 ( .A0(n1771), .A1(n1558), .B0(n1762), .B1(n1556), .Y(n1433)
         );
  AOI22X1TS U1723 ( .A0(n937), .A1(n1564), .B0(n1436), .B1(
        \dataoutbuffer[4][5] ), .Y(n1441) );
  AOI22X1TS U1724 ( .A0(n303), .A1(n1437), .B0(n1778), .B1(dataIn_EAST[5]), 
        .Y(n1440) );
  AOI22X1TS U1725 ( .A0(n1438), .A1(n1567), .B0(n1785), .B1(n1566), .Y(n1439)
         );
  AOI22X1TS U1726 ( .A0(n1733), .A1(n1520), .B0(n1448), .B1(
        \dataoutbuffer[5][0] ), .Y(n1447) );
  AOI22X1TS U1727 ( .A0(n1454), .A1(n1521), .B0(n927), .B1(n1472), .Y(n1446)
         );
  INVX2TS U1728 ( .A(n1443), .Y(n1739) );
  AOI22X1TS U1729 ( .A0(n1739), .A1(n1474), .B0(n1444), .B1(n1473), .Y(n1445)
         );
  AOI22X1TS U1730 ( .A0(n1744), .A1(n1530), .B0(n1448), .B1(
        \dataoutbuffer[5][1] ), .Y(n1452) );
  AOI22X1TS U1731 ( .A0(n260), .A1(n1531), .B0(n1735), .B1(n1480), .Y(n1451)
         );
  AOI22X1TS U1732 ( .A0(n1449), .A1(n1482), .B0(n263), .B1(n1481), .Y(n1450)
         );
  INVX2TS U1733 ( .A(n13), .Y(n1755) );
  INVX2TS U1734 ( .A(n1453), .Y(n1466) );
  AOI22X1TS U1735 ( .A0(n1755), .A1(n1538), .B0(n1466), .B1(
        \dataoutbuffer[5][2] ), .Y(n1457) );
  AOI22X1TS U1736 ( .A0(n1454), .A1(n1539), .B0(n1746), .B1(n1489), .Y(n1456)
         );
  AOI22X1TS U1737 ( .A0(n232), .A1(n1492), .B0(n1462), .B1(n1491), .Y(n1455)
         );
  AOI22X1TS U1738 ( .A0(n1733), .A1(n1545), .B0(n1466), .B1(
        \dataoutbuffer[5][3] ), .Y(n1461) );
  AOI22X1TS U1739 ( .A0(n1458), .A1(n1546), .B0(n222), .B1(n1497), .Y(n1460)
         );
  AOI22X1TS U1740 ( .A0(n1739), .A1(n1500), .B0(n1749), .B1(n1498), .Y(n1459)
         );
  AOI22X1TS U1741 ( .A0(n1744), .A1(n1553), .B0(n1466), .B1(
        \dataoutbuffer[5][4] ), .Y(n1465) );
  AOI22X1TS U1742 ( .A0(n1737), .A1(n1555), .B0(n1735), .B1(n1505), .Y(n1464)
         );
  AOI22X1TS U1743 ( .A0(n1750), .A1(n1507), .B0(n1462), .B1(n1506), .Y(n1463)
         );
  AOI22X1TS U1744 ( .A0(n1755), .A1(n1564), .B0(n1466), .B1(
        \dataoutbuffer[5][5] ), .Y(n1469) );
  AOI22X1TS U1745 ( .A0(n224), .A1(n1565), .B0(n1746), .B1(n1513), .Y(n1468)
         );
  AOI22X1TS U1746 ( .A0(n1729), .A1(n1516), .B0(n228), .B1(n1514), .Y(n1467)
         );
  AOI22X1TS U1747 ( .A0(n1702), .A1(n1470), .B0(n1478), .B1(
        \dataoutbuffer[6][0] ), .Y(n1477) );
  AOI22X1TS U1748 ( .A0(n1490), .A1(n1521), .B0(n911), .B1(n1472), .Y(n1476)
         );
  AOI22X1TS U1749 ( .A0(n92), .A1(n1474), .B0(n1499), .B1(n1473), .Y(n1475) );
  AOI22X1TS U1750 ( .A0(n87), .A1(n1479), .B0(n1478), .B1(
        \dataoutbuffer[6][1] ), .Y(n1485) );
  AOI22X1TS U1751 ( .A0(n1721), .A1(n1531), .B0(n1703), .B1(n1480), .Y(n1484)
         );
  AOI22X1TS U1752 ( .A0(n92), .A1(n1482), .B0(n94), .B1(n1481), .Y(n1483) );
  INVX2TS U1753 ( .A(n1486), .Y(n1720) );
  INVX2TS U1754 ( .A(n1487), .Y(n1511) );
  AOI22X1TS U1755 ( .A0(n1720), .A1(n1488), .B0(n1511), .B1(
        \dataoutbuffer[6][2] ), .Y(n1495) );
  AOI22X1TS U1756 ( .A0(n1490), .A1(n1539), .B0(n1712), .B1(n1489), .Y(n1494)
         );
  AOI22X1TS U1757 ( .A0(n92), .A1(n1492), .B0(n94), .B1(n1491), .Y(n1493) );
  AOI22X1TS U1758 ( .A0(n1702), .A1(n1496), .B0(n1511), .B1(
        \dataoutbuffer[6][3] ), .Y(n1503) );
  AOI22X1TS U1759 ( .A0(n109), .A1(n1546), .B0(n85), .B1(n1497), .Y(n1502) );
  AOI22X1TS U1760 ( .A0(n1715), .A1(n1500), .B0(n1499), .B1(n1498), .Y(n1501)
         );
  AOI22X1TS U1761 ( .A0(n900), .A1(n1504), .B0(n1511), .B1(
        \dataoutbuffer[6][4] ), .Y(n1510) );
  AOI22X1TS U1762 ( .A0(n1704), .A1(n1555), .B0(n1703), .B1(n1505), .Y(n1509)
         );
  AOI22X1TS U1763 ( .A0(n1698), .A1(n1507), .B0(n1515), .B1(n1506), .Y(n1508)
         );
  AOI22X1TS U1764 ( .A0(n1720), .A1(n1512), .B0(n1511), .B1(
        \dataoutbuffer[6][5] ), .Y(n1519) );
  AOI22X1TS U1765 ( .A0(n1721), .A1(n1565), .B0(n1712), .B1(n1513), .Y(n1518)
         );
  AOI22X1TS U1766 ( .A0(n104), .A1(n1516), .B0(n1515), .B1(n1514), .Y(n1517)
         );
  AOI22X1TS U1767 ( .A0(n1675), .A1(n1520), .B0(n1529), .B1(
        \dataoutbuffer[7][0] ), .Y(n1528) );
  AOI22X1TS U1768 ( .A0(n1522), .A1(n1521), .B0(n1669), .B1(dataIn_EAST[0]), 
        .Y(n1527) );
  AOI22X1TS U1769 ( .A0(n1559), .A1(n1525), .B0(n1524), .B1(n1523), .Y(n1526)
         );
  AOI22X1TS U1770 ( .A0(n36), .A1(n1530), .B0(n1529), .B1(
        \dataoutbuffer[7][1] ), .Y(n1536) );
  AOI22X1TS U1771 ( .A0(n1547), .A1(n1531), .B0(n1554), .B1(dataIn_EAST[1]), 
        .Y(n1535) );
  AOI22X1TS U1772 ( .A0(n1677), .A1(n1533), .B0(n1692), .B1(n1532), .Y(n1534)
         );
  INVX2TS U1773 ( .A(n1537), .Y(n1563) );
  AOI22X1TS U1774 ( .A0(n1691), .A1(n1538), .B0(n1563), .B1(
        \dataoutbuffer[7][2] ), .Y(n1544) );
  AOI22X1TS U1775 ( .A0(n1684), .A1(n1539), .B0(n1683), .B1(dataIn_EAST[2]), 
        .Y(n1543) );
  AOI22X1TS U1776 ( .A0(n1568), .A1(n1541), .B0(n46), .B1(n1540), .Y(n1542) );
  AOI22X1TS U1777 ( .A0(n1675), .A1(n1545), .B0(n1563), .B1(
        \dataoutbuffer[7][3] ), .Y(n1552) );
  AOI22X1TS U1778 ( .A0(n1547), .A1(n1546), .B0(n1669), .B1(dataIn_EAST[3]), 
        .Y(n1551) );
  AOI22X1TS U1779 ( .A0(n1693), .A1(n1549), .B0(n46), .B1(n1548), .Y(n1550) );
  AOI22X1TS U1780 ( .A0(n36), .A1(n1553), .B0(n1563), .B1(
        \dataoutbuffer[7][4] ), .Y(n1562) );
  AOI22X1TS U1781 ( .A0(n1670), .A1(n1555), .B0(n1554), .B1(dataIn_EAST[4]), 
        .Y(n1561) );
  AOI22X1TS U1782 ( .A0(n1559), .A1(n1558), .B0(n1557), .B1(n1556), .Y(n1560)
         );
  AOI22X1TS U1783 ( .A0(n1691), .A1(n1564), .B0(n1563), .B1(
        \dataoutbuffer[7][5] ), .Y(n1571) );
  AOI22X1TS U1784 ( .A0(n68), .A1(n1565), .B0(n34), .B1(dataIn_EAST[5]), .Y(
        n1570) );
  AOI22X1TS U1785 ( .A0(n1568), .A1(n1567), .B0(n1692), .B1(n1566), .Y(n1569)
         );
  CLKBUFX2TS U1786 ( .A(n1664), .Y(n1615) );
  INVX2TS U1787 ( .A(n1572), .Y(n1660) );
  AOI22X1TS U1788 ( .A0(n1574), .A1(n1597), .B0(n1596), .B1(n1573), .Y(n1576)
         );
  AOI22X1TS U1789 ( .A0(n1577), .A1(n1660), .B0(n1576), .B1(n1575), .Y(n1579)
         );
  AOI22X1TS U1790 ( .A0(n1580), .A1(n1615), .B0(n1579), .B1(n1578), .Y(n1583)
         );
  AOI32X1TS U1791 ( .A0(n1583), .A1(n1582), .A2(n1581), .B0(n1689), .B1(n1958), 
        .Y(n2085) );
  INVX2TS U1792 ( .A(n1572), .Y(n1633) );
  AOI22X1TS U1793 ( .A0(n1585), .A1(n1597), .B0(n1596), .B1(n1584), .Y(n1587)
         );
  AOI22X1TS U1794 ( .A0(n1588), .A1(n1633), .B0(n1587), .B1(n1586), .Y(n1590)
         );
  AOI22X1TS U1795 ( .A0(n1591), .A1(n1615), .B0(n1590), .B1(n1589), .Y(n1594)
         );
  AOI32X1TS U1796 ( .A0(n1594), .A1(n1593), .A2(n1592), .B0(n1719), .B1(n1959), 
        .Y(n2086) );
  AOI22X1TS U1797 ( .A0(n1598), .A1(n1597), .B0(n1596), .B1(n1595), .Y(n1600)
         );
  AOI22X1TS U1798 ( .A0(n1601), .A1(n1633), .B0(n1600), .B1(n1599), .Y(n1603)
         );
  AOI22X1TS U1799 ( .A0(n1604), .A1(n1615), .B0(n1603), .B1(n1602), .Y(n1607)
         );
  AOI32X1TS U1800 ( .A0(n1607), .A1(n1606), .A2(n1605), .B0(n1754), .B1(n1960), 
        .Y(n2087) );
  CLKBUFX2TS U1801 ( .A(n1656), .Y(n1643) );
  CLKBUFX2TS U1802 ( .A(n1655), .Y(n1642) );
  AOI22X1TS U1803 ( .A0(n1609), .A1(n1643), .B0(n1642), .B1(n1608), .Y(n1611)
         );
  AOI22X1TS U1804 ( .A0(n1612), .A1(n1660), .B0(n1611), .B1(n1610), .Y(n1614)
         );
  AOI22X1TS U1805 ( .A0(n1616), .A1(n1615), .B0(n1614), .B1(n1613), .Y(n1619)
         );
  AOI32X1TS U1806 ( .A0(n1619), .A1(n1618), .A2(n1617), .B0(n1783), .B1(n1961), 
        .Y(n2088) );
  AOI22X1TS U1807 ( .A0(n122), .A1(n1643), .B0(n1642), .B1(n28), .Y(n1621) );
  AOI22X1TS U1808 ( .A0(n1622), .A1(n1633), .B0(n1621), .B1(n1620), .Y(n1624)
         );
  AOI22X1TS U1809 ( .A0(n1625), .A1(n1664), .B0(n1624), .B1(n1623), .Y(n1628)
         );
  AOI32X1TS U1810 ( .A0(n1628), .A1(n1627), .A2(n1626), .B0(n1810), .B1(n1962), 
        .Y(n2089) );
  AOI22X1TS U1811 ( .A0(n1630), .A1(n1643), .B0(n1642), .B1(n1629), .Y(n1632)
         );
  AOI22X1TS U1812 ( .A0(n1634), .A1(n1633), .B0(n1632), .B1(n1631), .Y(n1636)
         );
  AOI22X1TS U1813 ( .A0(n1637), .A1(n1650), .B0(n1636), .B1(n1635), .Y(n1640)
         );
  AOI32X1TS U1814 ( .A0(n1640), .A1(n1639), .A2(n1638), .B0(n1839), .B1(n1963), 
        .Y(n2090) );
  AOI22X1TS U1815 ( .A0(n1644), .A1(n1643), .B0(n1642), .B1(n1641), .Y(n1646)
         );
  AOI22X1TS U1816 ( .A0(n1647), .A1(n1660), .B0(n1646), .B1(n1645), .Y(n1649)
         );
  AOI22X1TS U1817 ( .A0(n1651), .A1(n1650), .B0(n1649), .B1(n1648), .Y(n1653)
         );
  AOI32X1TS U1818 ( .A0(n1653), .A1(n359), .A2(n1652), .B0(n1879), .B1(n1964), 
        .Y(n2091) );
  AOI22X1TS U1819 ( .A0(n1657), .A1(n1656), .B0(n1655), .B1(n1654), .Y(n1659)
         );
  AOI22X1TS U1820 ( .A0(n1661), .A1(n1660), .B0(n1659), .B1(n1658), .Y(n1663)
         );
  AOI22X1TS U1821 ( .A0(n1665), .A1(n1664), .B0(n1663), .B1(n1662), .Y(n1667)
         );
  AOI32X1TS U1822 ( .A0(n1667), .A1(n429), .A2(n1666), .B0(n1919), .B1(n1965), 
        .Y(n2092) );
  AOI22X1TS U1823 ( .A0(n1846), .A1(n1668), .B0(n1681), .B1(
        \destinationAddressbuffer[7][0] ), .Y(n1673) );
  AOI22X1TS U1824 ( .A0(n1670), .A1(n1728), .B0(n1669), .B1(n1727), .Y(n1672)
         );
  CLKBUFX2TS U1825 ( .A(n1697), .Y(n1850) );
  AOI22X1TS U1826 ( .A0(n60), .A1(destinationAddressIn_SOUTH[0]), .B0(n1676), 
        .B1(n1850), .Y(n1671) );
  AOI22X1TS U1827 ( .A0(n1675), .A1(n1674), .B0(n1681), .B1(
        \destinationAddressbuffer[7][1] ), .Y(n1680) );
  AOI22X1TS U1828 ( .A0(n1684), .A1(n1736), .B0(n1683), .B1(n1734), .Y(n1679)
         );
  CLKBUFX2TS U1829 ( .A(n1705), .Y(n1861) );
  AOI22X1TS U1830 ( .A0(n1677), .A1(destinationAddressIn_SOUTH[1]), .B0(n1676), 
        .B1(n1861), .Y(n1678) );
  AOI22X1TS U1831 ( .A0(n1668), .A1(n1682), .B0(n1681), .B1(
        \destinationAddressbuffer[7][2] ), .Y(n1688) );
  AOI22X1TS U1832 ( .A0(n1684), .A1(n1747), .B0(n1683), .B1(n1745), .Y(n1687)
         );
  CLKBUFX2TS U1833 ( .A(n1713), .Y(n1874) );
  AOI22X1TS U1834 ( .A0(n1685), .A1(destinationAddressIn_SOUTH[2]), .B0(n888), 
        .B1(n1874), .Y(n1686) );
  AOI22X1TS U1835 ( .A0(n1691), .A1(n1690), .B0(n1689), .B1(
        \destinationAddressbuffer[7][3] ), .Y(n1696) );
  AOI22X1TS U1836 ( .A0(n44), .A1(n1757), .B0(n34), .B1(n1756), .Y(n1695) );
  CLKBUFX2TS U1837 ( .A(n1722), .Y(n1884) );
  AOI22X1TS U1838 ( .A0(n1693), .A1(destinationAddressIn_SOUTH[3]), .B0(n1692), 
        .B1(n1884), .Y(n1694) );
  AOI22X1TS U1839 ( .A0(n1889), .A1(n1720), .B0(n1711), .B1(
        \destinationAddressbuffer[6][0] ), .Y(n1701) );
  AOI22X1TS U1840 ( .A0(n89), .A1(n1728), .B0(n85), .B1(n1727), .Y(n1700) );
  CLKBUFX2TS U1841 ( .A(n1697), .Y(n1891) );
  CLKBUFX2TS U1842 ( .A(destinationAddressIn_SOUTH[0]), .Y(n1892) );
  CLKBUFX2TS U1843 ( .A(n1892), .Y(n1849) );
  AOI22X1TS U1844 ( .A0(n1698), .A1(n1891), .B0(n1714), .B1(n1849), .Y(n1699)
         );
  AOI22X1TS U1845 ( .A0(n1767), .A1(n1702), .B0(n1711), .B1(
        \destinationAddressbuffer[6][1] ), .Y(n1710) );
  AOI22X1TS U1846 ( .A0(n1704), .A1(n1736), .B0(n1703), .B1(n1734), .Y(n1709)
         );
  CLKBUFX2TS U1847 ( .A(n1705), .Y(n1901) );
  CLKBUFX2TS U1848 ( .A(destinationAddressIn_SOUTH[1]), .Y(n1903) );
  CLKBUFX2TS U1849 ( .A(n1903), .Y(n1860) );
  AOI22X1TS U1850 ( .A0(n1707), .A1(n1901), .B0(n1706), .B1(n1860), .Y(n1708)
         );
  AOI22X1TS U1851 ( .A0(n1777), .A1(n87), .B0(n1711), .B1(
        \destinationAddressbuffer[6][2] ), .Y(n1718) );
  AOI22X1TS U1852 ( .A0(n89), .A1(n1747), .B0(n1712), .B1(n1745), .Y(n1717) );
  CLKBUFX2TS U1853 ( .A(n1713), .Y(n1912) );
  CLKBUFX2TS U1854 ( .A(destinationAddressIn_SOUTH[2]), .Y(n1914) );
  CLKBUFX2TS U1855 ( .A(n1914), .Y(n1872) );
  AOI22X1TS U1856 ( .A0(n1715), .A1(n1912), .B0(n1714), .B1(n1872), .Y(n1716)
         );
  AOI22X1TS U1857 ( .A0(n1784), .A1(n1720), .B0(n1719), .B1(
        \destinationAddressbuffer[6][3] ), .Y(n1726) );
  AOI22X1TS U1858 ( .A0(n1721), .A1(n1757), .B0(n85), .B1(n1756), .Y(n1725) );
  CLKBUFX2TS U1859 ( .A(n1722), .Y(n1922) );
  CLKBUFX2TS U1860 ( .A(destinationAddressIn_SOUTH[3]), .Y(n1923) );
  CLKBUFX2TS U1861 ( .A(n1923), .Y(n1882) );
  AOI22X1TS U1862 ( .A0(n104), .A1(n1922), .B0(n1723), .B1(n1882), .Y(n1724)
         );
  AOI22X1TS U1863 ( .A0(n1889), .A1(n1755), .B0(n1743), .B1(
        \destinationAddressbuffer[5][0] ), .Y(n1732) );
  AOI22X1TS U1864 ( .A0(n1748), .A1(n1728), .B0(n222), .B1(n1727), .Y(n1731)
         );
  AOI22X1TS U1865 ( .A0(n1729), .A1(n1891), .B0(n1738), .B1(
        destinationAddressIn_SOUTH[0]), .Y(n1730) );
  AOI22X1TS U1866 ( .A0(readRequesterAddress[1]), .A1(n1733), .B0(n1743), .B1(
        \destinationAddressbuffer[5][1] ), .Y(n1742) );
  AOI22X1TS U1867 ( .A0(n1737), .A1(n1736), .B0(n1735), .B1(n1734), .Y(n1741)
         );
  AOI22X1TS U1868 ( .A0(n1739), .A1(n1901), .B0(n1738), .B1(
        destinationAddressIn_SOUTH[1]), .Y(n1740) );
  AOI22X1TS U1869 ( .A0(readRequesterAddress[2]), .A1(n1744), .B0(n1743), .B1(
        \destinationAddressbuffer[5][2] ), .Y(n1753) );
  AOI22X1TS U1870 ( .A0(n1748), .A1(n1747), .B0(n1746), .B1(n1745), .Y(n1752)
         );
  AOI22X1TS U1871 ( .A0(n1750), .A1(n1912), .B0(n1749), .B1(
        destinationAddressIn_SOUTH[2]), .Y(n1751) );
  AOI22X1TS U1872 ( .A0(readRequesterAddress[3]), .A1(n1755), .B0(n1754), .B1(
        \destinationAddressbuffer[5][3] ), .Y(n1760) );
  AOI22X1TS U1873 ( .A0(n224), .A1(n1757), .B0(n222), .B1(n1756), .Y(n1759) );
  AOI22X1TS U1874 ( .A0(n256), .A1(n1922), .B0(n1738), .B1(
        destinationAddressIn_SOUTH[3]), .Y(n1758) );
  AOI22X1TS U1875 ( .A0(n1790), .A1(n276), .B0(n1775), .B1(
        \destinationAddressbuffer[4][0] ), .Y(n1765) );
  AOI22X1TS U1876 ( .A0(n1761), .A1(n1791), .B0(n274), .B1(
        destinationAddressIn_EAST[0]), .Y(n1764) );
  AOI22X1TS U1877 ( .A0(n284), .A1(n1892), .B0(n1762), .B1(n1891), .Y(n1763)
         );
  AOI22X1TS U1878 ( .A0(n1767), .A1(n1766), .B0(n1775), .B1(
        \destinationAddressbuffer[4][1] ), .Y(n1774) );
  AOI22X1TS U1879 ( .A0(n1769), .A1(n1798), .B0(n1768), .B1(
        destinationAddressIn_EAST[1]), .Y(n1773) );
  AOI22X1TS U1880 ( .A0(n1771), .A1(n1903), .B0(n1770), .B1(n1901), .Y(n1772)
         );
  AOI22X1TS U1881 ( .A0(n1777), .A1(n1776), .B0(n1775), .B1(
        \destinationAddressbuffer[4][2] ), .Y(n1782) );
  AOI22X1TS U1882 ( .A0(n1779), .A1(n1805), .B0(n1778), .B1(
        destinationAddressIn_EAST[2]), .Y(n1781) );
  AOI22X1TS U1883 ( .A0(n284), .A1(n1914), .B0(n300), .B1(n1912), .Y(n1780) );
  AOI22X1TS U1884 ( .A0(n1784), .A1(n276), .B0(n1783), .B1(
        \destinationAddressbuffer[4][3] ), .Y(n1789) );
  AOI22X1TS U1885 ( .A0(n297), .A1(n1813), .B0(n274), .B1(
        destinationAddressIn_EAST[3]), .Y(n1788) );
  AOI22X1TS U1886 ( .A0(n1786), .A1(n1923), .B0(n1785), .B1(n1922), .Y(n1787)
         );
  AOI22X1TS U1887 ( .A0(n1790), .A1(n1811), .B0(n1804), .B1(
        \destinationAddressbuffer[3][0] ), .Y(n1795) );
  AOI22X1TS U1888 ( .A0(n1792), .A1(n1791), .B0(n1797), .B1(
        destinationAddressIn_EAST[0]), .Y(n1794) );
  AOI22X1TS U1889 ( .A0(n174), .A1(n1850), .B0(n1386), .B1(n1849), .Y(n1793)
         );
  AOI22X1TS U1890 ( .A0(n1856), .A1(n1796), .B0(n1804), .B1(
        \destinationAddressbuffer[3][1] ), .Y(n1803) );
  AOI22X1TS U1891 ( .A0(n1799), .A1(n1798), .B0(n1797), .B1(
        destinationAddressIn_EAST[1]), .Y(n1802) );
  AOI22X1TS U1892 ( .A0(n1800), .A1(n1861), .B0(n1815), .B1(n1860), .Y(n1801)
         );
  AOI22X1TS U1893 ( .A0(n1868), .A1(n132), .B0(n1804), .B1(
        \destinationAddressbuffer[3][2] ), .Y(n1809) );
  AOI22X1TS U1894 ( .A0(n149), .A1(n1805), .B0(n169), .B1(
        destinationAddressIn_EAST[2]), .Y(n1808) );
  AOI22X1TS U1895 ( .A0(n1806), .A1(n1874), .B0(n131), .B1(n1872), .Y(n1807)
         );
  AOI22X1TS U1896 ( .A0(n1880), .A1(n1811), .B0(n1810), .B1(
        \destinationAddressbuffer[3][3] ), .Y(n1818) );
  AOI22X1TS U1897 ( .A0(n1814), .A1(n1813), .B0(n1812), .B1(
        destinationAddressIn_EAST[3]), .Y(n1817) );
  AOI22X1TS U1898 ( .A0(n174), .A1(n1884), .B0(n1815), .B1(n1882), .Y(n1816)
         );
  AOI22X1TS U1899 ( .A0(n1846), .A1(n1840), .B0(n1830), .B1(
        \destinationAddressbuffer[2][0] ), .Y(n1822) );
  AOI22X1TS U1900 ( .A0(n1819), .A1(destinationAddressIn_WEST[0]), .B0(n1002), 
        .B1(n1847), .Y(n1821) );
  AOI22X1TS U1901 ( .A0(n184), .A1(n1850), .B0(n1834), .B1(n1849), .Y(n1820)
         );
  AOI22X1TS U1902 ( .A0(n1898), .A1(n1823), .B0(n1830), .B1(
        \destinationAddressbuffer[2][1] ), .Y(n1829) );
  AOI22X1TS U1903 ( .A0(n1825), .A1(destinationAddressIn_WEST[1]), .B0(n1824), 
        .B1(n1857), .Y(n1828) );
  AOI22X1TS U1904 ( .A0(n1826), .A1(n1861), .B0(n187), .B1(n1860), .Y(n1827)
         );
  AOI22X1TS U1905 ( .A0(n1909), .A1(n1831), .B0(n1830), .B1(
        \destinationAddressbuffer[2][2] ), .Y(n1838) );
  AOI22X1TS U1906 ( .A0(n1833), .A1(destinationAddressIn_WEST[2]), .B0(n1832), 
        .B1(n1869), .Y(n1837) );
  AOI22X1TS U1907 ( .A0(n1835), .A1(n1874), .B0(n1834), .B1(n1872), .Y(n1836)
         );
  AOI22X1TS U1908 ( .A0(n1921), .A1(n1840), .B0(n1839), .B1(
        \destinationAddressbuffer[2][3] ), .Y(n1845) );
  AOI22X1TS U1909 ( .A0(n213), .A1(destinationAddressIn_WEST[3]), .B0(n1), 
        .B1(n1881), .Y(n1844) );
  AOI22X1TS U1910 ( .A0(n1842), .A1(n1884), .B0(n1841), .B1(n1882), .Y(n1843)
         );
  AOI22X1TS U1911 ( .A0(n1846), .A1(n320), .B0(n1866), .B1(
        \destinationAddressbuffer[1][0] ), .Y(n1854) );
  AOI22X1TS U1912 ( .A0(n1848), .A1(destinationAddressIn_WEST[0]), .B0(n1029), 
        .B1(n1847), .Y(n1853) );
  AOI22X1TS U1913 ( .A0(n1851), .A1(n1850), .B0(n1873), .B1(n1849), .Y(n1852)
         );
  AOI22X1TS U1914 ( .A0(n1856), .A1(n1855), .B0(n1866), .B1(
        \destinationAddressbuffer[1][1] ), .Y(n1865) );
  AOI22X1TS U1915 ( .A0(n1859), .A1(destinationAddressIn_WEST[1]), .B0(n1858), 
        .B1(n1857), .Y(n1864) );
  AOI22X1TS U1916 ( .A0(n1862), .A1(n1861), .B0(n335), .B1(n1860), .Y(n1863)
         );
  AOI22X1TS U1917 ( .A0(n1868), .A1(n1867), .B0(n1866), .B1(
        \destinationAddressbuffer[1][2] ), .Y(n1878) );
  AOI22X1TS U1918 ( .A0(n1871), .A1(destinationAddressIn_WEST[2]), .B0(n1870), 
        .B1(n1869), .Y(n1877) );
  AOI22X1TS U1919 ( .A0(n1875), .A1(n1874), .B0(n1873), .B1(n1872), .Y(n1876)
         );
  AOI22X1TS U1920 ( .A0(n1880), .A1(n320), .B0(n1879), .B1(
        \destinationAddressbuffer[1][3] ), .Y(n1888) );
  AOI22X1TS U1921 ( .A0(n361), .A1(destinationAddressIn_WEST[3]), .B0(n318), 
        .B1(n1881), .Y(n1887) );
  AOI22X1TS U1922 ( .A0(n1885), .A1(n1884), .B0(n1883), .B1(n1882), .Y(n1886)
         );
  AOI22X1TS U1923 ( .A0(n1889), .A1(n1920), .B0(n1907), .B1(
        \destinationAddressbuffer[0][0] ), .Y(n1896) );
  AOI22X1TS U1924 ( .A0(n1890), .A1(destinationAddressIn_WEST[0]), .B0(n414), 
        .B1(destinationAddressIn_EAST[0]), .Y(n1895) );
  AOI22X1TS U1925 ( .A0(n1893), .A1(n1892), .B0(n1902), .B1(n1891), .Y(n1894)
         );
  AOI22X1TS U1926 ( .A0(n1898), .A1(n1897), .B0(n1907), .B1(
        \destinationAddressbuffer[0][1] ), .Y(n1906) );
  AOI22X1TS U1927 ( .A0(n1900), .A1(destinationAddressIn_WEST[1]), .B0(n1899), 
        .B1(destinationAddressIn_EAST[1]), .Y(n1905) );
  AOI22X1TS U1928 ( .A0(n439), .A1(n1903), .B0(n1902), .B1(n1901), .Y(n1904)
         );
  AOI22X1TS U1929 ( .A0(n1909), .A1(n1908), .B0(n1907), .B1(
        \destinationAddressbuffer[0][2] ), .Y(n1918) );
  AOI22X1TS U1930 ( .A0(n1911), .A1(destinationAddressIn_WEST[2]), .B0(n1910), 
        .B1(destinationAddressIn_EAST[2]), .Y(n1917) );
  AOI22X1TS U1931 ( .A0(n1915), .A1(n1914), .B0(n1913), .B1(n1912), .Y(n1916)
         );
  AOI22X1TS U1932 ( .A0(n1921), .A1(n1920), .B0(n1919), .B1(
        \destinationAddressbuffer[0][3] ), .Y(n1927) );
  AOI22X1TS U1933 ( .A0(n437), .A1(destinationAddressIn_WEST[3]), .B0(n1056), 
        .B1(destinationAddressIn_EAST[3]), .Y(n1926) );
  AOI22X1TS U1934 ( .A0(n1924), .A1(n1923), .B0(n411), .B1(n1922), .Y(n1925)
         );
endmodule


module outputPortArbiter_2 ( clk, reset, selectBit_NORTH, 
        destinationAddressIn_NORTH, requesterAddressIn_NORTH, readIn_NORTH, 
        writeIn_NORTH, dataIn_NORTH, selectBit_SOUTH, 
        destinationAddressIn_SOUTH, requesterAddressIn_SOUTH, readIn_SOUTH, 
        writeIn_SOUTH, dataIn_SOUTH, selectBit_EAST, destinationAddressIn_EAST, 
        requesterAddressIn_EAST, readIn_EAST, writeIn_EAST, dataIn_EAST, 
        selectBit_WEST, destinationAddressIn_WEST, requesterAddressIn_WEST, 
        readIn_WEST, writeIn_WEST, dataIn_WEST, readReady, 
        readRequesterAddress, cacheDataOut, destinationAddressOut, 
        requesterAddressOut, readOut, writeOut, dataOut );
  input [11:0] destinationAddressIn_NORTH;
  input [3:0] requesterAddressIn_NORTH;
  input [5:0] dataIn_NORTH;
  input [11:0] destinationAddressIn_SOUTH;
  input [3:0] requesterAddressIn_SOUTH;
  input [5:0] dataIn_SOUTH;
  input [11:0] destinationAddressIn_EAST;
  input [3:0] requesterAddressIn_EAST;
  input [5:0] dataIn_EAST;
  input [11:0] destinationAddressIn_WEST;
  input [3:0] requesterAddressIn_WEST;
  input [5:0] dataIn_WEST;
  input [3:0] readRequesterAddress;
  input [5:0] cacheDataOut;
  output [11:0] destinationAddressOut;
  output [3:0] requesterAddressOut;
  output [5:0] dataOut;
  input clk, reset, selectBit_NORTH, readIn_NORTH, writeIn_NORTH,
         selectBit_SOUTH, readIn_SOUTH, writeIn_SOUTH, selectBit_EAST,
         readIn_EAST, writeIn_EAST, selectBit_WEST, readIn_WEST, writeIn_WEST,
         readReady;
  output readOut, writeOut;
  wire   \requesterAddressbuffer[0][3] , \requesterAddressbuffer[0][2] ,
         \requesterAddressbuffer[0][1] , \requesterAddressbuffer[0][0] ,
         \requesterAddressbuffer[1][3] , \requesterAddressbuffer[1][2] ,
         \requesterAddressbuffer[1][1] , \requesterAddressbuffer[1][0] ,
         \requesterAddressbuffer[2][3] , \requesterAddressbuffer[2][2] ,
         \requesterAddressbuffer[2][1] , \requesterAddressbuffer[2][0] ,
         \requesterAddressbuffer[3][3] , \requesterAddressbuffer[3][2] ,
         \requesterAddressbuffer[3][1] , \requesterAddressbuffer[3][0] ,
         \requesterAddressbuffer[4][3] , \requesterAddressbuffer[4][2] ,
         \requesterAddressbuffer[4][1] , \requesterAddressbuffer[4][0] ,
         \requesterAddressbuffer[5][3] , \requesterAddressbuffer[5][2] ,
         \requesterAddressbuffer[5][1] , \requesterAddressbuffer[5][0] ,
         \requesterAddressbuffer[6][3] , \requesterAddressbuffer[6][2] ,
         \requesterAddressbuffer[6][1] , \requesterAddressbuffer[6][0] ,
         \requesterAddressbuffer[7][3] , \requesterAddressbuffer[7][2] ,
         \requesterAddressbuffer[7][1] , \requesterAddressbuffer[7][0] ,
         \destinationAddressbuffer[0][11] , \destinationAddressbuffer[0][10] ,
         \destinationAddressbuffer[0][9] , \destinationAddressbuffer[0][8] ,
         \destinationAddressbuffer[0][7] , \destinationAddressbuffer[0][6] ,
         \destinationAddressbuffer[0][5] , \destinationAddressbuffer[0][4] ,
         \destinationAddressbuffer[0][3] , \destinationAddressbuffer[0][2] ,
         \destinationAddressbuffer[0][1] , \destinationAddressbuffer[0][0] ,
         \destinationAddressbuffer[1][11] , \destinationAddressbuffer[1][10] ,
         \destinationAddressbuffer[1][9] , \destinationAddressbuffer[1][8] ,
         \destinationAddressbuffer[1][7] , \destinationAddressbuffer[1][6] ,
         \destinationAddressbuffer[1][5] , \destinationAddressbuffer[1][4] ,
         \destinationAddressbuffer[1][3] , \destinationAddressbuffer[1][2] ,
         \destinationAddressbuffer[1][1] , \destinationAddressbuffer[1][0] ,
         \destinationAddressbuffer[2][11] , \destinationAddressbuffer[2][10] ,
         \destinationAddressbuffer[2][9] , \destinationAddressbuffer[2][8] ,
         \destinationAddressbuffer[2][7] , \destinationAddressbuffer[2][6] ,
         \destinationAddressbuffer[2][5] , \destinationAddressbuffer[2][4] ,
         \destinationAddressbuffer[2][3] , \destinationAddressbuffer[2][2] ,
         \destinationAddressbuffer[2][1] , \destinationAddressbuffer[2][0] ,
         \destinationAddressbuffer[3][11] , \destinationAddressbuffer[3][10] ,
         \destinationAddressbuffer[3][9] , \destinationAddressbuffer[3][8] ,
         \destinationAddressbuffer[3][7] , \destinationAddressbuffer[3][6] ,
         \destinationAddressbuffer[3][5] , \destinationAddressbuffer[3][4] ,
         \destinationAddressbuffer[3][3] , \destinationAddressbuffer[3][2] ,
         \destinationAddressbuffer[3][1] , \destinationAddressbuffer[3][0] ,
         \destinationAddressbuffer[4][11] , \destinationAddressbuffer[4][10] ,
         \destinationAddressbuffer[4][9] , \destinationAddressbuffer[4][8] ,
         \destinationAddressbuffer[4][7] , \destinationAddressbuffer[4][6] ,
         \destinationAddressbuffer[4][5] , \destinationAddressbuffer[4][4] ,
         \destinationAddressbuffer[4][3] , \destinationAddressbuffer[4][2] ,
         \destinationAddressbuffer[4][1] , \destinationAddressbuffer[4][0] ,
         \destinationAddressbuffer[5][11] , \destinationAddressbuffer[5][10] ,
         \destinationAddressbuffer[5][9] , \destinationAddressbuffer[5][8] ,
         \destinationAddressbuffer[5][7] , \destinationAddressbuffer[5][6] ,
         \destinationAddressbuffer[5][5] , \destinationAddressbuffer[5][4] ,
         \destinationAddressbuffer[5][3] , \destinationAddressbuffer[5][2] ,
         \destinationAddressbuffer[5][1] , \destinationAddressbuffer[5][0] ,
         \destinationAddressbuffer[6][11] , \destinationAddressbuffer[6][10] ,
         \destinationAddressbuffer[6][9] , \destinationAddressbuffer[6][8] ,
         \destinationAddressbuffer[6][7] , \destinationAddressbuffer[6][6] ,
         \destinationAddressbuffer[6][5] , \destinationAddressbuffer[6][4] ,
         \destinationAddressbuffer[6][3] , \destinationAddressbuffer[6][2] ,
         \destinationAddressbuffer[6][1] , \destinationAddressbuffer[6][0] ,
         \destinationAddressbuffer[7][11] , \destinationAddressbuffer[7][10] ,
         \destinationAddressbuffer[7][9] , \destinationAddressbuffer[7][8] ,
         \destinationAddressbuffer[7][7] , \destinationAddressbuffer[7][6] ,
         \destinationAddressbuffer[7][5] , \destinationAddressbuffer[7][4] ,
         \destinationAddressbuffer[7][3] , \destinationAddressbuffer[7][2] ,
         \destinationAddressbuffer[7][1] , \destinationAddressbuffer[7][0] ,
         \dataoutbuffer[7][5] , \dataoutbuffer[7][4] , \dataoutbuffer[7][3] ,
         \dataoutbuffer[7][2] , \dataoutbuffer[7][1] , \dataoutbuffer[7][0] ,
         \dataoutbuffer[6][5] , \dataoutbuffer[6][4] , \dataoutbuffer[6][3] ,
         \dataoutbuffer[6][2] , \dataoutbuffer[6][1] , \dataoutbuffer[6][0] ,
         \dataoutbuffer[5][5] , \dataoutbuffer[5][4] , \dataoutbuffer[5][3] ,
         \dataoutbuffer[5][2] , \dataoutbuffer[5][1] , \dataoutbuffer[5][0] ,
         \dataoutbuffer[4][5] , \dataoutbuffer[4][4] , \dataoutbuffer[4][3] ,
         \dataoutbuffer[4][2] , \dataoutbuffer[4][1] , \dataoutbuffer[4][0] ,
         \dataoutbuffer[3][5] , \dataoutbuffer[3][4] , \dataoutbuffer[3][3] ,
         \dataoutbuffer[3][2] , \dataoutbuffer[3][1] , \dataoutbuffer[3][0] ,
         \dataoutbuffer[2][5] , \dataoutbuffer[2][4] , \dataoutbuffer[2][3] ,
         \dataoutbuffer[2][2] , \dataoutbuffer[2][1] , \dataoutbuffer[2][0] ,
         \dataoutbuffer[1][5] , \dataoutbuffer[1][4] , \dataoutbuffer[1][3] ,
         \dataoutbuffer[1][2] , \dataoutbuffer[1][1] , \dataoutbuffer[1][0] ,
         \dataoutbuffer[0][5] , \dataoutbuffer[0][4] , \dataoutbuffer[0][3] ,
         \dataoutbuffer[0][2] , \dataoutbuffer[0][1] , \dataoutbuffer[0][0] ,
         N2624, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167;
  wire   [0:7] writeOutbuffer;
  wire   [0:7] readOutbuffer;

  DFFNSRX1TS full_reg_reg ( .D(N2624), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(
        n1936) );
  DFFNSRX1TS \requesterAddressbuffer_reg[2][0]  ( .D(n1996), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[2][1]  ( .D(n1997), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[2][2]  ( .D(n1998), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[2][3]  ( .D(n1999), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][0]  ( .D(n2132), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][1]  ( .D(n2133), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][2]  ( .D(n2134), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][3]  ( .D(n2135), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][0]  ( .D(n2008), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][1]  ( .D(n2009), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][2]  ( .D(n2010), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][3]  ( .D(n2011), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][4]  ( .D(n2012), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][5]  ( .D(n2013), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][5] ) );
  DFFNSRX1TS \writeOutbuffer_reg[7]  ( .D(n2056), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[7]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][4]  ( .D(n2076), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][5]  ( .D(n2077), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][6]  ( .D(n2078), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][7]  ( .D(n2079), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][8]  ( .D(n2080), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][9]  ( .D(n2081), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][11]  ( .D(n2083), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[6]  ( .D(n2057), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[6]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][4]  ( .D(n2088), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][5]  ( .D(n2089), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][6]  ( .D(n2090), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][7]  ( .D(n2091), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][8]  ( .D(n2092), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][9]  ( .D(n2093), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][10]  ( .D(n2094), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][11]  ( .D(n2095), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[3]  ( .D(n2060), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[3]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][4]  ( .D(n2124), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][5]  ( .D(n2125), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][6]  ( .D(n2126), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][7]  ( .D(n2127), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][8]  ( .D(n2128), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][9]  ( .D(n2129), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][10]  ( .D(n2130), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][11]  ( .D(n2131), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[2]  ( .D(n2061), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[2]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][4]  ( .D(n2136), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][5]  ( .D(n2137), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][6]  ( .D(n2138), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][7]  ( .D(n2139), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][8]  ( .D(n2140), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][9]  ( .D(n2141), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][10]  ( .D(n2142), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][11]  ( .D(n2143), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][11] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][0]  ( .D(n2050), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][1]  ( .D(n2051), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][2]  ( .D(n2052), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][3]  ( .D(n2053), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][4]  ( .D(n2054), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][5]  ( .D(n2055), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][0]  ( .D(n2044), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][1]  ( .D(n2045), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][2]  ( .D(n2046), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][3]  ( .D(n2047), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][4]  ( .D(n2048), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][5]  ( .D(n2049), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][5] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[5][0]  ( .D(n1984), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[5][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[5][1]  ( .D(n1985), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[5][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[5][2]  ( .D(n1986), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[5][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[5][3]  ( .D(n1987), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[5][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][0]  ( .D(n2096), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][1]  ( .D(n2097), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][2]  ( .D(n2098), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][3]  ( .D(n2099), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[4][0]  ( .D(n1988), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[4][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[4][1]  ( .D(n1989), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[4][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[4][2]  ( .D(n1990), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[4][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[4][3]  ( .D(n1991), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[4][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][0]  ( .D(n2108), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][1]  ( .D(n2109), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][2]  ( .D(n2110), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][3]  ( .D(n2111), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][0]  ( .D(n2026), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][1]  ( .D(n2027), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][2]  ( .D(n2028), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][3]  ( .D(n2029), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][4]  ( .D(n2030), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][5]  ( .D(n2031), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][0]  ( .D(n2020), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][1]  ( .D(n2021), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][2]  ( .D(n2022), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][3]  ( .D(n2023), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][4]  ( .D(n2024), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][5]  ( .D(n2025), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][5] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[1][0]  ( .D(n2000), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[1][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[1][1]  ( .D(n2001), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[1][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[1][2]  ( .D(n2002), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[1][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[1][3]  ( .D(n2003), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[1][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][0]  ( .D(n2144), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][1]  ( .D(n2145), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][2]  ( .D(n2146), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][3]  ( .D(n2147), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[0][0]  ( .D(n2004), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[0][1]  ( .D(n2005), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[0][2]  ( .D(n2006), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[0][3]  ( .D(n2007), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][0]  ( .D(n2156), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][1]  ( .D(n2157), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][2]  ( .D(n2158), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][3]  ( .D(n2159), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[7][0]  ( .D(n1976), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[7][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[7][1]  ( .D(n1977), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[7][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[7][2]  ( .D(n1978), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[7][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[7][3]  ( .D(n1979), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[7][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][0]  ( .D(n2072), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][1]  ( .D(n2073), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][2]  ( .D(n2074), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][3]  ( .D(n2075), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[6][0]  ( .D(n1980), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[6][1]  ( .D(n1981), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[6][2]  ( .D(n1982), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[6][3]  ( .D(n1983), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][0]  ( .D(n2084), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][1]  ( .D(n2085), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][2]  ( .D(n2086), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][3]  ( .D(n2087), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][0]  ( .D(n2038), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][1]  ( .D(n2039), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][2]  ( .D(n2040), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][3]  ( .D(n2041), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][4]  ( .D(n2042), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][5]  ( .D(n2043), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][0]  ( .D(n2032), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][1]  ( .D(n2033), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][2]  ( .D(n2034), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][3]  ( .D(n2035), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][4]  ( .D(n2036), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][5]  ( .D(n2037), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][5] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[3][0]  ( .D(n1992), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[3][1]  ( .D(n1993), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[3][2]  ( .D(n1994), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[3][3]  ( .D(n1995), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][0]  ( .D(n2120), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][1]  ( .D(n2121), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][2]  ( .D(n2122), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][3]  ( .D(n2123), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][0]  ( .D(n2014), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][1]  ( .D(n2015), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][2]  ( .D(n2016), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][3]  ( .D(n2017), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][4]  ( .D(n2018), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][5]  ( .D(n2019), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][5] ) );
  DFFNSRX1TS \writeOutbuffer_reg[5]  ( .D(n2058), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[5]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][4]  ( .D(n2100), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][5]  ( .D(n2101), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][6]  ( .D(n2102), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][7]  ( .D(n2103), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][8]  ( .D(n2104), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][9]  ( .D(n2105), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][10]  ( .D(n2106), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][11]  ( .D(n2107), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[4]  ( .D(n2059), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[4]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][4]  ( .D(n2112), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][5]  ( .D(n2113), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][6]  ( .D(n2114), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][7]  ( .D(n2115), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][8]  ( .D(n2116), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][9]  ( .D(n2117), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][10]  ( .D(n2118), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][11]  ( .D(n2119), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[1]  ( .D(n2062), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[1]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][4]  ( .D(n2148), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][5]  ( .D(n2149), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][6]  ( .D(n2150), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][7]  ( .D(n2151), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][8]  ( .D(n2152), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][9]  ( .D(n2153), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][10]  ( .D(n2154), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][11]  ( .D(n2155), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[0]  ( .D(n2063), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[0]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][4]  ( .D(n2160), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][5]  ( .D(n2161), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][6]  ( .D(n2162), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][7]  ( .D(n2163), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][8]  ( .D(n2164), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][9]  ( .D(n2165), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][10]  ( .D(n2166), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][11]  ( .D(n2167), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][11] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][10]  ( .D(n2082), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][10] ) );
  DFFNSRX1TS writeOut_reg ( .D(n1953), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        writeOut) );
  DFFNSRX1TS \destinationAddressOut_reg[4]  ( .D(n1962), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[4]) );
  DFFNSRX1TS \destinationAddressOut_reg[5]  ( .D(n1963), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[5]) );
  DFFNSRX1TS \destinationAddressOut_reg[6]  ( .D(n1964), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[6]) );
  DFFNSRX1TS \destinationAddressOut_reg[7]  ( .D(n1965), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[7]) );
  DFFNSRX1TS \destinationAddressOut_reg[8]  ( .D(n1966), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[8]) );
  DFFNSRX1TS \destinationAddressOut_reg[9]  ( .D(n1967), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[9]) );
  DFFNSRX1TS \destinationAddressOut_reg[10]  ( .D(n1968), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[10]) );
  DFFNSRX1TS \destinationAddressOut_reg[11]  ( .D(n1969), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[11]) );
  DFFNSRX1TS readOut_reg ( .D(n1952), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        readOut) );
  DFFNSRX1TS \requesterAddressOut_reg[0]  ( .D(n1954), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[0]) );
  DFFNSRX1TS \requesterAddressOut_reg[1]  ( .D(n1955), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[1]) );
  DFFNSRX1TS \requesterAddressOut_reg[2]  ( .D(n1956), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[2]) );
  DFFNSRX1TS \requesterAddressOut_reg[3]  ( .D(n1957), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[3]) );
  DFFNSRX1TS \destinationAddressOut_reg[0]  ( .D(n1958), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[0]) );
  DFFNSRX1TS \destinationAddressOut_reg[1]  ( .D(n1959), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[1]) );
  DFFNSRX1TS \destinationAddressOut_reg[2]  ( .D(n1960), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[2]) );
  DFFNSRX1TS \destinationAddressOut_reg[3]  ( .D(n1961), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[3]) );
  DFFNSRX1TS \dataOut_reg[0]  ( .D(n1970), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[0]) );
  DFFNSRX1TS \dataOut_reg[1]  ( .D(n1971), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[1]) );
  DFFNSRX1TS \dataOut_reg[2]  ( .D(n1972), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[2]) );
  DFFNSRX1TS \dataOut_reg[3]  ( .D(n1973), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[3]) );
  DFFNSRX1TS \dataOut_reg[4]  ( .D(n1974), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[4]) );
  DFFNSRX1TS \dataOut_reg[5]  ( .D(n1975), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[5]) );
  DFFNSRX1TS \read_reg_reg[1]  ( .D(n1951), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1929), .QN(n1928) );
  DFFNSRX1TS \write_reg_reg[0]  ( .D(n1946), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1927), .QN(n1931) );
  DFFNSRX1TS \write_reg_reg[2]  ( .D(n1948), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1932), .QN(n1933) );
  DFFNSRX1TS \read_reg_reg[0]  ( .D(n1945), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1922), .QN(n1934) );
  DFFNSRX1TS \read_reg_reg[2]  ( .D(n1950), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1925), .QN(n1926) );
  DFFNSRX1TS empty_reg_reg ( .D(n1949), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        n1924), .QN(n1923) );
  DFFNSRX1TS \readOutbuffer_reg[7]  ( .D(n2064), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[7]), .QN(n1937) );
  DFFNSRX1TS \readOutbuffer_reg[4]  ( .D(n2067), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[4]), .QN(n1940) );
  DFFNSRX1TS \readOutbuffer_reg[6]  ( .D(n2065), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[6]), .QN(n1938) );
  DFFNSRX1TS \readOutbuffer_reg[5]  ( .D(n2066), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[5]), .QN(n1939) );
  DFFNSRX1TS \readOutbuffer_reg[0]  ( .D(n2071), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[0]), .QN(n1944) );
  DFFNSRX1TS \readOutbuffer_reg[2]  ( .D(n2069), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[2]), .QN(n1942) );
  DFFNSRX1TS \readOutbuffer_reg[1]  ( .D(n2070), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[1]), .QN(n1943) );
  DFFNSRX1TS \write_reg_reg[1]  ( .D(n1947), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1930), .QN(n1935) );
  DFFNSRX1TS \readOutbuffer_reg[3]  ( .D(n2068), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[3]), .QN(n1941) );
  CMPR32X2TS U3 ( .A(n475), .B(n483), .C(n474), .CO(n469), .S(n492) );
  CLKBUFX2TS U4 ( .A(n17), .Y(n219) );
  CMPR32X2TS U5 ( .A(n529), .B(n452), .C(n455), .CO(n445), .S(n457) );
  CMPR32X2TS U6 ( .A(n451), .B(n513), .C(n450), .CO(n453), .S(n466) );
  CMPR32X2TS U7 ( .A(n454), .B(n85), .C(n19), .CO(n20), .S(n17) );
  CLKBUFX2TS U8 ( .A(n23), .Y(n83) );
  CMPR32X2TS U9 ( .A(selectBit_SOUTH), .B(selectBit_NORTH), .C(selectBit_EAST), 
        .CO(n454), .S(n450) );
  NOR3XLTS U10 ( .A(n511), .B(selectBit_EAST), .C(n513), .Y(n506) );
  NOR2XLTS U11 ( .A(n1561), .B(n41), .Y(n45) );
  NOR2XLTS U12 ( .A(n129), .B(n381), .Y(n1610) );
  ADDHXLTS U13 ( .A(n442), .B(n450), .CO(n19), .S(n18) );
  INVX2TS U14 ( .A(n1635), .Y(n1633) );
  INVX2TS U15 ( .A(n1576), .Y(n1574) );
  NOR2XLTS U16 ( .A(selectBit_NORTH), .B(selectBit_SOUTH), .Y(n537) );
  NOR2XLTS U17 ( .A(n314), .B(n1640), .Y(n315) );
  NOR2XLTS U18 ( .A(n314), .B(n1614), .Y(n134) );
  NOR2XLTS U19 ( .A(n386), .B(n1605), .Y(n274) );
  NOR3XLTS U20 ( .A(n1592), .B(n1587), .C(n226), .Y(n222) );
  NOR2XLTS U21 ( .A(n481), .B(n1580), .Y(n88) );
  NOR2XLTS U22 ( .A(n1569), .B(n386), .Y(n36) );
  NOR2XLTS U23 ( .A(n1619), .B(n189), .Y(n187) );
  CLKBUFX2TS U24 ( .A(n1355), .Y(n1349) );
  INVX2TS U25 ( .A(reset), .Y(n490) );
  AOI211XLTS U26 ( .A0(n479), .A1(n524), .B0(n478), .C0(n477), .Y(n480) );
  NOR2X1TS U27 ( .A(n1572), .B(n93), .Y(n94) );
  NAND2BXLTS U28 ( .AN(n137), .B(n132), .Y(n136) );
  OAI2BB2XLTS U29 ( .B0(n1936), .B1(n502), .A0N(n495), .A1N(n480), .Y(N2624)
         );
  NAND2BXLTS U30 ( .AN(n91), .B(n90), .Y(n93) );
  NAND2BXLTS U31 ( .AN(n394), .B(n393), .Y(n396) );
  NAND2BXLTS U32 ( .AN(n277), .B(n276), .Y(n279) );
  INVX1TS U33 ( .A(n1589), .Y(n1587) );
  NOR2X1TS U34 ( .A(n1613), .B(n1610), .Y(n132) );
  NAND2BX1TS U35 ( .AN(n128), .B(selectBit_EAST), .Y(n381) );
  XOR2XLTS U36 ( .A(n523), .B(n491), .Y(n478) );
  NAND3X1TS U37 ( .A(n85), .B(n32), .C(n220), .Y(n1561) );
  NAND3X1TS U38 ( .A(n27), .B(n220), .C(n269), .Y(n1583) );
  NOR2X1TS U39 ( .A(n220), .B(n82), .Y(n309) );
  INVX1TS U40 ( .A(n1579), .Y(n1577) );
  INVX1TS U41 ( .A(n1604), .Y(n1601) );
  NOR3X1TS U42 ( .A(n179), .B(n81), .C(n379), .Y(n1613) );
  NAND2BX1TS U43 ( .AN(n127), .B(n511), .Y(n379) );
  INVX1TS U44 ( .A(n25), .Y(n130) );
  AND2X2TS U45 ( .A(n522), .B(n1936), .Y(n273) );
  NOR2X1TS U46 ( .A(n449), .B(n503), .Y(n21) );
  INVX1TS U47 ( .A(n1933), .Y(n497) );
  NOR2XLTS U48 ( .A(n1592), .B(n1589), .Y(n225) );
  NOR3BXLTS U49 ( .AN(readReady), .B(n511), .C(n510), .Y(n536) );
  INVX2TS U50 ( .A(n322), .Y(n361) );
  OR2X1TS U51 ( .A(n275), .B(n931), .Y(n1407) );
  OR2X1TS U52 ( .A(n223), .B(n912), .Y(n1438) );
  OR2X1TS U53 ( .A(n184), .B(n983), .Y(n1345) );
  OR2X1TS U54 ( .A(n135), .B(n956), .Y(n1379) );
  OR2X1TS U55 ( .A(n89), .B(n894), .Y(n1475) );
  OR2X1TS U56 ( .A(n37), .B(n1653), .Y(n1527) );
  NAND4XLTS U57 ( .A(n486), .B(n473), .C(n509), .D(n485), .Y(n1614) );
  CLKBUFX2TS U58 ( .A(n1379), .Y(n1615) );
  CLKAND2X2TS U59 ( .A(n468), .B(n467), .Y(n474) );
  NAND4XLTS U60 ( .A(n442), .B(n508), .C(n482), .D(n384), .Y(n1640) );
  NOR3X1TS U61 ( .A(n126), .B(n179), .C(n379), .Y(n1626) );
  INVX2TS U62 ( .A(n1623), .Y(n1620) );
  CLKBUFX2TS U63 ( .A(n1345), .Y(n1628) );
  NOR3X1TS U64 ( .A(n219), .B(n18), .C(n379), .Y(n1650) );
  INVX2TS U65 ( .A(n1647), .Y(n1644) );
  NOR3X1TS U66 ( .A(n219), .B(n81), .C(n266), .Y(n1592) );
  CLKBUFX2TS U67 ( .A(n1438), .Y(n1594) );
  NAND4XLTS U68 ( .A(n85), .B(n497), .C(n508), .D(n389), .Y(n1580) );
  NOR3XLTS U69 ( .A(n18), .B(n179), .C(n266), .Y(n1579) );
  INVX2TS U70 ( .A(n1573), .Y(n1572) );
  CLKBUFX2TS U71 ( .A(n1475), .Y(n1581) );
  NAND4XLTS U72 ( .A(n271), .B(n509), .C(n389), .D(n384), .Y(n1605) );
  NOR3XLTS U73 ( .A(n219), .B(n18), .C(n266), .Y(n1604) );
  INVX2TS U74 ( .A(n1600), .Y(n1598) );
  CLKBUFX2TS U75 ( .A(n1407), .Y(n1606) );
  NAND4XLTS U76 ( .A(n1927), .B(n493), .C(n497), .D(n508), .Y(n1569) );
  INVX2TS U77 ( .A(n1565), .Y(n1563) );
  CLKBUFX2TS U78 ( .A(n1527), .Y(n1570) );
  NAND3XLTS U79 ( .A(n537), .B(n1924), .C(n536), .Y(n559) );
  CLKAND2X2TS U80 ( .A(n522), .B(n520), .Y(n550) );
  INVX2TS U81 ( .A(selectBit_NORTH), .Y(n503) );
  NOR2XLTS U82 ( .A(n1604), .B(n1600), .Y(n276) );
  NOR2XLTS U83 ( .A(n1568), .B(n1565), .Y(n39) );
  NOR2XLTS U84 ( .A(n1650), .B(n1647), .Y(n393) );
  AO21X1TS U85 ( .A0(n449), .A1(n503), .B0(n311), .Y(n24) );
  OAI21XLTS U86 ( .A0(n31), .A1(n28), .B0(n30), .Y(n128) );
  NAND3XLTS U87 ( .A(selectBit_NORTH), .B(n506), .C(n505), .Y(n517) );
  NAND3XLTS U88 ( .A(n504), .B(n506), .C(n503), .Y(n516) );
  NOR2XLTS U89 ( .A(n1639), .B(n1635), .Y(n319) );
  NAND2BXLTS U90 ( .AN(n226), .B(n225), .Y(n227) );
  NAND3XLTS U91 ( .A(n311), .B(n444), .C(n388), .Y(n221) );
  NOR2XLTS U92 ( .A(n1579), .B(n1576), .Y(n90) );
  NAND2X1TS U93 ( .A(n135), .B(n1614), .Y(n137) );
  NAND2BXLTS U94 ( .AN(n40), .B(n39), .Y(n41) );
  XOR2XLTS U95 ( .A(n445), .B(n447), .Y(n463) );
  OAI21XLTS U96 ( .A0(n486), .A1(n1928), .B0(n447), .Y(n448) );
  NOR2X1TS U97 ( .A(n12), .B(n82), .Y(n31) );
  INVX2TS U98 ( .A(n269), .Y(n383) );
  XOR2X1TS U99 ( .A(n497), .B(n20), .Y(n127) );
  NAND2BXLTS U100 ( .AN(n320), .B(n319), .Y(n323) );
  NAND2BXLTS U101 ( .AN(n186), .B(n185), .Y(n189) );
  XOR2XLTS U102 ( .A(n471), .B(n470), .Y(n494) );
  INVX2TS U103 ( .A(n1613), .Y(n1611) );
  INVX2TS U104 ( .A(n1610), .Y(n1608) );
  NOR2XLTS U105 ( .A(n87), .B(reset), .Y(n496) );
  NOR3XLTS U106 ( .A(n32), .B(n383), .C(n12), .Y(n1632) );
  INVX2TS U107 ( .A(n1632), .Y(n1630) );
  INVX2TS U108 ( .A(n1639), .Y(n1636) );
  NOR3XLTS U109 ( .A(n310), .B(n309), .C(n381), .Y(n1635) );
  NAND4XLTS U110 ( .A(n483), .B(readReady), .C(n389), .D(n485), .Y(n1627) );
  NOR3XLTS U111 ( .A(n32), .B(n83), .C(n269), .Y(n1619) );
  INVX2TS U112 ( .A(n1619), .Y(n1617) );
  INVX2TS U113 ( .A(n1626), .Y(n1624) );
  NAND4XLTS U114 ( .A(n513), .B(n389), .C(n388), .D(n485), .Y(n1651) );
  NOR3XLTS U115 ( .A(n32), .B(n383), .C(n83), .Y(n1643) );
  INVX2TS U116 ( .A(n1650), .Y(n1648) );
  INVX2TS U117 ( .A(n1643), .Y(n1642) );
  NOR3BXLTS U118 ( .AN(n382), .B(n381), .C(n380), .Y(n1647) );
  NAND4XLTS U119 ( .A(n473), .B(n271), .C(readReady), .D(n384), .Y(n1593) );
  INVX2TS U120 ( .A(n1592), .Y(n1590) );
  INVX2TS U121 ( .A(n1583), .Y(n1586) );
  NOR3XLTS U122 ( .A(n310), .B(n309), .C(n268), .Y(n1589) );
  NOR3XLTS U123 ( .A(n383), .B(n23), .C(n26), .Y(n1597) );
  INVX2TS U124 ( .A(n1597), .Y(n1596) );
  NOR3BXLTS U125 ( .AN(n382), .B(n268), .C(n267), .Y(n1600) );
  NAND4XLTS U126 ( .A(n17), .B(n126), .C(n127), .D(n451), .Y(n1566) );
  INVX2TS U127 ( .A(n1561), .Y(n1562) );
  NOR2XLTS U128 ( .A(n129), .B(n268), .Y(n1565) );
  INVX2TS U129 ( .A(destinationAddressIn_SOUTH[11]), .Y(n144) );
  INVX2TS U130 ( .A(destinationAddressIn_SOUTH[10]), .Y(n148) );
  INVX2TS U131 ( .A(destinationAddressIn_SOUTH[9]), .Y(n154) );
  INVX2TS U132 ( .A(destinationAddressIn_SOUTH[8]), .Y(n140) );
  CLKAND2X2TS U133 ( .A(n468), .B(n466), .Y(n472) );
  AO22XLTS U134 ( .A0(n497), .A1(n496), .B0(n495), .B1(n494), .Y(n1948) );
  AO22XLTS U135 ( .A0(n1927), .A1(n496), .B0(n495), .B1(n491), .Y(n1946) );
  AO22XLTS U136 ( .A0(n493), .A1(n496), .B0(n495), .B1(n492), .Y(n1947) );
  OAI21XLTS U137 ( .A0(n87), .A1(n489), .B0(n490), .Y(n1949) );
  NAND4XLTS U138 ( .A(n872), .B(n871), .C(n870), .D(n869), .Y(n1975) );
  NAND4XLTS U139 ( .A(n848), .B(n847), .C(n846), .D(n845), .Y(n1974) );
  NAND4XLTS U140 ( .A(n836), .B(n835), .C(n834), .D(n833), .Y(n1973) );
  NAND4XLTS U141 ( .A(n824), .B(n823), .C(n822), .D(n821), .Y(n1972) );
  NAND4XLTS U142 ( .A(n805), .B(n804), .C(n803), .D(n802), .Y(n1971) );
  NAND4XLTS U143 ( .A(n785), .B(n784), .C(n783), .D(n782), .Y(n1970) );
  NAND4XLTS U144 ( .A(n655), .B(n654), .C(n653), .D(n652), .Y(n1961) );
  NAND4XLTS U145 ( .A(n643), .B(n642), .C(n641), .D(n640), .Y(n1960) );
  NAND4XLTS U146 ( .A(n624), .B(n623), .C(n622), .D(n621), .Y(n1959) );
  NAND4XLTS U147 ( .A(n609), .B(n608), .C(n607), .D(n606), .Y(n1958) );
  NAND4XLTS U148 ( .A(n598), .B(n597), .C(n596), .D(n652), .Y(n1957) );
  NAND4XLTS U149 ( .A(n587), .B(n586), .C(n585), .D(n640), .Y(n1956) );
  NAND4XLTS U150 ( .A(n579), .B(n578), .C(n577), .D(n621), .Y(n1955) );
  NAND4XLTS U151 ( .A(n562), .B(n561), .C(n560), .D(n606), .Y(n1954) );
  NAND4XLTS U152 ( .A(n540), .B(n539), .C(n538), .D(n559), .Y(n1952) );
  NAND3XLTS U153 ( .A(n775), .B(n774), .C(n773), .Y(n1969) );
  NAND3XLTS U154 ( .A(n761), .B(n760), .C(n759), .Y(n1968) );
  NAND3XLTS U155 ( .A(n746), .B(n745), .C(n744), .Y(n1967) );
  NAND3XLTS U156 ( .A(n728), .B(n727), .C(n726), .Y(n1966) );
  NAND3XLTS U157 ( .A(n714), .B(n713), .C(n712), .Y(n1965) );
  NAND3XLTS U158 ( .A(n703), .B(n702), .C(n701), .Y(n1964) );
  NAND3XLTS U159 ( .A(n688), .B(n687), .C(n686), .Y(n1963) );
  NAND3XLTS U160 ( .A(n666), .B(n665), .C(n664), .Y(n1962) );
  NAND3XLTS U161 ( .A(n553), .B(n552), .C(n551), .Y(n1953) );
  NAND3XLTS U162 ( .A(n1110), .B(n1109), .C(n1108), .Y(n2019) );
  NAND3XLTS U163 ( .A(n1105), .B(n1104), .C(n1103), .Y(n2018) );
  NAND3XLTS U164 ( .A(n1100), .B(n1099), .C(n1098), .Y(n2017) );
  NAND3XLTS U165 ( .A(n1095), .B(n1094), .C(n1093), .Y(n2016) );
  NAND3XLTS U166 ( .A(n1087), .B(n1086), .C(n1085), .Y(n2015) );
  NAND3XLTS U167 ( .A(n1082), .B(n1081), .C(n1080), .Y(n2014) );
  NAND3XLTS U168 ( .A(n1799), .B(n1798), .C(n1797), .Y(n2123) );
  NAND3XLTS U169 ( .A(n1790), .B(n1789), .C(n1788), .Y(n2122) );
  NAND3XLTS U170 ( .A(n1783), .B(n1782), .C(n1781), .Y(n2121) );
  NAND3XLTS U171 ( .A(n1776), .B(n1775), .C(n1774), .Y(n2120) );
  NAND3XLTS U172 ( .A(n978), .B(n977), .C(n976), .Y(n1995) );
  NAND3XLTS U173 ( .A(n971), .B(n970), .C(n969), .Y(n1994) );
  NAND3XLTS U174 ( .A(n963), .B(n962), .C(n961), .Y(n1993) );
  NAND3XLTS U175 ( .A(n954), .B(n953), .C(n952), .Y(n1992) );
  NAND3XLTS U176 ( .A(n1428), .B(n1427), .C(n1426), .Y(n2037) );
  NAND3XLTS U177 ( .A(n1422), .B(n1421), .C(n1420), .Y(n2036) );
  NAND3XLTS U178 ( .A(n1418), .B(n1417), .C(n1416), .Y(n2035) );
  NAND3XLTS U179 ( .A(n1414), .B(n1413), .C(n1412), .Y(n2034) );
  NAND3XLTS U180 ( .A(n1405), .B(n1404), .C(n1403), .Y(n2033) );
  NAND3XLTS U181 ( .A(n1400), .B(n1399), .C(n1398), .Y(n2032) );
  NAND3XLTS U182 ( .A(n1457), .B(n1456), .C(n1455), .Y(n2043) );
  NAND3XLTS U183 ( .A(n1453), .B(n1452), .C(n1451), .Y(n2042) );
  NAND3XLTS U184 ( .A(n1449), .B(n1448), .C(n1447), .Y(n2041) );
  NAND3XLTS U185 ( .A(n1443), .B(n1442), .C(n1441), .Y(n2040) );
  NAND3XLTS U186 ( .A(n1437), .B(n1436), .C(n1435), .Y(n2039) );
  NAND3XLTS U187 ( .A(n1433), .B(n1432), .C(n1431), .Y(n2038) );
  NAND3XLTS U188 ( .A(n1706), .B(n1705), .C(n1704), .Y(n2087) );
  NAND3XLTS U189 ( .A(n1700), .B(n1699), .C(n1698), .Y(n2086) );
  NAND3XLTS U190 ( .A(n1693), .B(n1692), .C(n1691), .Y(n2085) );
  NAND3XLTS U191 ( .A(n1685), .B(n1684), .C(n1683), .Y(n2084) );
  NAND3XLTS U192 ( .A(n907), .B(n906), .C(n905), .Y(n1983) );
  NAND3XLTS U193 ( .A(n901), .B(n900), .C(n899), .Y(n1982) );
  NAND3XLTS U194 ( .A(n898), .B(n897), .C(n896), .Y(n1981) );
  NAND3XLTS U195 ( .A(n893), .B(n892), .C(n891), .Y(n1980) );
  NAND3XLTS U196 ( .A(n1681), .B(n1680), .C(n1679), .Y(n2075) );
  NAND3XLTS U197 ( .A(n1673), .B(n1672), .C(n1671), .Y(n2074) );
  NAND3XLTS U198 ( .A(n1665), .B(n1664), .C(n1663), .Y(n2073) );
  NAND3XLTS U199 ( .A(n1658), .B(n1657), .C(n1656), .Y(n2072) );
  NAND3XLTS U200 ( .A(n890), .B(n889), .C(n888), .Y(n1979) );
  NAND3XLTS U201 ( .A(n885), .B(n884), .C(n883), .Y(n1978) );
  NAND3XLTS U202 ( .A(n880), .B(n879), .C(n878), .Y(n1977) );
  NAND3XLTS U203 ( .A(n877), .B(n876), .C(n875), .Y(n1976) );
  NAND3XLTS U204 ( .A(n1906), .B(n1905), .C(n1904), .Y(n2159) );
  NAND3XLTS U205 ( .A(n1897), .B(n1896), .C(n1895), .Y(n2158) );
  NAND3XLTS U206 ( .A(n1885), .B(n1884), .C(n1883), .Y(n2157) );
  NAND3XLTS U207 ( .A(n1875), .B(n1874), .C(n1873), .Y(n2156) );
  NAND3XLTS U208 ( .A(n1051), .B(n1050), .C(n1049), .Y(n2007) );
  NAND3XLTS U209 ( .A(n1044), .B(n1043), .C(n1042), .Y(n2006) );
  NAND3XLTS U210 ( .A(n1039), .B(n1038), .C(n1037), .Y(n2005) );
  NAND3XLTS U211 ( .A(n1033), .B(n1032), .C(n1031), .Y(n2004) );
  NAND3XLTS U212 ( .A(n1867), .B(n1866), .C(n1865), .Y(n2147) );
  NAND3XLTS U213 ( .A(n1859), .B(n1858), .C(n1857), .Y(n2146) );
  NAND3XLTS U214 ( .A(n1846), .B(n1845), .C(n1844), .Y(n2145) );
  NAND3XLTS U215 ( .A(n1835), .B(n1834), .C(n1833), .Y(n2144) );
  NAND3XLTS U216 ( .A(n1026), .B(n1025), .C(n1024), .Y(n2003) );
  NAND3XLTS U217 ( .A(n1017), .B(n1016), .C(n1015), .Y(n2002) );
  NAND3XLTS U218 ( .A(n1009), .B(n1008), .C(n1007), .Y(n2001) );
  NAND3XLTS U219 ( .A(n1002), .B(n1001), .C(n1000), .Y(n2000) );
  NAND3XLTS U220 ( .A(n1367), .B(n1366), .C(n1365), .Y(n2025) );
  NAND3XLTS U221 ( .A(n1362), .B(n1361), .C(n1360), .Y(n2024) );
  NAND3XLTS U222 ( .A(n1358), .B(n1357), .C(n1356), .Y(n2023) );
  NAND3XLTS U223 ( .A(n1352), .B(n1351), .C(n1350), .Y(n2022) );
  NAND3XLTS U224 ( .A(n1344), .B(n1343), .C(n1342), .Y(n2021) );
  NAND3XLTS U225 ( .A(n1339), .B(n1338), .C(n1337), .Y(n2020) );
  NAND3XLTS U226 ( .A(n1395), .B(n1394), .C(n1393), .Y(n2031) );
  NAND3XLTS U227 ( .A(n1390), .B(n1389), .C(n1388), .Y(n2030) );
  NAND3XLTS U228 ( .A(n1385), .B(n1384), .C(n1383), .Y(n2029) );
  NAND3XLTS U229 ( .A(n1382), .B(n1381), .C(n1380), .Y(n2028) );
  NAND3XLTS U230 ( .A(n1377), .B(n1376), .C(n1375), .Y(n2027) );
  NAND3XLTS U231 ( .A(n1371), .B(n1370), .C(n1369), .Y(n2026) );
  NAND3XLTS U232 ( .A(n1769), .B(n1768), .C(n1767), .Y(n2111) );
  NAND3XLTS U233 ( .A(n1763), .B(n1762), .C(n1761), .Y(n2110) );
  NAND3XLTS U234 ( .A(n1753), .B(n1752), .C(n1751), .Y(n2109) );
  NAND3XLTS U235 ( .A(n1745), .B(n1744), .C(n1743), .Y(n2108) );
  NAND3XLTS U236 ( .A(n948), .B(n947), .C(n946), .Y(n1991) );
  NAND3XLTS U237 ( .A(n941), .B(n940), .C(n939), .Y(n1990) );
  NAND3XLTS U238 ( .A(n936), .B(n935), .C(n934), .Y(n1989) );
  NAND3XLTS U239 ( .A(n930), .B(n929), .C(n928), .Y(n1988) );
  NAND3XLTS U240 ( .A(n1740), .B(n1739), .C(n1738), .Y(n2099) );
  NAND3XLTS U241 ( .A(n1732), .B(n1731), .C(n1730), .Y(n2098) );
  NAND3XLTS U242 ( .A(n1722), .B(n1721), .C(n1720), .Y(n2097) );
  NAND3XLTS U243 ( .A(n1713), .B(n1712), .C(n1711), .Y(n2096) );
  NAND3XLTS U244 ( .A(n923), .B(n922), .C(n921), .Y(n1987) );
  NAND3XLTS U245 ( .A(n918), .B(n917), .C(n916), .Y(n1986) );
  NAND3XLTS U246 ( .A(n915), .B(n914), .C(n913), .Y(n1985) );
  NAND3XLTS U247 ( .A(n911), .B(n910), .C(n909), .Y(n1984) );
  NAND3XLTS U248 ( .A(n1509), .B(n1508), .C(n1507), .Y(n2049) );
  NAND3XLTS U249 ( .A(n1500), .B(n1499), .C(n1498), .Y(n2048) );
  NAND3XLTS U250 ( .A(n1493), .B(n1492), .C(n1491), .Y(n2047) );
  NAND3XLTS U251 ( .A(n1485), .B(n1484), .C(n1483), .Y(n2046) );
  NAND3XLTS U252 ( .A(n1473), .B(n1472), .C(n1471), .Y(n2045) );
  NAND3XLTS U253 ( .A(n1465), .B(n1464), .C(n1463), .Y(n2044) );
  NAND3XLTS U254 ( .A(n1560), .B(n1559), .C(n1558), .Y(n2055) );
  NAND3XLTS U255 ( .A(n1551), .B(n1550), .C(n1549), .Y(n2054) );
  NAND3XLTS U256 ( .A(n1541), .B(n1540), .C(n1539), .Y(n2053) );
  NAND3XLTS U257 ( .A(n1534), .B(n1533), .C(n1532), .Y(n2052) );
  NAND3XLTS U258 ( .A(n1526), .B(n1525), .C(n1524), .Y(n2051) );
  NAND3XLTS U259 ( .A(n1518), .B(n1517), .C(n1516), .Y(n2050) );
  NAND3XLTS U260 ( .A(n1077), .B(n1076), .C(n1075), .Y(n2013) );
  NAND3XLTS U261 ( .A(n1073), .B(n1072), .C(n1071), .Y(n2012) );
  NAND3XLTS U262 ( .A(n1069), .B(n1068), .C(n1067), .Y(n2011) );
  NAND3XLTS U263 ( .A(n1066), .B(n1065), .C(n1064), .Y(n2010) );
  NAND3XLTS U264 ( .A(n1060), .B(n1059), .C(n1058), .Y(n2009) );
  NAND3XLTS U265 ( .A(n1055), .B(n1054), .C(n1053), .Y(n2008) );
  NAND3XLTS U266 ( .A(n1826), .B(n1825), .C(n1824), .Y(n2135) );
  NAND3XLTS U267 ( .A(n1821), .B(n1820), .C(n1819), .Y(n2134) );
  NAND3XLTS U268 ( .A(n1812), .B(n1811), .C(n1810), .Y(n2133) );
  NAND3XLTS U269 ( .A(n1805), .B(n1804), .C(n1803), .Y(n2132) );
  NAND3XLTS U270 ( .A(n994), .B(n993), .C(n992), .Y(n1999) );
  NAND3XLTS U271 ( .A(n989), .B(n988), .C(n987), .Y(n1998) );
  NAND3XLTS U272 ( .A(n986), .B(n985), .C(n984), .Y(n1997) );
  NAND3XLTS U273 ( .A(n982), .B(n981), .C(n980), .Y(n1996) );
  NOR2XLTS U274 ( .A(n1626), .B(n1623), .Y(n185) );
  INVX2TS U275 ( .A(n188), .Y(n215) );
  OR2X1TS U276 ( .A(n316), .B(n1003), .Y(n353) );
  CLKBUFX2TS U277 ( .A(n321), .Y(n322) );
  NOR2XLTS U278 ( .A(n1632), .B(n323), .Y(n321) );
  NAND2X1TS U279 ( .A(n31), .B(n28), .Y(n29) );
  OR2X1TS U280 ( .A(n1586), .B(n227), .Y(n2) );
  OR2X1TS U281 ( .A(n1596), .B(n279), .Y(n3) );
  OR2X1TS U282 ( .A(n1642), .B(n396), .Y(n4) );
  OR2X1TS U283 ( .A(n1573), .B(n93), .Y(n5) );
  OR2X1TS U284 ( .A(n1611), .B(n137), .Y(n6) );
  OR2X1TS U285 ( .A(n1617), .B(n189), .Y(n7) );
  OR2X1TS U286 ( .A(n1630), .B(n323), .Y(n8) );
  OR2X1TS U287 ( .A(n1597), .B(n279), .Y(n9) );
  OR2X1TS U288 ( .A(n1643), .B(n396), .Y(n10) );
  OA21XLTS U289 ( .A0(n311), .A1(n493), .B0(n25), .Y(n11) );
  OR2X1TS U290 ( .A(n24), .B(n505), .Y(n12) );
  NOR2XLTS U291 ( .A(n29), .B(n136), .Y(n133) );
  CLKBUFX2TS U292 ( .A(n187), .Y(n188) );
  OR2X1TS U293 ( .A(n481), .B(n1627), .Y(n13) );
  OR2X1TS U294 ( .A(n391), .B(n1034), .Y(n422) );
  NOR3XLTS U295 ( .A(n1639), .B(n1633), .C(n320), .Y(n313) );
  NOR3XLTS U296 ( .A(n1650), .B(n1644), .C(n394), .Y(n390) );
  NOR3XLTS U297 ( .A(n1579), .B(n1574), .C(n91), .Y(n86) );
  NOR3XLTS U298 ( .A(n1604), .B(n1598), .C(n277), .Y(n272) );
  NOR3XLTS U299 ( .A(n1626), .B(n1620), .C(n186), .Y(n183) );
  NOR3XLTS U300 ( .A(n1568), .B(n1563), .C(n40), .Y(n34) );
  OR2X1TS U301 ( .A(n440), .B(n1593), .Y(n14) );
  OR2X1TS U302 ( .A(n481), .B(n1651), .Y(n15) );
  NOR2XLTS U303 ( .A(n843), .B(n517), .Y(n690) );
  NOR2XLTS U304 ( .A(n843), .B(n516), .Y(n542) );
  INVX2TS U305 ( .A(destinationAddressIn_EAST[5]), .Y(n64) );
  INVX2TS U306 ( .A(destinationAddressIn_EAST[6]), .Y(n75) );
  INVX2TS U307 ( .A(destinationAddressIn_EAST[4]), .Y(n72) );
  INVX2TS U308 ( .A(destinationAddressIn_EAST[7]), .Y(n67) );
  INVX2TS U309 ( .A(destinationAddressIn_EAST[9]), .Y(n44) );
  INVX2TS U310 ( .A(destinationAddressIn_EAST[8]), .Y(n49) );
  INVX2TS U311 ( .A(destinationAddressIn_EAST[10]), .Y(n52) );
  INVX2TS U312 ( .A(destinationAddressIn_EAST[11]), .Y(n35) );
  INVX2TS U313 ( .A(writeIn_EAST), .Y(n57) );
  CLKBUFX2TS U314 ( .A(n1928), .Y(n16) );
  INVX2TS U330 ( .A(n1935), .Y(n85) );
  INVX2TS U331 ( .A(n1931), .Y(n442) );
  INVX2TS U332 ( .A(n18), .Y(n81) );
  INVX2TS U333 ( .A(n81), .Y(n126) );
  INVX2TS U334 ( .A(selectBit_WEST), .Y(n446) );
  INVX2TS U335 ( .A(n1566), .Y(n1568) );
  INVX2TS U336 ( .A(n1927), .Y(n449) );
  INVX2TS U337 ( .A(n21), .Y(n22) );
  INVX2TS U338 ( .A(n22), .Y(n311) );
  INVX2TS U339 ( .A(selectBit_SOUTH), .Y(n505) );
  INVX2TS U340 ( .A(n12), .Y(n220) );
  INVX2TS U341 ( .A(n1935), .Y(n493) );
  INVX2TS U342 ( .A(n1935), .Y(n483) );
  NAND2X1TS U343 ( .A(n21), .B(n483), .Y(n25) );
  INVX2TS U344 ( .A(n11), .Y(n82) );
  INVX2TS U345 ( .A(n505), .Y(n504) );
  NAND2X1TS U346 ( .A(n504), .B(n24), .Y(n23) );
  OAI21XLTS U347 ( .A0(selectBit_SOUTH), .A1(n24), .B0(n83), .Y(n267) );
  NAND2X1TS U348 ( .A(n309), .B(n267), .Y(n129) );
  INVX2TS U349 ( .A(selectBit_EAST), .Y(n512) );
  INVX2TS U350 ( .A(n512), .Y(n510) );
  INVX2TS U351 ( .A(n1933), .Y(n271) );
  INVX2TS U352 ( .A(n1932), .Y(n443) );
  AOI22X1TS U353 ( .A0(n271), .A1(n25), .B0(n130), .B1(n443), .Y(n26) );
  INVX2TS U354 ( .A(n26), .Y(n27) );
  INVX2TS U355 ( .A(n27), .Y(n28) );
  INVX2TS U356 ( .A(n29), .Y(n125) );
  INVX2TS U357 ( .A(n125), .Y(n30) );
  NAND2X1TS U358 ( .A(n510), .B(n128), .Y(n268) );
  NAND2X1TS U359 ( .A(n444), .B(n130), .Y(n33) );
  INVX2TS U360 ( .A(n28), .Y(n32) );
  INVX2TS U361 ( .A(n446), .Y(n511) );
  INVX2TS U362 ( .A(readReady), .Y(n182) );
  INVX2TS U363 ( .A(n182), .Y(n513) );
  NAND2X1TS U364 ( .A(n537), .B(n506), .Y(n522) );
  INVX2TS U365 ( .A(n273), .Y(n314) );
  INVX2TS U366 ( .A(n314), .Y(n87) );
  INVX2TS U367 ( .A(n87), .Y(n180) );
  AOI31XLTS U368 ( .A0(n39), .A1(n33), .A2(n1561), .B0(n180), .Y(n37) );
  INVX2TS U369 ( .A(n182), .Y(n508) );
  NAND2X1TS U370 ( .A(n37), .B(n1569), .Y(n40) );
  INVX2TS U371 ( .A(n34), .Y(n887) );
  INVX2TS U372 ( .A(n887), .Y(n1668) );
  CLKBUFX2TS U373 ( .A(n1668), .Y(n48) );
  INVX2TS U374 ( .A(n48), .Y(n71) );
  INVX2TS U375 ( .A(destinationAddressIn_EAST[11]), .Y(n244) );
  INVX2TS U376 ( .A(n36), .Y(n886) );
  INVX2TS U377 ( .A(n886), .Y(n1653) );
  INVX2TS U378 ( .A(n1527), .Y(n53) );
  OR2X1TS U379 ( .A(n1566), .B(n40), .Y(n58) );
  INVX2TS U380 ( .A(n58), .Y(n1669) );
  INVX2TS U381 ( .A(n1669), .Y(n881) );
  INVX2TS U382 ( .A(n881), .Y(n38) );
  CLKBUFX2TS U383 ( .A(destinationAddressIn_WEST[11]), .Y(n410) );
  CLKBUFX2TS U384 ( .A(n410), .Y(n762) );
  AOI22X1TS U385 ( .A0(n53), .A1(\destinationAddressbuffer[7][11] ), .B0(n38), 
        .B1(n762), .Y(n43) );
  INVX2TS U386 ( .A(n45), .Y(n60) );
  INVX2TS U387 ( .A(n60), .Y(n1548) );
  INVX2TS U388 ( .A(n144), .Y(n765) );
  OR2X1TS U389 ( .A(n1562), .B(n41), .Y(n68) );
  INVX2TS U390 ( .A(n68), .Y(n1514) );
  CLKBUFX2TS U391 ( .A(destinationAddressIn_NORTH[11]), .Y(n766) );
  CLKBUFX2TS U392 ( .A(n766), .Y(n337) );
  AOI22X1TS U393 ( .A0(n1548), .A1(n765), .B0(n1514), .B1(n337), .Y(n42) );
  OAI211XLTS U394 ( .A0(n71), .A1(n244), .B0(n43), .C0(n42), .Y(n2083) );
  INVX2TS U395 ( .A(destinationAddressIn_EAST[9]), .Y(n234) );
  INVX2TS U396 ( .A(n881), .Y(n76) );
  CLKBUFX2TS U397 ( .A(destinationAddressIn_WEST[9]), .Y(n392) );
  CLKBUFX2TS U398 ( .A(n392), .Y(n730) );
  AOI22X1TS U399 ( .A0(n53), .A1(\destinationAddressbuffer[7][9] ), .B0(n76), 
        .B1(n730), .Y(n47) );
  INVX2TS U400 ( .A(n45), .Y(n873) );
  INVX2TS U401 ( .A(n873), .Y(n1662) );
  INVX2TS U402 ( .A(n154), .Y(n731) );
  INVX2TS U403 ( .A(n1514), .Y(n874) );
  INVX2TS U404 ( .A(n874), .Y(n882) );
  CLKBUFX2TS U405 ( .A(destinationAddressIn_NORTH[9]), .Y(n733) );
  CLKBUFX2TS U406 ( .A(n733), .Y(n344) );
  AOI22X1TS U407 ( .A0(n1662), .A1(n731), .B0(n882), .B1(n344), .Y(n46) );
  OAI211XLTS U408 ( .A0(n71), .A1(n234), .B0(n47), .C0(n46), .Y(n2081) );
  INVX2TS U409 ( .A(n48), .Y(n80) );
  INVX2TS U410 ( .A(destinationAddressIn_EAST[8]), .Y(n231) );
  INVX2TS U411 ( .A(n58), .Y(n1655) );
  CLKBUFX2TS U412 ( .A(destinationAddressIn_WEST[8]), .Y(n400) );
  CLKBUFX2TS U413 ( .A(n400), .Y(n715) );
  AOI22X1TS U414 ( .A0(n53), .A1(\destinationAddressbuffer[7][8] ), .B0(n1655), 
        .B1(n715), .Y(n51) );
  INVX2TS U415 ( .A(n60), .Y(n1670) );
  INVX2TS U416 ( .A(n140), .Y(n716) );
  INVX2TS U417 ( .A(n68), .Y(n1546) );
  CLKBUFX2TS U418 ( .A(destinationAddressIn_NORTH[8]), .Y(n717) );
  CLKBUFX2TS U419 ( .A(n717), .Y(n325) );
  AOI22X1TS U420 ( .A0(n1670), .A1(n716), .B0(n1546), .B1(n325), .Y(n50) );
  OAI211XLTS U421 ( .A0(n80), .A1(n231), .B0(n51), .C0(n50), .Y(n2080) );
  INVX2TS U422 ( .A(destinationAddressIn_EAST[10]), .Y(n238) );
  INVX2TS U423 ( .A(n58), .Y(n1512) );
  CLKBUFX2TS U424 ( .A(destinationAddressIn_WEST[10]), .Y(n405) );
  CLKBUFX2TS U425 ( .A(n405), .Y(n747) );
  AOI22X1TS U426 ( .A0(n53), .A1(\destinationAddressbuffer[7][10] ), .B0(n1512), .B1(n747), .Y(n56) );
  INVX2TS U427 ( .A(n60), .Y(n54) );
  INVX2TS U428 ( .A(n148), .Y(n750) );
  CLKBUFX2TS U429 ( .A(destinationAddressIn_NORTH[10]), .Y(n751) );
  CLKBUFX2TS U430 ( .A(n751), .Y(n330) );
  AOI22X1TS U431 ( .A0(n54), .A1(n750), .B0(n1546), .B1(n330), .Y(n55) );
  OAI211XLTS U432 ( .A0(n71), .A1(n238), .B0(n56), .C0(n55), .Y(n2082) );
  INVX2TS U433 ( .A(writeIn_EAST), .Y(n249) );
  INVX2TS U434 ( .A(n1570), .Y(n1674) );
  INVX2TS U435 ( .A(n58), .Y(n59) );
  CLKBUFX2TS U436 ( .A(writeIn_WEST), .Y(n418) );
  CLKBUFX2TS U437 ( .A(n418), .Y(n541) );
  AOI22X1TS U438 ( .A0(n1674), .A1(writeOutbuffer[7]), .B0(n59), .B1(n541), 
        .Y(n63) );
  INVX2TS U439 ( .A(n60), .Y(n1678) );
  INVX2TS U440 ( .A(writeIn_SOUTH), .Y(n157) );
  INVX2TS U441 ( .A(n157), .Y(n543) );
  INVX2TS U442 ( .A(n68), .Y(n61) );
  CLKBUFX2TS U443 ( .A(writeIn_NORTH), .Y(n544) );
  CLKBUFX2TS U444 ( .A(n544), .Y(n350) );
  AOI22X1TS U445 ( .A0(n1678), .A1(n543), .B0(n61), .B1(n350), .Y(n62) );
  OAI211XLTS U446 ( .A0(n80), .A1(n249), .B0(n63), .C0(n62), .Y(n2056) );
  INVX2TS U447 ( .A(destinationAddressIn_EAST[5]), .Y(n260) );
  INVX2TS U448 ( .A(n1527), .Y(n77) );
  AOI22X1TS U449 ( .A0(n77), .A1(\destinationAddressbuffer[7][5] ), .B0(n59), 
        .B1(destinationAddressIn_WEST[5]), .Y(n66) );
  INVX2TS U450 ( .A(destinationAddressIn_SOUTH[5]), .Y(n160) );
  INVX2TS U451 ( .A(n160), .Y(n671) );
  AOI22X1TS U452 ( .A0(n1678), .A1(n671), .B0(n61), .B1(
        destinationAddressIn_NORTH[5]), .Y(n65) );
  OAI211XLTS U453 ( .A0(n80), .A1(n260), .B0(n66), .C0(n65), .Y(n2077) );
  INVX2TS U454 ( .A(destinationAddressIn_EAST[7]), .Y(n252) );
  AOI22X1TS U455 ( .A0(n77), .A1(\destinationAddressbuffer[7][7] ), .B0(n1655), 
        .B1(destinationAddressIn_WEST[7]), .Y(n70) );
  INVX2TS U456 ( .A(destinationAddressIn_SOUTH[7]), .Y(n165) );
  INVX2TS U457 ( .A(n165), .Y(n705) );
  INVX2TS U458 ( .A(n68), .Y(n1661) );
  AOI22X1TS U459 ( .A0(n54), .A1(n705), .B0(n1661), .B1(
        destinationAddressIn_NORTH[7]), .Y(n69) );
  OAI211XLTS U460 ( .A0(n71), .A1(n252), .B0(n70), .C0(n69), .Y(n2079) );
  INVX2TS U461 ( .A(destinationAddressIn_EAST[4]), .Y(n256) );
  AOI22X1TS U462 ( .A0(n77), .A1(\destinationAddressbuffer[7][4] ), .B0(n1512), 
        .B1(destinationAddressIn_WEST[4]), .Y(n74) );
  INVX2TS U463 ( .A(destinationAddressIn_SOUTH[4]), .Y(n178) );
  INVX2TS U464 ( .A(n178), .Y(n658) );
  AOI22X1TS U465 ( .A0(n1548), .A1(n658), .B0(n1661), .B1(
        destinationAddressIn_NORTH[4]), .Y(n73) );
  OAI211XLTS U466 ( .A0(n887), .A1(n256), .B0(n74), .C0(n73), .Y(n2076) );
  INVX2TS U467 ( .A(destinationAddressIn_EAST[6]), .Y(n264) );
  AOI22X1TS U468 ( .A0(n77), .A1(\destinationAddressbuffer[7][6] ), .B0(n76), 
        .B1(destinationAddressIn_WEST[6]), .Y(n79) );
  INVX2TS U469 ( .A(destinationAddressIn_SOUTH[6]), .Y(n170) );
  INVX2TS U470 ( .A(n170), .Y(n691) );
  AOI22X1TS U471 ( .A0(n1670), .A1(n691), .B0(n882), .B1(
        destinationAddressIn_NORTH[6]), .Y(n78) );
  OAI211XLTS U472 ( .A0(n80), .A1(n264), .B0(n79), .C0(n78), .Y(n2078) );
  INVX2TS U473 ( .A(n17), .Y(n179) );
  NAND2X1TS U474 ( .A(n127), .B(n451), .Y(n266) );
  AOI21X1TS U475 ( .A0(n220), .A1(n82), .B0(n309), .Y(n382) );
  NOR3XLTS U476 ( .A(n382), .B(n268), .C(n267), .Y(n1576) );
  INVX2TS U477 ( .A(n1935), .Y(n486) );
  NOR2XLTS U478 ( .A(n442), .B(n503), .Y(n385) );
  INVX2TS U479 ( .A(n11), .Y(n269) );
  NOR3XLTS U480 ( .A(n26), .B(n83), .C(n269), .Y(n1573) );
  AOI31XLTS U481 ( .A0(n271), .A1(n486), .A2(n385), .B0(n1573), .Y(n84) );
  AOI21X1TS U482 ( .A0(n90), .A1(n84), .B0(n314), .Y(n89) );
  INVX2TS U483 ( .A(n1927), .Y(n389) );
  NAND2X1TS U484 ( .A(n89), .B(n1580), .Y(n91) );
  INVX2TS U485 ( .A(n86), .Y(n1459) );
  INVX2TS U486 ( .A(n1459), .Y(n903) );
  CLKBUFX2TS U487 ( .A(n903), .Y(n100) );
  INVX2TS U488 ( .A(n100), .Y(n118) );
  INVX2TS U489 ( .A(n87), .Y(n481) );
  INVX2TS U490 ( .A(n88), .Y(n1474) );
  INVX2TS U491 ( .A(n1474), .Y(n894) );
  INVX2TS U492 ( .A(n1475), .Y(n103) );
  OR2X1TS U493 ( .A(n1577), .B(n91), .Y(n108) );
  INVX2TS U494 ( .A(n108), .Y(n1478) );
  AOI22X1TS U495 ( .A0(n103), .A1(\destinationAddressbuffer[6][11] ), .B0(n115), .B1(n762), .Y(n97) );
  INVX2TS U496 ( .A(n5), .Y(n92) );
  INVX2TS U497 ( .A(n92), .Y(n104) );
  INVX2TS U498 ( .A(n104), .Y(n1482) );
  CLKBUFX2TS U499 ( .A(n766), .Y(n412) );
  INVX2TS U500 ( .A(n94), .Y(n105) );
  INVX2TS U501 ( .A(n105), .Y(n95) );
  INVX2TS U502 ( .A(n95), .Y(n904) );
  INVX2TS U503 ( .A(n904), .Y(n112) );
  INVX2TS U504 ( .A(n144), .Y(n336) );
  AOI22X1TS U505 ( .A0(n1482), .A1(n412), .B0(n112), .B1(n336), .Y(n96) );
  OAI211XLTS U506 ( .A0(n118), .A1(n244), .B0(n97), .C0(n96), .Y(n2095) );
  INVX2TS U507 ( .A(n108), .Y(n1488) );
  AOI22X1TS U508 ( .A0(n103), .A1(\destinationAddressbuffer[6][8] ), .B0(n1488), .B1(n715), .Y(n99) );
  INVX2TS U509 ( .A(n5), .Y(n1682) );
  CLKBUFX2TS U510 ( .A(n717), .Y(n401) );
  INVX2TS U511 ( .A(n105), .Y(n1505) );
  INVX2TS U512 ( .A(n140), .Y(n324) );
  AOI22X1TS U513 ( .A0(n1682), .A1(n401), .B0(n1505), .B1(n324), .Y(n98) );
  OAI211XLTS U514 ( .A0(n118), .A1(n231), .B0(n99), .C0(n98), .Y(n2092) );
  INVX2TS U515 ( .A(n100), .Y(n124) );
  AOI22X1TS U516 ( .A0(n103), .A1(\destinationAddressbuffer[6][9] ), .B0(n109), 
        .B1(n730), .Y(n102) );
  CLKBUFX2TS U517 ( .A(n733), .Y(n397) );
  INVX2TS U518 ( .A(n105), .Y(n1689) );
  INVX2TS U519 ( .A(n154), .Y(n343) );
  AOI22X1TS U520 ( .A0(n1482), .A1(n397), .B0(n1689), .B1(n343), .Y(n101) );
  OAI211XLTS U521 ( .A0(n124), .A1(n234), .B0(n102), .C0(n101), .Y(n2093) );
  INVX2TS U522 ( .A(n108), .Y(n1688) );
  AOI22X1TS U523 ( .A0(n103), .A1(\destinationAddressbuffer[6][10] ), .B0(
        n1688), .B1(n747), .Y(n107) );
  INVX2TS U524 ( .A(n104), .Y(n895) );
  CLKBUFX2TS U525 ( .A(n751), .Y(n407) );
  INVX2TS U526 ( .A(n105), .Y(n1703) );
  INVX2TS U527 ( .A(n148), .Y(n329) );
  AOI22X1TS U528 ( .A0(n895), .A1(n407), .B0(n112), .B1(n329), .Y(n106) );
  OAI211XLTS U529 ( .A0(n118), .A1(n238), .B0(n107), .C0(n106), .Y(n2094) );
  INVX2TS U530 ( .A(n1581), .Y(n1701) );
  INVX2TS U531 ( .A(n108), .Y(n109) );
  INVX2TS U532 ( .A(n109), .Y(n902) );
  INVX2TS U533 ( .A(n902), .Y(n115) );
  AOI22X1TS U534 ( .A0(n1701), .A1(writeOutbuffer[6]), .B0(n115), .B1(n541), 
        .Y(n111) );
  INVX2TS U535 ( .A(n5), .Y(n1697) );
  CLKBUFX2TS U536 ( .A(n544), .Y(n419) );
  INVX2TS U537 ( .A(n157), .Y(n348) );
  AOI22X1TS U538 ( .A0(n1697), .A1(n419), .B0(n1505), .B1(n348), .Y(n110) );
  OAI211XLTS U539 ( .A0(n124), .A1(n249), .B0(n111), .C0(n110), .Y(n2057) );
  INVX2TS U540 ( .A(n1581), .Y(n121) );
  AOI22X1TS U541 ( .A0(n121), .A1(\destinationAddressbuffer[6][6] ), .B0(n1478), .B1(destinationAddressIn_WEST[6]), .Y(n114) );
  CLKBUFX2TS U542 ( .A(destinationAddressIn_NORTH[6]), .Y(n356) );
  CLKBUFX2TS U543 ( .A(n356), .Y(n428) );
  INVX2TS U544 ( .A(n170), .Y(n355) );
  AOI22X1TS U545 ( .A0(n895), .A1(n428), .B0(n112), .B1(n355), .Y(n113) );
  OAI211XLTS U546 ( .A0(n124), .A1(n264), .B0(n114), .C0(n113), .Y(n2090) );
  AOI22X1TS U547 ( .A0(n121), .A1(\destinationAddressbuffer[6][5] ), .B0(n115), 
        .B1(destinationAddressIn_WEST[5]), .Y(n117) );
  INVX2TS U548 ( .A(n5), .Y(n1690) );
  CLKBUFX2TS U549 ( .A(destinationAddressIn_NORTH[5]), .Y(n375) );
  CLKBUFX2TS U550 ( .A(n375), .Y(n424) );
  INVX2TS U551 ( .A(n160), .Y(n374) );
  AOI22X1TS U552 ( .A0(n1690), .A1(n424), .B0(n1703), .B1(n374), .Y(n116) );
  OAI211XLTS U553 ( .A0(n118), .A1(n260), .B0(n117), .C0(n116), .Y(n2089) );
  AOI22X1TS U554 ( .A0(n121), .A1(\destinationAddressbuffer[6][7] ), .B0(n1488), .B1(destinationAddressIn_WEST[7]), .Y(n120) );
  CLKBUFX2TS U555 ( .A(destinationAddressIn_NORTH[7]), .Y(n369) );
  CLKBUFX2TS U556 ( .A(n369), .Y(n436) );
  INVX2TS U557 ( .A(n165), .Y(n368) );
  AOI22X1TS U558 ( .A0(n1690), .A1(n436), .B0(n1703), .B1(n368), .Y(n119) );
  OAI211XLTS U559 ( .A0(n1459), .A1(n252), .B0(n120), .C0(n119), .Y(n2091) );
  AOI22X1TS U560 ( .A0(n121), .A1(\destinationAddressbuffer[6][4] ), .B0(n1688), .B1(destinationAddressIn_WEST[4]), .Y(n123) );
  CLKBUFX2TS U561 ( .A(destinationAddressIn_NORTH[4]), .Y(n363) );
  CLKBUFX2TS U562 ( .A(n363), .Y(n432) );
  INVX2TS U563 ( .A(n178), .Y(n362) );
  AOI22X1TS U564 ( .A0(n1682), .A1(n432), .B0(n1689), .B1(n362), .Y(n122) );
  OAI211XLTS U565 ( .A0(n124), .A1(n256), .B0(n123), .C0(n122), .Y(n2088) );
  INVX2TS U566 ( .A(n1932), .Y(n482) );
  NAND2X1TS U567 ( .A(n130), .B(n482), .Y(n131) );
  AOI31XLTS U568 ( .A0(n132), .A1(n30), .A2(n131), .B0(n481), .Y(n135) );
  INVX2TS U569 ( .A(n1931), .Y(n473) );
  INVX2TS U570 ( .A(n182), .Y(n509) );
  INVX2TS U571 ( .A(n1932), .Y(n485) );
  INVX2TS U572 ( .A(n133), .Y(n966) );
  INVX2TS U573 ( .A(n966), .Y(n1374) );
  CLKBUFX2TS U574 ( .A(n1374), .Y(n145) );
  INVX2TS U575 ( .A(n145), .Y(n166) );
  INVX2TS U576 ( .A(n134), .Y(n1378) );
  INVX2TS U577 ( .A(n1378), .Y(n956) );
  INVX2TS U578 ( .A(n1615), .Y(n150) );
  NOR3XLTS U579 ( .A(n1613), .B(n1608), .C(n137), .Y(n149) );
  INVX2TS U580 ( .A(n149), .Y(n172) );
  INVX2TS U581 ( .A(n172), .Y(n1368) );
  AOI22X1TS U582 ( .A0(n150), .A1(\destinationAddressbuffer[3][8] ), .B0(n1368), .B1(destinationAddressIn_EAST[8]), .Y(n139) );
  NOR2XLTS U583 ( .A(n125), .B(n136), .Y(n151) );
  INVX2TS U584 ( .A(n151), .Y(n161) );
  INVX2TS U585 ( .A(n161), .Y(n1787) );
  INVX2TS U586 ( .A(n6), .Y(n1387) );
  CLKBUFX2TS U587 ( .A(n400), .Y(n318) );
  AOI22X1TS U588 ( .A0(n1787), .A1(n325), .B0(n1387), .B1(n318), .Y(n138) );
  OAI211XLTS U589 ( .A0(n166), .A1(n140), .B0(n139), .C0(n138), .Y(n2128) );
  INVX2TS U590 ( .A(n145), .Y(n171) );
  INVX2TS U591 ( .A(n172), .Y(n1778) );
  AOI22X1TS U592 ( .A0(n150), .A1(\destinationAddressbuffer[3][11] ), .B0(
        n1778), .B1(destinationAddressIn_EAST[11]), .Y(n143) );
  INVX2TS U593 ( .A(n161), .Y(n1773) );
  INVX2TS U594 ( .A(n6), .Y(n141) );
  CLKBUFX2TS U595 ( .A(n410), .Y(n334) );
  AOI22X1TS U596 ( .A0(n1773), .A1(n337), .B0(n141), .B1(n334), .Y(n142) );
  OAI211XLTS U597 ( .A0(n171), .A1(n144), .B0(n143), .C0(n142), .Y(n2131) );
  AOI22X1TS U598 ( .A0(n150), .A1(\destinationAddressbuffer[3][10] ), .B0(
        n1368), .B1(destinationAddressIn_EAST[10]), .Y(n147) );
  INVX2TS U599 ( .A(n161), .Y(n1780) );
  INVX2TS U600 ( .A(n6), .Y(n1772) );
  CLKBUFX2TS U601 ( .A(n405), .Y(n328) );
  AOI22X1TS U602 ( .A0(n1780), .A1(n330), .B0(n1772), .B1(n328), .Y(n146) );
  OAI211XLTS U603 ( .A0(n966), .A1(n148), .B0(n147), .C0(n146), .Y(n2130) );
  INVX2TS U604 ( .A(n149), .Y(n957) );
  INVX2TS U605 ( .A(n957), .Y(n167) );
  AOI22X1TS U606 ( .A0(n150), .A1(\destinationAddressbuffer[3][9] ), .B0(n167), 
        .B1(destinationAddressIn_EAST[9]), .Y(n153) );
  INVX2TS U607 ( .A(n151), .Y(n1373) );
  INVX2TS U608 ( .A(n1373), .Y(n967) );
  INVX2TS U609 ( .A(n1387), .Y(n973) );
  INVX2TS U610 ( .A(n973), .Y(n958) );
  CLKBUFX2TS U611 ( .A(n392), .Y(n341) );
  AOI22X1TS U612 ( .A0(n967), .A1(n344), .B0(n958), .B1(n341), .Y(n152) );
  OAI211XLTS U613 ( .A0(n166), .A1(n154), .B0(n153), .C0(n152), .Y(n2129) );
  INVX2TS U614 ( .A(n1615), .Y(n1791) );
  INVX2TS U615 ( .A(n172), .Y(n1386) );
  AOI22X1TS U616 ( .A0(n1791), .A1(writeOutbuffer[3]), .B0(n1386), .B1(
        writeIn_EAST), .Y(n156) );
  INVX2TS U617 ( .A(n6), .Y(n1795) );
  CLKBUFX2TS U618 ( .A(n418), .Y(n347) );
  AOI22X1TS U619 ( .A0(n1780), .A1(n350), .B0(n1795), .B1(n347), .Y(n155) );
  OAI211XLTS U620 ( .A0(n171), .A1(n157), .B0(n156), .C0(n155), .Y(n2060) );
  INVX2TS U621 ( .A(n1379), .Y(n174) );
  AOI22X1TS U622 ( .A0(n174), .A1(\destinationAddressbuffer[3][5] ), .B0(n1778), .B1(destinationAddressIn_EAST[5]), .Y(n159) );
  CLKBUFX2TS U623 ( .A(destinationAddressIn_WEST[5]), .Y(n669) );
  CLKBUFX2TS U624 ( .A(n669), .Y(n372) );
  AOI22X1TS U625 ( .A0(n967), .A1(n375), .B0(n141), .B1(n372), .Y(n158) );
  OAI211XLTS U626 ( .A0(n166), .A1(n160), .B0(n159), .C0(n158), .Y(n2125) );
  AOI22X1TS U627 ( .A0(n174), .A1(\destinationAddressbuffer[3][7] ), .B0(n1386), .B1(destinationAddressIn_EAST[7]), .Y(n164) );
  INVX2TS U628 ( .A(n161), .Y(n162) );
  CLKBUFX2TS U629 ( .A(destinationAddressIn_WEST[7]), .Y(n704) );
  CLKBUFX2TS U630 ( .A(n704), .Y(n367) );
  AOI22X1TS U631 ( .A0(n162), .A1(n369), .B0(n1795), .B1(n367), .Y(n163) );
  OAI211XLTS U632 ( .A0(n166), .A1(n165), .B0(n164), .C0(n163), .Y(n2127) );
  AOI22X1TS U633 ( .A0(n174), .A1(\destinationAddressbuffer[3][6] ), .B0(n167), 
        .B1(destinationAddressIn_EAST[6]), .Y(n169) );
  CLKBUFX2TS U634 ( .A(destinationAddressIn_WEST[6]), .Y(n689) );
  CLKBUFX2TS U635 ( .A(n689), .Y(n354) );
  AOI22X1TS U636 ( .A0(n162), .A1(n356), .B0(n1772), .B1(n354), .Y(n168) );
  OAI211XLTS U637 ( .A0(n171), .A1(n170), .B0(n169), .C0(n168), .Y(n2126) );
  INVX2TS U638 ( .A(n172), .Y(n173) );
  AOI22X1TS U639 ( .A0(n174), .A1(\destinationAddressbuffer[3][4] ), .B0(n167), 
        .B1(destinationAddressIn_EAST[4]), .Y(n177) );
  INVX2TS U640 ( .A(n973), .Y(n175) );
  CLKBUFX2TS U641 ( .A(destinationAddressIn_WEST[4]), .Y(n656) );
  CLKBUFX2TS U642 ( .A(n656), .Y(n359) );
  AOI22X1TS U643 ( .A0(n1773), .A1(n363), .B0(n175), .B1(n359), .Y(n176) );
  OAI211XLTS U644 ( .A0(n171), .A1(n178), .B0(n177), .C0(n176), .Y(n2124) );
  INVX2TS U645 ( .A(n267), .Y(n310) );
  INVX2TS U646 ( .A(n310), .Y(n380) );
  NOR3XLTS U647 ( .A(n382), .B(n380), .C(n381), .Y(n1623) );
  AOI31XLTS U648 ( .A0(n493), .A1(n385), .A2(n443), .B0(n1619), .Y(n181) );
  AOI21X1TS U649 ( .A0(n185), .A1(n181), .B0(n180), .Y(n184) );
  NAND2X1TS U650 ( .A(n184), .B(n1627), .Y(n186) );
  INVX2TS U651 ( .A(n183), .Y(n1346) );
  INVX2TS U652 ( .A(n1346), .Y(n991) );
  CLKBUFX2TS U653 ( .A(n991), .Y(n195) );
  INVX2TS U654 ( .A(n195), .Y(n211) );
  INVX2TS U655 ( .A(n13), .Y(n983) );
  INVX2TS U656 ( .A(n1345), .Y(n200) );
  OR2X1TS U657 ( .A(n1624), .B(n186), .Y(n198) );
  INVX2TS U658 ( .A(n198), .Y(n1816) );
  AOI22X1TS U659 ( .A0(n200), .A1(\destinationAddressbuffer[2][11] ), .B0(
        n1816), .B1(n334), .Y(n192) );
  INVX2TS U660 ( .A(n215), .Y(n1355) );
  INVX2TS U661 ( .A(n7), .Y(n190) );
  INVX2TS U662 ( .A(n190), .Y(n979) );
  INVX2TS U663 ( .A(n979), .Y(n203) );
  AOI22X1TS U664 ( .A0(n1355), .A1(n337), .B0(n203), .B1(n336), .Y(n191) );
  OAI211XLTS U665 ( .A0(n211), .A1(n244), .B0(n192), .C0(n191), .Y(n2143) );
  INVX2TS U666 ( .A(n198), .Y(n1800) );
  AOI22X1TS U667 ( .A0(n200), .A1(\destinationAddressbuffer[2][9] ), .B0(n1800), .B1(n341), .Y(n194) );
  INVX2TS U668 ( .A(n7), .Y(n1354) );
  AOI22X1TS U669 ( .A0(n187), .A1(n344), .B0(n1354), .B1(n343), .Y(n193) );
  OAI211XLTS U670 ( .A0(n211), .A1(n234), .B0(n194), .C0(n193), .Y(n2141) );
  INVX2TS U671 ( .A(n195), .Y(n218) );
  INVX2TS U672 ( .A(n198), .Y(n1808) );
  AOI22X1TS U673 ( .A0(n200), .A1(\destinationAddressbuffer[2][10] ), .B0(
        n1808), .B1(n328), .Y(n197) );
  INVX2TS U674 ( .A(n215), .Y(n1112) );
  INVX2TS U675 ( .A(n7), .Y(n1801) );
  AOI22X1TS U676 ( .A0(n1112), .A1(n330), .B0(n1801), .B1(n329), .Y(n196) );
  OAI211XLTS U677 ( .A0(n218), .A1(n238), .B0(n197), .C0(n196), .Y(n2142) );
  INVX2TS U678 ( .A(n198), .Y(n199) );
  INVX2TS U679 ( .A(n199), .Y(n990) );
  INVX2TS U680 ( .A(n990), .Y(n208) );
  AOI22X1TS U681 ( .A0(n200), .A1(\destinationAddressbuffer[2][8] ), .B0(n208), 
        .B1(n318), .Y(n202) );
  INVX2TS U682 ( .A(n7), .Y(n1809) );
  AOI22X1TS U683 ( .A0(n1112), .A1(n325), .B0(n1809), .B1(n324), .Y(n201) );
  OAI211XLTS U684 ( .A0(n211), .A1(n231), .B0(n202), .C0(n201), .Y(n2140) );
  INVX2TS U685 ( .A(n1628), .Y(n1822) );
  AOI22X1TS U686 ( .A0(n1822), .A1(writeOutbuffer[2]), .B0(n208), .B1(n347), 
        .Y(n205) );
  AOI22X1TS U687 ( .A0(n187), .A1(n350), .B0(n203), .B1(n348), .Y(n204) );
  OAI211XLTS U688 ( .A0(n218), .A1(n249), .B0(n205), .C0(n204), .Y(n2061) );
  INVX2TS U689 ( .A(n1345), .Y(n214) );
  AOI22X1TS U690 ( .A0(n214), .A1(\destinationAddressbuffer[2][6] ), .B0(n199), 
        .B1(n354), .Y(n207) );
  AOI22X1TS U691 ( .A0(n1355), .A1(destinationAddressIn_NORTH[6]), .B0(n190), 
        .B1(n355), .Y(n206) );
  OAI211XLTS U692 ( .A0(n218), .A1(n264), .B0(n207), .C0(n206), .Y(n2138) );
  AOI22X1TS U693 ( .A0(n214), .A1(\destinationAddressbuffer[2][4] ), .B0(n208), 
        .B1(n359), .Y(n210) );
  INVX2TS U694 ( .A(n215), .Y(n1802) );
  AOI22X1TS U695 ( .A0(n1802), .A1(destinationAddressIn_NORTH[4]), .B0(n1801), 
        .B1(n362), .Y(n209) );
  OAI211XLTS U696 ( .A0(n211), .A1(n256), .B0(n210), .C0(n209), .Y(n2136) );
  AOI22X1TS U697 ( .A0(n214), .A1(\destinationAddressbuffer[2][5] ), .B0(n1808), .B1(n372), .Y(n213) );
  AOI22X1TS U698 ( .A0(n1818), .A1(destinationAddressIn_NORTH[5]), .B0(n203), 
        .B1(n374), .Y(n212) );
  OAI211XLTS U699 ( .A0(n1346), .A1(n260), .B0(n213), .C0(n212), .Y(n2137) );
  AOI22X1TS U700 ( .A0(n214), .A1(\destinationAddressbuffer[2][7] ), .B0(n1816), .B1(n367), .Y(n217) );
  INVX2TS U701 ( .A(n215), .Y(n1818) );
  AOI22X1TS U702 ( .A0(n1818), .A1(destinationAddressIn_NORTH[7]), .B0(n1809), 
        .B1(n368), .Y(n216) );
  OAI211XLTS U703 ( .A0(n218), .A1(n252), .B0(n217), .C0(n216), .Y(n2139) );
  INVX2TS U704 ( .A(n1930), .Y(n388) );
  INVX2TS U705 ( .A(n273), .Y(n440) );
  AOI31XLTS U706 ( .A0(n225), .A1(n1583), .A2(n221), .B0(n440), .Y(n223) );
  INVX2TS U707 ( .A(n1930), .Y(n384) );
  NAND2X1TS U708 ( .A(n223), .B(n1593), .Y(n226) );
  INVX2TS U709 ( .A(n222), .Y(n1429) );
  INVX2TS U710 ( .A(n1429), .Y(n920) );
  CLKBUFX2TS U711 ( .A(n920), .Y(n235) );
  INVX2TS U712 ( .A(n235), .Y(n257) );
  INVX2TS U713 ( .A(n14), .Y(n912) );
  INVX2TS U714 ( .A(n1438), .Y(n240) );
  OR2X1TS U715 ( .A(n1590), .B(n226), .Y(n239) );
  INVX2TS U716 ( .A(n239), .Y(n224) );
  INVX2TS U717 ( .A(n224), .Y(n919) );
  INVX2TS U718 ( .A(n919), .Y(n253) );
  AOI22X1TS U719 ( .A0(n240), .A1(\destinationAddressbuffer[5][8] ), .B0(n253), 
        .B1(n715), .Y(n230) );
  INVX2TS U720 ( .A(n2), .Y(n1430) );
  OR2X1TS U721 ( .A(n1583), .B(n227), .Y(n245) );
  INVX2TS U722 ( .A(n245), .Y(n228) );
  INVX2TS U723 ( .A(n228), .Y(n908) );
  INVX2TS U724 ( .A(n908), .Y(n241) );
  AOI22X1TS U725 ( .A0(n1430), .A1(n401), .B0(n241), .B1(n324), .Y(n229) );
  OAI211XLTS U726 ( .A0(n257), .A1(n231), .B0(n230), .C0(n229), .Y(n2104) );
  INVX2TS U727 ( .A(n239), .Y(n1439) );
  AOI22X1TS U728 ( .A0(n240), .A1(\destinationAddressbuffer[5][9] ), .B0(n1439), .B1(n730), .Y(n233) );
  INVX2TS U729 ( .A(n2), .Y(n1446) );
  INVX2TS U730 ( .A(n1446), .Y(n1450) );
  INVX2TS U731 ( .A(n1450), .Y(n246) );
  INVX2TS U732 ( .A(n245), .Y(n1729) );
  AOI22X1TS U733 ( .A0(n246), .A1(n397), .B0(n241), .B1(n343), .Y(n232) );
  OAI211XLTS U734 ( .A0(n257), .A1(n234), .B0(n233), .C0(n232), .Y(n2105) );
  INVX2TS U735 ( .A(n235), .Y(n265) );
  INVX2TS U736 ( .A(n239), .Y(n1444) );
  AOI22X1TS U737 ( .A0(n240), .A1(\destinationAddressbuffer[5][10] ), .B0(
        n1444), .B1(n747), .Y(n237) );
  INVX2TS U738 ( .A(n245), .Y(n1719) );
  AOI22X1TS U739 ( .A0(n1440), .A1(n407), .B0(n1719), .B1(n329), .Y(n236) );
  OAI211XLTS U740 ( .A0(n265), .A1(n238), .B0(n237), .C0(n236), .Y(n2106) );
  INVX2TS U741 ( .A(n239), .Y(n1718) );
  AOI22X1TS U742 ( .A0(n240), .A1(\destinationAddressbuffer[5][11] ), .B0(
        n1718), .B1(n762), .Y(n243) );
  AOI22X1TS U743 ( .A0(n1446), .A1(n412), .B0(n241), .B1(n336), .Y(n242) );
  OAI211XLTS U744 ( .A0(n257), .A1(n244), .B0(n243), .C0(n242), .Y(n2107) );
  INVX2TS U745 ( .A(n1594), .Y(n1733) );
  AOI22X1TS U746 ( .A0(n1733), .A1(writeOutbuffer[5]), .B0(n253), .B1(n541), 
        .Y(n248) );
  INVX2TS U747 ( .A(n245), .Y(n1445) );
  AOI22X1TS U748 ( .A0(n246), .A1(n419), .B0(n1445), .B1(n348), .Y(n247) );
  OAI211XLTS U749 ( .A0(n265), .A1(n249), .B0(n248), .C0(n247), .Y(n2058) );
  INVX2TS U750 ( .A(n1594), .Y(n261) );
  AOI22X1TS U751 ( .A0(n261), .A1(\destinationAddressbuffer[5][7] ), .B0(n1718), .B1(n704), .Y(n251) );
  INVX2TS U752 ( .A(n2), .Y(n1710) );
  AOI22X1TS U753 ( .A0(n1710), .A1(n436), .B0(n1445), .B1(n368), .Y(n250) );
  OAI211XLTS U754 ( .A0(n265), .A1(n252), .B0(n251), .C0(n250), .Y(n2103) );
  AOI22X1TS U755 ( .A0(n261), .A1(\destinationAddressbuffer[5][4] ), .B0(n253), 
        .B1(n656), .Y(n255) );
  INVX2TS U756 ( .A(n2), .Y(n1440) );
  AOI22X1TS U757 ( .A0(n1440), .A1(n432), .B0(n241), .B1(n362), .Y(n254) );
  OAI211XLTS U758 ( .A0(n257), .A1(n256), .B0(n255), .C0(n254), .Y(n2100) );
  AOI22X1TS U759 ( .A0(n261), .A1(\destinationAddressbuffer[5][5] ), .B0(n1444), .B1(n669), .Y(n259) );
  AOI22X1TS U760 ( .A0(n246), .A1(n424), .B0(n1719), .B1(n374), .Y(n258) );
  OAI211XLTS U761 ( .A0(n1429), .A1(n260), .B0(n259), .C0(n258), .Y(n2101) );
  AOI22X1TS U762 ( .A0(n261), .A1(\destinationAddressbuffer[5][6] ), .B0(n224), 
        .B1(n689), .Y(n263) );
  AOI22X1TS U763 ( .A0(n1446), .A1(n428), .B0(n1709), .B1(n355), .Y(n262) );
  OAI211XLTS U764 ( .A0(n265), .A1(n264), .B0(n263), .C0(n262), .Y(n2102) );
  AOI31XLTS U765 ( .A0(n444), .A1(n385), .A2(n388), .B0(n1597), .Y(n270) );
  AOI21X1TS U766 ( .A0(n276), .A1(n270), .B0(n440), .Y(n275) );
  NAND2X1TS U767 ( .A(n275), .B(n1605), .Y(n277) );
  INVX2TS U768 ( .A(n272), .Y(n1396) );
  INVX2TS U769 ( .A(n1396), .Y(n943) );
  CLKBUFX2TS U770 ( .A(n943), .Y(n285) );
  INVX2TS U771 ( .A(n285), .Y(n301) );
  INVX2TS U772 ( .A(n273), .Y(n386) );
  INVX2TS U773 ( .A(n274), .Y(n1406) );
  INVX2TS U774 ( .A(n1406), .Y(n931) );
  INVX2TS U775 ( .A(n1407), .Y(n291) );
  OR2X1TS U776 ( .A(n1601), .B(n277), .Y(n289) );
  INVX2TS U777 ( .A(n289), .Y(n1741) );
  AOI22X1TS U778 ( .A0(n291), .A1(\destinationAddressbuffer[4][9] ), .B0(n1741), .B1(n341), .Y(n281) );
  INVX2TS U779 ( .A(n3), .Y(n278) );
  INVX2TS U780 ( .A(n278), .Y(n926) );
  INVX2TS U781 ( .A(n926), .Y(n298) );
  INVX2TS U782 ( .A(n9), .Y(n1742) );
  AOI22X1TS U783 ( .A0(n298), .A1(n731), .B0(n282), .B1(n397), .Y(n280) );
  OAI211XLTS U784 ( .A0(n301), .A1(n44), .B0(n281), .C0(n280), .Y(n2117) );
  INVX2TS U785 ( .A(n289), .Y(n1758) );
  AOI22X1TS U786 ( .A0(n291), .A1(\destinationAddressbuffer[4][11] ), .B0(
        n1758), .B1(n334), .Y(n284) );
  INVX2TS U787 ( .A(n3), .Y(n1411) );
  INVX2TS U788 ( .A(n9), .Y(n282) );
  INVX2TS U789 ( .A(n282), .Y(n286) );
  INVX2TS U790 ( .A(n286), .Y(n1410) );
  AOI22X1TS U791 ( .A0(n1411), .A1(n765), .B0(n1410), .B1(n412), .Y(n283) );
  OAI211XLTS U792 ( .A0(n301), .A1(n35), .B0(n284), .C0(n283), .Y(n2119) );
  INVX2TS U793 ( .A(n285), .Y(n308) );
  INVX2TS U794 ( .A(n289), .Y(n1749) );
  AOI22X1TS U795 ( .A0(n291), .A1(\destinationAddressbuffer[4][10] ), .B0(
        n1749), .B1(n328), .Y(n288) );
  INVX2TS U796 ( .A(n286), .Y(n927) );
  AOI22X1TS U797 ( .A0(n1760), .A1(n750), .B0(n927), .B1(n407), .Y(n287) );
  OAI211XLTS U798 ( .A0(n308), .A1(n52), .B0(n288), .C0(n287), .Y(n2118) );
  INVX2TS U799 ( .A(n289), .Y(n290) );
  INVX2TS U800 ( .A(n290), .Y(n942) );
  INVX2TS U801 ( .A(n942), .Y(n302) );
  AOI22X1TS U802 ( .A0(n291), .A1(\destinationAddressbuffer[4][8] ), .B0(n302), 
        .B1(n318), .Y(n293) );
  INVX2TS U803 ( .A(n3), .Y(n1766) );
  INVX2TS U804 ( .A(n9), .Y(n1759) );
  AOI22X1TS U805 ( .A0(n1766), .A1(n716), .B0(n1759), .B1(n401), .Y(n292) );
  OAI211XLTS U806 ( .A0(n301), .A1(n49), .B0(n293), .C0(n292), .Y(n2116) );
  INVX2TS U807 ( .A(n1606), .Y(n1764) );
  AOI22X1TS U808 ( .A0(n1764), .A1(writeOutbuffer[4]), .B0(n302), .B1(n347), 
        .Y(n295) );
  INVX2TS U809 ( .A(n9), .Y(n1750) );
  AOI22X1TS U810 ( .A0(n1766), .A1(n543), .B0(n1750), .B1(n419), .Y(n294) );
  OAI211XLTS U811 ( .A0(n308), .A1(n57), .B0(n295), .C0(n294), .Y(n2059) );
  INVX2TS U812 ( .A(n1606), .Y(n305) );
  AOI22X1TS U813 ( .A0(n305), .A1(\destinationAddressbuffer[4][6] ), .B0(n290), 
        .B1(n354), .Y(n297) );
  INVX2TS U814 ( .A(n3), .Y(n1425) );
  AOI22X1TS U815 ( .A0(n1425), .A1(n691), .B0(n282), .B1(n428), .Y(n296) );
  OAI211XLTS U816 ( .A0(n308), .A1(n75), .B0(n297), .C0(n296), .Y(n2114) );
  AOI22X1TS U817 ( .A0(n305), .A1(\destinationAddressbuffer[4][5] ), .B0(n1749), .B1(n372), .Y(n300) );
  AOI22X1TS U818 ( .A0(n298), .A1(n671), .B0(n927), .B1(n424), .Y(n299) );
  OAI211XLTS U819 ( .A0(n301), .A1(n64), .B0(n300), .C0(n299), .Y(n2113) );
  AOI22X1TS U820 ( .A0(n305), .A1(\destinationAddressbuffer[4][4] ), .B0(n302), 
        .B1(n359), .Y(n304) );
  AOI22X1TS U821 ( .A0(n278), .A1(n658), .B0(n1759), .B1(n432), .Y(n303) );
  OAI211XLTS U822 ( .A0(n1396), .A1(n72), .B0(n304), .C0(n303), .Y(n2112) );
  AOI22X1TS U823 ( .A0(n305), .A1(\destinationAddressbuffer[4][7] ), .B0(n1758), .B1(n367), .Y(n307) );
  AOI22X1TS U824 ( .A0(n278), .A1(n705), .B0(n1750), .B1(n436), .Y(n306) );
  OAI211XLTS U825 ( .A0(n308), .A1(n67), .B0(n307), .C0(n306), .Y(n2115) );
  NOR3X1TS U826 ( .A(n219), .B(n81), .C(n379), .Y(n1639) );
  AOI31XLTS U827 ( .A0(n311), .A1(n388), .A2(n443), .B0(n1632), .Y(n312) );
  AOI21X1TS U828 ( .A0(n319), .A1(n312), .B0(n386), .Y(n316) );
  NAND2X1TS U829 ( .A(n316), .B(n1640), .Y(n320) );
  INVX2TS U830 ( .A(n313), .Y(n1090) );
  INVX2TS U831 ( .A(n1090), .Y(n1019) );
  CLKBUFX2TS U832 ( .A(n1019), .Y(n333) );
  INVX2TS U833 ( .A(n333), .Y(n366) );
  INVX2TS U834 ( .A(n315), .Y(n1088) );
  INVX2TS U835 ( .A(n1088), .Y(n1003) );
  CLKBUFX2TS U836 ( .A(n353), .Y(n1010) );
  INVX2TS U837 ( .A(n1010), .Y(n342) );
  OR2X1TS U838 ( .A(n1636), .B(n320), .Y(n340) );
  INVX2TS U839 ( .A(n340), .Y(n317) );
  INVX2TS U840 ( .A(n317), .Y(n1018) );
  INVX2TS U841 ( .A(n1018), .Y(n360) );
  AOI22X1TS U842 ( .A0(n342), .A1(\destinationAddressbuffer[1][8] ), .B0(n360), 
        .B1(n318), .Y(n327) );
  INVX2TS U843 ( .A(n361), .Y(n1832) );
  INVX2TS U844 ( .A(n8), .Y(n1842) );
  AOI22X1TS U845 ( .A0(n1832), .A1(n325), .B0(n1842), .B1(n324), .Y(n326) );
  OAI211XLTS U846 ( .A0(n366), .A1(n49), .B0(n327), .C0(n326), .Y(n2152) );
  INVX2TS U847 ( .A(n340), .Y(n1840) );
  AOI22X1TS U848 ( .A0(n342), .A1(\destinationAddressbuffer[1][10] ), .B0(
        n1840), .B1(n328), .Y(n332) );
  INVX2TS U849 ( .A(n1092), .Y(n1012) );
  INVX2TS U850 ( .A(n8), .Y(n1102) );
  AOI22X1TS U851 ( .A0(n1012), .A1(n330), .B0(n1102), .B1(n329), .Y(n331) );
  OAI211XLTS U852 ( .A0(n366), .A1(n52), .B0(n332), .C0(n331), .Y(n2154) );
  INVX2TS U853 ( .A(n333), .Y(n378) );
  INVX2TS U854 ( .A(n340), .Y(n1852) );
  AOI22X1TS U855 ( .A0(n342), .A1(\destinationAddressbuffer[1][11] ), .B0(
        n1852), .B1(n334), .Y(n339) );
  INVX2TS U856 ( .A(n361), .Y(n1856) );
  INVX2TS U857 ( .A(n8), .Y(n335) );
  INVX2TS U858 ( .A(n335), .Y(n997) );
  INVX2TS U859 ( .A(n997), .Y(n349) );
  AOI22X1TS U860 ( .A0(n1856), .A1(n337), .B0(n349), .B1(n336), .Y(n338) );
  OAI211XLTS U861 ( .A0(n378), .A1(n35), .B0(n339), .C0(n338), .Y(n2155) );
  INVX2TS U862 ( .A(n340), .Y(n1829) );
  AOI22X1TS U863 ( .A0(n342), .A1(\destinationAddressbuffer[1][9] ), .B0(n1829), .B1(n341), .Y(n346) );
  INVX2TS U864 ( .A(n1856), .Y(n1092) );
  INVX2TS U865 ( .A(n8), .Y(n1097) );
  AOI22X1TS U866 ( .A0(n321), .A1(n344), .B0(n1097), .B1(n343), .Y(n345) );
  OAI211XLTS U867 ( .A0(n366), .A1(n44), .B0(n346), .C0(n345), .Y(n2153) );
  INVX2TS U868 ( .A(n353), .Y(n1860) );
  AOI22X1TS U869 ( .A0(n1860), .A1(writeOutbuffer[1]), .B0(n360), .B1(n347), 
        .Y(n352) );
  INVX2TS U870 ( .A(n361), .Y(n1021) );
  AOI22X1TS U871 ( .A0(n1021), .A1(n350), .B0(n349), .B1(n348), .Y(n351) );
  OAI211XLTS U872 ( .A0(n378), .A1(n57), .B0(n352), .C0(n351), .Y(n2062) );
  INVX2TS U873 ( .A(n353), .Y(n373) );
  AOI22X1TS U874 ( .A0(n373), .A1(\destinationAddressbuffer[1][6] ), .B0(n317), 
        .B1(n354), .Y(n358) );
  AOI22X1TS U875 ( .A0(n1856), .A1(n356), .B0(n335), .B1(n355), .Y(n357) );
  OAI211XLTS U876 ( .A0(n378), .A1(n75), .B0(n358), .C0(n357), .Y(n2150) );
  AOI22X1TS U877 ( .A0(n373), .A1(\destinationAddressbuffer[1][4] ), .B0(n360), 
        .B1(n359), .Y(n365) );
  INVX2TS U878 ( .A(n361), .Y(n1079) );
  AOI22X1TS U879 ( .A0(n1079), .A1(n363), .B0(n1102), .B1(n362), .Y(n364) );
  OAI211XLTS U880 ( .A0(n366), .A1(n72), .B0(n365), .C0(n364), .Y(n2148) );
  AOI22X1TS U881 ( .A0(n373), .A1(\destinationAddressbuffer[1][7] ), .B0(n1852), .B1(n367), .Y(n371) );
  AOI22X1TS U882 ( .A0(n1021), .A1(n369), .B0(n1842), .B1(n368), .Y(n370) );
  OAI211XLTS U883 ( .A0(n1090), .A1(n67), .B0(n371), .C0(n370), .Y(n2151) );
  AOI22X1TS U884 ( .A0(n373), .A1(\destinationAddressbuffer[1][5] ), .B0(n1840), .B1(n372), .Y(n377) );
  AOI22X1TS U885 ( .A0(n1012), .A1(n375), .B0(n349), .B1(n374), .Y(n376) );
  OAI211XLTS U886 ( .A0(n378), .A1(n64), .B0(n377), .C0(n376), .Y(n2149) );
  AOI31XLTS U887 ( .A0(n385), .A1(n384), .A2(n482), .B0(n1643), .Y(n387) );
  AOI21X1TS U888 ( .A0(n393), .A1(n387), .B0(n386), .Y(n391) );
  NAND2X1TS U889 ( .A(n391), .B(n1651), .Y(n394) );
  INVX2TS U890 ( .A(n390), .Y(n1062) );
  INVX2TS U891 ( .A(n1062), .Y(n1046) );
  CLKBUFX2TS U892 ( .A(n1046), .Y(n404) );
  INVX2TS U893 ( .A(n404), .Y(n431) );
  INVX2TS U894 ( .A(n15), .Y(n1034) );
  INVX2TS U895 ( .A(n422), .Y(n411) );
  OR2X1TS U896 ( .A(n1648), .B(n394), .Y(n416) );
  INVX2TS U897 ( .A(n416), .Y(n1869) );
  AOI22X1TS U898 ( .A0(n411), .A1(\destinationAddressbuffer[0][9] ), .B0(n417), 
        .B1(n392), .Y(n399) );
  INVX2TS U899 ( .A(n4), .Y(n395) );
  INVX2TS U900 ( .A(n395), .Y(n1028) );
  INVX2TS U901 ( .A(n1028), .Y(n425) );
  INVX2TS U902 ( .A(n10), .Y(n1881) );
  AOI22X1TS U903 ( .A0(n425), .A1(n731), .B0(n406), .B1(n397), .Y(n398) );
  OAI211XLTS U904 ( .A0(n431), .A1(n44), .B0(n399), .C0(n398), .Y(n2165) );
  INVX2TS U905 ( .A(n416), .Y(n1879) );
  AOI22X1TS U906 ( .A0(n411), .A1(\destinationAddressbuffer[0][8] ), .B0(n1879), .B1(n400), .Y(n403) );
  INVX2TS U907 ( .A(n4), .Y(n1057) );
  INVX2TS U908 ( .A(n10), .Y(n1892) );
  AOI22X1TS U909 ( .A0(n1057), .A1(n716), .B0(n1892), .B1(n401), .Y(n402) );
  OAI211XLTS U910 ( .A0(n431), .A1(n49), .B0(n403), .C0(n402), .Y(n2164) );
  INVX2TS U911 ( .A(n404), .Y(n439) );
  INVX2TS U912 ( .A(n416), .Y(n1890) );
  AOI22X1TS U913 ( .A0(n411), .A1(\destinationAddressbuffer[0][10] ), .B0(
        n1890), .B1(n405), .Y(n409) );
  INVX2TS U914 ( .A(n10), .Y(n406) );
  INVX2TS U915 ( .A(n406), .Y(n1029) );
  INVX2TS U916 ( .A(n1029), .Y(n413) );
  AOI22X1TS U917 ( .A0(n395), .A1(n750), .B0(n413), .B1(n407), .Y(n408) );
  OAI211XLTS U918 ( .A0(n439), .A1(n52), .B0(n409), .C0(n408), .Y(n2166) );
  AOI22X1TS U919 ( .A0(n411), .A1(\destinationAddressbuffer[0][11] ), .B0(n423), .B1(n410), .Y(n415) );
  INVX2TS U920 ( .A(n4), .Y(n1894) );
  AOI22X1TS U921 ( .A0(n1894), .A1(n765), .B0(n413), .B1(n412), .Y(n414) );
  OAI211XLTS U922 ( .A0(n431), .A1(n35), .B0(n415), .C0(n414), .Y(n2167) );
  INVX2TS U923 ( .A(n422), .Y(n1898) );
  INVX2TS U924 ( .A(n416), .Y(n417) );
  INVX2TS U925 ( .A(n417), .Y(n1045) );
  INVX2TS U926 ( .A(n1045), .Y(n423) );
  AOI22X1TS U927 ( .A0(n1898), .A1(writeOutbuffer[0]), .B0(n423), .B1(n418), 
        .Y(n421) );
  INVX2TS U928 ( .A(n10), .Y(n1052) );
  AOI22X1TS U929 ( .A0(n1057), .A1(n543), .B0(n1052), .B1(n419), .Y(n420) );
  OAI211XLTS U930 ( .A0(n439), .A1(n57), .B0(n421), .C0(n420), .Y(n2063) );
  CLKBUFX2TS U931 ( .A(n422), .Y(n1061) );
  INVX2TS U932 ( .A(n1061), .Y(n435) );
  AOI22X1TS U933 ( .A0(n435), .A1(\destinationAddressbuffer[0][5] ), .B0(n423), 
        .B1(destinationAddressIn_WEST[5]), .Y(n427) );
  AOI22X1TS U934 ( .A0(n425), .A1(n671), .B0(n413), .B1(n424), .Y(n426) );
  OAI211XLTS U935 ( .A0(n439), .A1(n64), .B0(n427), .C0(n426), .Y(n2161) );
  AOI22X1TS U936 ( .A0(n435), .A1(\destinationAddressbuffer[0][6] ), .B0(n1869), .B1(destinationAddressIn_WEST[6]), .Y(n430) );
  INVX2TS U937 ( .A(n4), .Y(n1872) );
  AOI22X1TS U938 ( .A0(n1872), .A1(n691), .B0(n406), .B1(n428), .Y(n429) );
  OAI211XLTS U939 ( .A0(n431), .A1(n75), .B0(n430), .C0(n429), .Y(n2162) );
  AOI22X1TS U940 ( .A0(n435), .A1(\destinationAddressbuffer[0][4] ), .B0(n1890), .B1(destinationAddressIn_WEST[4]), .Y(n434) );
  AOI22X1TS U941 ( .A0(n395), .A1(n658), .B0(n1892), .B1(n432), .Y(n433) );
  OAI211XLTS U942 ( .A0(n1062), .A1(n72), .B0(n434), .C0(n433), .Y(n2160) );
  AOI22X1TS U943 ( .A0(n435), .A1(\destinationAddressbuffer[0][7] ), .B0(n1879), .B1(destinationAddressIn_WEST[7]), .Y(n438) );
  AOI22X1TS U944 ( .A0(n395), .A1(n705), .B0(n1052), .B1(n436), .Y(n437) );
  OAI211XLTS U945 ( .A0(n439), .A1(n67), .B0(n438), .C0(n437), .Y(n2163) );
  NAND2X1TS U946 ( .A(n490), .B(n1924), .Y(n502) );
  NOR2XLTS U947 ( .A(reset), .B(n440), .Y(n495) );
  INVX2TS U948 ( .A(n1928), .Y(n529) );
  INVX2TS U949 ( .A(n1930), .Y(n452) );
  INVX2TS U950 ( .A(n1922), .Y(n441) );
  NAND2X1TS U951 ( .A(n442), .B(n441), .Y(n455) );
  INVX2TS U952 ( .A(n1933), .Y(n444) );
  INVX2TS U953 ( .A(n1925), .Y(n525) );
  INVX2TS U954 ( .A(n1926), .Y(n528) );
  AOI22X1TS U955 ( .A0(n444), .A1(n525), .B0(n528), .B1(n443), .Y(n447) );
  INVX2TS U956 ( .A(n446), .Y(n451) );
  INVX2TS U957 ( .A(n465), .Y(n462) );
  INVX2TS U958 ( .A(n1934), .Y(n526) );
  AOI21X1TS U959 ( .A0(n526), .A1(n449), .B0(n448), .Y(n461) );
  ADDHX1TS U960 ( .A(n454), .B(n453), .CO(n465), .S(n467) );
  INVX2TS U961 ( .A(n467), .Y(n456) );
  OAI21XLTS U962 ( .A0(n473), .A1(n1934), .B0(n455), .Y(n487) );
  AOI21X1TS U963 ( .A0(n457), .A1(n456), .B0(n487), .Y(n459) );
  OAI22X1TS U964 ( .A0(n457), .A1(n456), .B0(n463), .B1(n462), .Y(n458) );
  AOI21X1TS U965 ( .A0(n466), .A1(n459), .B0(n458), .Y(n460) );
  AOI211X1TS U966 ( .A0(n463), .A1(n462), .B0(n461), .C0(n460), .Y(n464) );
  INVX2TS U967 ( .A(n464), .Y(n468) );
  NAND2X1TS U968 ( .A(n468), .B(n465), .Y(n471) );
  XNOR2X1TS U969 ( .A(n1932), .B(n469), .Y(n470) );
  INVX2TS U970 ( .A(n494), .Y(n479) );
  INVX2TS U971 ( .A(n1926), .Y(n524) );
  INVX2TS U972 ( .A(n1934), .Y(n523) );
  ADDHXLTS U973 ( .A(n473), .B(n472), .CO(n475), .S(n491) );
  XNOR2X1TS U974 ( .A(n1929), .B(n492), .Y(n476) );
  OAI21X1TS U975 ( .A0(n479), .A1(n524), .B0(n476), .Y(n477) );
  NAND2X1TS U976 ( .A(n523), .B(n529), .Y(n527) );
  OAI21XLTS U977 ( .A0(n526), .A1(n1929), .B0(n527), .Y(n501) );
  INVX2TS U978 ( .A(n1925), .Y(n530) );
  NOR2XLTS U979 ( .A(n527), .B(n525), .Y(n837) );
  CLKBUFX2TS U980 ( .A(n837), .Y(n795) );
  CLKBUFX2TS U981 ( .A(n795), .Y(n814) );
  AOI21X1TS U982 ( .A0(n527), .A1(n530), .B0(n814), .Y(n498) );
  OAI22X1TS U983 ( .A0(n483), .A1(n501), .B0(n482), .B1(n498), .Y(n484) );
  AOI221XLTS U984 ( .A0(n501), .A1(n486), .B0(n485), .B1(n498), .C0(n484), .Y(
        n488) );
  AOI21X1TS U985 ( .A0(n488), .A1(n487), .B0(n1924), .Y(n489) );
  NAND2X1TS U986 ( .A(n490), .B(n1923), .Y(n500) );
  AOI22X1TS U987 ( .A0(n1922), .A1(n502), .B0(n500), .B1(n441), .Y(n1945) );
  INVX2TS U988 ( .A(n498), .Y(n499) );
  OAI22X1TS U989 ( .A0(n530), .A1(n502), .B0(n499), .B1(n500), .Y(n1950) );
  OAI22X1TS U990 ( .A0(n16), .A1(n502), .B0(n501), .B1(n500), .Y(n1951) );
  CLKBUFX2TS U991 ( .A(readIn_SOUTH), .Y(n1585) );
  CLKBUFX2TS U992 ( .A(n1923), .Y(n843) );
  CLKBUFX2TS U993 ( .A(n542), .Y(n852) );
  CLKBUFX2TS U994 ( .A(readIn_WEST), .Y(n1603) );
  CLKBUFX2TS U995 ( .A(n1603), .Y(n1638) );
  INVX2TS U996 ( .A(n1923), .Y(n519) );
  NAND2X1TS U997 ( .A(n537), .B(n519), .Y(n507) );
  NOR4XLTS U998 ( .A(n509), .B(n510), .C(n446), .D(n507), .Y(n611) );
  CLKBUFX2TS U999 ( .A(n611), .Y(n626) );
  CLKBUFX2TS U1000 ( .A(n626), .Y(n806) );
  CLKBUFX2TS U1001 ( .A(n806), .Y(n564) );
  AOI22X1TS U1002 ( .A0(n1585), .A1(n852), .B0(n1638), .B1(n564), .Y(n540) );
  CLKBUFX2TS U1003 ( .A(readIn_NORTH), .Y(n1618) );
  CLKBUFX2TS U1004 ( .A(n1618), .Y(n1584) );
  CLKBUFX2TS U1005 ( .A(n690), .Y(n625) );
  CLKBUFX2TS U1006 ( .A(n625), .Y(n563) );
  NOR4XLTS U1007 ( .A(selectBit_WEST), .B(n508), .C(n512), .D(n507), .Y(n644)
         );
  CLKBUFX2TS U1008 ( .A(n644), .Y(n776) );
  CLKBUFX2TS U1009 ( .A(n776), .Y(n667) );
  CLKBUFX2TS U1010 ( .A(n667), .Y(n825) );
  AOI22X1TS U1011 ( .A0(n1584), .A1(n563), .B0(readIn_EAST), .B1(n825), .Y(
        n539) );
  NOR3XLTS U1012 ( .A(n510), .B(n509), .C(n446), .Y(n515) );
  NOR3XLTS U1013 ( .A(selectBit_WEST), .B(n513), .C(n512), .Y(n514) );
  OAI31X1TS U1014 ( .A0(n515), .A1(n536), .A2(n514), .B0(n537), .Y(n518) );
  NAND4XLTS U1015 ( .A(n519), .B(n518), .C(n517), .D(n516), .Y(n673) );
  INVX2TS U1016 ( .A(n673), .Y(n520) );
  INVX2TS U1017 ( .A(n520), .Y(n627) );
  INVX2TS U1018 ( .A(n627), .Y(n521) );
  CLKBUFX2TS U1019 ( .A(n1923), .Y(n599) );
  NOR3XLTS U1020 ( .A(n523), .B(n524), .C(n1928), .Y(n718) );
  CLKBUFX2TS U1021 ( .A(n718), .Y(n628) );
  CLKBUFX2TS U1022 ( .A(n628), .Y(n566) );
  NOR3XLTS U1023 ( .A(n526), .B(n1929), .C(n524), .Y(n692) );
  CLKBUFX2TS U1024 ( .A(n692), .Y(n629) );
  CLKBUFX2TS U1025 ( .A(n629), .Y(n565) );
  AOI22X1TS U1026 ( .A0(readOutbuffer[2]), .A1(n566), .B0(readOutbuffer[0]), 
        .B1(n565), .Y(n534) );
  NOR3XLTS U1027 ( .A(n523), .B(n16), .C(n525), .Y(n719) );
  CLKBUFX2TS U1028 ( .A(n719), .Y(n630) );
  CLKBUFX2TS U1029 ( .A(n630), .Y(n568) );
  NOR3XLTS U1030 ( .A(n526), .B(n529), .C(n530), .Y(n693) );
  CLKBUFX2TS U1031 ( .A(n693), .Y(n631) );
  CLKBUFX2TS U1032 ( .A(n631), .Y(n567) );
  AOI22X1TS U1033 ( .A0(readOutbuffer[6]), .A1(n568), .B0(readOutbuffer[4]), 
        .B1(n567), .Y(n533) );
  NOR2XLTS U1034 ( .A(n528), .B(n527), .Y(n720) );
  CLKBUFX2TS U1035 ( .A(n720), .Y(n632) );
  CLKBUFX2TS U1036 ( .A(n632), .Y(n570) );
  NOR3XLTS U1037 ( .A(n529), .B(n528), .C(n1934), .Y(n694) );
  CLKBUFX2TS U1038 ( .A(n694), .Y(n633) );
  CLKBUFX2TS U1039 ( .A(n633), .Y(n569) );
  AOI22X1TS U1040 ( .A0(readOutbuffer[3]), .A1(n570), .B0(readOutbuffer[1]), 
        .B1(n569), .Y(n532) );
  CLKBUFX2TS U1041 ( .A(n837), .Y(n859) );
  NOR3XLTS U1042 ( .A(n1929), .B(n441), .C(n530), .Y(n860) );
  CLKBUFX2TS U1043 ( .A(n860), .Y(n634) );
  CLKBUFX2TS U1044 ( .A(n634), .Y(n571) );
  AOI22X1TS U1045 ( .A0(readOutbuffer[7]), .A1(n859), .B0(readOutbuffer[5]), 
        .B1(n571), .Y(n531) );
  NAND4XLTS U1046 ( .A(n534), .B(n533), .C(n532), .D(n531), .Y(n535) );
  AOI22X1TS U1047 ( .A0(readOut), .A1(n550), .B0(n599), .B1(n535), .Y(n538) );
  CLKBUFX2TS U1048 ( .A(n667), .Y(n748) );
  AOI22X1TS U1049 ( .A0(writeIn_EAST), .A1(n748), .B0(n541), .B1(n564), .Y(
        n553) );
  CLKBUFX2TS U1050 ( .A(n542), .Y(n670) );
  CLKBUFX2TS U1051 ( .A(n670), .Y(n764) );
  AOI22X1TS U1052 ( .A0(n544), .A1(n563), .B0(n543), .B1(n764), .Y(n552) );
  AOI22X1TS U1053 ( .A0(writeOutbuffer[2]), .A1(n566), .B0(writeOutbuffer[0]), 
        .B1(n565), .Y(n548) );
  AOI22X1TS U1054 ( .A0(writeOutbuffer[6]), .A1(n568), .B0(writeOutbuffer[4]), 
        .B1(n567), .Y(n547) );
  AOI22X1TS U1055 ( .A0(writeOutbuffer[3]), .A1(n570), .B0(writeOutbuffer[1]), 
        .B1(n569), .Y(n546) );
  AOI22X1TS U1056 ( .A0(writeOutbuffer[7]), .A1(n859), .B0(writeOutbuffer[5]), 
        .B1(n571), .Y(n545) );
  NAND4XLTS U1057 ( .A(n548), .B(n547), .C(n546), .D(n545), .Y(n549) );
  AOI22X1TS U1058 ( .A0(writeOut), .A1(n550), .B0(n599), .B1(n549), .Y(n551)
         );
  CLKBUFX2TS U1059 ( .A(requesterAddressIn_NORTH[0]), .Y(n998) );
  CLKBUFX2TS U1060 ( .A(requesterAddressIn_EAST[0]), .Y(n1027) );
  CLKBUFX2TS U1061 ( .A(n1027), .Y(n996) );
  CLKBUFX2TS U1062 ( .A(n667), .Y(n588) );
  AOI22X1TS U1063 ( .A0(n998), .A1(n563), .B0(n996), .B1(n588), .Y(n562) );
  CLKBUFX2TS U1064 ( .A(requesterAddressIn_SOUTH[0]), .Y(n999) );
  CLKBUFX2TS U1065 ( .A(n670), .Y(n657) );
  CLKBUFX2TS U1066 ( .A(requesterAddressIn_WEST[0]), .Y(n925) );
  CLKBUFX2TS U1067 ( .A(n925), .Y(n950) );
  AOI22X1TS U1068 ( .A0(n999), .A1(n657), .B0(n950), .B1(n564), .Y(n561) );
  INVX2TS U1069 ( .A(n673), .Y(n700) );
  CLKBUFX2TS U1070 ( .A(n599), .Y(n594) );
  AOI22X1TS U1071 ( .A0(\requesterAddressbuffer[2][0] ), .A1(n566), .B0(
        \requesterAddressbuffer[0][0] ), .B1(n565), .Y(n557) );
  AOI22X1TS U1072 ( .A0(\requesterAddressbuffer[6][0] ), .A1(n568), .B0(
        \requesterAddressbuffer[4][0] ), .B1(n567), .Y(n556) );
  AOI22X1TS U1073 ( .A0(\requesterAddressbuffer[3][0] ), .A1(n570), .B0(
        \requesterAddressbuffer[1][0] ), .B1(n569), .Y(n555) );
  CLKBUFX2TS U1074 ( .A(n795), .Y(n752) );
  CLKBUFX2TS U1075 ( .A(n752), .Y(n600) );
  AOI22X1TS U1076 ( .A0(\requesterAddressbuffer[7][0] ), .A1(n600), .B0(
        \requesterAddressbuffer[5][0] ), .B1(n571), .Y(n554) );
  NAND4XLTS U1077 ( .A(n557), .B(n556), .C(n555), .D(n554), .Y(n558) );
  AOI22X1TS U1078 ( .A0(requesterAddressOut[0]), .A1(n700), .B0(n594), .B1(
        n558), .Y(n560) );
  INVX2TS U1079 ( .A(readRequesterAddress[0]), .Y(n949) );
  INVX2TS U1080 ( .A(n949), .Y(n995) );
  INVX2TS U1081 ( .A(n559), .Y(n595) );
  NAND2X1TS U1082 ( .A(n995), .B(n595), .Y(n606) );
  CLKBUFX2TS U1083 ( .A(requesterAddressIn_NORTH[1]), .Y(n1005) );
  CLKBUFX2TS U1084 ( .A(requesterAddressIn_EAST[1]), .Y(n1035) );
  CLKBUFX2TS U1085 ( .A(n1035), .Y(n1004) );
  AOI22X1TS U1086 ( .A0(n1005), .A1(n563), .B0(n1004), .B1(n588), .Y(n579) );
  CLKBUFX2TS U1087 ( .A(requesterAddressIn_SOUTH[1]), .Y(n1006) );
  CLKBUFX2TS U1088 ( .A(n542), .Y(n807) );
  CLKBUFX2TS U1089 ( .A(requesterAddressIn_WEST[1]), .Y(n933) );
  CLKBUFX2TS U1090 ( .A(n933), .Y(n959) );
  AOI22X1TS U1091 ( .A0(n1006), .A1(n807), .B0(n959), .B1(n564), .Y(n578) );
  AOI22X1TS U1092 ( .A0(\requesterAddressbuffer[2][1] ), .A1(n566), .B0(
        \requesterAddressbuffer[0][1] ), .B1(n565), .Y(n575) );
  AOI22X1TS U1093 ( .A0(\requesterAddressbuffer[6][1] ), .A1(n568), .B0(
        \requesterAddressbuffer[4][1] ), .B1(n567), .Y(n574) );
  AOI22X1TS U1094 ( .A0(\requesterAddressbuffer[3][1] ), .A1(n570), .B0(
        \requesterAddressbuffer[1][1] ), .B1(n569), .Y(n573) );
  AOI22X1TS U1095 ( .A0(\requesterAddressbuffer[7][1] ), .A1(n600), .B0(
        \requesterAddressbuffer[5][1] ), .B1(n571), .Y(n572) );
  NAND4XLTS U1096 ( .A(n575), .B(n574), .C(n573), .D(n572), .Y(n576) );
  AOI22X1TS U1097 ( .A0(requesterAddressOut[1]), .A1(n521), .B0(n594), .B1(
        n576), .Y(n577) );
  INVX2TS U1098 ( .A(readRequesterAddress[1]), .Y(n955) );
  INVX2TS U1099 ( .A(n955), .Y(n1659) );
  NAND2X1TS U1100 ( .A(n1659), .B(n595), .Y(n621) );
  CLKBUFX2TS U1101 ( .A(requesterAddressIn_NORTH[2]), .Y(n1013) );
  CLKBUFX2TS U1102 ( .A(n625), .Y(n610) );
  CLKBUFX2TS U1103 ( .A(requesterAddressIn_EAST[2]), .Y(n1040) );
  CLKBUFX2TS U1104 ( .A(n1040), .Y(n1011) );
  AOI22X1TS U1105 ( .A0(n1013), .A1(n610), .B0(n1011), .B1(n588), .Y(n587) );
  CLKBUFX2TS U1106 ( .A(requesterAddressIn_SOUTH[2]), .Y(n1014) );
  CLKBUFX2TS U1107 ( .A(requesterAddressIn_WEST[2]), .Y(n938) );
  CLKBUFX2TS U1108 ( .A(n938), .Y(n965) );
  AOI22X1TS U1109 ( .A0(n1014), .A1(n657), .B0(n965), .B1(n626), .Y(n586) );
  INVX2TS U1110 ( .A(n673), .Y(n743) );
  CLKBUFX2TS U1111 ( .A(n628), .Y(n612) );
  AOI22X1TS U1112 ( .A0(\requesterAddressbuffer[2][2] ), .A1(n612), .B0(
        \requesterAddressbuffer[0][2] ), .B1(n692), .Y(n583) );
  CLKBUFX2TS U1113 ( .A(n630), .Y(n613) );
  AOI22X1TS U1114 ( .A0(\requesterAddressbuffer[6][2] ), .A1(n613), .B0(
        \requesterAddressbuffer[4][2] ), .B1(n693), .Y(n582) );
  CLKBUFX2TS U1115 ( .A(n632), .Y(n614) );
  AOI22X1TS U1116 ( .A0(\requesterAddressbuffer[3][2] ), .A1(n614), .B0(
        \requesterAddressbuffer[1][2] ), .B1(n694), .Y(n581) );
  CLKBUFX2TS U1117 ( .A(n634), .Y(n615) );
  AOI22X1TS U1118 ( .A0(\requesterAddressbuffer[7][2] ), .A1(n600), .B0(
        \requesterAddressbuffer[5][2] ), .B1(n615), .Y(n580) );
  NAND4XLTS U1119 ( .A(n583), .B(n582), .C(n581), .D(n580), .Y(n584) );
  AOI22X1TS U1120 ( .A0(requesterAddressOut[2]), .A1(n743), .B0(n594), .B1(
        n584), .Y(n585) );
  INVX2TS U1121 ( .A(readRequesterAddress[2]), .Y(n964) );
  INVX2TS U1122 ( .A(n964), .Y(n1667) );
  NAND2X1TS U1123 ( .A(n1667), .B(n595), .Y(n640) );
  CLKBUFX2TS U1124 ( .A(requesterAddressIn_NORTH[3]), .Y(n1022) );
  CLKBUFX2TS U1125 ( .A(requesterAddressIn_EAST[3]), .Y(n1047) );
  CLKBUFX2TS U1126 ( .A(n1047), .Y(n1020) );
  AOI22X1TS U1127 ( .A0(n1022), .A1(n610), .B0(n1020), .B1(n588), .Y(n598) );
  CLKBUFX2TS U1128 ( .A(requesterAddressIn_SOUTH[3]), .Y(n1023) );
  CLKBUFX2TS U1129 ( .A(requesterAddressIn_WEST[3]), .Y(n945) );
  CLKBUFX2TS U1130 ( .A(n945), .Y(n974) );
  AOI22X1TS U1131 ( .A0(n1023), .A1(n807), .B0(n974), .B1(n611), .Y(n597) );
  AOI22X1TS U1132 ( .A0(\requesterAddressbuffer[2][3] ), .A1(n612), .B0(
        \requesterAddressbuffer[0][3] ), .B1(n692), .Y(n592) );
  AOI22X1TS U1133 ( .A0(\requesterAddressbuffer[6][3] ), .A1(n613), .B0(
        \requesterAddressbuffer[4][3] ), .B1(n693), .Y(n591) );
  AOI22X1TS U1134 ( .A0(\requesterAddressbuffer[3][3] ), .A1(n614), .B0(
        \requesterAddressbuffer[1][3] ), .B1(n694), .Y(n590) );
  CLKBUFX2TS U1135 ( .A(n752), .Y(n645) );
  AOI22X1TS U1136 ( .A0(\requesterAddressbuffer[7][3] ), .A1(n645), .B0(
        \requesterAddressbuffer[5][3] ), .B1(n615), .Y(n589) );
  NAND4XLTS U1137 ( .A(n592), .B(n591), .C(n590), .D(n589), .Y(n593) );
  AOI22X1TS U1138 ( .A0(requesterAddressOut[3]), .A1(n743), .B0(n594), .B1(
        n593), .Y(n596) );
  INVX2TS U1139 ( .A(readRequesterAddress[3]), .Y(n972) );
  INVX2TS U1140 ( .A(n972), .Y(n1675) );
  NAND2X1TS U1141 ( .A(n1675), .B(n595), .Y(n652) );
  CLKBUFX2TS U1142 ( .A(destinationAddressIn_EAST[0]), .Y(n1828) );
  CLKBUFX2TS U1143 ( .A(n1828), .Y(n1707) );
  AOI22X1TS U1144 ( .A0(destinationAddressIn_NORTH[0]), .A1(n610), .B0(n1707), 
        .B1(n776), .Y(n609) );
  CLKBUFX2TS U1145 ( .A(destinationAddressIn_WEST[0]), .Y(n1708) );
  CLKBUFX2TS U1146 ( .A(n1708), .Y(n1771) );
  AOI22X1TS U1147 ( .A0(destinationAddressIn_SOUTH[0]), .A1(n657), .B0(n1771), 
        .B1(n611), .Y(n608) );
  CLKBUFX2TS U1148 ( .A(n599), .Y(n651) );
  AOI22X1TS U1149 ( .A0(\destinationAddressbuffer[2][0] ), .A1(n612), .B0(
        \destinationAddressbuffer[0][0] ), .B1(n629), .Y(n604) );
  AOI22X1TS U1150 ( .A0(\destinationAddressbuffer[6][0] ), .A1(n613), .B0(
        \destinationAddressbuffer[4][0] ), .B1(n631), .Y(n603) );
  AOI22X1TS U1151 ( .A0(\destinationAddressbuffer[3][0] ), .A1(n614), .B0(
        \destinationAddressbuffer[1][0] ), .B1(n633), .Y(n602) );
  AOI22X1TS U1152 ( .A0(\destinationAddressbuffer[7][0] ), .A1(n600), .B0(
        \destinationAddressbuffer[5][0] ), .B1(n615), .Y(n601) );
  NAND4XLTS U1153 ( .A(n604), .B(n603), .C(n602), .D(n601), .Y(n605) );
  AOI22X1TS U1154 ( .A0(destinationAddressOut[0]), .A1(n743), .B0(n651), .B1(
        n605), .Y(n607) );
  CLKBUFX2TS U1155 ( .A(destinationAddressIn_EAST[1]), .Y(n1838) );
  CLKBUFX2TS U1156 ( .A(n1838), .Y(n1715) );
  AOI22X1TS U1157 ( .A0(destinationAddressIn_NORTH[1]), .A1(n610), .B0(n1715), 
        .B1(n644), .Y(n624) );
  CLKBUFX2TS U1158 ( .A(destinationAddressIn_WEST[1]), .Y(n1717) );
  CLKBUFX2TS U1159 ( .A(n1717), .Y(n1779) );
  AOI22X1TS U1160 ( .A0(destinationAddressIn_SOUTH[1]), .A1(n807), .B0(n1779), 
        .B1(n611), .Y(n623) );
  AOI22X1TS U1161 ( .A0(\destinationAddressbuffer[2][1] ), .A1(n612), .B0(
        \destinationAddressbuffer[0][1] ), .B1(n629), .Y(n619) );
  AOI22X1TS U1162 ( .A0(\destinationAddressbuffer[6][1] ), .A1(n613), .B0(
        \destinationAddressbuffer[4][1] ), .B1(n631), .Y(n618) );
  AOI22X1TS U1163 ( .A0(\destinationAddressbuffer[3][1] ), .A1(n614), .B0(
        \destinationAddressbuffer[1][1] ), .B1(n633), .Y(n617) );
  AOI22X1TS U1164 ( .A0(\destinationAddressbuffer[7][1] ), .A1(n645), .B0(
        \destinationAddressbuffer[5][1] ), .B1(n615), .Y(n616) );
  NAND4XLTS U1165 ( .A(n619), .B(n618), .C(n617), .D(n616), .Y(n620) );
  AOI22X1TS U1166 ( .A0(destinationAddressOut[1]), .A1(n700), .B0(n651), .B1(
        n620), .Y(n622) );
  CLKBUFX2TS U1167 ( .A(n625), .Y(n672) );
  CLKBUFX2TS U1168 ( .A(destinationAddressIn_EAST[2]), .Y(n1850) );
  CLKBUFX2TS U1169 ( .A(n1850), .Y(n1725) );
  AOI22X1TS U1170 ( .A0(destinationAddressIn_NORTH[2]), .A1(n672), .B0(n1725), 
        .B1(n644), .Y(n643) );
  CLKBUFX2TS U1171 ( .A(n542), .Y(n788) );
  CLKBUFX2TS U1172 ( .A(destinationAddressIn_WEST[2]), .Y(n1727) );
  CLKBUFX2TS U1173 ( .A(n1727), .Y(n1785) );
  CLKBUFX2TS U1174 ( .A(n626), .Y(n668) );
  AOI22X1TS U1175 ( .A0(destinationAddressIn_SOUTH[2]), .A1(n788), .B0(n1785), 
        .B1(n668), .Y(n642) );
  INVX2TS U1176 ( .A(n627), .Y(n867) );
  CLKBUFX2TS U1177 ( .A(n628), .Y(n675) );
  CLKBUFX2TS U1178 ( .A(n629), .Y(n674) );
  AOI22X1TS U1179 ( .A0(\destinationAddressbuffer[2][2] ), .A1(n675), .B0(
        \destinationAddressbuffer[0][2] ), .B1(n674), .Y(n638) );
  CLKBUFX2TS U1180 ( .A(n630), .Y(n677) );
  CLKBUFX2TS U1181 ( .A(n631), .Y(n676) );
  AOI22X1TS U1182 ( .A0(\destinationAddressbuffer[6][2] ), .A1(n677), .B0(
        \destinationAddressbuffer[4][2] ), .B1(n676), .Y(n637) );
  CLKBUFX2TS U1183 ( .A(n632), .Y(n679) );
  CLKBUFX2TS U1184 ( .A(n633), .Y(n678) );
  AOI22X1TS U1185 ( .A0(\destinationAddressbuffer[3][2] ), .A1(n679), .B0(
        \destinationAddressbuffer[1][2] ), .B1(n678), .Y(n636) );
  CLKBUFX2TS U1186 ( .A(n634), .Y(n680) );
  AOI22X1TS U1187 ( .A0(\destinationAddressbuffer[7][2] ), .A1(n645), .B0(
        \destinationAddressbuffer[5][2] ), .B1(n680), .Y(n635) );
  NAND4XLTS U1188 ( .A(n638), .B(n637), .C(n636), .D(n635), .Y(n639) );
  AOI22X1TS U1189 ( .A0(destinationAddressOut[2]), .A1(n867), .B0(n651), .B1(
        n639), .Y(n641) );
  CLKBUFX2TS U1190 ( .A(destinationAddressIn_EAST[3]), .Y(n1862) );
  CLKBUFX2TS U1191 ( .A(n1862), .Y(n1735) );
  AOI22X1TS U1192 ( .A0(destinationAddressIn_NORTH[3]), .A1(n672), .B0(n1735), 
        .B1(n644), .Y(n655) );
  CLKBUFX2TS U1193 ( .A(destinationAddressIn_WEST[3]), .Y(n1736) );
  CLKBUFX2TS U1194 ( .A(n1736), .Y(n1794) );
  AOI22X1TS U1195 ( .A0(destinationAddressIn_SOUTH[3]), .A1(n788), .B0(n1794), 
        .B1(n668), .Y(n654) );
  AOI22X1TS U1196 ( .A0(\destinationAddressbuffer[2][3] ), .A1(n675), .B0(
        \destinationAddressbuffer[0][3] ), .B1(n674), .Y(n649) );
  AOI22X1TS U1197 ( .A0(\destinationAddressbuffer[6][3] ), .A1(n677), .B0(
        \destinationAddressbuffer[4][3] ), .B1(n676), .Y(n648) );
  AOI22X1TS U1198 ( .A0(\destinationAddressbuffer[3][3] ), .A1(n679), .B0(
        \destinationAddressbuffer[1][3] ), .B1(n678), .Y(n647) );
  AOI22X1TS U1199 ( .A0(\destinationAddressbuffer[7][3] ), .A1(n645), .B0(
        \destinationAddressbuffer[5][3] ), .B1(n680), .Y(n646) );
  NAND4XLTS U1200 ( .A(n649), .B(n648), .C(n647), .D(n646), .Y(n650) );
  AOI22X1TS U1201 ( .A0(destinationAddressOut[3]), .A1(n521), .B0(n651), .B1(
        n650), .Y(n653) );
  AOI22X1TS U1202 ( .A0(destinationAddressIn_EAST[4]), .A1(n748), .B0(n656), 
        .B1(n668), .Y(n666) );
  AOI22X1TS U1203 ( .A0(destinationAddressIn_NORTH[4]), .A1(n672), .B0(n658), 
        .B1(n657), .Y(n665) );
  INVX2TS U1204 ( .A(n1924), .Y(n767) );
  CLKBUFX2TS U1205 ( .A(n767), .Y(n866) );
  AOI22X1TS U1206 ( .A0(\destinationAddressbuffer[2][4] ), .A1(n675), .B0(
        \destinationAddressbuffer[0][4] ), .B1(n674), .Y(n662) );
  AOI22X1TS U1207 ( .A0(\destinationAddressbuffer[6][4] ), .A1(n677), .B0(
        \destinationAddressbuffer[4][4] ), .B1(n676), .Y(n661) );
  AOI22X1TS U1208 ( .A0(\destinationAddressbuffer[3][4] ), .A1(n679), .B0(
        \destinationAddressbuffer[1][4] ), .B1(n678), .Y(n660) );
  CLKBUFX2TS U1209 ( .A(n752), .Y(n706) );
  AOI22X1TS U1210 ( .A0(\destinationAddressbuffer[7][4] ), .A1(n706), .B0(
        \destinationAddressbuffer[5][4] ), .B1(n680), .Y(n659) );
  NAND4XLTS U1211 ( .A(n662), .B(n661), .C(n660), .D(n659), .Y(n663) );
  AOI22X1TS U1212 ( .A0(destinationAddressOut[4]), .A1(n700), .B0(n866), .B1(
        n663), .Y(n664) );
  CLKBUFX2TS U1213 ( .A(n667), .Y(n763) );
  AOI22X1TS U1214 ( .A0(destinationAddressIn_EAST[5]), .A1(n763), .B0(n669), 
        .B1(n668), .Y(n688) );
  CLKBUFX2TS U1215 ( .A(n670), .Y(n749) );
  AOI22X1TS U1216 ( .A0(destinationAddressIn_NORTH[5]), .A1(n672), .B0(n671), 
        .B1(n749), .Y(n687) );
  INVX2TS U1217 ( .A(n673), .Y(n832) );
  AOI22X1TS U1218 ( .A0(\destinationAddressbuffer[2][5] ), .A1(n675), .B0(
        \destinationAddressbuffer[0][5] ), .B1(n674), .Y(n684) );
  AOI22X1TS U1219 ( .A0(\destinationAddressbuffer[6][5] ), .A1(n677), .B0(
        \destinationAddressbuffer[4][5] ), .B1(n676), .Y(n683) );
  AOI22X1TS U1220 ( .A0(\destinationAddressbuffer[3][5] ), .A1(n679), .B0(
        \destinationAddressbuffer[1][5] ), .B1(n678), .Y(n682) );
  AOI22X1TS U1221 ( .A0(\destinationAddressbuffer[7][5] ), .A1(n706), .B0(
        \destinationAddressbuffer[5][5] ), .B1(n680), .Y(n681) );
  NAND4XLTS U1222 ( .A(n684), .B(n683), .C(n682), .D(n681), .Y(n685) );
  AOI22X1TS U1223 ( .A0(destinationAddressOut[5]), .A1(n832), .B0(n866), .B1(
        n685), .Y(n686) );
  CLKBUFX2TS U1224 ( .A(n806), .Y(n729) );
  AOI22X1TS U1225 ( .A0(destinationAddressIn_EAST[6]), .A1(n763), .B0(n689), 
        .B1(n729), .Y(n703) );
  CLKBUFX2TS U1226 ( .A(n690), .Y(n732) );
  AOI22X1TS U1227 ( .A0(destinationAddressIn_NORTH[6]), .A1(n732), .B0(n691), 
        .B1(n749), .Y(n702) );
  CLKBUFX2TS U1228 ( .A(n692), .Y(n808) );
  CLKBUFX2TS U1229 ( .A(n808), .Y(n734) );
  AOI22X1TS U1230 ( .A0(\destinationAddressbuffer[2][6] ), .A1(n718), .B0(
        \destinationAddressbuffer[0][6] ), .B1(n734), .Y(n698) );
  CLKBUFX2TS U1231 ( .A(n693), .Y(n810) );
  CLKBUFX2TS U1232 ( .A(n810), .Y(n735) );
  AOI22X1TS U1233 ( .A0(\destinationAddressbuffer[6][6] ), .A1(n719), .B0(
        \destinationAddressbuffer[4][6] ), .B1(n735), .Y(n697) );
  CLKBUFX2TS U1234 ( .A(n694), .Y(n812) );
  CLKBUFX2TS U1235 ( .A(n812), .Y(n736) );
  AOI22X1TS U1236 ( .A0(\destinationAddressbuffer[3][6] ), .A1(n720), .B0(
        \destinationAddressbuffer[1][6] ), .B1(n736), .Y(n696) );
  CLKBUFX2TS U1237 ( .A(n860), .Y(n826) );
  CLKBUFX2TS U1238 ( .A(n826), .Y(n737) );
  AOI22X1TS U1239 ( .A0(\destinationAddressbuffer[7][6] ), .A1(n706), .B0(
        \destinationAddressbuffer[5][6] ), .B1(n737), .Y(n695) );
  NAND4XLTS U1240 ( .A(n698), .B(n697), .C(n696), .D(n695), .Y(n699) );
  AOI22X1TS U1241 ( .A0(destinationAddressOut[6]), .A1(n700), .B0(n866), .B1(
        n699), .Y(n701) );
  AOI22X1TS U1242 ( .A0(destinationAddressIn_EAST[7]), .A1(n825), .B0(n704), 
        .B1(n729), .Y(n714) );
  AOI22X1TS U1243 ( .A0(destinationAddressIn_NORTH[7]), .A1(n732), .B0(n705), 
        .B1(n764), .Y(n713) );
  CLKBUFX2TS U1244 ( .A(n767), .Y(n758) );
  AOI22X1TS U1245 ( .A0(\destinationAddressbuffer[2][7] ), .A1(n718), .B0(
        \destinationAddressbuffer[0][7] ), .B1(n734), .Y(n710) );
  AOI22X1TS U1246 ( .A0(\destinationAddressbuffer[6][7] ), .A1(n719), .B0(
        \destinationAddressbuffer[4][7] ), .B1(n735), .Y(n709) );
  AOI22X1TS U1247 ( .A0(\destinationAddressbuffer[3][7] ), .A1(n720), .B0(
        \destinationAddressbuffer[1][7] ), .B1(n736), .Y(n708) );
  AOI22X1TS U1248 ( .A0(\destinationAddressbuffer[7][7] ), .A1(n706), .B0(
        \destinationAddressbuffer[5][7] ), .B1(n737), .Y(n707) );
  NAND4XLTS U1249 ( .A(n710), .B(n709), .C(n708), .D(n707), .Y(n711) );
  AOI22X1TS U1250 ( .A0(destinationAddressOut[7]), .A1(n520), .B0(n758), .B1(
        n711), .Y(n712) );
  AOI22X1TS U1251 ( .A0(destinationAddressIn_EAST[8]), .A1(n748), .B0(n715), 
        .B1(n729), .Y(n728) );
  AOI22X1TS U1252 ( .A0(n717), .A1(n732), .B0(n716), .B1(n749), .Y(n727) );
  CLKBUFX2TS U1253 ( .A(n718), .Y(n809) );
  AOI22X1TS U1254 ( .A0(\destinationAddressbuffer[2][8] ), .A1(n809), .B0(
        \destinationAddressbuffer[0][8] ), .B1(n734), .Y(n724) );
  CLKBUFX2TS U1255 ( .A(n719), .Y(n811) );
  AOI22X1TS U1256 ( .A0(\destinationAddressbuffer[6][8] ), .A1(n811), .B0(
        \destinationAddressbuffer[4][8] ), .B1(n735), .Y(n723) );
  CLKBUFX2TS U1257 ( .A(n720), .Y(n813) );
  AOI22X1TS U1258 ( .A0(\destinationAddressbuffer[3][8] ), .A1(n813), .B0(
        \destinationAddressbuffer[1][8] ), .B1(n736), .Y(n722) );
  AOI22X1TS U1259 ( .A0(\destinationAddressbuffer[7][8] ), .A1(n814), .B0(
        \destinationAddressbuffer[5][8] ), .B1(n737), .Y(n721) );
  NAND4XLTS U1260 ( .A(n724), .B(n723), .C(n722), .D(n721), .Y(n725) );
  AOI22X1TS U1261 ( .A0(destinationAddressOut[8]), .A1(n867), .B0(n758), .B1(
        n725), .Y(n726) );
  AOI22X1TS U1262 ( .A0(destinationAddressIn_EAST[9]), .A1(n763), .B0(n730), 
        .B1(n729), .Y(n746) );
  AOI22X1TS U1263 ( .A0(n733), .A1(n732), .B0(n731), .B1(n764), .Y(n745) );
  AOI22X1TS U1264 ( .A0(\destinationAddressbuffer[2][9] ), .A1(n809), .B0(
        \destinationAddressbuffer[0][9] ), .B1(n734), .Y(n741) );
  AOI22X1TS U1265 ( .A0(\destinationAddressbuffer[6][9] ), .A1(n811), .B0(
        \destinationAddressbuffer[4][9] ), .B1(n735), .Y(n740) );
  AOI22X1TS U1266 ( .A0(\destinationAddressbuffer[3][9] ), .A1(n813), .B0(
        \destinationAddressbuffer[1][9] ), .B1(n736), .Y(n739) );
  AOI22X1TS U1267 ( .A0(\destinationAddressbuffer[7][9] ), .A1(n814), .B0(
        \destinationAddressbuffer[5][9] ), .B1(n737), .Y(n738) );
  NAND4XLTS U1268 ( .A(n741), .B(n740), .C(n739), .D(n738), .Y(n742) );
  AOI22X1TS U1269 ( .A0(destinationAddressOut[9]), .A1(n743), .B0(n758), .B1(
        n742), .Y(n744) );
  CLKBUFX2TS U1270 ( .A(n806), .Y(n787) );
  AOI22X1TS U1271 ( .A0(destinationAddressIn_EAST[10]), .A1(n748), .B0(n747), 
        .B1(n787), .Y(n761) );
  CLKBUFX2TS U1272 ( .A(n690), .Y(n786) );
  AOI22X1TS U1273 ( .A0(n751), .A1(n786), .B0(n750), .B1(n749), .Y(n760) );
  CLKBUFX2TS U1274 ( .A(n809), .Y(n789) );
  CLKBUFX2TS U1275 ( .A(n808), .Y(n790) );
  AOI22X1TS U1276 ( .A0(\destinationAddressbuffer[2][10] ), .A1(n789), .B0(
        \destinationAddressbuffer[0][10] ), .B1(n790), .Y(n756) );
  CLKBUFX2TS U1277 ( .A(n811), .Y(n791) );
  CLKBUFX2TS U1278 ( .A(n810), .Y(n792) );
  AOI22X1TS U1279 ( .A0(\destinationAddressbuffer[6][10] ), .A1(n791), .B0(
        \destinationAddressbuffer[4][10] ), .B1(n792), .Y(n755) );
  CLKBUFX2TS U1280 ( .A(n813), .Y(n793) );
  CLKBUFX2TS U1281 ( .A(n812), .Y(n794) );
  AOI22X1TS U1282 ( .A0(\destinationAddressbuffer[3][10] ), .A1(n793), .B0(
        \destinationAddressbuffer[1][10] ), .B1(n794), .Y(n754) );
  CLKBUFX2TS U1283 ( .A(n826), .Y(n796) );
  AOI22X1TS U1284 ( .A0(\destinationAddressbuffer[7][10] ), .A1(n752), .B0(
        \destinationAddressbuffer[5][10] ), .B1(n796), .Y(n753) );
  NAND4XLTS U1285 ( .A(n756), .B(n755), .C(n754), .D(n753), .Y(n757) );
  AOI22X1TS U1286 ( .A0(destinationAddressOut[10]), .A1(n867), .B0(n758), .B1(
        n757), .Y(n759) );
  AOI22X1TS U1287 ( .A0(destinationAddressIn_EAST[11]), .A1(n763), .B0(n762), 
        .B1(n787), .Y(n775) );
  AOI22X1TS U1288 ( .A0(n766), .A1(n786), .B0(n765), .B1(n764), .Y(n774) );
  CLKBUFX2TS U1289 ( .A(n767), .Y(n820) );
  AOI22X1TS U1290 ( .A0(\destinationAddressbuffer[2][11] ), .A1(n789), .B0(
        \destinationAddressbuffer[0][11] ), .B1(n790), .Y(n771) );
  AOI22X1TS U1291 ( .A0(\destinationAddressbuffer[6][11] ), .A1(n791), .B0(
        \destinationAddressbuffer[4][11] ), .B1(n792), .Y(n770) );
  AOI22X1TS U1292 ( .A0(\destinationAddressbuffer[3][11] ), .A1(n793), .B0(
        \destinationAddressbuffer[1][11] ), .B1(n794), .Y(n769) );
  AOI22X1TS U1293 ( .A0(\destinationAddressbuffer[7][11] ), .A1(n795), .B0(
        \destinationAddressbuffer[5][11] ), .B1(n796), .Y(n768) );
  NAND4XLTS U1294 ( .A(n771), .B(n770), .C(n769), .D(n768), .Y(n772) );
  AOI22X1TS U1295 ( .A0(destinationAddressOut[11]), .A1(n520), .B0(n820), .B1(
        n772), .Y(n773) );
  CLKBUFX2TS U1296 ( .A(dataIn_EAST[0]), .Y(n1460) );
  CLKBUFX2TS U1297 ( .A(n1460), .Y(n1111) );
  CLKBUFX2TS U1298 ( .A(n776), .Y(n849) );
  AOI22X1TS U1299 ( .A0(dataIn_NORTH[0]), .A1(n786), .B0(n1111), .B1(n849), 
        .Y(n785) );
  CLKBUFX2TS U1300 ( .A(dataIn_WEST[0]), .Y(n1511) );
  CLKBUFX2TS U1301 ( .A(n1511), .Y(n1397) );
  AOI22X1TS U1302 ( .A0(dataIn_SOUTH[0]), .A1(n788), .B0(n1397), .B1(n787), 
        .Y(n784) );
  AOI22X1TS U1303 ( .A0(\dataoutbuffer[0][0] ), .A1(n790), .B0(
        \dataoutbuffer[2][0] ), .B1(n789), .Y(n780) );
  AOI22X1TS U1304 ( .A0(\dataoutbuffer[4][0] ), .A1(n792), .B0(
        \dataoutbuffer[6][0] ), .B1(n791), .Y(n779) );
  AOI22X1TS U1305 ( .A0(\dataoutbuffer[1][0] ), .A1(n794), .B0(
        \dataoutbuffer[3][0] ), .B1(n793), .Y(n778) );
  AOI22X1TS U1306 ( .A0(\dataoutbuffer[5][0] ), .A1(n796), .B0(
        \dataoutbuffer[7][0] ), .B1(n859), .Y(n777) );
  NAND4XLTS U1307 ( .A(n780), .B(n779), .C(n778), .D(n777), .Y(n781) );
  AOI22X1TS U1308 ( .A0(dataOut[0]), .A1(n521), .B0(n820), .B1(n781), .Y(n783)
         );
  INVX2TS U1309 ( .A(cacheDataOut[0]), .Y(n1078) );
  INVX2TS U1310 ( .A(n559), .Y(n844) );
  NAND2X1TS U1311 ( .A(cacheDataOut[0]), .B(n844), .Y(n782) );
  CLKBUFX2TS U1312 ( .A(dataIn_EAST[1]), .Y(n1468) );
  CLKBUFX2TS U1313 ( .A(n1468), .Y(n1341) );
  AOI22X1TS U1314 ( .A0(dataIn_NORTH[1]), .A1(n786), .B0(n1341), .B1(n825), 
        .Y(n805) );
  CLKBUFX2TS U1315 ( .A(dataIn_WEST[1]), .Y(n1521) );
  CLKBUFX2TS U1316 ( .A(n1521), .Y(n1402) );
  AOI22X1TS U1317 ( .A0(dataIn_SOUTH[1]), .A1(n788), .B0(n1402), .B1(n787), 
        .Y(n804) );
  AOI22X1TS U1318 ( .A0(\dataoutbuffer[0][1] ), .A1(n790), .B0(
        \dataoutbuffer[2][1] ), .B1(n789), .Y(n800) );
  AOI22X1TS U1319 ( .A0(\dataoutbuffer[4][1] ), .A1(n792), .B0(
        \dataoutbuffer[6][1] ), .B1(n791), .Y(n799) );
  AOI22X1TS U1320 ( .A0(\dataoutbuffer[1][1] ), .A1(n794), .B0(
        \dataoutbuffer[3][1] ), .B1(n793), .Y(n798) );
  AOI22X1TS U1321 ( .A0(\dataoutbuffer[5][1] ), .A1(n796), .B0(
        \dataoutbuffer[7][1] ), .B1(n795), .Y(n797) );
  NAND4XLTS U1322 ( .A(n800), .B(n799), .C(n798), .D(n797), .Y(n801) );
  AOI22X1TS U1323 ( .A0(dataOut[1]), .A1(n832), .B0(n820), .B1(n801), .Y(n803)
         );
  INVX2TS U1324 ( .A(cacheDataOut[1]), .Y(n1083) );
  INVX2TS U1325 ( .A(n559), .Y(n868) );
  NAND2X1TS U1326 ( .A(cacheDataOut[1]), .B(n868), .Y(n802) );
  CLKBUFX2TS U1327 ( .A(n690), .Y(n850) );
  CLKBUFX2TS U1328 ( .A(dataIn_EAST[2]), .Y(n1477) );
  CLKBUFX2TS U1329 ( .A(n1477), .Y(n1347) );
  AOI22X1TS U1330 ( .A0(dataIn_NORTH[2]), .A1(n850), .B0(n1347), .B1(n849), 
        .Y(n824) );
  CLKBUFX2TS U1331 ( .A(dataIn_WEST[2]), .Y(n1529) );
  CLKBUFX2TS U1332 ( .A(n1529), .Y(n1408) );
  CLKBUFX2TS U1333 ( .A(n806), .Y(n851) );
  AOI22X1TS U1334 ( .A0(dataIn_SOUTH[2]), .A1(n807), .B0(n1408), .B1(n851), 
        .Y(n823) );
  CLKBUFX2TS U1335 ( .A(n808), .Y(n854) );
  CLKBUFX2TS U1336 ( .A(n809), .Y(n853) );
  AOI22X1TS U1337 ( .A0(\dataoutbuffer[0][2] ), .A1(n854), .B0(
        \dataoutbuffer[2][2] ), .B1(n853), .Y(n818) );
  CLKBUFX2TS U1338 ( .A(n810), .Y(n856) );
  CLKBUFX2TS U1339 ( .A(n811), .Y(n855) );
  AOI22X1TS U1340 ( .A0(\dataoutbuffer[4][2] ), .A1(n856), .B0(
        \dataoutbuffer[6][2] ), .B1(n855), .Y(n817) );
  CLKBUFX2TS U1341 ( .A(n812), .Y(n858) );
  CLKBUFX2TS U1342 ( .A(n813), .Y(n857) );
  AOI22X1TS U1343 ( .A0(\dataoutbuffer[1][2] ), .A1(n858), .B0(
        \dataoutbuffer[3][2] ), .B1(n857), .Y(n816) );
  AOI22X1TS U1344 ( .A0(\dataoutbuffer[5][2] ), .A1(n826), .B0(
        \dataoutbuffer[7][2] ), .B1(n814), .Y(n815) );
  NAND4XLTS U1345 ( .A(n818), .B(n817), .C(n816), .D(n815), .Y(n819) );
  AOI22X1TS U1346 ( .A0(dataOut[2]), .A1(n832), .B0(n820), .B1(n819), .Y(n822)
         );
  INVX2TS U1347 ( .A(cacheDataOut[2]), .Y(n1089) );
  NAND2X1TS U1348 ( .A(cacheDataOut[2]), .B(n844), .Y(n821) );
  CLKBUFX2TS U1349 ( .A(dataIn_EAST[3]), .Y(n1487) );
  CLKBUFX2TS U1350 ( .A(n1487), .Y(n1353) );
  AOI22X1TS U1351 ( .A0(dataIn_NORTH[3]), .A1(n850), .B0(n1353), .B1(n825), 
        .Y(n836) );
  CLKBUFX2TS U1352 ( .A(dataIn_WEST[3]), .Y(n1536) );
  CLKBUFX2TS U1353 ( .A(n1536), .Y(n1415) );
  AOI22X1TS U1354 ( .A0(dataIn_SOUTH[3]), .A1(n852), .B0(n1415), .B1(n851), 
        .Y(n835) );
  AOI22X1TS U1355 ( .A0(\dataoutbuffer[0][3] ), .A1(n854), .B0(
        \dataoutbuffer[2][3] ), .B1(n853), .Y(n830) );
  AOI22X1TS U1356 ( .A0(\dataoutbuffer[4][3] ), .A1(n856), .B0(
        \dataoutbuffer[6][3] ), .B1(n855), .Y(n829) );
  AOI22X1TS U1357 ( .A0(\dataoutbuffer[1][3] ), .A1(n858), .B0(
        \dataoutbuffer[3][3] ), .B1(n857), .Y(n828) );
  AOI22X1TS U1358 ( .A0(\dataoutbuffer[5][3] ), .A1(n826), .B0(
        \dataoutbuffer[7][3] ), .B1(n837), .Y(n827) );
  NAND4XLTS U1359 ( .A(n830), .B(n829), .C(n828), .D(n827), .Y(n831) );
  AOI22X1TS U1360 ( .A0(dataOut[3]), .A1(n832), .B0(n843), .B1(n831), .Y(n834)
         );
  INVX2TS U1361 ( .A(cacheDataOut[3]), .Y(n1096) );
  NAND2X1TS U1362 ( .A(cacheDataOut[3]), .B(n868), .Y(n833) );
  CLKBUFX2TS U1363 ( .A(dataIn_EAST[4]), .Y(n1495) );
  CLKBUFX2TS U1364 ( .A(n1495), .Y(n1359) );
  AOI22X1TS U1365 ( .A0(dataIn_NORTH[4]), .A1(n850), .B0(n1359), .B1(n849), 
        .Y(n848) );
  CLKBUFX2TS U1366 ( .A(dataIn_WEST[4]), .Y(n1544) );
  CLKBUFX2TS U1367 ( .A(n1544), .Y(n1419) );
  AOI22X1TS U1368 ( .A0(dataIn_SOUTH[4]), .A1(n852), .B0(n1419), .B1(n851), 
        .Y(n847) );
  AOI22X1TS U1369 ( .A0(\dataoutbuffer[0][4] ), .A1(n854), .B0(
        \dataoutbuffer[2][4] ), .B1(n853), .Y(n841) );
  AOI22X1TS U1370 ( .A0(\dataoutbuffer[4][4] ), .A1(n856), .B0(
        \dataoutbuffer[6][4] ), .B1(n855), .Y(n840) );
  AOI22X1TS U1371 ( .A0(\dataoutbuffer[1][4] ), .A1(n858), .B0(
        \dataoutbuffer[3][4] ), .B1(n857), .Y(n839) );
  AOI22X1TS U1372 ( .A0(\dataoutbuffer[5][4] ), .A1(n860), .B0(
        \dataoutbuffer[7][4] ), .B1(n837), .Y(n838) );
  NAND4XLTS U1373 ( .A(n841), .B(n840), .C(n839), .D(n838), .Y(n842) );
  AOI22X1TS U1374 ( .A0(dataOut[4]), .A1(n521), .B0(n843), .B1(n842), .Y(n846)
         );
  INVX2TS U1375 ( .A(cacheDataOut[4]), .Y(n1101) );
  NAND2X1TS U1376 ( .A(cacheDataOut[4]), .B(n844), .Y(n845) );
  CLKBUFX2TS U1377 ( .A(dataIn_EAST[5]), .Y(n1503) );
  CLKBUFX2TS U1378 ( .A(n1503), .Y(n1364) );
  AOI22X1TS U1379 ( .A0(dataIn_NORTH[5]), .A1(n850), .B0(n1364), .B1(n849), 
        .Y(n872) );
  CLKBUFX2TS U1380 ( .A(dataIn_WEST[5]), .Y(n1554) );
  CLKBUFX2TS U1381 ( .A(n1554), .Y(n1424) );
  AOI22X1TS U1382 ( .A0(dataIn_SOUTH[5]), .A1(n852), .B0(n1424), .B1(n851), 
        .Y(n871) );
  AOI22X1TS U1383 ( .A0(\dataoutbuffer[0][5] ), .A1(n854), .B0(
        \dataoutbuffer[2][5] ), .B1(n853), .Y(n864) );
  AOI22X1TS U1384 ( .A0(\dataoutbuffer[4][5] ), .A1(n856), .B0(
        \dataoutbuffer[6][5] ), .B1(n855), .Y(n863) );
  AOI22X1TS U1385 ( .A0(\dataoutbuffer[1][5] ), .A1(n858), .B0(
        \dataoutbuffer[3][5] ), .B1(n857), .Y(n862) );
  AOI22X1TS U1386 ( .A0(\dataoutbuffer[5][5] ), .A1(n860), .B0(
        \dataoutbuffer[7][5] ), .B1(n859), .Y(n861) );
  NAND4XLTS U1387 ( .A(n864), .B(n863), .C(n862), .D(n861), .Y(n865) );
  AOI22X1TS U1388 ( .A0(dataOut[5]), .A1(n867), .B0(n866), .B1(n865), .Y(n870)
         );
  INVX2TS U1389 ( .A(cacheDataOut[5]), .Y(n1106) );
  NAND2X1TS U1390 ( .A(cacheDataOut[5]), .B(n868), .Y(n869) );
  INVX2TS U1391 ( .A(n949), .Y(n1770) );
  INVX2TS U1392 ( .A(n1570), .Y(n1666) );
  AOI22X1TS U1393 ( .A0(n1770), .A1(n1653), .B0(n1666), .B1(
        \requesterAddressbuffer[7][0] ), .Y(n877) );
  INVX2TS U1394 ( .A(n887), .Y(n1543) );
  CLKBUFX2TS U1395 ( .A(n1027), .Y(n924) );
  AOI22X1TS U1396 ( .A0(n59), .A1(n950), .B0(n1543), .B1(n924), .Y(n876) );
  INVX2TS U1397 ( .A(n873), .Y(n1557) );
  CLKBUFX2TS U1398 ( .A(requesterAddressIn_SOUTH[0]), .Y(n1030) );
  INVX2TS U1399 ( .A(n874), .Y(n1677) );
  CLKBUFX2TS U1400 ( .A(n998), .Y(n951) );
  AOI22X1TS U1401 ( .A0(n1557), .A1(n1030), .B0(n1677), .B1(n951), .Y(n875) );
  INVX2TS U1402 ( .A(n886), .Y(n1660) );
  AOI22X1TS U1403 ( .A0(n1660), .A1(n1659), .B0(n1674), .B1(
        \requesterAddressbuffer[7][1] ), .Y(n880) );
  INVX2TS U1404 ( .A(n887), .Y(n1654) );
  CLKBUFX2TS U1405 ( .A(n1035), .Y(n932) );
  AOI22X1TS U1406 ( .A0(n59), .A1(n959), .B0(n1654), .B1(n932), .Y(n879) );
  CLKBUFX2TS U1407 ( .A(requesterAddressIn_SOUTH[1]), .Y(n1036) );
  CLKBUFX2TS U1408 ( .A(n1005), .Y(n960) );
  AOI22X1TS U1409 ( .A0(n1662), .A1(n1036), .B0(n1514), .B1(n960), .Y(n878) );
  INVX2TS U1410 ( .A(n1570), .Y(n1519) );
  AOI22X1TS U1411 ( .A0(n36), .A1(n1667), .B0(n1519), .B1(
        \requesterAddressbuffer[7][2] ), .Y(n885) );
  CLKBUFX2TS U1412 ( .A(n1040), .Y(n937) );
  AOI22X1TS U1413 ( .A0(n38), .A1(n965), .B0(n1543), .B1(n937), .Y(n884) );
  CLKBUFX2TS U1414 ( .A(requesterAddressIn_SOUTH[2]), .Y(n1041) );
  CLKBUFX2TS U1415 ( .A(n1013), .Y(n968) );
  AOI22X1TS U1416 ( .A0(n1557), .A1(n1041), .B0(n882), .B1(n968), .Y(n883) );
  INVX2TS U1417 ( .A(n886), .Y(n1676) );
  AOI22X1TS U1418 ( .A0(n1676), .A1(n1675), .B0(n1519), .B1(
        \requesterAddressbuffer[7][3] ), .Y(n890) );
  CLKBUFX2TS U1419 ( .A(n1047), .Y(n944) );
  AOI22X1TS U1420 ( .A0(n1512), .A1(n974), .B0(n34), .B1(n944), .Y(n889) );
  CLKBUFX2TS U1421 ( .A(requesterAddressIn_SOUTH[3]), .Y(n1048) );
  CLKBUFX2TS U1422 ( .A(n1022), .Y(n975) );
  AOI22X1TS U1423 ( .A0(n1670), .A1(n1048), .B0(n1546), .B1(n975), .Y(n888) );
  INVX2TS U1424 ( .A(n949), .Y(n1827) );
  INVX2TS U1425 ( .A(n1475), .Y(n1694) );
  AOI22X1TS U1426 ( .A0(n1827), .A1(n894), .B0(n1694), .B1(
        \requesterAddressbuffer[6][0] ), .Y(n893) );
  INVX2TS U1427 ( .A(n1459), .Y(n1687) );
  AOI22X1TS U1428 ( .A0(n925), .A1(n1478), .B0(n924), .B1(n1687), .Y(n892) );
  AOI22X1TS U1429 ( .A0(requesterAddressIn_SOUTH[0]), .A1(n1703), .B0(n951), 
        .B1(n1690), .Y(n891) );
  INVX2TS U1430 ( .A(n955), .Y(n1747) );
  AOI22X1TS U1431 ( .A0(n1747), .A1(n894), .B0(n1701), .B1(
        \requesterAddressbuffer[6][1] ), .Y(n898) );
  INVX2TS U1432 ( .A(n1459), .Y(n1695) );
  AOI22X1TS U1433 ( .A0(n933), .A1(n1696), .B0(n932), .B1(n1695), .Y(n897) );
  AOI22X1TS U1434 ( .A0(requesterAddressIn_SOUTH[1]), .A1(n95), .B0(n960), 
        .B1(n895), .Y(n896) );
  INVX2TS U1435 ( .A(n964), .Y(n1756) );
  INVX2TS U1436 ( .A(n1474), .Y(n1686) );
  INVX2TS U1437 ( .A(n1581), .Y(n1466) );
  AOI22X1TS U1438 ( .A0(n1756), .A1(n1686), .B0(n1466), .B1(
        \requesterAddressbuffer[6][2] ), .Y(n901) );
  AOI22X1TS U1439 ( .A0(n938), .A1(n1488), .B0(n937), .B1(n903), .Y(n900) );
  AOI22X1TS U1440 ( .A0(requesterAddressIn_SOUTH[2]), .A1(n1689), .B0(n968), 
        .B1(n895), .Y(n899) );
  INVX2TS U1441 ( .A(n972), .Y(n1765) );
  AOI22X1TS U1442 ( .A0(n1765), .A1(n88), .B0(n1466), .B1(
        \requesterAddressbuffer[6][3] ), .Y(n907) );
  INVX2TS U1443 ( .A(n902), .Y(n1696) );
  AOI22X1TS U1444 ( .A0(n945), .A1(n1696), .B0(n944), .B1(n903), .Y(n906) );
  INVX2TS U1445 ( .A(n904), .Y(n1480) );
  AOI22X1TS U1446 ( .A0(requesterAddressIn_SOUTH[3]), .A1(n1480), .B0(n975), 
        .B1(n1697), .Y(n905) );
  INVX2TS U1447 ( .A(n1438), .Y(n1723) );
  AOI22X1TS U1448 ( .A0(n995), .A1(n912), .B0(n1723), .B1(
        \requesterAddressbuffer[5][0] ), .Y(n911) );
  INVX2TS U1449 ( .A(n1429), .Y(n1716) );
  AOI22X1TS U1450 ( .A0(n925), .A1(n1439), .B0(n924), .B1(n1716), .Y(n910) );
  INVX2TS U1451 ( .A(n908), .Y(n1709) );
  AOI22X1TS U1452 ( .A0(n1030), .A1(n1709), .B0(requesterAddressIn_NORTH[0]), 
        .B1(n1440), .Y(n909) );
  AOI22X1TS U1453 ( .A0(n1659), .A1(n912), .B0(n1733), .B1(
        \requesterAddressbuffer[5][1] ), .Y(n915) );
  INVX2TS U1454 ( .A(n1429), .Y(n1726) );
  AOI22X1TS U1455 ( .A0(n933), .A1(n1728), .B0(n932), .B1(n1726), .Y(n914) );
  AOI22X1TS U1456 ( .A0(n1036), .A1(n1729), .B0(requesterAddressIn_NORTH[1]), 
        .B1(n1430), .Y(n913) );
  INVX2TS U1457 ( .A(n14), .Y(n1714) );
  INVX2TS U1458 ( .A(n1594), .Y(n1434) );
  AOI22X1TS U1459 ( .A0(n1667), .A1(n1714), .B0(n1434), .B1(
        \requesterAddressbuffer[5][2] ), .Y(n918) );
  AOI22X1TS U1460 ( .A0(n938), .A1(n1444), .B0(n937), .B1(n920), .Y(n917) );
  AOI22X1TS U1461 ( .A0(n1041), .A1(n1445), .B0(requesterAddressIn_NORTH[2]), 
        .B1(n1430), .Y(n916) );
  INVX2TS U1462 ( .A(n14), .Y(n1724) );
  AOI22X1TS U1463 ( .A0(n1675), .A1(n1724), .B0(n1434), .B1(
        \requesterAddressbuffer[5][3] ), .Y(n923) );
  INVX2TS U1464 ( .A(n919), .Y(n1728) );
  AOI22X1TS U1465 ( .A0(n945), .A1(n1728), .B0(n944), .B1(n920), .Y(n922) );
  AOI22X1TS U1466 ( .A0(n1048), .A1(n228), .B0(requesterAddressIn_NORTH[3]), 
        .B1(n1710), .Y(n921) );
  INVX2TS U1467 ( .A(n1407), .Y(n1754) );
  AOI22X1TS U1468 ( .A0(n995), .A1(n931), .B0(n1754), .B1(
        \requesterAddressbuffer[4][0] ), .Y(n930) );
  INVX2TS U1469 ( .A(n1396), .Y(n1748) );
  AOI22X1TS U1470 ( .A0(n925), .A1(n1741), .B0(n924), .B1(n1748), .Y(n929) );
  INVX2TS U1471 ( .A(n926), .Y(n1760) );
  AOI22X1TS U1472 ( .A0(n1030), .A1(n1760), .B0(requesterAddressIn_NORTH[0]), 
        .B1(n927), .Y(n928) );
  INVX2TS U1473 ( .A(n955), .Y(n1877) );
  AOI22X1TS U1474 ( .A0(n1877), .A1(n931), .B0(n1764), .B1(
        \requesterAddressbuffer[4][1] ), .Y(n936) );
  INVX2TS U1475 ( .A(n1396), .Y(n1757) );
  AOI22X1TS U1476 ( .A0(n933), .A1(n1409), .B0(n932), .B1(n1757), .Y(n935) );
  AOI22X1TS U1477 ( .A0(n1036), .A1(n1766), .B0(requesterAddressIn_NORTH[1]), 
        .B1(n1742), .Y(n934) );
  INVX2TS U1478 ( .A(n964), .Y(n1888) );
  INVX2TS U1479 ( .A(n1406), .Y(n1746) );
  INVX2TS U1480 ( .A(n1606), .Y(n1401) );
  AOI22X1TS U1481 ( .A0(n1888), .A1(n1746), .B0(n1401), .B1(
        \requesterAddressbuffer[4][2] ), .Y(n941) );
  AOI22X1TS U1482 ( .A0(n938), .A1(n1749), .B0(n937), .B1(n943), .Y(n940) );
  AOI22X1TS U1483 ( .A0(n1041), .A1(n1425), .B0(requesterAddressIn_NORTH[2]), 
        .B1(n1742), .Y(n939) );
  INVX2TS U1484 ( .A(n972), .Y(n1900) );
  INVX2TS U1485 ( .A(n1406), .Y(n1755) );
  AOI22X1TS U1486 ( .A0(n1900), .A1(n1755), .B0(n1401), .B1(
        \requesterAddressbuffer[4][3] ), .Y(n948) );
  INVX2TS U1487 ( .A(n942), .Y(n1409) );
  AOI22X1TS U1488 ( .A0(n945), .A1(n1409), .B0(n944), .B1(n943), .Y(n947) );
  AOI22X1TS U1489 ( .A0(n1048), .A1(n1411), .B0(requesterAddressIn_NORTH[3]), 
        .B1(n1750), .Y(n946) );
  INVX2TS U1490 ( .A(n949), .Y(n1868) );
  INVX2TS U1491 ( .A(n1379), .Y(n1784) );
  AOI22X1TS U1492 ( .A0(n1868), .A1(n956), .B0(n1784), .B1(
        \requesterAddressbuffer[3][0] ), .Y(n954) );
  AOI22X1TS U1493 ( .A0(n950), .A1(n175), .B0(n996), .B1(n173), .Y(n953) );
  INVX2TS U1494 ( .A(n966), .Y(n1392) );
  AOI22X1TS U1495 ( .A0(n999), .A1(n1392), .B0(n951), .B1(n1796), .Y(n952) );
  INVX2TS U1496 ( .A(n955), .Y(n1837) );
  AOI22X1TS U1497 ( .A0(n1837), .A1(n956), .B0(n1791), .B1(
        \requesterAddressbuffer[3][1] ), .Y(n963) );
  INVX2TS U1498 ( .A(n957), .Y(n1793) );
  AOI22X1TS U1499 ( .A0(n959), .A1(n958), .B0(n1004), .B1(n1793), .Y(n962) );
  INVX2TS U1500 ( .A(n966), .Y(n1786) );
  AOI22X1TS U1501 ( .A0(n1006), .A1(n1786), .B0(n960), .B1(n1780), .Y(n961) );
  INVX2TS U1502 ( .A(n964), .Y(n1849) );
  INVX2TS U1503 ( .A(n1378), .Y(n1777) );
  INVX2TS U1504 ( .A(n1615), .Y(n1372) );
  AOI22X1TS U1505 ( .A0(n1849), .A1(n1777), .B0(n1372), .B1(
        \requesterAddressbuffer[3][2] ), .Y(n971) );
  AOI22X1TS U1506 ( .A0(n965), .A1(n1772), .B0(n1011), .B1(n1368), .Y(n970) );
  AOI22X1TS U1507 ( .A0(n1014), .A1(n133), .B0(n968), .B1(n967), .Y(n969) );
  INVX2TS U1508 ( .A(n972), .Y(n1861) );
  AOI22X1TS U1509 ( .A0(n1861), .A1(n134), .B0(n1372), .B1(
        \requesterAddressbuffer[3][3] ), .Y(n978) );
  AOI22X1TS U1510 ( .A0(n974), .A1(n175), .B0(n1020), .B1(n1386), .Y(n977) );
  AOI22X1TS U1511 ( .A0(n1023), .A1(n1392), .B0(n975), .B1(n1787), .Y(n976) );
  INVX2TS U1512 ( .A(n1628), .Y(n1813) );
  AOI22X1TS U1513 ( .A0(n1770), .A1(n983), .B0(n1813), .B1(
        \requesterAddressbuffer[2][0] ), .Y(n982) );
  INVX2TS U1514 ( .A(n1346), .Y(n1807) );
  AOI22X1TS U1515 ( .A0(requesterAddressIn_WEST[0]), .A1(n1800), .B0(n996), 
        .B1(n1807), .Y(n981) );
  INVX2TS U1516 ( .A(n979), .Y(n1817) );
  AOI22X1TS U1517 ( .A0(n999), .A1(n1817), .B0(n998), .B1(n1802), .Y(n980) );
  AOI22X1TS U1518 ( .A0(n1877), .A1(n983), .B0(n1822), .B1(
        \requesterAddressbuffer[2][1] ), .Y(n986) );
  INVX2TS U1519 ( .A(n1346), .Y(n1815) );
  AOI22X1TS U1520 ( .A0(requesterAddressIn_WEST[1]), .A1(n1348), .B0(n1004), 
        .B1(n1815), .Y(n985) );
  AOI22X1TS U1521 ( .A0(n1006), .A1(n1354), .B0(n1005), .B1(n1112), .Y(n984)
         );
  INVX2TS U1522 ( .A(n13), .Y(n1806) );
  INVX2TS U1523 ( .A(n1628), .Y(n1340) );
  AOI22X1TS U1524 ( .A0(n1888), .A1(n1806), .B0(n1340), .B1(
        \requesterAddressbuffer[2][2] ), .Y(n989) );
  AOI22X1TS U1525 ( .A0(requesterAddressIn_WEST[2]), .A1(n1808), .B0(n1011), 
        .B1(n991), .Y(n988) );
  AOI22X1TS U1526 ( .A0(n1014), .A1(n1809), .B0(n1013), .B1(n1802), .Y(n987)
         );
  INVX2TS U1527 ( .A(n13), .Y(n1814) );
  AOI22X1TS U1528 ( .A0(n1900), .A1(n1814), .B0(n1340), .B1(
        \requesterAddressbuffer[2][3] ), .Y(n994) );
  INVX2TS U1529 ( .A(n990), .Y(n1348) );
  AOI22X1TS U1530 ( .A0(requesterAddressIn_WEST[3]), .A1(n1348), .B0(n1020), 
        .B1(n991), .Y(n993) );
  AOI22X1TS U1531 ( .A0(n1023), .A1(n190), .B0(n1022), .B1(n1818), .Y(n992) );
  INVX2TS U1532 ( .A(n1010), .Y(n1847) );
  AOI22X1TS U1533 ( .A0(n995), .A1(n1003), .B0(n1847), .B1(
        \requesterAddressbuffer[1][0] ), .Y(n1002) );
  INVX2TS U1534 ( .A(n1090), .Y(n1839) );
  AOI22X1TS U1535 ( .A0(requesterAddressIn_WEST[0]), .A1(n1829), .B0(n996), 
        .B1(n1839), .Y(n1001) );
  INVX2TS U1536 ( .A(n997), .Y(n1854) );
  AOI22X1TS U1537 ( .A0(n999), .A1(n1854), .B0(n998), .B1(n1079), .Y(n1000) );
  AOI22X1TS U1538 ( .A0(n1747), .A1(n1003), .B0(n1860), .B1(
        \requesterAddressbuffer[1][1] ), .Y(n1009) );
  INVX2TS U1539 ( .A(n1090), .Y(n1851) );
  AOI22X1TS U1540 ( .A0(requesterAddressIn_WEST[1]), .A1(n1091), .B0(n1004), 
        .B1(n1851), .Y(n1008) );
  AOI22X1TS U1541 ( .A0(n1006), .A1(n1097), .B0(n1005), .B1(n1832), .Y(n1007)
         );
  INVX2TS U1542 ( .A(n1088), .Y(n1836) );
  INVX2TS U1543 ( .A(n1010), .Y(n1084) );
  AOI22X1TS U1544 ( .A0(n1756), .A1(n1836), .B0(n1084), .B1(
        \requesterAddressbuffer[1][2] ), .Y(n1017) );
  AOI22X1TS U1545 ( .A0(requesterAddressIn_WEST[2]), .A1(n1840), .B0(n1011), 
        .B1(n1019), .Y(n1016) );
  AOI22X1TS U1546 ( .A0(n1014), .A1(n1842), .B0(n1013), .B1(n1012), .Y(n1015)
         );
  INVX2TS U1547 ( .A(n1088), .Y(n1848) );
  AOI22X1TS U1548 ( .A0(n1765), .A1(n1848), .B0(n1084), .B1(
        \requesterAddressbuffer[1][3] ), .Y(n1026) );
  INVX2TS U1549 ( .A(n1018), .Y(n1091) );
  AOI22X1TS U1550 ( .A0(requesterAddressIn_WEST[3]), .A1(n1091), .B0(n1020), 
        .B1(n1019), .Y(n1025) );
  AOI22X1TS U1551 ( .A0(n1023), .A1(n335), .B0(n1022), .B1(n1021), .Y(n1024)
         );
  INVX2TS U1552 ( .A(n1061), .Y(n1886) );
  AOI22X1TS U1553 ( .A0(readRequesterAddress[0]), .A1(n1034), .B0(n1886), .B1(
        \requesterAddressbuffer[0][0] ), .Y(n1033) );
  INVX2TS U1554 ( .A(n1062), .Y(n1878) );
  AOI22X1TS U1555 ( .A0(requesterAddressIn_WEST[0]), .A1(n1869), .B0(n1027), 
        .B1(n1878), .Y(n1032) );
  INVX2TS U1556 ( .A(n1028), .Y(n1903) );
  INVX2TS U1557 ( .A(n1029), .Y(n1070) );
  AOI22X1TS U1558 ( .A0(n1030), .A1(n1903), .B0(requesterAddressIn_NORTH[0]), 
        .B1(n1070), .Y(n1031) );
  AOI22X1TS U1559 ( .A0(n1837), .A1(n1034), .B0(n1898), .B1(
        \requesterAddressbuffer[0][1] ), .Y(n1039) );
  INVX2TS U1560 ( .A(n1062), .Y(n1889) );
  AOI22X1TS U1561 ( .A0(requesterAddressIn_WEST[1]), .A1(n1063), .B0(n1035), 
        .B1(n1889), .Y(n1038) );
  AOI22X1TS U1562 ( .A0(n1036), .A1(n1057), .B0(requesterAddressIn_NORTH[1]), 
        .B1(n1881), .Y(n1037) );
  INVX2TS U1563 ( .A(n15), .Y(n1876) );
  INVX2TS U1564 ( .A(n1061), .Y(n1056) );
  AOI22X1TS U1565 ( .A0(n1849), .A1(n1876), .B0(n1056), .B1(
        \requesterAddressbuffer[0][2] ), .Y(n1044) );
  AOI22X1TS U1566 ( .A0(requesterAddressIn_WEST[2]), .A1(n1879), .B0(n1040), 
        .B1(n1046), .Y(n1043) );
  AOI22X1TS U1567 ( .A0(n1041), .A1(n1872), .B0(requesterAddressIn_NORTH[2]), 
        .B1(n1881), .Y(n1042) );
  INVX2TS U1568 ( .A(n15), .Y(n1887) );
  AOI22X1TS U1569 ( .A0(n1861), .A1(n1887), .B0(n1056), .B1(
        \requesterAddressbuffer[0][3] ), .Y(n1051) );
  INVX2TS U1570 ( .A(n1045), .Y(n1063) );
  AOI22X1TS U1571 ( .A0(requesterAddressIn_WEST[3]), .A1(n1063), .B0(n1047), 
        .B1(n1046), .Y(n1050) );
  AOI22X1TS U1572 ( .A0(n1048), .A1(n1894), .B0(requesterAddressIn_NORTH[3]), 
        .B1(n1052), .Y(n1049) );
  INVX2TS U1573 ( .A(n1078), .Y(n1458) );
  AOI22X1TS U1574 ( .A0(n1876), .A1(n1458), .B0(n1056), .B1(
        \dataoutbuffer[0][0] ), .Y(n1055) );
  AOI22X1TS U1575 ( .A0(n1063), .A1(n1397), .B0(n1878), .B1(n1111), .Y(n1054)
         );
  CLKBUFX2TS U1576 ( .A(dataIn_NORTH[0]), .Y(n1462) );
  AOI22X1TS U1577 ( .A0(n1903), .A1(dataIn_SOUTH[0]), .B0(n1052), .B1(n1462), 
        .Y(n1053) );
  INVX2TS U1578 ( .A(n1083), .Y(n1467) );
  AOI22X1TS U1579 ( .A0(n1887), .A1(n1467), .B0(n1056), .B1(
        \dataoutbuffer[0][1] ), .Y(n1060) );
  AOI22X1TS U1580 ( .A0(n417), .A1(n1402), .B0(n1889), .B1(n1341), .Y(n1059)
         );
  CLKBUFX2TS U1581 ( .A(dataIn_NORTH[1]), .Y(n1470) );
  AOI22X1TS U1582 ( .A0(n1057), .A1(dataIn_SOUTH[1]), .B0(n413), .B1(n1470), 
        .Y(n1058) );
  INVX2TS U1583 ( .A(n15), .Y(n1899) );
  INVX2TS U1584 ( .A(n1089), .Y(n1476) );
  INVX2TS U1585 ( .A(n1061), .Y(n1074) );
  AOI22X1TS U1586 ( .A0(n1899), .A1(n1476), .B0(n1074), .B1(
        \dataoutbuffer[0][2] ), .Y(n1066) );
  AOI22X1TS U1587 ( .A0(n1063), .A1(n1408), .B0(n390), .B1(n1347), .Y(n1065)
         );
  CLKBUFX2TS U1588 ( .A(dataIn_NORTH[2]), .Y(n1481) );
  AOI22X1TS U1589 ( .A0(n1903), .A1(dataIn_SOUTH[2]), .B0(n1070), .B1(n1481), 
        .Y(n1064) );
  INVX2TS U1590 ( .A(n1096), .Y(n1486) );
  AOI22X1TS U1591 ( .A0(n1876), .A1(n1486), .B0(n1074), .B1(
        \dataoutbuffer[0][3] ), .Y(n1069) );
  AOI22X1TS U1592 ( .A0(n1890), .A1(n1415), .B0(n1878), .B1(n1353), .Y(n1068)
         );
  CLKBUFX2TS U1593 ( .A(dataIn_NORTH[3]), .Y(n1490) );
  AOI22X1TS U1594 ( .A0(n425), .A1(dataIn_SOUTH[3]), .B0(n1892), .B1(n1490), 
        .Y(n1067) );
  INVX2TS U1595 ( .A(n1101), .Y(n1494) );
  AOI22X1TS U1596 ( .A0(n1887), .A1(n1494), .B0(n1074), .B1(
        \dataoutbuffer[0][4] ), .Y(n1073) );
  AOI22X1TS U1597 ( .A0(n1869), .A1(n1419), .B0(n1889), .B1(n1359), .Y(n1072)
         );
  CLKBUFX2TS U1598 ( .A(dataIn_NORTH[4]), .Y(n1497) );
  AOI22X1TS U1599 ( .A0(n1894), .A1(dataIn_SOUTH[4]), .B0(n1070), .B1(n1497), 
        .Y(n1071) );
  INVX2TS U1600 ( .A(n1106), .Y(n1502) );
  AOI22X1TS U1601 ( .A0(n1899), .A1(n1502), .B0(n1074), .B1(
        \dataoutbuffer[0][5] ), .Y(n1077) );
  AOI22X1TS U1602 ( .A0(n417), .A1(n1424), .B0(n390), .B1(n1364), .Y(n1076) );
  CLKBUFX2TS U1603 ( .A(dataIn_NORTH[5]), .Y(n1506) );
  AOI22X1TS U1604 ( .A0(n1872), .A1(dataIn_SOUTH[5]), .B0(n406), .B1(n1506), 
        .Y(n1075) );
  INVX2TS U1605 ( .A(n1078), .Y(n1510) );
  AOI22X1TS U1606 ( .A0(n1836), .A1(n1510), .B0(n1084), .B1(
        \dataoutbuffer[1][0] ), .Y(n1082) );
  AOI22X1TS U1607 ( .A0(n1091), .A1(dataIn_WEST[0]), .B0(n1839), .B1(n1111), 
        .Y(n1081) );
  CLKBUFX2TS U1608 ( .A(dataIn_NORTH[0]), .Y(n1513) );
  CLKBUFX2TS U1609 ( .A(dataIn_SOUTH[0]), .Y(n1515) );
  CLKBUFX2TS U1610 ( .A(n1515), .Y(n1461) );
  AOI22X1TS U1611 ( .A0(n1079), .A1(n1513), .B0(n1097), .B1(n1461), .Y(n1080)
         );
  INVX2TS U1612 ( .A(n1083), .Y(n1520) );
  AOI22X1TS U1613 ( .A0(n1848), .A1(n1520), .B0(n1084), .B1(
        \dataoutbuffer[1][1] ), .Y(n1087) );
  AOI22X1TS U1614 ( .A0(n317), .A1(dataIn_WEST[1]), .B0(n1851), .B1(n1341), 
        .Y(n1086) );
  CLKBUFX2TS U1615 ( .A(dataIn_NORTH[1]), .Y(n1522) );
  CLKBUFX2TS U1616 ( .A(dataIn_SOUTH[1]), .Y(n1523) );
  CLKBUFX2TS U1617 ( .A(n1523), .Y(n1469) );
  AOI22X1TS U1618 ( .A0(n1832), .A1(n1522), .B0(n1854), .B1(n1469), .Y(n1085)
         );
  INVX2TS U1619 ( .A(n1089), .Y(n1528) );
  INVX2TS U1620 ( .A(n1010), .Y(n1107) );
  AOI22X1TS U1621 ( .A0(n315), .A1(n1528), .B0(n1107), .B1(
        \dataoutbuffer[1][2] ), .Y(n1095) );
  AOI22X1TS U1622 ( .A0(n1091), .A1(dataIn_WEST[2]), .B0(n313), .B1(n1347), 
        .Y(n1094) );
  CLKBUFX2TS U1623 ( .A(dataIn_NORTH[2]), .Y(n1530) );
  CLKBUFX2TS U1624 ( .A(dataIn_SOUTH[2]), .Y(n1531) );
  CLKBUFX2TS U1625 ( .A(n1531), .Y(n1479) );
  AOI22X1TS U1626 ( .A0(n1012), .A1(n1530), .B0(n1102), .B1(n1479), .Y(n1093)
         );
  INVX2TS U1627 ( .A(n1096), .Y(n1535) );
  AOI22X1TS U1628 ( .A0(n1836), .A1(n1535), .B0(n1107), .B1(
        \dataoutbuffer[1][3] ), .Y(n1100) );
  AOI22X1TS U1629 ( .A0(n1852), .A1(dataIn_WEST[3]), .B0(n1839), .B1(n1353), 
        .Y(n1099) );
  CLKBUFX2TS U1630 ( .A(dataIn_NORTH[3]), .Y(n1537) );
  CLKBUFX2TS U1631 ( .A(dataIn_SOUTH[3]), .Y(n1538) );
  CLKBUFX2TS U1632 ( .A(n1538), .Y(n1489) );
  AOI22X1TS U1633 ( .A0(n322), .A1(n1537), .B0(n1097), .B1(n1489), .Y(n1098)
         );
  INVX2TS U1634 ( .A(n1101), .Y(n1542) );
  AOI22X1TS U1635 ( .A0(n1848), .A1(n1542), .B0(n1107), .B1(
        \dataoutbuffer[1][4] ), .Y(n1105) );
  AOI22X1TS U1636 ( .A0(n1829), .A1(dataIn_WEST[4]), .B0(n1851), .B1(n1359), 
        .Y(n1104) );
  CLKBUFX2TS U1637 ( .A(dataIn_NORTH[4]), .Y(n1545) );
  CLKBUFX2TS U1638 ( .A(dataIn_SOUTH[4]), .Y(n1547) );
  CLKBUFX2TS U1639 ( .A(n1547), .Y(n1496) );
  AOI22X1TS U1640 ( .A0(n322), .A1(n1545), .B0(n1102), .B1(n1496), .Y(n1103)
         );
  INVX2TS U1641 ( .A(n1106), .Y(n1553) );
  AOI22X1TS U1642 ( .A0(n1003), .A1(n1553), .B0(n1107), .B1(
        \dataoutbuffer[1][5] ), .Y(n1110) );
  AOI22X1TS U1643 ( .A0(n317), .A1(dataIn_WEST[5]), .B0(n313), .B1(n1364), .Y(
        n1109) );
  CLKBUFX2TS U1644 ( .A(dataIn_NORTH[5]), .Y(n1555) );
  CLKBUFX2TS U1645 ( .A(dataIn_SOUTH[5]), .Y(n1556) );
  CLKBUFX2TS U1646 ( .A(n1556), .Y(n1504) );
  AOI22X1TS U1647 ( .A0(n1021), .A1(n1555), .B0(n349), .B1(n1504), .Y(n1108)
         );
  AOI22X1TS U1648 ( .A0(n1806), .A1(n1458), .B0(n1340), .B1(
        \dataoutbuffer[2][0] ), .Y(n1339) );
  AOI22X1TS U1649 ( .A0(n1348), .A1(dataIn_WEST[0]), .B0(n1807), .B1(n1111), 
        .Y(n1338) );
  AOI22X1TS U1650 ( .A0(n1112), .A1(n1513), .B0(n1354), .B1(dataIn_SOUTH[0]), 
        .Y(n1337) );
  AOI22X1TS U1651 ( .A0(n1814), .A1(n1467), .B0(n1340), .B1(
        \dataoutbuffer[2][1] ), .Y(n1344) );
  AOI22X1TS U1652 ( .A0(n199), .A1(dataIn_WEST[1]), .B0(n1815), .B1(n1341), 
        .Y(n1343) );
  AOI22X1TS U1653 ( .A0(n1349), .A1(n1522), .B0(n1817), .B1(dataIn_SOUTH[1]), 
        .Y(n1342) );
  INVX2TS U1654 ( .A(n13), .Y(n1823) );
  INVX2TS U1655 ( .A(n1345), .Y(n1363) );
  AOI22X1TS U1656 ( .A0(n1823), .A1(n1476), .B0(n1363), .B1(
        \dataoutbuffer[2][2] ), .Y(n1352) );
  AOI22X1TS U1657 ( .A0(n1348), .A1(dataIn_WEST[2]), .B0(n183), .B1(n1347), 
        .Y(n1351) );
  AOI22X1TS U1658 ( .A0(n1349), .A1(n1530), .B0(n1817), .B1(dataIn_SOUTH[2]), 
        .Y(n1350) );
  AOI22X1TS U1659 ( .A0(n1806), .A1(n1486), .B0(n1363), .B1(
        \dataoutbuffer[2][3] ), .Y(n1358) );
  AOI22X1TS U1660 ( .A0(n1816), .A1(dataIn_WEST[3]), .B0(n1807), .B1(n1353), 
        .Y(n1357) );
  AOI22X1TS U1661 ( .A0(n1355), .A1(n1537), .B0(n1354), .B1(dataIn_SOUTH[3]), 
        .Y(n1356) );
  AOI22X1TS U1662 ( .A0(n1814), .A1(n1494), .B0(n1363), .B1(
        \dataoutbuffer[2][4] ), .Y(n1362) );
  AOI22X1TS U1663 ( .A0(n1800), .A1(dataIn_WEST[4]), .B0(n1815), .B1(n1359), 
        .Y(n1361) );
  AOI22X1TS U1664 ( .A0(n1349), .A1(n1545), .B0(n1801), .B1(dataIn_SOUTH[4]), 
        .Y(n1360) );
  AOI22X1TS U1665 ( .A0(n1823), .A1(n1502), .B0(n1363), .B1(
        \dataoutbuffer[2][5] ), .Y(n1367) );
  AOI22X1TS U1666 ( .A0(n199), .A1(dataIn_WEST[5]), .B0(n183), .B1(n1364), .Y(
        n1366) );
  AOI22X1TS U1667 ( .A0(n188), .A1(n1555), .B0(n203), .B1(dataIn_SOUTH[5]), 
        .Y(n1365) );
  AOI22X1TS U1668 ( .A0(n1777), .A1(n1458), .B0(n1372), .B1(
        \dataoutbuffer[3][0] ), .Y(n1371) );
  AOI22X1TS U1669 ( .A0(n1387), .A1(dataIn_WEST[0]), .B0(n1368), .B1(
        dataIn_EAST[0]), .Y(n1370) );
  AOI22X1TS U1670 ( .A0(n967), .A1(n1462), .B0(n1374), .B1(n1461), .Y(n1369)
         );
  AOI22X1TS U1671 ( .A0(n134), .A1(n1467), .B0(n1372), .B1(
        \dataoutbuffer[3][1] ), .Y(n1377) );
  AOI22X1TS U1672 ( .A0(n1795), .A1(dataIn_WEST[1]), .B0(n1793), .B1(
        dataIn_EAST[1]), .Y(n1376) );
  INVX2TS U1673 ( .A(n1373), .Y(n1796) );
  AOI22X1TS U1674 ( .A0(n1796), .A1(n1470), .B0(n1374), .B1(n1469), .Y(n1375)
         );
  INVX2TS U1675 ( .A(n1378), .Y(n1792) );
  INVX2TS U1676 ( .A(n1379), .Y(n1391) );
  AOI22X1TS U1677 ( .A0(n1792), .A1(n1476), .B0(n1391), .B1(
        \dataoutbuffer[3][2] ), .Y(n1382) );
  AOI22X1TS U1678 ( .A0(n958), .A1(dataIn_WEST[2]), .B0(n173), .B1(
        dataIn_EAST[2]), .Y(n1381) );
  AOI22X1TS U1679 ( .A0(n162), .A1(n1481), .B0(n1392), .B1(n1479), .Y(n1380)
         );
  AOI22X1TS U1680 ( .A0(n1777), .A1(n1486), .B0(n1391), .B1(
        \dataoutbuffer[3][3] ), .Y(n1385) );
  AOI22X1TS U1681 ( .A0(n141), .A1(dataIn_WEST[3]), .B0(n167), .B1(
        dataIn_EAST[3]), .Y(n1384) );
  AOI22X1TS U1682 ( .A0(n1787), .A1(n1490), .B0(n1786), .B1(n1489), .Y(n1383)
         );
  AOI22X1TS U1683 ( .A0(n956), .A1(n1494), .B0(n1391), .B1(
        \dataoutbuffer[3][4] ), .Y(n1390) );
  AOI22X1TS U1684 ( .A0(n1387), .A1(dataIn_WEST[4]), .B0(n1386), .B1(
        dataIn_EAST[4]), .Y(n1389) );
  AOI22X1TS U1685 ( .A0(n1773), .A1(n1497), .B0(n145), .B1(n1496), .Y(n1388)
         );
  AOI22X1TS U1686 ( .A0(n1792), .A1(n1502), .B0(n1391), .B1(
        \dataoutbuffer[3][5] ), .Y(n1395) );
  AOI22X1TS U1687 ( .A0(n175), .A1(dataIn_WEST[5]), .B0(n1793), .B1(
        dataIn_EAST[5]), .Y(n1394) );
  AOI22X1TS U1688 ( .A0(n1796), .A1(n1506), .B0(n1392), .B1(n1504), .Y(n1393)
         );
  AOI22X1TS U1689 ( .A0(n1746), .A1(n1510), .B0(n1401), .B1(
        \dataoutbuffer[4][0] ), .Y(n1400) );
  AOI22X1TS U1690 ( .A0(n1409), .A1(n1397), .B0(n943), .B1(dataIn_EAST[0]), 
        .Y(n1399) );
  AOI22X1TS U1691 ( .A0(n1411), .A1(n1515), .B0(n1410), .B1(n1513), .Y(n1398)
         );
  AOI22X1TS U1692 ( .A0(n1755), .A1(n1520), .B0(n1401), .B1(
        \dataoutbuffer[4][1] ), .Y(n1405) );
  AOI22X1TS U1693 ( .A0(n302), .A1(n1402), .B0(n1748), .B1(dataIn_EAST[1]), 
        .Y(n1404) );
  AOI22X1TS U1694 ( .A0(n278), .A1(n1523), .B0(n927), .B1(n1522), .Y(n1403) );
  INVX2TS U1695 ( .A(n1407), .Y(n1423) );
  AOI22X1TS U1696 ( .A0(n274), .A1(n1528), .B0(n1423), .B1(
        \dataoutbuffer[4][2] ), .Y(n1414) );
  AOI22X1TS U1697 ( .A0(n1409), .A1(n1408), .B0(n1757), .B1(dataIn_EAST[2]), 
        .Y(n1413) );
  AOI22X1TS U1698 ( .A0(n1411), .A1(n1531), .B0(n1410), .B1(n1530), .Y(n1412)
         );
  AOI22X1TS U1699 ( .A0(n1746), .A1(n1535), .B0(n1423), .B1(
        \dataoutbuffer[4][3] ), .Y(n1418) );
  AOI22X1TS U1700 ( .A0(n1758), .A1(n1415), .B0(n272), .B1(dataIn_EAST[3]), 
        .Y(n1417) );
  AOI22X1TS U1701 ( .A0(n1425), .A1(n1538), .B0(n1759), .B1(n1537), .Y(n1416)
         );
  AOI22X1TS U1702 ( .A0(n1755), .A1(n1542), .B0(n1423), .B1(
        \dataoutbuffer[4][4] ), .Y(n1422) );
  AOI22X1TS U1703 ( .A0(n1741), .A1(n1419), .B0(n1748), .B1(dataIn_EAST[4]), 
        .Y(n1421) );
  AOI22X1TS U1704 ( .A0(n298), .A1(n1547), .B0(n1742), .B1(n1545), .Y(n1420)
         );
  AOI22X1TS U1705 ( .A0(n931), .A1(n1553), .B0(n1423), .B1(
        \dataoutbuffer[4][5] ), .Y(n1428) );
  AOI22X1TS U1706 ( .A0(n290), .A1(n1424), .B0(n1757), .B1(dataIn_EAST[5]), 
        .Y(n1427) );
  AOI22X1TS U1707 ( .A0(n1425), .A1(n1556), .B0(n1410), .B1(n1555), .Y(n1426)
         );
  AOI22X1TS U1708 ( .A0(n1714), .A1(n1510), .B0(n1434), .B1(
        \dataoutbuffer[5][0] ), .Y(n1433) );
  AOI22X1TS U1709 ( .A0(n1439), .A1(n1511), .B0(n920), .B1(n1460), .Y(n1432)
         );
  AOI22X1TS U1710 ( .A0(n1430), .A1(n1462), .B0(n1709), .B1(n1461), .Y(n1431)
         );
  AOI22X1TS U1711 ( .A0(n1724), .A1(n1520), .B0(n1434), .B1(
        \dataoutbuffer[5][1] ), .Y(n1437) );
  AOI22X1TS U1712 ( .A0(n253), .A1(n1521), .B0(n1716), .B1(n1468), .Y(n1436)
         );
  AOI22X1TS U1713 ( .A0(n246), .A1(n1470), .B0(n228), .B1(n1469), .Y(n1435) );
  INVX2TS U1714 ( .A(n14), .Y(n1734) );
  INVX2TS U1715 ( .A(n1438), .Y(n1454) );
  AOI22X1TS U1716 ( .A0(n1734), .A1(n1528), .B0(n1454), .B1(
        \dataoutbuffer[5][2] ), .Y(n1443) );
  AOI22X1TS U1717 ( .A0(n1439), .A1(n1529), .B0(n1726), .B1(n1477), .Y(n1442)
         );
  AOI22X1TS U1718 ( .A0(n1440), .A1(n1481), .B0(n1719), .B1(n1479), .Y(n1441)
         );
  AOI22X1TS U1719 ( .A0(n1714), .A1(n1535), .B0(n1454), .B1(
        \dataoutbuffer[5][3] ), .Y(n1449) );
  AOI22X1TS U1720 ( .A0(n1444), .A1(n1536), .B0(n222), .B1(n1487), .Y(n1448)
         );
  AOI22X1TS U1721 ( .A0(n1446), .A1(n1490), .B0(n1445), .B1(n1489), .Y(n1447)
         );
  AOI22X1TS U1722 ( .A0(n1724), .A1(n1542), .B0(n1454), .B1(
        \dataoutbuffer[5][4] ), .Y(n1453) );
  AOI22X1TS U1723 ( .A0(n1718), .A1(n1544), .B0(n1716), .B1(n1495), .Y(n1452)
         );
  INVX2TS U1724 ( .A(n1450), .Y(n1737) );
  AOI22X1TS U1725 ( .A0(n1737), .A1(n1497), .B0(n1729), .B1(n1496), .Y(n1451)
         );
  AOI22X1TS U1726 ( .A0(n1734), .A1(n1553), .B0(n1454), .B1(
        \dataoutbuffer[5][5] ), .Y(n1457) );
  AOI22X1TS U1727 ( .A0(n224), .A1(n1554), .B0(n1726), .B1(n1503), .Y(n1456)
         );
  AOI22X1TS U1728 ( .A0(n1737), .A1(n1506), .B0(n228), .B1(n1504), .Y(n1455)
         );
  AOI22X1TS U1729 ( .A0(n1686), .A1(n1458), .B0(n1466), .B1(
        \dataoutbuffer[6][0] ), .Y(n1465) );
  AOI22X1TS U1730 ( .A0(n1478), .A1(n1511), .B0(n903), .B1(n1460), .Y(n1464)
         );
  AOI22X1TS U1731 ( .A0(n1482), .A1(n1462), .B0(n94), .B1(n1461), .Y(n1463) );
  AOI22X1TS U1732 ( .A0(n88), .A1(n1467), .B0(n1466), .B1(
        \dataoutbuffer[6][1] ), .Y(n1473) );
  AOI22X1TS U1733 ( .A0(n115), .A1(n1521), .B0(n1687), .B1(n1468), .Y(n1472)
         );
  AOI22X1TS U1734 ( .A0(n92), .A1(n1470), .B0(n1480), .B1(n1469), .Y(n1471) );
  INVX2TS U1735 ( .A(n1474), .Y(n1702) );
  INVX2TS U1736 ( .A(n1475), .Y(n1501) );
  AOI22X1TS U1737 ( .A0(n1702), .A1(n1476), .B0(n1501), .B1(
        \dataoutbuffer[6][2] ), .Y(n1485) );
  AOI22X1TS U1738 ( .A0(n1478), .A1(n1529), .B0(n1695), .B1(n1477), .Y(n1484)
         );
  AOI22X1TS U1739 ( .A0(n1482), .A1(n1481), .B0(n1480), .B1(n1479), .Y(n1483)
         );
  AOI22X1TS U1740 ( .A0(n1686), .A1(n1486), .B0(n1501), .B1(
        \dataoutbuffer[6][3] ), .Y(n1493) );
  AOI22X1TS U1741 ( .A0(n1488), .A1(n1536), .B0(n86), .B1(n1487), .Y(n1492) );
  AOI22X1TS U1742 ( .A0(n1697), .A1(n1490), .B0(n94), .B1(n1489), .Y(n1491) );
  AOI22X1TS U1743 ( .A0(n894), .A1(n1494), .B0(n1501), .B1(
        \dataoutbuffer[6][4] ), .Y(n1500) );
  AOI22X1TS U1744 ( .A0(n1688), .A1(n1544), .B0(n1687), .B1(n1495), .Y(n1499)
         );
  AOI22X1TS U1745 ( .A0(n1682), .A1(n1497), .B0(n1505), .B1(n1496), .Y(n1498)
         );
  AOI22X1TS U1746 ( .A0(n1702), .A1(n1502), .B0(n1501), .B1(
        \dataoutbuffer[6][5] ), .Y(n1509) );
  AOI22X1TS U1747 ( .A0(n109), .A1(n1554), .B0(n1695), .B1(n1503), .Y(n1508)
         );
  AOI22X1TS U1748 ( .A0(n92), .A1(n1506), .B0(n1505), .B1(n1504), .Y(n1507) );
  AOI22X1TS U1749 ( .A0(n1660), .A1(n1510), .B0(n1519), .B1(
        \dataoutbuffer[7][0] ), .Y(n1518) );
  AOI22X1TS U1750 ( .A0(n1512), .A1(n1511), .B0(n1654), .B1(dataIn_EAST[0]), 
        .Y(n1517) );
  AOI22X1TS U1751 ( .A0(n1548), .A1(n1515), .B0(n1514), .B1(n1513), .Y(n1516)
         );
  AOI22X1TS U1752 ( .A0(n36), .A1(n1520), .B0(n1519), .B1(
        \dataoutbuffer[7][1] ), .Y(n1526) );
  AOI22X1TS U1753 ( .A0(n76), .A1(n1521), .B0(n1543), .B1(dataIn_EAST[1]), .Y(
        n1525) );
  AOI22X1TS U1754 ( .A0(n1662), .A1(n1523), .B0(n1677), .B1(n1522), .Y(n1524)
         );
  INVX2TS U1755 ( .A(n1527), .Y(n1552) );
  AOI22X1TS U1756 ( .A0(n1676), .A1(n1528), .B0(n1552), .B1(
        \dataoutbuffer[7][2] ), .Y(n1534) );
  AOI22X1TS U1757 ( .A0(n1669), .A1(n1529), .B0(n1668), .B1(dataIn_EAST[2]), 
        .Y(n1533) );
  AOI22X1TS U1758 ( .A0(n1557), .A1(n1531), .B0(n61), .B1(n1530), .Y(n1532) );
  AOI22X1TS U1759 ( .A0(n1660), .A1(n1535), .B0(n1552), .B1(
        \dataoutbuffer[7][3] ), .Y(n1541) );
  AOI22X1TS U1760 ( .A0(n38), .A1(n1536), .B0(n1654), .B1(dataIn_EAST[3]), .Y(
        n1540) );
  AOI22X1TS U1761 ( .A0(n1678), .A1(n1538), .B0(n61), .B1(n1537), .Y(n1539) );
  AOI22X1TS U1762 ( .A0(n36), .A1(n1542), .B0(n1552), .B1(
        \dataoutbuffer[7][4] ), .Y(n1551) );
  AOI22X1TS U1763 ( .A0(n1655), .A1(n1544), .B0(n1543), .B1(dataIn_EAST[4]), 
        .Y(n1550) );
  AOI22X1TS U1764 ( .A0(n1548), .A1(n1547), .B0(n1546), .B1(n1545), .Y(n1549)
         );
  AOI22X1TS U1765 ( .A0(n1676), .A1(n1553), .B0(n1552), .B1(
        \dataoutbuffer[7][5] ), .Y(n1560) );
  AOI22X1TS U1766 ( .A0(n38), .A1(n1554), .B0(n34), .B1(dataIn_EAST[5]), .Y(
        n1559) );
  AOI22X1TS U1767 ( .A0(n1557), .A1(n1556), .B0(n1677), .B1(n1555), .Y(n1558)
         );
  INVX2TS U1768 ( .A(readIn_EAST), .Y(n1646) );
  AOI22X1TS U1769 ( .A0(n1562), .A1(n1585), .B0(n1584), .B1(n1561), .Y(n1564)
         );
  AOI22X1TS U1770 ( .A0(n1565), .A1(n1646), .B0(n1564), .B1(n1563), .Y(n1567)
         );
  AOI22X1TS U1771 ( .A0(n1568), .A1(n1638), .B0(n1567), .B1(n1566), .Y(n1571)
         );
  AOI32X1TS U1772 ( .A0(n1571), .A1(n1570), .A2(n1569), .B0(n1674), .B1(n1937), 
        .Y(n2064) );
  INVX2TS U1773 ( .A(readIn_EAST), .Y(n1622) );
  AOI22X1TS U1774 ( .A0(n1573), .A1(n1585), .B0(n1584), .B1(n1572), .Y(n1575)
         );
  AOI22X1TS U1775 ( .A0(n1576), .A1(n1622), .B0(n1575), .B1(n1574), .Y(n1578)
         );
  AOI22X1TS U1776 ( .A0(n1579), .A1(n1603), .B0(n1578), .B1(n1577), .Y(n1582)
         );
  AOI32X1TS U1777 ( .A0(n1582), .A1(n1581), .A2(n1580), .B0(n1701), .B1(n1938), 
        .Y(n2065) );
  AOI22X1TS U1778 ( .A0(n1586), .A1(n1585), .B0(n1584), .B1(n1583), .Y(n1588)
         );
  AOI22X1TS U1779 ( .A0(n1589), .A1(n1622), .B0(n1588), .B1(n1587), .Y(n1591)
         );
  AOI22X1TS U1780 ( .A0(n1592), .A1(n1603), .B0(n1591), .B1(n1590), .Y(n1595)
         );
  AOI32X1TS U1781 ( .A0(n1595), .A1(n1594), .A2(n1593), .B0(n1733), .B1(n1939), 
        .Y(n2066) );
  CLKBUFX2TS U1782 ( .A(readIn_SOUTH), .Y(n1631) );
  AOI22X1TS U1783 ( .A0(n1597), .A1(n1631), .B0(n1618), .B1(n1596), .Y(n1599)
         );
  AOI22X1TS U1784 ( .A0(n1600), .A1(n1646), .B0(n1599), .B1(n1598), .Y(n1602)
         );
  AOI22X1TS U1785 ( .A0(n1604), .A1(n1603), .B0(n1602), .B1(n1601), .Y(n1607)
         );
  AOI32X1TS U1786 ( .A0(n1607), .A1(n1606), .A2(n1605), .B0(n1764), .B1(n1940), 
        .Y(n2067) );
  AOI22X1TS U1787 ( .A0(n125), .A1(n1631), .B0(readIn_NORTH), .B1(n29), .Y(
        n1609) );
  AOI22X1TS U1788 ( .A0(n1610), .A1(n1622), .B0(n1609), .B1(n1608), .Y(n1612)
         );
  AOI22X1TS U1789 ( .A0(n1613), .A1(readIn_WEST), .B0(n1612), .B1(n1611), .Y(
        n1616) );
  AOI32X1TS U1790 ( .A0(n1616), .A1(n1615), .A2(n1614), .B0(n1791), .B1(n1941), 
        .Y(n2068) );
  AOI22X1TS U1791 ( .A0(n1619), .A1(n1631), .B0(n1618), .B1(n1617), .Y(n1621)
         );
  AOI22X1TS U1792 ( .A0(n1623), .A1(n1622), .B0(n1621), .B1(n1620), .Y(n1625)
         );
  AOI22X1TS U1793 ( .A0(n1626), .A1(readIn_WEST), .B0(n1625), .B1(n1624), .Y(
        n1629) );
  AOI32X1TS U1794 ( .A0(n1629), .A1(n1628), .A2(n1627), .B0(n1822), .B1(n1942), 
        .Y(n2069) );
  AOI22X1TS U1795 ( .A0(n1632), .A1(n1631), .B0(readIn_NORTH), .B1(n1630), .Y(
        n1634) );
  AOI22X1TS U1796 ( .A0(n1635), .A1(n1646), .B0(n1634), .B1(n1633), .Y(n1637)
         );
  AOI22X1TS U1797 ( .A0(n1639), .A1(n1638), .B0(n1637), .B1(n1636), .Y(n1641)
         );
  AOI32X1TS U1798 ( .A0(n1641), .A1(n353), .A2(n1640), .B0(n1860), .B1(n1943), 
        .Y(n2070) );
  AOI22X1TS U1799 ( .A0(n1643), .A1(readIn_SOUTH), .B0(readIn_NORTH), .B1(
        n1642), .Y(n1645) );
  AOI22X1TS U1800 ( .A0(n1647), .A1(n1646), .B0(n1645), .B1(n1644), .Y(n1649)
         );
  AOI22X1TS U1801 ( .A0(n1650), .A1(readIn_WEST), .B0(n1649), .B1(n1648), .Y(
        n1652) );
  AOI32X1TS U1802 ( .A0(n1652), .A1(n422), .A2(n1651), .B0(n1898), .B1(n1944), 
        .Y(n2071) );
  AOI22X1TS U1803 ( .A0(n1827), .A1(n1653), .B0(n1666), .B1(
        \destinationAddressbuffer[7][0] ), .Y(n1658) );
  AOI22X1TS U1804 ( .A0(n1655), .A1(n1708), .B0(n1654), .B1(n1707), .Y(n1657)
         );
  CLKBUFX2TS U1805 ( .A(destinationAddressIn_NORTH[0]), .Y(n1831) );
  AOI22X1TS U1806 ( .A0(n54), .A1(destinationAddressIn_SOUTH[0]), .B0(n1661), 
        .B1(n1831), .Y(n1656) );
  AOI22X1TS U1807 ( .A0(n1660), .A1(n1659), .B0(n1666), .B1(
        \destinationAddressbuffer[7][1] ), .Y(n1665) );
  AOI22X1TS U1808 ( .A0(n1669), .A1(n1717), .B0(n1668), .B1(n1715), .Y(n1664)
         );
  CLKBUFX2TS U1809 ( .A(destinationAddressIn_NORTH[1]), .Y(n1843) );
  AOI22X1TS U1810 ( .A0(n1662), .A1(destinationAddressIn_SOUTH[1]), .B0(n1661), 
        .B1(n1843), .Y(n1663) );
  AOI22X1TS U1811 ( .A0(n1653), .A1(n1667), .B0(n1666), .B1(
        \destinationAddressbuffer[7][2] ), .Y(n1673) );
  AOI22X1TS U1812 ( .A0(n1669), .A1(n1727), .B0(n1668), .B1(n1725), .Y(n1672)
         );
  CLKBUFX2TS U1813 ( .A(destinationAddressIn_NORTH[2]), .Y(n1855) );
  AOI22X1TS U1814 ( .A0(n1670), .A1(destinationAddressIn_SOUTH[2]), .B0(n882), 
        .B1(n1855), .Y(n1671) );
  AOI22X1TS U1815 ( .A0(n1676), .A1(n1675), .B0(n1674), .B1(
        \destinationAddressbuffer[7][3] ), .Y(n1681) );
  AOI22X1TS U1816 ( .A0(n76), .A1(n1736), .B0(n34), .B1(n1735), .Y(n1680) );
  CLKBUFX2TS U1817 ( .A(destinationAddressIn_NORTH[3]), .Y(n1864) );
  AOI22X1TS U1818 ( .A0(n1678), .A1(destinationAddressIn_SOUTH[3]), .B0(n1677), 
        .B1(n1864), .Y(n1679) );
  AOI22X1TS U1819 ( .A0(n1868), .A1(n1702), .B0(n1694), .B1(
        \destinationAddressbuffer[6][0] ), .Y(n1685) );
  AOI22X1TS U1820 ( .A0(n1696), .A1(n1708), .B0(n86), .B1(n1707), .Y(n1684) );
  CLKBUFX2TS U1821 ( .A(destinationAddressIn_NORTH[0]), .Y(n1870) );
  CLKBUFX2TS U1822 ( .A(destinationAddressIn_SOUTH[0]), .Y(n1871) );
  CLKBUFX2TS U1823 ( .A(n1871), .Y(n1830) );
  AOI22X1TS U1824 ( .A0(n1682), .A1(n1870), .B0(n1480), .B1(n1830), .Y(n1683)
         );
  AOI22X1TS U1825 ( .A0(n1747), .A1(n1686), .B0(n1694), .B1(
        \destinationAddressbuffer[6][1] ), .Y(n1693) );
  AOI22X1TS U1826 ( .A0(n1688), .A1(n1717), .B0(n1687), .B1(n1715), .Y(n1692)
         );
  CLKBUFX2TS U1827 ( .A(destinationAddressIn_NORTH[1]), .Y(n1880) );
  CLKBUFX2TS U1828 ( .A(destinationAddressIn_SOUTH[1]), .Y(n1882) );
  CLKBUFX2TS U1829 ( .A(n1882), .Y(n1841) );
  AOI22X1TS U1830 ( .A0(n1690), .A1(n1880), .B0(n1689), .B1(n1841), .Y(n1691)
         );
  AOI22X1TS U1831 ( .A0(n1756), .A1(n88), .B0(n1694), .B1(
        \destinationAddressbuffer[6][2] ), .Y(n1700) );
  AOI22X1TS U1832 ( .A0(n1696), .A1(n1727), .B0(n1695), .B1(n1725), .Y(n1699)
         );
  CLKBUFX2TS U1833 ( .A(destinationAddressIn_NORTH[2]), .Y(n1891) );
  CLKBUFX2TS U1834 ( .A(destinationAddressIn_SOUTH[2]), .Y(n1893) );
  CLKBUFX2TS U1835 ( .A(n1893), .Y(n1853) );
  AOI22X1TS U1836 ( .A0(n1697), .A1(n1891), .B0(n112), .B1(n1853), .Y(n1698)
         );
  AOI22X1TS U1837 ( .A0(n1765), .A1(n1702), .B0(n1701), .B1(
        \destinationAddressbuffer[6][3] ), .Y(n1706) );
  AOI22X1TS U1838 ( .A0(n109), .A1(n1736), .B0(n86), .B1(n1735), .Y(n1705) );
  CLKBUFX2TS U1839 ( .A(destinationAddressIn_NORTH[3]), .Y(n1901) );
  CLKBUFX2TS U1840 ( .A(destinationAddressIn_SOUTH[3]), .Y(n1902) );
  CLKBUFX2TS U1841 ( .A(n1902), .Y(n1863) );
  AOI22X1TS U1842 ( .A0(n92), .A1(n1901), .B0(n1703), .B1(n1863), .Y(n1704) );
  AOI22X1TS U1843 ( .A0(n1868), .A1(n1734), .B0(n1723), .B1(
        \destinationAddressbuffer[5][0] ), .Y(n1713) );
  AOI22X1TS U1844 ( .A0(n1728), .A1(n1708), .B0(n222), .B1(n1707), .Y(n1712)
         );
  AOI22X1TS U1845 ( .A0(n1710), .A1(n1870), .B0(n1709), .B1(
        destinationAddressIn_SOUTH[0]), .Y(n1711) );
  AOI22X1TS U1846 ( .A0(readRequesterAddress[1]), .A1(n1714), .B0(n1723), .B1(
        \destinationAddressbuffer[5][1] ), .Y(n1722) );
  AOI22X1TS U1847 ( .A0(n1718), .A1(n1717), .B0(n1716), .B1(n1715), .Y(n1721)
         );
  AOI22X1TS U1848 ( .A0(n1710), .A1(n1880), .B0(n1719), .B1(
        destinationAddressIn_SOUTH[1]), .Y(n1720) );
  AOI22X1TS U1849 ( .A0(readRequesterAddress[2]), .A1(n1724), .B0(n1723), .B1(
        \destinationAddressbuffer[5][2] ), .Y(n1732) );
  AOI22X1TS U1850 ( .A0(n1728), .A1(n1727), .B0(n1726), .B1(n1725), .Y(n1731)
         );
  AOI22X1TS U1851 ( .A0(n1737), .A1(n1891), .B0(n1729), .B1(
        destinationAddressIn_SOUTH[2]), .Y(n1730) );
  AOI22X1TS U1852 ( .A0(readRequesterAddress[3]), .A1(n1734), .B0(n1733), .B1(
        \destinationAddressbuffer[5][3] ), .Y(n1740) );
  AOI22X1TS U1853 ( .A0(n224), .A1(n1736), .B0(n222), .B1(n1735), .Y(n1739) );
  AOI22X1TS U1854 ( .A0(n1737), .A1(n1901), .B0(n1729), .B1(
        destinationAddressIn_SOUTH[3]), .Y(n1738) );
  AOI22X1TS U1855 ( .A0(n1770), .A1(n274), .B0(n1754), .B1(
        \destinationAddressbuffer[4][0] ), .Y(n1745) );
  AOI22X1TS U1856 ( .A0(n1741), .A1(n1771), .B0(n272), .B1(
        destinationAddressIn_EAST[0]), .Y(n1744) );
  AOI22X1TS U1857 ( .A0(n1760), .A1(n1871), .B0(n1742), .B1(n1870), .Y(n1743)
         );
  AOI22X1TS U1858 ( .A0(n1747), .A1(n1746), .B0(n1754), .B1(
        \destinationAddressbuffer[4][1] ), .Y(n1753) );
  AOI22X1TS U1859 ( .A0(n1749), .A1(n1779), .B0(n1748), .B1(
        destinationAddressIn_EAST[1]), .Y(n1752) );
  AOI22X1TS U1860 ( .A0(n298), .A1(n1882), .B0(n1750), .B1(n1880), .Y(n1751)
         );
  AOI22X1TS U1861 ( .A0(n1756), .A1(n1755), .B0(n1754), .B1(
        \destinationAddressbuffer[4][2] ), .Y(n1763) );
  AOI22X1TS U1862 ( .A0(n1758), .A1(n1785), .B0(n1757), .B1(
        destinationAddressIn_EAST[2]), .Y(n1762) );
  AOI22X1TS U1863 ( .A0(n1760), .A1(n1893), .B0(n1759), .B1(n1891), .Y(n1761)
         );
  AOI22X1TS U1864 ( .A0(n1765), .A1(n274), .B0(n1764), .B1(
        \destinationAddressbuffer[4][3] ), .Y(n1769) );
  AOI22X1TS U1865 ( .A0(n290), .A1(n1794), .B0(n272), .B1(
        destinationAddressIn_EAST[3]), .Y(n1768) );
  AOI22X1TS U1866 ( .A0(n1766), .A1(n1902), .B0(n282), .B1(n1901), .Y(n1767)
         );
  AOI22X1TS U1867 ( .A0(n1770), .A1(n1792), .B0(n1784), .B1(
        \destinationAddressbuffer[3][0] ), .Y(n1776) );
  AOI22X1TS U1868 ( .A0(n1772), .A1(n1771), .B0(n1778), .B1(
        destinationAddressIn_EAST[0]), .Y(n1775) );
  AOI22X1TS U1869 ( .A0(n1773), .A1(n1831), .B0(n1786), .B1(n1830), .Y(n1774)
         );
  AOI22X1TS U1870 ( .A0(n1837), .A1(n1777), .B0(n1784), .B1(
        \destinationAddressbuffer[3][1] ), .Y(n1783) );
  AOI22X1TS U1871 ( .A0(n141), .A1(n1779), .B0(n1778), .B1(
        destinationAddressIn_EAST[1]), .Y(n1782) );
  AOI22X1TS U1872 ( .A0(n1780), .A1(n1843), .B0(n1374), .B1(n1841), .Y(n1781)
         );
  AOI22X1TS U1873 ( .A0(n1849), .A1(n134), .B0(n1784), .B1(
        \destinationAddressbuffer[3][2] ), .Y(n1790) );
  AOI22X1TS U1874 ( .A0(n958), .A1(n1785), .B0(n173), .B1(
        destinationAddressIn_EAST[2]), .Y(n1789) );
  AOI22X1TS U1875 ( .A0(n1787), .A1(n1855), .B0(n1786), .B1(n1853), .Y(n1788)
         );
  AOI22X1TS U1876 ( .A0(n1861), .A1(n1792), .B0(n1791), .B1(
        \destinationAddressbuffer[3][3] ), .Y(n1799) );
  AOI22X1TS U1877 ( .A0(n1795), .A1(n1794), .B0(n1793), .B1(
        destinationAddressIn_EAST[3]), .Y(n1798) );
  AOI22X1TS U1878 ( .A0(n1796), .A1(n1864), .B0(n133), .B1(n1863), .Y(n1797)
         );
  AOI22X1TS U1879 ( .A0(n1827), .A1(n1823), .B0(n1813), .B1(
        \destinationAddressbuffer[2][0] ), .Y(n1805) );
  AOI22X1TS U1880 ( .A0(n1800), .A1(destinationAddressIn_WEST[0]), .B0(n991), 
        .B1(n1828), .Y(n1804) );
  AOI22X1TS U1881 ( .A0(n1802), .A1(n1831), .B0(n1801), .B1(n1830), .Y(n1803)
         );
  AOI22X1TS U1882 ( .A0(n1877), .A1(n1806), .B0(n1813), .B1(
        \destinationAddressbuffer[2][1] ), .Y(n1812) );
  AOI22X1TS U1883 ( .A0(n1808), .A1(destinationAddressIn_WEST[1]), .B0(n1807), 
        .B1(n1838), .Y(n1811) );
  AOI22X1TS U1884 ( .A0(n1349), .A1(n1843), .B0(n1809), .B1(n1841), .Y(n1810)
         );
  AOI22X1TS U1885 ( .A0(n1888), .A1(n1814), .B0(n1813), .B1(
        \destinationAddressbuffer[2][2] ), .Y(n1821) );
  AOI22X1TS U1886 ( .A0(n1816), .A1(destinationAddressIn_WEST[2]), .B0(n1815), 
        .B1(n1850), .Y(n1820) );
  AOI22X1TS U1887 ( .A0(n1818), .A1(n1855), .B0(n1817), .B1(n1853), .Y(n1819)
         );
  AOI22X1TS U1888 ( .A0(n1900), .A1(n1823), .B0(n1822), .B1(
        \destinationAddressbuffer[2][3] ), .Y(n1826) );
  AOI22X1TS U1889 ( .A0(n208), .A1(destinationAddressIn_WEST[3]), .B0(n183), 
        .B1(n1862), .Y(n1825) );
  AOI22X1TS U1890 ( .A0(n188), .A1(n1864), .B0(n190), .B1(n1863), .Y(n1824) );
  AOI22X1TS U1891 ( .A0(n1827), .A1(n315), .B0(n1847), .B1(
        \destinationAddressbuffer[1][0] ), .Y(n1835) );
  AOI22X1TS U1892 ( .A0(n1829), .A1(destinationAddressIn_WEST[0]), .B0(n333), 
        .B1(n1828), .Y(n1834) );
  AOI22X1TS U1893 ( .A0(n1832), .A1(n1831), .B0(n1854), .B1(n1830), .Y(n1833)
         );
  AOI22X1TS U1894 ( .A0(n1837), .A1(n1836), .B0(n1847), .B1(
        \destinationAddressbuffer[1][1] ), .Y(n1846) );
  AOI22X1TS U1895 ( .A0(n1840), .A1(destinationAddressIn_WEST[1]), .B0(n1839), 
        .B1(n1838), .Y(n1845) );
  AOI22X1TS U1896 ( .A0(n322), .A1(n1843), .B0(n1842), .B1(n1841), .Y(n1844)
         );
  AOI22X1TS U1897 ( .A0(n1849), .A1(n1848), .B0(n1847), .B1(
        \destinationAddressbuffer[1][2] ), .Y(n1859) );
  AOI22X1TS U1898 ( .A0(n1852), .A1(destinationAddressIn_WEST[2]), .B0(n1851), 
        .B1(n1850), .Y(n1858) );
  AOI22X1TS U1899 ( .A0(n1856), .A1(n1855), .B0(n1854), .B1(n1853), .Y(n1857)
         );
  AOI22X1TS U1900 ( .A0(n1861), .A1(n315), .B0(n1860), .B1(
        \destinationAddressbuffer[1][3] ), .Y(n1867) );
  AOI22X1TS U1901 ( .A0(n360), .A1(destinationAddressIn_WEST[3]), .B0(n1019), 
        .B1(n1862), .Y(n1866) );
  AOI22X1TS U1902 ( .A0(n1079), .A1(n1864), .B0(n335), .B1(n1863), .Y(n1865)
         );
  AOI22X1TS U1903 ( .A0(n1868), .A1(n1899), .B0(n1886), .B1(
        \destinationAddressbuffer[0][0] ), .Y(n1875) );
  AOI22X1TS U1904 ( .A0(n1869), .A1(destinationAddressIn_WEST[0]), .B0(n1046), 
        .B1(destinationAddressIn_EAST[0]), .Y(n1874) );
  AOI22X1TS U1905 ( .A0(n1872), .A1(n1871), .B0(n1881), .B1(n1870), .Y(n1873)
         );
  AOI22X1TS U1906 ( .A0(n1877), .A1(n1876), .B0(n1886), .B1(
        \destinationAddressbuffer[0][1] ), .Y(n1885) );
  AOI22X1TS U1907 ( .A0(n1879), .A1(destinationAddressIn_WEST[1]), .B0(n1878), 
        .B1(destinationAddressIn_EAST[1]), .Y(n1884) );
  AOI22X1TS U1908 ( .A0(n425), .A1(n1882), .B0(n1881), .B1(n1880), .Y(n1883)
         );
  AOI22X1TS U1909 ( .A0(n1888), .A1(n1887), .B0(n1886), .B1(
        \destinationAddressbuffer[0][2] ), .Y(n1897) );
  AOI22X1TS U1910 ( .A0(n1890), .A1(destinationAddressIn_WEST[2]), .B0(n1889), 
        .B1(destinationAddressIn_EAST[2]), .Y(n1896) );
  AOI22X1TS U1911 ( .A0(n1894), .A1(n1893), .B0(n1892), .B1(n1891), .Y(n1895)
         );
  AOI22X1TS U1912 ( .A0(n1900), .A1(n1899), .B0(n1898), .B1(
        \destinationAddressbuffer[0][3] ), .Y(n1906) );
  AOI22X1TS U1913 ( .A0(n423), .A1(destinationAddressIn_WEST[3]), .B0(n390), 
        .B1(destinationAddressIn_EAST[3]), .Y(n1905) );
  AOI22X1TS U1914 ( .A0(n1903), .A1(n1902), .B0(n1070), .B1(n1901), .Y(n1904)
         );
endmodule


module outputPortArbiter_3 ( clk, reset, selectBit_NORTH, 
        destinationAddressIn_NORTH, requesterAddressIn_NORTH, readIn_NORTH, 
        writeIn_NORTH, dataIn_NORTH, selectBit_SOUTH, 
        destinationAddressIn_SOUTH, requesterAddressIn_SOUTH, readIn_SOUTH, 
        writeIn_SOUTH, dataIn_SOUTH, selectBit_EAST, destinationAddressIn_EAST, 
        requesterAddressIn_EAST, readIn_EAST, writeIn_EAST, dataIn_EAST, 
        selectBit_WEST, destinationAddressIn_WEST, requesterAddressIn_WEST, 
        readIn_WEST, writeIn_WEST, dataIn_WEST, readReady, 
        readRequesterAddress, cacheDataOut, destinationAddressOut, 
        requesterAddressOut, readOut, writeOut, dataOut );
  input [11:0] destinationAddressIn_NORTH;
  input [3:0] requesterAddressIn_NORTH;
  input [5:0] dataIn_NORTH;
  input [11:0] destinationAddressIn_SOUTH;
  input [3:0] requesterAddressIn_SOUTH;
  input [5:0] dataIn_SOUTH;
  input [11:0] destinationAddressIn_EAST;
  input [3:0] requesterAddressIn_EAST;
  input [5:0] dataIn_EAST;
  input [11:0] destinationAddressIn_WEST;
  input [3:0] requesterAddressIn_WEST;
  input [5:0] dataIn_WEST;
  input [3:0] readRequesterAddress;
  input [5:0] cacheDataOut;
  output [11:0] destinationAddressOut;
  output [3:0] requesterAddressOut;
  output [5:0] dataOut;
  input clk, reset, selectBit_NORTH, readIn_NORTH, writeIn_NORTH,
         selectBit_SOUTH, readIn_SOUTH, writeIn_SOUTH, selectBit_EAST,
         readIn_EAST, writeIn_EAST, selectBit_WEST, readIn_WEST, writeIn_WEST,
         readReady;
  output readOut, writeOut;
  wire   \requesterAddressbuffer[0][3] , \requesterAddressbuffer[0][2] ,
         \requesterAddressbuffer[0][1] , \requesterAddressbuffer[0][0] ,
         \requesterAddressbuffer[1][3] , \requesterAddressbuffer[1][2] ,
         \requesterAddressbuffer[1][1] , \requesterAddressbuffer[1][0] ,
         \requesterAddressbuffer[2][3] , \requesterAddressbuffer[2][2] ,
         \requesterAddressbuffer[2][1] , \requesterAddressbuffer[2][0] ,
         \requesterAddressbuffer[3][3] , \requesterAddressbuffer[3][2] ,
         \requesterAddressbuffer[3][1] , \requesterAddressbuffer[3][0] ,
         \requesterAddressbuffer[4][3] , \requesterAddressbuffer[4][2] ,
         \requesterAddressbuffer[4][1] , \requesterAddressbuffer[4][0] ,
         \requesterAddressbuffer[5][3] , \requesterAddressbuffer[5][2] ,
         \requesterAddressbuffer[5][1] , \requesterAddressbuffer[5][0] ,
         \requesterAddressbuffer[6][3] , \requesterAddressbuffer[6][2] ,
         \requesterAddressbuffer[6][1] , \requesterAddressbuffer[6][0] ,
         \requesterAddressbuffer[7][3] , \requesterAddressbuffer[7][2] ,
         \requesterAddressbuffer[7][1] , \requesterAddressbuffer[7][0] ,
         \destinationAddressbuffer[0][11] , \destinationAddressbuffer[0][10] ,
         \destinationAddressbuffer[0][9] , \destinationAddressbuffer[0][8] ,
         \destinationAddressbuffer[0][7] , \destinationAddressbuffer[0][6] ,
         \destinationAddressbuffer[0][5] , \destinationAddressbuffer[0][4] ,
         \destinationAddressbuffer[0][3] , \destinationAddressbuffer[0][2] ,
         \destinationAddressbuffer[0][1] , \destinationAddressbuffer[0][0] ,
         \destinationAddressbuffer[1][11] , \destinationAddressbuffer[1][10] ,
         \destinationAddressbuffer[1][9] , \destinationAddressbuffer[1][8] ,
         \destinationAddressbuffer[1][7] , \destinationAddressbuffer[1][6] ,
         \destinationAddressbuffer[1][5] , \destinationAddressbuffer[1][4] ,
         \destinationAddressbuffer[1][3] , \destinationAddressbuffer[1][2] ,
         \destinationAddressbuffer[1][1] , \destinationAddressbuffer[1][0] ,
         \destinationAddressbuffer[2][11] , \destinationAddressbuffer[2][10] ,
         \destinationAddressbuffer[2][9] , \destinationAddressbuffer[2][8] ,
         \destinationAddressbuffer[2][7] , \destinationAddressbuffer[2][6] ,
         \destinationAddressbuffer[2][5] , \destinationAddressbuffer[2][4] ,
         \destinationAddressbuffer[2][3] , \destinationAddressbuffer[2][2] ,
         \destinationAddressbuffer[2][1] , \destinationAddressbuffer[2][0] ,
         \destinationAddressbuffer[3][11] , \destinationAddressbuffer[3][10] ,
         \destinationAddressbuffer[3][9] , \destinationAddressbuffer[3][8] ,
         \destinationAddressbuffer[3][7] , \destinationAddressbuffer[3][6] ,
         \destinationAddressbuffer[3][5] , \destinationAddressbuffer[3][4] ,
         \destinationAddressbuffer[3][3] , \destinationAddressbuffer[3][2] ,
         \destinationAddressbuffer[3][1] , \destinationAddressbuffer[3][0] ,
         \destinationAddressbuffer[4][11] , \destinationAddressbuffer[4][10] ,
         \destinationAddressbuffer[4][9] , \destinationAddressbuffer[4][8] ,
         \destinationAddressbuffer[4][7] , \destinationAddressbuffer[4][6] ,
         \destinationAddressbuffer[4][5] , \destinationAddressbuffer[4][4] ,
         \destinationAddressbuffer[4][3] , \destinationAddressbuffer[4][2] ,
         \destinationAddressbuffer[4][1] , \destinationAddressbuffer[4][0] ,
         \destinationAddressbuffer[5][11] , \destinationAddressbuffer[5][10] ,
         \destinationAddressbuffer[5][9] , \destinationAddressbuffer[5][8] ,
         \destinationAddressbuffer[5][7] , \destinationAddressbuffer[5][6] ,
         \destinationAddressbuffer[5][5] , \destinationAddressbuffer[5][4] ,
         \destinationAddressbuffer[5][3] , \destinationAddressbuffer[5][2] ,
         \destinationAddressbuffer[5][1] , \destinationAddressbuffer[5][0] ,
         \destinationAddressbuffer[6][11] , \destinationAddressbuffer[6][10] ,
         \destinationAddressbuffer[6][9] , \destinationAddressbuffer[6][8] ,
         \destinationAddressbuffer[6][7] , \destinationAddressbuffer[6][6] ,
         \destinationAddressbuffer[6][5] , \destinationAddressbuffer[6][4] ,
         \destinationAddressbuffer[6][3] , \destinationAddressbuffer[6][2] ,
         \destinationAddressbuffer[6][1] , \destinationAddressbuffer[6][0] ,
         \destinationAddressbuffer[7][11] , \destinationAddressbuffer[7][10] ,
         \destinationAddressbuffer[7][9] , \destinationAddressbuffer[7][8] ,
         \destinationAddressbuffer[7][7] , \destinationAddressbuffer[7][6] ,
         \destinationAddressbuffer[7][5] , \destinationAddressbuffer[7][4] ,
         \destinationAddressbuffer[7][3] , \destinationAddressbuffer[7][2] ,
         \destinationAddressbuffer[7][1] , \destinationAddressbuffer[7][0] ,
         \dataoutbuffer[7][5] , \dataoutbuffer[7][4] , \dataoutbuffer[7][3] ,
         \dataoutbuffer[7][2] , \dataoutbuffer[7][1] , \dataoutbuffer[7][0] ,
         \dataoutbuffer[6][5] , \dataoutbuffer[6][4] , \dataoutbuffer[6][3] ,
         \dataoutbuffer[6][2] , \dataoutbuffer[6][1] , \dataoutbuffer[6][0] ,
         \dataoutbuffer[5][5] , \dataoutbuffer[5][4] , \dataoutbuffer[5][3] ,
         \dataoutbuffer[5][2] , \dataoutbuffer[5][1] , \dataoutbuffer[5][0] ,
         \dataoutbuffer[4][5] , \dataoutbuffer[4][4] , \dataoutbuffer[4][3] ,
         \dataoutbuffer[4][2] , \dataoutbuffer[4][1] , \dataoutbuffer[4][0] ,
         \dataoutbuffer[3][5] , \dataoutbuffer[3][4] , \dataoutbuffer[3][3] ,
         \dataoutbuffer[3][2] , \dataoutbuffer[3][1] , \dataoutbuffer[3][0] ,
         \dataoutbuffer[2][5] , \dataoutbuffer[2][4] , \dataoutbuffer[2][3] ,
         \dataoutbuffer[2][2] , \dataoutbuffer[2][1] , \dataoutbuffer[2][0] ,
         \dataoutbuffer[1][5] , \dataoutbuffer[1][4] , \dataoutbuffer[1][3] ,
         \dataoutbuffer[1][2] , \dataoutbuffer[1][1] , \dataoutbuffer[1][0] ,
         \dataoutbuffer[0][5] , \dataoutbuffer[0][4] , \dataoutbuffer[0][3] ,
         \dataoutbuffer[0][2] , \dataoutbuffer[0][1] , \dataoutbuffer[0][0] ,
         N2624, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182;
  wire   [0:7] writeOutbuffer;
  wire   [0:7] readOutbuffer;

  DFFNSRX1TS full_reg_reg ( .D(N2624), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(
        n1951) );
  DFFNSRX1TS \requesterAddressbuffer_reg[2][0]  ( .D(n2011), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[2][1]  ( .D(n2012), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[2][2]  ( .D(n2013), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[2][3]  ( .D(n2014), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][0]  ( .D(n2147), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][1]  ( .D(n2148), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][2]  ( .D(n2149), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][3]  ( .D(n2150), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][0]  ( .D(n2023), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][1]  ( .D(n2024), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][2]  ( .D(n2025), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][3]  ( .D(n2026), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][4]  ( .D(n2027), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[0][5]  ( .D(n2028), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[0][5] ) );
  DFFNSRX1TS \writeOutbuffer_reg[7]  ( .D(n2071), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[7]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][4]  ( .D(n2091), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][5]  ( .D(n2092), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][6]  ( .D(n2093), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][7]  ( .D(n2094), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][8]  ( .D(n2095), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][9]  ( .D(n2096), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][11]  ( .D(n2098), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[6]  ( .D(n2072), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[6]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][4]  ( .D(n2103), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][5]  ( .D(n2104), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][6]  ( .D(n2105), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][7]  ( .D(n2106), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][8]  ( .D(n2107), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][9]  ( .D(n2108), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][10]  ( .D(n2109), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][11]  ( .D(n2110), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[3]  ( .D(n2075), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[3]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][4]  ( .D(n2139), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][5]  ( .D(n2140), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][6]  ( .D(n2141), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][7]  ( .D(n2142), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][8]  ( .D(n2143), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][9]  ( .D(n2144), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][10]  ( .D(n2145), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][11]  ( .D(n2146), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[2]  ( .D(n2076), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[2]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][4]  ( .D(n2151), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][5]  ( .D(n2152), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][6]  ( .D(n2153), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][7]  ( .D(n2154), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][8]  ( .D(n2155), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][9]  ( .D(n2156), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][10]  ( .D(n2157), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[2][11]  ( .D(n2158), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[2][11] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][0]  ( .D(n2065), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][1]  ( .D(n2066), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][2]  ( .D(n2067), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][3]  ( .D(n2068), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][4]  ( .D(n2069), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[7][5]  ( .D(n2070), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[7][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][0]  ( .D(n2059), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][1]  ( .D(n2060), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][2]  ( .D(n2061), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][3]  ( .D(n2062), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][4]  ( .D(n2063), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[6][5]  ( .D(n2064), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[6][5] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[5][0]  ( .D(n1999), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[5][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[5][1]  ( .D(n2000), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[5][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[5][2]  ( .D(n2001), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[5][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[5][3]  ( .D(n2002), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[5][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][0]  ( .D(n2111), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][1]  ( .D(n2112), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][2]  ( .D(n2113), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][3]  ( .D(n2114), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[4][0]  ( .D(n2003), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[4][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[4][1]  ( .D(n2004), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[4][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[4][2]  ( .D(n2005), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[4][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[4][3]  ( .D(n2006), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[4][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][0]  ( .D(n2123), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][1]  ( .D(n2124), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][2]  ( .D(n2125), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][3]  ( .D(n2126), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][0]  ( .D(n2041), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][1]  ( .D(n2042), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][2]  ( .D(n2043), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][3]  ( .D(n2044), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][4]  ( .D(n2045), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[3][5]  ( .D(n2046), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[3][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][0]  ( .D(n2035), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][1]  ( .D(n2036), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][2]  ( .D(n2037), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][3]  ( .D(n2038), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][4]  ( .D(n2039), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[2][5]  ( .D(n2040), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[2][5] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[1][0]  ( .D(n2015), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[1][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[1][1]  ( .D(n2016), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[1][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[1][2]  ( .D(n2017), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[1][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[1][3]  ( .D(n2018), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[1][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][0]  ( .D(n2159), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][1]  ( .D(n2160), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][2]  ( .D(n2161), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][3]  ( .D(n2162), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[0][0]  ( .D(n2019), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[0][1]  ( .D(n2020), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[0][2]  ( .D(n2021), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[0][3]  ( .D(n2022), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][0]  ( .D(n2171), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][1]  ( .D(n2172), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][2]  ( .D(n2173), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][3]  ( .D(n2174), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[7][0]  ( .D(n1991), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[7][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[7][1]  ( .D(n1992), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[7][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[7][2]  ( .D(n1993), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[7][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[7][3]  ( .D(n1994), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[7][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][0]  ( .D(n2087), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][1]  ( .D(n2088), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][2]  ( .D(n2089), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][3]  ( .D(n2090), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][3] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[6][0]  ( .D(n1995), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[6][1]  ( .D(n1996), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[6][2]  ( .D(n1997), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[6][3]  ( .D(n1998), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][0]  ( .D(n2099), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][1]  ( .D(n2100), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][2]  ( .D(n2101), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[6][3]  ( .D(n2102), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[6][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][0]  ( .D(n2053), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][1]  ( .D(n2054), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][2]  ( .D(n2055), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][3]  ( .D(n2056), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][4]  ( .D(n2057), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[5][5]  ( .D(n2058), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[5][5] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][0]  ( .D(n2047), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][1]  ( .D(n2048), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][2]  ( .D(n2049), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][3]  ( .D(n2050), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][4]  ( .D(n2051), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[4][5]  ( .D(n2052), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[4][5] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[3][0]  ( .D(n2007), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][0] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[3][1]  ( .D(n2008), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][1] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[3][2]  ( .D(n2009), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][2] ) );
  DFFNSRX1TS \requesterAddressbuffer_reg[3][3]  ( .D(n2010), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][3] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][0]  ( .D(n2135), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][0] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][1]  ( .D(n2136), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][1] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][2]  ( .D(n2137), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][2] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[3][3]  ( .D(n2138), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[3][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][0]  ( .D(n2029), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][0] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][1]  ( .D(n2030), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][1] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][2]  ( .D(n2031), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][2] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][3]  ( .D(n2032), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][3] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][4]  ( .D(n2033), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][4] ) );
  DFFNSRX1TS \dataoutbuffer_reg[1][5]  ( .D(n2034), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\dataoutbuffer[1][5] ) );
  DFFNSRX1TS \writeOutbuffer_reg[5]  ( .D(n2073), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[5]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][4]  ( .D(n2115), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][5]  ( .D(n2116), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][6]  ( .D(n2117), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][7]  ( .D(n2118), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][8]  ( .D(n2119), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][9]  ( .D(n2120), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][10]  ( .D(n2121), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[5][11]  ( .D(n2122), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[5][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[4]  ( .D(n2074), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[4]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][4]  ( .D(n2127), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][5]  ( .D(n2128), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][6]  ( .D(n2129), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][7]  ( .D(n2130), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][8]  ( .D(n2131), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][9]  ( .D(n2132), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][10]  ( .D(n2133), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[4][11]  ( .D(n2134), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[4][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[1]  ( .D(n2077), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[1]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][4]  ( .D(n2163), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][5]  ( .D(n2164), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][6]  ( .D(n2165), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][7]  ( .D(n2166), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][8]  ( .D(n2167), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][9]  ( .D(n2168), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][10]  ( .D(n2169), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[1][11]  ( .D(n2170), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[1][11] ) );
  DFFNSRX1TS \writeOutbuffer_reg[0]  ( .D(n2078), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(writeOutbuffer[0]) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][4]  ( .D(n2175), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][4] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][5]  ( .D(n2176), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][5] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][6]  ( .D(n2177), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][6] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][7]  ( .D(n2178), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][7] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][8]  ( .D(n2179), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][8] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][9]  ( .D(n2180), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][9] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][10]  ( .D(n2181), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][10] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[0][11]  ( .D(n2182), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[0][11] ) );
  DFFNSRX1TS \destinationAddressbuffer_reg[7][10]  ( .D(n2097), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(\destinationAddressbuffer[7][10] ) );
  DFFNSRX1TS writeOut_reg ( .D(n1968), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        writeOut) );
  DFFNSRX1TS \destinationAddressOut_reg[4]  ( .D(n1977), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[4]) );
  DFFNSRX1TS \destinationAddressOut_reg[5]  ( .D(n1978), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[5]) );
  DFFNSRX1TS \destinationAddressOut_reg[6]  ( .D(n1979), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[6]) );
  DFFNSRX1TS \destinationAddressOut_reg[7]  ( .D(n1980), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[7]) );
  DFFNSRX1TS \destinationAddressOut_reg[8]  ( .D(n1981), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[8]) );
  DFFNSRX1TS \destinationAddressOut_reg[9]  ( .D(n1982), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[9]) );
  DFFNSRX1TS \destinationAddressOut_reg[10]  ( .D(n1983), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[10]) );
  DFFNSRX1TS \destinationAddressOut_reg[11]  ( .D(n1984), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[11]) );
  DFFNSRX1TS readOut_reg ( .D(n1967), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        readOut) );
  DFFNSRX1TS \requesterAddressOut_reg[0]  ( .D(n1969), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[0]) );
  DFFNSRX1TS \requesterAddressOut_reg[1]  ( .D(n1970), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[1]) );
  DFFNSRX1TS \requesterAddressOut_reg[2]  ( .D(n1971), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[2]) );
  DFFNSRX1TS \requesterAddressOut_reg[3]  ( .D(n1972), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[3]) );
  DFFNSRX1TS \destinationAddressOut_reg[0]  ( .D(n1973), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[0]) );
  DFFNSRX1TS \destinationAddressOut_reg[1]  ( .D(n1974), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[1]) );
  DFFNSRX1TS \destinationAddressOut_reg[2]  ( .D(n1975), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[2]) );
  DFFNSRX1TS \destinationAddressOut_reg[3]  ( .D(n1976), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[3]) );
  DFFNSRX1TS \dataOut_reg[0]  ( .D(n1985), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[0]) );
  DFFNSRX1TS \dataOut_reg[1]  ( .D(n1986), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[1]) );
  DFFNSRX1TS \dataOut_reg[2]  ( .D(n1987), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[2]) );
  DFFNSRX1TS \dataOut_reg[3]  ( .D(n1988), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[3]) );
  DFFNSRX1TS \dataOut_reg[4]  ( .D(n1989), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[4]) );
  DFFNSRX1TS \dataOut_reg[5]  ( .D(n1990), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[5]) );
  DFFNSRX1TS \read_reg_reg[1]  ( .D(n1966), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1944), .QN(n1943) );
  DFFNSRX1TS \write_reg_reg[0]  ( .D(n1961), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1942), .QN(n1946) );
  DFFNSRX1TS \write_reg_reg[2]  ( .D(n1963), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1947), .QN(n1948) );
  DFFNSRX1TS \read_reg_reg[0]  ( .D(n1960), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1937), .QN(n1949) );
  DFFNSRX1TS \read_reg_reg[2]  ( .D(n1965), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1940), .QN(n1941) );
  DFFNSRX1TS empty_reg_reg ( .D(n1964), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        n1939), .QN(n1938) );
  DFFNSRX1TS \readOutbuffer_reg[7]  ( .D(n2079), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[7]), .QN(n1952) );
  DFFNSRX1TS \readOutbuffer_reg[4]  ( .D(n2082), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[4]), .QN(n1955) );
  DFFNSRX1TS \readOutbuffer_reg[6]  ( .D(n2080), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[6]), .QN(n1953) );
  DFFNSRX1TS \readOutbuffer_reg[5]  ( .D(n2081), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[5]), .QN(n1954) );
  DFFNSRX1TS \readOutbuffer_reg[1]  ( .D(n2085), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[1]), .QN(n1958) );
  DFFNSRX1TS \readOutbuffer_reg[2]  ( .D(n2084), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[2]), .QN(n1957) );
  DFFNSRX1TS \readOutbuffer_reg[0]  ( .D(n2086), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[0]), .QN(n1959) );
  DFFNSRX1TS \readOutbuffer_reg[3]  ( .D(n2083), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer[3]), .QN(n1956) );
  DFFNSRX1TS \write_reg_reg[1]  ( .D(n1962), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1945), .QN(n1950) );
  CMPR32X2TS U3 ( .A(n493), .B(n492), .C(n491), .CO(n486), .S(n501) );
  CLKBUFX2TS U4 ( .A(n13), .Y(n209) );
  CMPR32X2TS U5 ( .A(n471), .B(n502), .C(n15), .CO(n16), .S(n13) );
  ADDHXLTS U6 ( .A(n453), .B(n466), .CO(n15), .S(n14) );
  CMPR32X2TS U7 ( .A(n537), .B(n469), .C(n468), .CO(n460), .S(n474) );
  CMPR32X2TS U8 ( .A(n467), .B(n521), .C(n466), .CO(n470), .S(n483) );
  NOR2XLTS U9 ( .A(n465), .B(n511), .Y(n17) );
  CLKBUFX2TS U10 ( .A(n19), .Y(n71) );
  CLKBUFX2TS U11 ( .A(n17), .Y(n18) );
  NOR3XLTS U12 ( .A(n519), .B(selectBit_EAST), .C(n521), .Y(n514) );
  NOR2XLTS U13 ( .A(n1605), .B(n272), .Y(n276) );
  NOR2XLTS U14 ( .A(n1570), .B(n37), .Y(n41) );
  NOR2XLTS U15 ( .A(n116), .B(n381), .Y(n1619) );
  INVX2TS U16 ( .A(n1609), .Y(n1607) );
  INVX2TS U17 ( .A(n1598), .Y(n1596) );
  INVX2TS U18 ( .A(n1585), .Y(n1583) );
  INVX2TS U19 ( .A(n1574), .Y(n1572) );
  INVX2TS U20 ( .A(n1648), .Y(n1645) );
  INVX2TS U21 ( .A(n1588), .Y(n1586) );
  NOR2XLTS U22 ( .A(selectBit_NORTH), .B(n512), .Y(n545) );
  NOR2XLTS U23 ( .A(n1638), .B(n317), .Y(n318) );
  NOR2XLTS U24 ( .A(n1620), .B(n125), .Y(n126) );
  NOR2XLTS U25 ( .A(n310), .B(n1649), .Y(n311) );
  NOR2XLTS U26 ( .A(n310), .B(n1623), .Y(n122) );
  NOR3XLTS U27 ( .A(n1613), .B(n1607), .C(n271), .Y(n266) );
  NOR3XLTS U28 ( .A(n1601), .B(n1596), .C(n217), .Y(n213) );
  NOR2XLTS U29 ( .A(n448), .B(n1589), .Y(n76) );
  NOR2XLTS U30 ( .A(n1578), .B(n29), .Y(n32) );
  NOR2XLTS U31 ( .A(n1626), .B(n175), .Y(n176) );
  NOR2XLTS U32 ( .A(n25), .B(n124), .Y(n121) );
  OAI21XLTS U33 ( .A0(n497), .A1(n532), .B0(n494), .Y(n495) );
  AOI211XLTS U34 ( .A0(n497), .A1(n532), .B0(n496), .C0(n495), .Y(n498) );
  NOR2X1TS U35 ( .A(n1595), .B(n219), .Y(n227) );
  NOR2X1TS U36 ( .A(n1628), .B(n175), .Y(n179) );
  NOR2X1TS U37 ( .A(n1640), .B(n317), .Y(n339) );
  NAND2BXLTS U38 ( .AN(n315), .B(n314), .Y(n317) );
  NAND2BXLTS U39 ( .AN(n174), .B(n173), .Y(n175) );
  NAND2BXLTS U40 ( .AN(n393), .B(n392), .Y(n394) );
  NAND2BXLTS U41 ( .AN(n271), .B(n270), .Y(n272) );
  NAND2BXLTS U42 ( .AN(n79), .B(n78), .Y(n80) );
  XOR2XLTS U43 ( .A(n531), .B(n500), .Y(n496) );
  OAI21X1TS U44 ( .A0(n27), .A1(n24), .B0(n26), .Y(n115) );
  NAND3X1TS U45 ( .A(n73), .B(n28), .C(n210), .Y(n1570) );
  OAI21X1TS U46 ( .A0(selectBit_SOUTH), .A1(n20), .B0(n71), .Y(n261) );
  NOR2X1TS U47 ( .A(n210), .B(n70), .Y(n306) );
  NAND3X1TS U48 ( .A(n23), .B(n210), .C(n263), .Y(n1592) );
  INVX1TS U49 ( .A(n1634), .Y(n1632) );
  NOR2X1TS U50 ( .A(n267), .B(n1614), .Y(n268) );
  INVX1TS U51 ( .A(n1613), .Y(n1610) );
  INVX1TS U52 ( .A(n1660), .Y(n1658) );
  AND2X2TS U53 ( .A(n530), .B(n1951), .Y(n211) );
  CLKBUFX2TS U54 ( .A(readIn_EAST), .Y(n1569) );
  INVX1TS U55 ( .A(n1948), .Y(n487) );
  NAND2BX1TS U56 ( .AN(n114), .B(n467), .Y(n379) );
  OR3X1TS U57 ( .A(n1648), .B(n1641), .C(n315), .Y(n1) );
  INVX2TS U58 ( .A(n1), .Y(n309) );
  NOR2X1TS U59 ( .A(n8), .B(n70), .Y(n27) );
  NAND2BX1TS U60 ( .AN(n115), .B(selectBit_EAST), .Y(n381) );
  NOR3X1TS U61 ( .A(n307), .B(n306), .C(n262), .Y(n1598) );
  NOR2X1TS U62 ( .A(n116), .B(n262), .Y(n1574) );
  NOR2XLTS U63 ( .A(n1601), .B(n1598), .Y(n216) );
  NOR3BXLTS U64 ( .AN(readReady), .B(n519), .C(n518), .Y(n544) );
  NAND2BXLTS U65 ( .AN(n125), .B(n120), .Y(n124) );
  NAND2X1TS U66 ( .A(n123), .B(n1623), .Y(n125) );
  OR2X1TS U67 ( .A(n269), .B(n937), .Y(n1420) );
  OR2X1TS U68 ( .A(n215), .B(n920), .Y(n1451) );
  OR2X1TS U69 ( .A(n172), .B(n989), .Y(n1356) );
  OR2X1TS U70 ( .A(n123), .B(n964), .Y(n1389) );
  OR2X1TS U71 ( .A(n77), .B(n902), .Y(n1485) );
  OR2X1TS U72 ( .A(n33), .B(n1663), .Y(n1538) );
  CLKAND2X2TS U73 ( .A(n485), .B(n484), .Y(n491) );
  NAND4XLTS U74 ( .A(n463), .B(n453), .C(n516), .D(n449), .Y(n1623) );
  INVX2TS U75 ( .A(n1622), .Y(n1620) );
  CLKBUFX2TS U76 ( .A(n1389), .Y(n1624) );
  NOR3XLTS U77 ( .A(n13), .B(n113), .C(n379), .Y(n1660) );
  INVX2TS U78 ( .A(n1657), .Y(n1654) );
  NOR3XLTS U79 ( .A(n14), .B(n169), .C(n379), .Y(n1634) );
  INVX2TS U80 ( .A(n1631), .Y(n1629) );
  CLKBUFX2TS U81 ( .A(n1356), .Y(n1636) );
  NAND4XLTS U82 ( .A(n454), .B(n516), .C(n451), .D(n387), .Y(n1649) );
  NOR3XLTS U83 ( .A(n13), .B(n69), .C(n379), .Y(n1648) );
  INVX2TS U84 ( .A(n1644), .Y(n1641) );
  NOR3X1TS U85 ( .A(n209), .B(n69), .C(n260), .Y(n1601) );
  CLKBUFX2TS U86 ( .A(n1451), .Y(n1603) );
  NAND4XLTS U87 ( .A(n73), .B(n459), .C(n517), .D(n388), .Y(n1589) );
  NOR3XLTS U88 ( .A(n14), .B(n169), .C(n260), .Y(n1588) );
  CLKBUFX2TS U89 ( .A(n1485), .Y(n1590) );
  NAND4XLTS U90 ( .A(n265), .B(n516), .C(n388), .D(n384), .Y(n1614) );
  NOR3XLTS U91 ( .A(n209), .B(n14), .C(n260), .Y(n1613) );
  CLKBUFX2TS U92 ( .A(n1420), .Y(n1615) );
  NAND4XLTS U93 ( .A(n1942), .B(n502), .C(n487), .D(n521), .Y(n1578) );
  CLKBUFX2TS U94 ( .A(n1538), .Y(n1579) );
  NAND3XLTS U95 ( .A(n545), .B(n1939), .C(n544), .Y(n567) );
  CLKAND2X2TS U96 ( .A(n530), .B(n528), .Y(n558) );
  NOR3XLTS U97 ( .A(n1634), .B(n1629), .C(n174), .Y(n171) );
  INVX2TS U98 ( .A(selectBit_NORTH), .Y(n511) );
  NOR2XLTS U99 ( .A(n1613), .B(n1609), .Y(n270) );
  NOR2XLTS U100 ( .A(n1588), .B(n1585), .Y(n78) );
  NOR2XLTS U101 ( .A(n1577), .B(n1574), .Y(n35) );
  NOR2XLTS U102 ( .A(n1660), .B(n1657), .Y(n392) );
  AO21X1TS U103 ( .A0(n465), .A1(n511), .B0(n18), .Y(n20) );
  NAND3XLTS U104 ( .A(selectBit_NORTH), .B(n514), .C(n513), .Y(n525) );
  NAND3XLTS U105 ( .A(n512), .B(n514), .C(n511), .Y(n524) );
  NOR2XLTS U106 ( .A(n1648), .B(n1644), .Y(n314) );
  NOR2XLTS U107 ( .A(n1622), .B(n1619), .Y(n120) );
  NAND2BXLTS U108 ( .AN(n217), .B(n216), .Y(n219) );
  NAND3XLTS U109 ( .A(n18), .B(n459), .C(n387), .Y(n212) );
  NOR2XLTS U110 ( .A(n1634), .B(n1631), .Y(n173) );
  NAND2BXLTS U111 ( .AN(n36), .B(n35), .Y(n37) );
  XOR2XLTS U112 ( .A(n460), .B(n462), .Y(n480) );
  OAI21XLTS U113 ( .A0(n463), .A1(n1943), .B0(n462), .Y(n464) );
  INVX2TS U114 ( .A(n263), .Y(n383) );
  XOR2X1TS U115 ( .A(n487), .B(n16), .Y(n114) );
  NOR2XLTS U116 ( .A(n75), .B(reset), .Y(n505) );
  NOR3X1TS U117 ( .A(n169), .B(n69), .C(n379), .Y(n1622) );
  INVX2TS U118 ( .A(n1619), .Y(n1617) );
  NAND4XLTS U119 ( .A(n517), .B(n388), .C(n387), .D(n449), .Y(n1661) );
  NOR3XLTS U120 ( .A(n28), .B(n383), .C(n71), .Y(n1653) );
  INVX2TS U121 ( .A(n1653), .Y(n1651) );
  NOR3BXLTS U122 ( .AN(n382), .B(n381), .C(n380), .Y(n1657) );
  NAND4XLTS U123 ( .A(n492), .B(n517), .C(n388), .D(n451), .Y(n1635) );
  NOR3XLTS U124 ( .A(n28), .B(n71), .C(n263), .Y(n1628) );
  INVX2TS U125 ( .A(n1628), .Y(n1626) );
  NOR3XLTS U126 ( .A(n28), .B(n383), .C(n8), .Y(n1640) );
  INVX2TS U127 ( .A(n1640), .Y(n1638) );
  NOR3XLTS U128 ( .A(n307), .B(n306), .C(n381), .Y(n1644) );
  NAND4XLTS U129 ( .A(n454), .B(n459), .C(readReady), .D(n384), .Y(n1602) );
  INVX2TS U130 ( .A(n1592), .Y(n1595) );
  INVX2TS U131 ( .A(n1601), .Y(n1599) );
  INVX2TS U132 ( .A(n1582), .Y(n1581) );
  NOR3XLTS U133 ( .A(n383), .B(n19), .C(n22), .Y(n1606) );
  INVX2TS U134 ( .A(n1606), .Y(n1605) );
  NOR3BXLTS U135 ( .AN(n382), .B(n262), .C(n261), .Y(n1609) );
  NAND4XLTS U136 ( .A(n209), .B(n113), .C(n114), .D(n467), .Y(n1575) );
  INVX2TS U137 ( .A(n1570), .Y(n1571) );
  INVX2TS U138 ( .A(destinationAddressIn_SOUTH[11]), .Y(n138) );
  INVX2TS U139 ( .A(destinationAddressIn_SOUTH[10]), .Y(n142) );
  INVX2TS U140 ( .A(destinationAddressIn_SOUTH[9]), .Y(n133) );
  INVX2TS U141 ( .A(destinationAddressIn_SOUTH[8]), .Y(n129) );
  CLKAND2X2TS U142 ( .A(n485), .B(n483), .Y(n490) );
  AO22XLTS U143 ( .A0(n1947), .A1(n505), .B0(n504), .B1(n503), .Y(n1963) );
  AO22XLTS U144 ( .A0(n1942), .A1(n505), .B0(n504), .B1(n500), .Y(n1961) );
  AO22XLTS U145 ( .A0(n502), .A1(n505), .B0(n504), .B1(n501), .Y(n1962) );
  OAI21XLTS U146 ( .A0(n75), .A1(n456), .B0(n499), .Y(n1964) );
  NAND4XLTS U147 ( .A(n880), .B(n879), .C(n878), .D(n877), .Y(n1990) );
  NAND4XLTS U148 ( .A(n856), .B(n855), .C(n854), .D(n853), .Y(n1989) );
  NAND4XLTS U149 ( .A(n844), .B(n843), .C(n842), .D(n841), .Y(n1988) );
  NAND4XLTS U150 ( .A(n832), .B(n831), .C(n830), .D(n829), .Y(n1987) );
  NAND4XLTS U151 ( .A(n813), .B(n812), .C(n811), .D(n810), .Y(n1986) );
  NAND4XLTS U152 ( .A(n793), .B(n792), .C(n791), .D(n790), .Y(n1985) );
  NAND4XLTS U153 ( .A(n664), .B(n663), .C(n662), .D(n661), .Y(n1976) );
  NAND4XLTS U154 ( .A(n652), .B(n651), .C(n650), .D(n649), .Y(n1975) );
  NAND4XLTS U155 ( .A(n632), .B(n631), .C(n630), .D(n629), .Y(n1974) );
  NAND4XLTS U156 ( .A(n617), .B(n616), .C(n615), .D(n614), .Y(n1973) );
  NAND4XLTS U157 ( .A(n606), .B(n605), .C(n604), .D(n661), .Y(n1972) );
  NAND4XLTS U158 ( .A(n595), .B(n594), .C(n593), .D(n649), .Y(n1971) );
  NAND4XLTS U159 ( .A(n587), .B(n586), .C(n585), .D(n629), .Y(n1970) );
  NAND4XLTS U160 ( .A(n570), .B(n569), .C(n568), .D(n614), .Y(n1969) );
  NAND4XLTS U161 ( .A(n548), .B(n547), .C(n546), .D(n567), .Y(n1967) );
  NAND3XLTS U162 ( .A(n783), .B(n782), .C(n781), .Y(n1984) );
  NAND3XLTS U163 ( .A(n769), .B(n768), .C(n767), .Y(n1983) );
  NAND3XLTS U164 ( .A(n754), .B(n753), .C(n752), .Y(n1982) );
  NAND3XLTS U165 ( .A(n736), .B(n735), .C(n734), .Y(n1981) );
  NAND3XLTS U166 ( .A(n722), .B(n721), .C(n720), .Y(n1980) );
  NAND3XLTS U167 ( .A(n711), .B(n710), .C(n709), .Y(n1979) );
  NAND3XLTS U168 ( .A(n696), .B(n695), .C(n694), .Y(n1978) );
  NAND3XLTS U169 ( .A(n675), .B(n674), .C(n673), .Y(n1977) );
  NAND3XLTS U170 ( .A(n561), .B(n560), .C(n559), .Y(n1968) );
  NAND3XLTS U171 ( .A(n1345), .B(n1344), .C(n1343), .Y(n2034) );
  NAND3XLTS U172 ( .A(n1339), .B(n1338), .C(n1337), .Y(n2033) );
  NAND3XLTS U173 ( .A(n1110), .B(n1109), .C(n1108), .Y(n2032) );
  NAND3XLTS U174 ( .A(n1104), .B(n1103), .C(n1102), .Y(n2031) );
  NAND3XLTS U175 ( .A(n1096), .B(n1095), .C(n1094), .Y(n2030) );
  NAND3XLTS U176 ( .A(n1090), .B(n1089), .C(n1088), .Y(n2029) );
  NAND3XLTS U177 ( .A(n1813), .B(n1812), .C(n1811), .Y(n2138) );
  NAND3XLTS U178 ( .A(n1804), .B(n1803), .C(n1802), .Y(n2137) );
  NAND3XLTS U179 ( .A(n1798), .B(n1797), .C(n1796), .Y(n2136) );
  NAND3XLTS U180 ( .A(n1790), .B(n1789), .C(n1788), .Y(n2135) );
  NAND3XLTS U181 ( .A(n985), .B(n984), .C(n983), .Y(n2010) );
  NAND3XLTS U182 ( .A(n979), .B(n978), .C(n977), .Y(n2009) );
  NAND3XLTS U183 ( .A(n971), .B(n970), .C(n969), .Y(n2008) );
  NAND3XLTS U184 ( .A(n962), .B(n961), .C(n960), .Y(n2007) );
  NAND3XLTS U185 ( .A(n1439), .B(n1438), .C(n1437), .Y(n2052) );
  NAND3XLTS U186 ( .A(n1433), .B(n1432), .C(n1431), .Y(n2051) );
  NAND3XLTS U187 ( .A(n1429), .B(n1428), .C(n1427), .Y(n2050) );
  NAND3XLTS U188 ( .A(n1425), .B(n1424), .C(n1423), .Y(n2049) );
  NAND3XLTS U189 ( .A(n1418), .B(n1417), .C(n1416), .Y(n2048) );
  NAND3XLTS U190 ( .A(n1411), .B(n1410), .C(n1409), .Y(n2047) );
  NAND3XLTS U191 ( .A(n1467), .B(n1466), .C(n1465), .Y(n2058) );
  NAND3XLTS U192 ( .A(n1463), .B(n1462), .C(n1461), .Y(n2057) );
  NAND3XLTS U193 ( .A(n1459), .B(n1458), .C(n1457), .Y(n2056) );
  NAND3XLTS U194 ( .A(n1455), .B(n1454), .C(n1453), .Y(n2055) );
  NAND3XLTS U195 ( .A(n1450), .B(n1449), .C(n1448), .Y(n2054) );
  NAND3XLTS U196 ( .A(n1445), .B(n1444), .C(n1443), .Y(n2053) );
  NAND3XLTS U197 ( .A(n1721), .B(n1720), .C(n1719), .Y(n2102) );
  NAND3XLTS U198 ( .A(n1713), .B(n1712), .C(n1711), .Y(n2101) );
  NAND3XLTS U199 ( .A(n1706), .B(n1705), .C(n1704), .Y(n2100) );
  NAND3XLTS U200 ( .A(n1697), .B(n1696), .C(n1695), .Y(n2099) );
  NAND3XLTS U201 ( .A(n915), .B(n914), .C(n913), .Y(n1998) );
  NAND3XLTS U202 ( .A(n911), .B(n910), .C(n909), .Y(n1997) );
  NAND3XLTS U203 ( .A(n908), .B(n907), .C(n906), .Y(n1996) );
  NAND3XLTS U204 ( .A(n901), .B(n900), .C(n899), .Y(n1995) );
  NAND3XLTS U205 ( .A(n1692), .B(n1691), .C(n1690), .Y(n2090) );
  NAND3XLTS U206 ( .A(n1683), .B(n1682), .C(n1681), .Y(n2089) );
  NAND3XLTS U207 ( .A(n1676), .B(n1675), .C(n1674), .Y(n2088) );
  NAND3XLTS U208 ( .A(n1668), .B(n1667), .C(n1666), .Y(n2087) );
  NAND3XLTS U209 ( .A(n898), .B(n897), .C(n896), .Y(n1994) );
  NAND3XLTS U210 ( .A(n893), .B(n892), .C(n891), .Y(n1993) );
  NAND3XLTS U211 ( .A(n888), .B(n887), .C(n886), .Y(n1992) );
  NAND3XLTS U212 ( .A(n885), .B(n884), .C(n883), .Y(n1991) );
  NAND3XLTS U213 ( .A(n1921), .B(n1920), .C(n1919), .Y(n2174) );
  NAND3XLTS U214 ( .A(n1912), .B(n1911), .C(n1910), .Y(n2173) );
  NAND3XLTS U215 ( .A(n1901), .B(n1900), .C(n1899), .Y(n2172) );
  NAND3XLTS U216 ( .A(n1890), .B(n1889), .C(n1888), .Y(n2171) );
  NAND3XLTS U217 ( .A(n1058), .B(n1057), .C(n1056), .Y(n2022) );
  NAND3XLTS U218 ( .A(n1051), .B(n1050), .C(n1049), .Y(n2021) );
  NAND3XLTS U219 ( .A(n1046), .B(n1045), .C(n1044), .Y(n2020) );
  NAND3XLTS U220 ( .A(n1040), .B(n1039), .C(n1038), .Y(n2019) );
  NAND3XLTS U221 ( .A(n1883), .B(n1882), .C(n1881), .Y(n2162) );
  NAND3XLTS U222 ( .A(n1873), .B(n1872), .C(n1871), .Y(n2161) );
  NAND3XLTS U223 ( .A(n1860), .B(n1859), .C(n1858), .Y(n2160) );
  NAND3XLTS U224 ( .A(n1849), .B(n1848), .C(n1847), .Y(n2159) );
  NAND3XLTS U225 ( .A(n1033), .B(n1032), .C(n1031), .Y(n2018) );
  NAND3XLTS U226 ( .A(n1024), .B(n1023), .C(n1022), .Y(n2017) );
  NAND3XLTS U227 ( .A(n1016), .B(n1015), .C(n1014), .Y(n2016) );
  NAND3XLTS U228 ( .A(n1009), .B(n1008), .C(n1007), .Y(n2015) );
  NAND3XLTS U229 ( .A(n1378), .B(n1377), .C(n1376), .Y(n2040) );
  NAND3XLTS U230 ( .A(n1373), .B(n1372), .C(n1371), .Y(n2039) );
  NAND3XLTS U231 ( .A(n1369), .B(n1368), .C(n1367), .Y(n2038) );
  NAND3XLTS U232 ( .A(n1364), .B(n1363), .C(n1362), .Y(n2037) );
  NAND3XLTS U233 ( .A(n1355), .B(n1354), .C(n1353), .Y(n2036) );
  NAND3XLTS U234 ( .A(n1349), .B(n1348), .C(n1347), .Y(n2035) );
  NAND3XLTS U235 ( .A(n1406), .B(n1405), .C(n1404), .Y(n2046) );
  NAND3XLTS U236 ( .A(n1401), .B(n1400), .C(n1399), .Y(n2045) );
  NAND3XLTS U237 ( .A(n1395), .B(n1394), .C(n1393), .Y(n2044) );
  NAND3XLTS U238 ( .A(n1392), .B(n1391), .C(n1390), .Y(n2043) );
  NAND3XLTS U239 ( .A(n1387), .B(n1386), .C(n1385), .Y(n2042) );
  NAND3XLTS U240 ( .A(n1382), .B(n1381), .C(n1380), .Y(n2041) );
  NAND3XLTS U241 ( .A(n1784), .B(n1783), .C(n1782), .Y(n2126) );
  NAND3XLTS U242 ( .A(n1777), .B(n1776), .C(n1775), .Y(n2125) );
  NAND3XLTS U243 ( .A(n1769), .B(n1768), .C(n1767), .Y(n2124) );
  NAND3XLTS U244 ( .A(n1760), .B(n1759), .C(n1758), .Y(n2123) );
  NAND3XLTS U245 ( .A(n955), .B(n954), .C(n953), .Y(n2006) );
  NAND3XLTS U246 ( .A(n949), .B(n948), .C(n947), .Y(n2005) );
  NAND3XLTS U247 ( .A(n944), .B(n943), .C(n942), .Y(n2004) );
  NAND3XLTS U248 ( .A(n936), .B(n935), .C(n934), .Y(n2003) );
  NAND3XLTS U249 ( .A(n1755), .B(n1754), .C(n1753), .Y(n2114) );
  NAND3XLTS U250 ( .A(n1748), .B(n1747), .C(n1746), .Y(n2113) );
  NAND3XLTS U251 ( .A(n1737), .B(n1736), .C(n1735), .Y(n2112) );
  NAND3XLTS U252 ( .A(n1727), .B(n1726), .C(n1725), .Y(n2111) );
  NAND3XLTS U253 ( .A(n931), .B(n930), .C(n929), .Y(n2002) );
  NAND3XLTS U254 ( .A(n926), .B(n925), .C(n924), .Y(n2001) );
  NAND3XLTS U255 ( .A(n923), .B(n922), .C(n921), .Y(n2000) );
  NAND3XLTS U256 ( .A(n919), .B(n918), .C(n917), .Y(n1999) );
  NAND3XLTS U257 ( .A(n1518), .B(n1517), .C(n1516), .Y(n2064) );
  NAND3XLTS U258 ( .A(n1509), .B(n1508), .C(n1507), .Y(n2063) );
  NAND3XLTS U259 ( .A(n1502), .B(n1501), .C(n1500), .Y(n2062) );
  NAND3XLTS U260 ( .A(n1494), .B(n1493), .C(n1492), .Y(n2061) );
  NAND3XLTS U261 ( .A(n1483), .B(n1482), .C(n1481), .Y(n2060) );
  NAND3XLTS U262 ( .A(n1475), .B(n1474), .C(n1473), .Y(n2059) );
  NAND3XLTS U263 ( .A(n1568), .B(n1567), .C(n1566), .Y(n2070) );
  NAND3XLTS U264 ( .A(n1560), .B(n1559), .C(n1558), .Y(n2069) );
  NAND3XLTS U265 ( .A(n1552), .B(n1551), .C(n1550), .Y(n2068) );
  NAND3XLTS U266 ( .A(n1545), .B(n1544), .C(n1543), .Y(n2067) );
  NAND3XLTS U267 ( .A(n1537), .B(n1536), .C(n1535), .Y(n2066) );
  NAND3XLTS U268 ( .A(n1527), .B(n1526), .C(n1525), .Y(n2065) );
  NAND3XLTS U269 ( .A(n1085), .B(n1084), .C(n1083), .Y(n2028) );
  NAND3XLTS U270 ( .A(n1080), .B(n1079), .C(n1078), .Y(n2027) );
  NAND3XLTS U271 ( .A(n1076), .B(n1075), .C(n1074), .Y(n2026) );
  NAND3XLTS U272 ( .A(n1073), .B(n1072), .C(n1071), .Y(n2025) );
  NAND3XLTS U273 ( .A(n1066), .B(n1065), .C(n1064), .Y(n2024) );
  NAND3XLTS U274 ( .A(n1062), .B(n1061), .C(n1060), .Y(n2023) );
  NAND3XLTS U275 ( .A(n1840), .B(n1839), .C(n1838), .Y(n2150) );
  NAND3XLTS U276 ( .A(n1833), .B(n1832), .C(n1831), .Y(n2149) );
  NAND3XLTS U277 ( .A(n1824), .B(n1823), .C(n1822), .Y(n2148) );
  NAND3XLTS U278 ( .A(n1817), .B(n1816), .C(n1815), .Y(n2147) );
  NAND3XLTS U279 ( .A(n1002), .B(n1001), .C(n1000), .Y(n2014) );
  NAND3XLTS U280 ( .A(n997), .B(n996), .C(n995), .Y(n2013) );
  NAND3XLTS U281 ( .A(n992), .B(n991), .C(n990), .Y(n2012) );
  NAND3XLTS U282 ( .A(n988), .B(n987), .C(n986), .Y(n2011) );
  OR2X1TS U283 ( .A(n312), .B(n1010), .Y(n350) );
  NAND2X1TS U284 ( .A(n27), .B(n24), .Y(n25) );
  OR2X1TS U285 ( .A(n1651), .B(n394), .Y(n2) );
  OR2X1TS U286 ( .A(n1582), .B(n80), .Y(n3) );
  OR2X1TS U287 ( .A(n1581), .B(n80), .Y(n4) );
  OR2X1TS U288 ( .A(n1653), .B(n394), .Y(n5) );
  OR2X1TS U289 ( .A(n1606), .B(n272), .Y(n6) );
  OA21XLTS U290 ( .A0(n18), .A1(n73), .B0(n21), .Y(n7) );
  OR2X1TS U291 ( .A(n20), .B(n513), .Y(n8) );
  OR2X1TS U292 ( .A(n448), .B(n1635), .Y(n9) );
  OR2X1TS U293 ( .A(n390), .B(n1041), .Y(n425) );
  NOR3XLTS U294 ( .A(n1660), .B(n1654), .C(n393), .Y(n389) );
  NOR3XLTS U295 ( .A(n1577), .B(n1572), .C(n36), .Y(n31) );
  NOR3XLTS U296 ( .A(n1588), .B(n1583), .C(n79), .Y(n74) );
  OR2X1TS U297 ( .A(n457), .B(n1602), .Y(n10) );
  OR2X1TS U298 ( .A(n448), .B(n1661), .Y(n11) );
  NOR2XLTS U299 ( .A(n851), .B(n525), .Y(n698) );
  NOR2XLTS U300 ( .A(n851), .B(n524), .Y(n550) );
  CLKBUFX2TS U301 ( .A(n1943), .Y(n12) );
  INVX2TS U317 ( .A(n1950), .Y(n502) );
  INVX2TS U318 ( .A(n1946), .Y(n453) );
  ADDFHX1TS U319 ( .A(selectBit_SOUTH), .B(selectBit_NORTH), .CI(
        selectBit_EAST), .CO(n471), .S(n466) );
  INVX2TS U320 ( .A(n14), .Y(n69) );
  INVX2TS U321 ( .A(n69), .Y(n113) );
  INVX2TS U322 ( .A(selectBit_WEST), .Y(n461) );
  INVX2TS U323 ( .A(n1575), .Y(n1577) );
  INVX2TS U324 ( .A(n1942), .Y(n465) );
  INVX2TS U325 ( .A(selectBit_SOUTH), .Y(n513) );
  INVX2TS U326 ( .A(n8), .Y(n210) );
  INVX2TS U327 ( .A(n1950), .Y(n73) );
  INVX2TS U328 ( .A(n1950), .Y(n492) );
  NAND2X1TS U329 ( .A(n17), .B(n492), .Y(n21) );
  INVX2TS U330 ( .A(n7), .Y(n70) );
  NAND2X1TS U331 ( .A(selectBit_SOUTH), .B(n20), .Y(n19) );
  NAND2X1TS U332 ( .A(n306), .B(n261), .Y(n116) );
  INVX2TS U333 ( .A(selectBit_EAST), .Y(n520) );
  INVX2TS U334 ( .A(n520), .Y(n518) );
  INVX2TS U335 ( .A(n1948), .Y(n265) );
  INVX2TS U336 ( .A(n21), .Y(n117) );
  INVX2TS U337 ( .A(n1947), .Y(n458) );
  AOI22X1TS U338 ( .A0(n265), .A1(n21), .B0(n117), .B1(n458), .Y(n22) );
  INVX2TS U339 ( .A(n22), .Y(n23) );
  INVX2TS U340 ( .A(n23), .Y(n24) );
  INVX2TS U341 ( .A(n25), .Y(n112) );
  INVX2TS U342 ( .A(n112), .Y(n26) );
  NAND2X1TS U343 ( .A(n518), .B(n115), .Y(n262) );
  NAND2X1TS U344 ( .A(n265), .B(n117), .Y(n30) );
  INVX2TS U345 ( .A(n24), .Y(n28) );
  INVX2TS U346 ( .A(n513), .Y(n512) );
  INVX2TS U347 ( .A(n461), .Y(n519) );
  INVX2TS U348 ( .A(readReady), .Y(n119) );
  INVX2TS U349 ( .A(n119), .Y(n521) );
  NAND2X1TS U350 ( .A(n545), .B(n514), .Y(n530) );
  INVX2TS U351 ( .A(n211), .Y(n310) );
  INVX2TS U352 ( .A(n310), .Y(n75) );
  INVX2TS U353 ( .A(n75), .Y(n29) );
  AOI31XLTS U354 ( .A0(n35), .A1(n30), .A2(n1570), .B0(n29), .Y(n33) );
  NAND2X1TS U355 ( .A(n33), .B(n1578), .Y(n36) );
  INVX2TS U356 ( .A(n31), .Y(n1530) );
  INVX2TS U357 ( .A(n1530), .Y(n889) );
  CLKBUFX2TS U358 ( .A(n889), .Y(n44) );
  INVX2TS U359 ( .A(n44), .Y(n60) );
  INVX2TS U360 ( .A(destinationAddressIn_EAST[11]), .Y(n222) );
  INVX2TS U361 ( .A(n32), .Y(n894) );
  INVX2TS U362 ( .A(n894), .Y(n1663) );
  INVX2TS U363 ( .A(n1538), .Y(n48) );
  OR2X1TS U364 ( .A(n1575), .B(n36), .Y(n47) );
  INVX2TS U365 ( .A(n47), .Y(n34) );
  INVX2TS U366 ( .A(n34), .Y(n881) );
  INVX2TS U367 ( .A(n881), .Y(n63) );
  CLKBUFX2TS U368 ( .A(destinationAddressIn_WEST[11]), .Y(n391) );
  CLKBUFX2TS U369 ( .A(n391), .Y(n770) );
  AOI22X1TS U370 ( .A0(n48), .A1(\destinationAddressbuffer[7][11] ), .B0(n63), 
        .B1(n770), .Y(n40) );
  INVX2TS U371 ( .A(n41), .Y(n1532) );
  INVX2TS U372 ( .A(n1532), .Y(n895) );
  INVX2TS U373 ( .A(n138), .Y(n773) );
  OR2X1TS U374 ( .A(n1571), .B(n37), .Y(n54) );
  INVX2TS U375 ( .A(n54), .Y(n38) );
  CLKBUFX2TS U376 ( .A(destinationAddressIn_NORTH[11]), .Y(n774) );
  CLKBUFX2TS U377 ( .A(n774), .Y(n326) );
  AOI22X1TS U378 ( .A0(n895), .A1(n773), .B0(n38), .B1(n326), .Y(n39) );
  OAI211XLTS U379 ( .A0(n60), .A1(n222), .B0(n40), .C0(n39), .Y(n2098) );
  INVX2TS U380 ( .A(destinationAddressIn_EAST[10]), .Y(n214) );
  INVX2TS U381 ( .A(n47), .Y(n1521) );
  CLKBUFX2TS U382 ( .A(destinationAddressIn_WEST[10]), .Y(n406) );
  CLKBUFX2TS U383 ( .A(n406), .Y(n755) );
  AOI22X1TS U384 ( .A0(n48), .A1(\destinationAddressbuffer[7][10] ), .B0(n1521), .B1(n755), .Y(n43) );
  INVX2TS U385 ( .A(n41), .Y(n57) );
  INVX2TS U386 ( .A(n142), .Y(n758) );
  INVX2TS U387 ( .A(n54), .Y(n1556) );
  CLKBUFX2TS U388 ( .A(destinationAddressIn_NORTH[10]), .Y(n759) );
  CLKBUFX2TS U389 ( .A(n759), .Y(n321) );
  AOI22X1TS U390 ( .A0(n49), .A1(n758), .B0(n1556), .B1(n321), .Y(n42) );
  OAI211XLTS U391 ( .A0(n60), .A1(n214), .B0(n43), .C0(n42), .Y(n2097) );
  INVX2TS U392 ( .A(n44), .Y(n68) );
  INVX2TS U393 ( .A(destinationAddressIn_EAST[8]), .Y(n230) );
  INVX2TS U394 ( .A(n47), .Y(n1664) );
  CLKBUFX2TS U395 ( .A(destinationAddressIn_WEST[8]), .Y(n400) );
  CLKBUFX2TS U396 ( .A(n400), .Y(n723) );
  AOI22X1TS U397 ( .A0(n48), .A1(\destinationAddressbuffer[7][8] ), .B0(n1664), 
        .B1(n723), .Y(n46) );
  INVX2TS U398 ( .A(n129), .Y(n724) );
  INVX2TS U399 ( .A(n54), .Y(n1523) );
  CLKBUFX2TS U400 ( .A(destinationAddressIn_NORTH[8]), .Y(n725) );
  CLKBUFX2TS U401 ( .A(n725), .Y(n333) );
  AOI22X1TS U402 ( .A0(n895), .A1(n724), .B0(n1523), .B1(n333), .Y(n45) );
  OAI211XLTS U403 ( .A0(n68), .A1(n230), .B0(n46), .C0(n45), .Y(n2095) );
  INVX2TS U404 ( .A(destinationAddressIn_EAST[9]), .Y(n226) );
  INVX2TS U405 ( .A(n47), .Y(n1672) );
  CLKBUFX2TS U406 ( .A(destinationAddressIn_WEST[9]), .Y(n412) );
  CLKBUFX2TS U407 ( .A(n412), .Y(n738) );
  AOI22X1TS U408 ( .A0(n48), .A1(\destinationAddressbuffer[7][9] ), .B0(n34), 
        .B1(n738), .Y(n51) );
  INVX2TS U409 ( .A(n57), .Y(n49) );
  INVX2TS U410 ( .A(n57), .Y(n65) );
  INVX2TS U411 ( .A(n133), .Y(n739) );
  INVX2TS U412 ( .A(n1523), .Y(n882) );
  INVX2TS U413 ( .A(n882), .Y(n890) );
  CLKBUFX2TS U414 ( .A(destinationAddressIn_NORTH[9]), .Y(n741) );
  CLKBUFX2TS U415 ( .A(n741), .Y(n342) );
  AOI22X1TS U416 ( .A0(n65), .A1(n739), .B0(n890), .B1(n342), .Y(n50) );
  OAI211XLTS U417 ( .A0(n60), .A1(n226), .B0(n51), .C0(n50), .Y(n2096) );
  INVX2TS U418 ( .A(writeIn_EAST), .Y(n237) );
  INVX2TS U419 ( .A(n1579), .Y(n1684) );
  CLKBUFX2TS U420 ( .A(writeIn_WEST), .Y(n420) );
  CLKBUFX2TS U421 ( .A(n420), .Y(n549) );
  AOI22X1TS U422 ( .A0(n1684), .A1(writeOutbuffer[7]), .B0(n63), .B1(n549), 
        .Y(n53) );
  INVX2TS U423 ( .A(n57), .Y(n1680) );
  INVX2TS U424 ( .A(writeIn_SOUTH), .Y(n146) );
  INVX2TS U425 ( .A(n146), .Y(n551) );
  CLKBUFX2TS U426 ( .A(writeIn_NORTH), .Y(n552) );
  CLKBUFX2TS U427 ( .A(n552), .Y(n347) );
  AOI22X1TS U428 ( .A0(n1680), .A1(n551), .B0(n1556), .B1(n347), .Y(n52) );
  OAI211XLTS U429 ( .A0(n68), .A1(n237), .B0(n53), .C0(n52), .Y(n2071) );
  INVX2TS U430 ( .A(destinationAddressIn_EAST[7]), .Y(n255) );
  INVX2TS U431 ( .A(n1538), .Y(n64) );
  AOI22X1TS U432 ( .A0(n64), .A1(\destinationAddressbuffer[7][7] ), .B0(n1664), 
        .B1(destinationAddressIn_WEST[7]), .Y(n56) );
  INVX2TS U433 ( .A(destinationAddressIn_SOUTH[7]), .Y(n161) );
  INVX2TS U434 ( .A(n161), .Y(n713) );
  INVX2TS U435 ( .A(n54), .Y(n1673) );
  AOI22X1TS U436 ( .A0(n1680), .A1(n713), .B0(n1673), .B1(
        destinationAddressIn_NORTH[7]), .Y(n55) );
  OAI211XLTS U437 ( .A0(n68), .A1(n255), .B0(n56), .C0(n55), .Y(n2094) );
  INVX2TS U438 ( .A(destinationAddressIn_EAST[6]), .Y(n240) );
  AOI22X1TS U439 ( .A0(n64), .A1(\destinationAddressbuffer[7][6] ), .B0(n1672), 
        .B1(destinationAddressIn_WEST[6]), .Y(n59) );
  INVX2TS U440 ( .A(destinationAddressIn_SOUTH[6]), .Y(n156) );
  INVX2TS U441 ( .A(n156), .Y(n699) );
  AOI22X1TS U442 ( .A0(n895), .A1(n699), .B0(n890), .B1(
        destinationAddressIn_NORTH[6]), .Y(n58) );
  OAI211XLTS U443 ( .A0(n60), .A1(n240), .B0(n59), .C0(n58), .Y(n2093) );
  INVX2TS U444 ( .A(destinationAddressIn_EAST[4]), .Y(n249) );
  AOI22X1TS U445 ( .A0(n64), .A1(\destinationAddressbuffer[7][4] ), .B0(n1521), 
        .B1(destinationAddressIn_WEST[4]), .Y(n62) );
  INVX2TS U446 ( .A(destinationAddressIn_SOUTH[4]), .Y(n167) );
  INVX2TS U447 ( .A(n167), .Y(n667) );
  AOI22X1TS U448 ( .A0(n49), .A1(n667), .B0(n1673), .B1(
        destinationAddressIn_NORTH[4]), .Y(n61) );
  OAI211XLTS U449 ( .A0(n1530), .A1(n249), .B0(n62), .C0(n61), .Y(n2091) );
  INVX2TS U450 ( .A(destinationAddressIn_EAST[5]), .Y(n244) );
  AOI22X1TS U451 ( .A0(n64), .A1(\destinationAddressbuffer[7][5] ), .B0(n63), 
        .B1(destinationAddressIn_WEST[5]), .Y(n67) );
  INVX2TS U452 ( .A(destinationAddressIn_SOUTH[5]), .Y(n150) );
  INVX2TS U453 ( .A(n150), .Y(n679) );
  AOI22X1TS U454 ( .A0(n65), .A1(n679), .B0(n38), .B1(
        destinationAddressIn_NORTH[5]), .Y(n66) );
  OAI211XLTS U455 ( .A0(n68), .A1(n244), .B0(n67), .C0(n66), .Y(n2092) );
  INVX2TS U456 ( .A(n209), .Y(n169) );
  NAND2X1TS U457 ( .A(n114), .B(n519), .Y(n260) );
  AOI21X1TS U458 ( .A0(n210), .A1(n70), .B0(n306), .Y(n382) );
  NOR3XLTS U459 ( .A(n382), .B(n262), .C(n261), .Y(n1585) );
  INVX2TS U460 ( .A(n1950), .Y(n463) );
  INVX2TS U461 ( .A(n1946), .Y(n454) );
  NOR2XLTS U462 ( .A(n454), .B(n511), .Y(n385) );
  INVX2TS U463 ( .A(n7), .Y(n263) );
  NOR3XLTS U464 ( .A(n24), .B(n71), .C(n263), .Y(n1582) );
  AOI31XLTS U465 ( .A0(n265), .A1(n463), .A2(n385), .B0(n1582), .Y(n72) );
  AOI21X1TS U466 ( .A0(n78), .A1(n72), .B0(n267), .Y(n77) );
  INVX2TS U467 ( .A(n119), .Y(n517) );
  INVX2TS U468 ( .A(n1942), .Y(n388) );
  NAND2X1TS U469 ( .A(n77), .B(n1589), .Y(n79) );
  INVX2TS U470 ( .A(n74), .Y(n1469) );
  INVX2TS U471 ( .A(n1469), .Y(n912) );
  CLKBUFX2TS U472 ( .A(n912), .Y(n86) );
  INVX2TS U473 ( .A(n86), .Y(n103) );
  INVX2TS U474 ( .A(n75), .Y(n448) );
  INVX2TS U475 ( .A(n76), .Y(n1484) );
  INVX2TS U476 ( .A(n1484), .Y(n902) );
  INVX2TS U477 ( .A(n1485), .Y(n91) );
  OR2X1TS U478 ( .A(n1586), .B(n79), .Y(n89) );
  INVX2TS U479 ( .A(n89), .Y(n1488) );
  INVX2TS U480 ( .A(n1488), .Y(n903) );
  INVX2TS U481 ( .A(n903), .Y(n104) );
  AOI22X1TS U482 ( .A0(n91), .A1(\destinationAddressbuffer[6][9] ), .B0(n104), 
        .B1(n738), .Y(n82) );
  CLKBUFX2TS U483 ( .A(n741), .Y(n414) );
  INVX2TS U484 ( .A(n4), .Y(n1718) );
  INVX2TS U485 ( .A(n1718), .Y(n904) );
  INVX2TS U486 ( .A(n904), .Y(n1498) );
  INVX2TS U487 ( .A(n133), .Y(n341) );
  AOI22X1TS U488 ( .A0(n97), .A1(n414), .B0(n1498), .B1(n341), .Y(n81) );
  OAI211XLTS U489 ( .A0(n103), .A1(n226), .B0(n82), .C0(n81), .Y(n2108) );
  INVX2TS U490 ( .A(n86), .Y(n108) );
  INVX2TS U491 ( .A(n89), .Y(n1700) );
  AOI22X1TS U492 ( .A0(n91), .A1(\destinationAddressbuffer[6][10] ), .B0(n1700), .B1(n755), .Y(n85) );
  INVX2TS U493 ( .A(n3), .Y(n1703) );
  CLKBUFX2TS U494 ( .A(n759), .Y(n407) );
  INVX2TS U495 ( .A(n4), .Y(n83) );
  INVX2TS U496 ( .A(n142), .Y(n319) );
  AOI22X1TS U497 ( .A0(n1703), .A1(n407), .B0(n83), .B1(n319), .Y(n84) );
  OAI211XLTS U498 ( .A0(n108), .A1(n214), .B0(n85), .C0(n84), .Y(n2109) );
  AOI22X1TS U499 ( .A0(n91), .A1(\destinationAddressbuffer[6][8] ), .B0(n94), 
        .B1(n723), .Y(n88) );
  INVX2TS U500 ( .A(n3), .Y(n1710) );
  CLKBUFX2TS U501 ( .A(n725), .Y(n401) );
  INVX2TS U502 ( .A(n4), .Y(n1702) );
  INVX2TS U503 ( .A(n129), .Y(n332) );
  AOI22X1TS U504 ( .A0(n1710), .A1(n401), .B0(n1702), .B1(n332), .Y(n87) );
  OAI211XLTS U505 ( .A0(n103), .A1(n230), .B0(n88), .C0(n87), .Y(n2107) );
  INVX2TS U506 ( .A(n89), .Y(n90) );
  AOI22X1TS U507 ( .A0(n91), .A1(\destinationAddressbuffer[6][11] ), .B0(n90), 
        .B1(n770), .Y(n93) );
  INVX2TS U508 ( .A(n3), .Y(n1694) );
  CLKBUFX2TS U509 ( .A(n774), .Y(n396) );
  INVX2TS U510 ( .A(n138), .Y(n325) );
  AOI22X1TS U511 ( .A0(n1694), .A1(n396), .B0(n1718), .B1(n325), .Y(n92) );
  OAI211XLTS U512 ( .A0(n103), .A1(n222), .B0(n93), .C0(n92), .Y(n2110) );
  INVX2TS U513 ( .A(n1590), .Y(n1714) );
  INVX2TS U514 ( .A(n903), .Y(n94) );
  AOI22X1TS U515 ( .A0(n1714), .A1(writeOutbuffer[6]), .B0(n94), .B1(n549), 
        .Y(n96) );
  CLKBUFX2TS U516 ( .A(n552), .Y(n421) );
  INVX2TS U517 ( .A(n4), .Y(n1514) );
  INVX2TS U518 ( .A(n146), .Y(n346) );
  AOI22X1TS U519 ( .A0(n1703), .A1(n421), .B0(n1514), .B1(n346), .Y(n95) );
  OAI211XLTS U520 ( .A0(n108), .A1(n237), .B0(n96), .C0(n95), .Y(n2072) );
  INVX2TS U521 ( .A(n1590), .Y(n109) );
  AOI22X1TS U522 ( .A0(n109), .A1(\destinationAddressbuffer[6][7] ), .B0(n104), 
        .B1(destinationAddressIn_WEST[7]), .Y(n99) );
  INVX2TS U523 ( .A(n3), .Y(n97) );
  INVX2TS U524 ( .A(n97), .Y(n905) );
  INVX2TS U525 ( .A(n905), .Y(n100) );
  CLKBUFX2TS U526 ( .A(destinationAddressIn_NORTH[7]), .Y(n359) );
  CLKBUFX2TS U527 ( .A(n359), .Y(n442) );
  INVX2TS U528 ( .A(n161), .Y(n358) );
  AOI22X1TS U529 ( .A0(n100), .A1(n442), .B0(n83), .B1(n358), .Y(n98) );
  OAI211XLTS U530 ( .A0(n108), .A1(n255), .B0(n99), .C0(n98), .Y(n2106) );
  AOI22X1TS U531 ( .A0(n109), .A1(\destinationAddressbuffer[6][4] ), .B0(n1700), .B1(destinationAddressIn_WEST[4]), .Y(n102) );
  CLKBUFX2TS U532 ( .A(destinationAddressIn_NORTH[4]), .Y(n375) );
  CLKBUFX2TS U533 ( .A(n375), .Y(n437) );
  INVX2TS U534 ( .A(n167), .Y(n374) );
  AOI22X1TS U535 ( .A0(n100), .A1(n437), .B0(n1514), .B1(n374), .Y(n101) );
  OAI211XLTS U536 ( .A0(n103), .A1(n249), .B0(n102), .C0(n101), .Y(n2103) );
  AOI22X1TS U537 ( .A0(n109), .A1(\destinationAddressbuffer[6][6] ), .B0(n104), 
        .B1(destinationAddressIn_WEST[6]), .Y(n107) );
  CLKBUFX2TS U538 ( .A(destinationAddressIn_NORTH[6]), .Y(n367) );
  CLKBUFX2TS U539 ( .A(n367), .Y(n432) );
  INVX2TS U540 ( .A(n904), .Y(n105) );
  INVX2TS U541 ( .A(n156), .Y(n365) );
  AOI22X1TS U542 ( .A0(n97), .A1(n432), .B0(n105), .B1(n365), .Y(n106) );
  OAI211XLTS U543 ( .A0(n108), .A1(n240), .B0(n107), .C0(n106), .Y(n2105) );
  AOI22X1TS U544 ( .A0(n109), .A1(\destinationAddressbuffer[6][5] ), .B0(n90), 
        .B1(destinationAddressIn_WEST[5]), .Y(n111) );
  CLKBUFX2TS U545 ( .A(destinationAddressIn_NORTH[5]), .Y(n354) );
  CLKBUFX2TS U546 ( .A(n354), .Y(n427) );
  INVX2TS U547 ( .A(n150), .Y(n353) );
  AOI22X1TS U548 ( .A0(n1694), .A1(n427), .B0(n1702), .B1(n353), .Y(n110) );
  OAI211XLTS U549 ( .A0(n1469), .A1(n244), .B0(n111), .C0(n110), .Y(n2104) );
  INVX2TS U550 ( .A(n1947), .Y(n451) );
  NAND2X1TS U551 ( .A(n117), .B(n451), .Y(n118) );
  INVX2TS U552 ( .A(n211), .Y(n457) );
  AOI31XLTS U553 ( .A0(n120), .A1(n26), .A2(n118), .B0(n457), .Y(n123) );
  INVX2TS U554 ( .A(n119), .Y(n516) );
  INVX2TS U555 ( .A(n1947), .Y(n449) );
  INVX2TS U556 ( .A(n121), .Y(n974) );
  INVX2TS U557 ( .A(n974), .Y(n1384) );
  CLKBUFX2TS U558 ( .A(n1384), .Y(n134) );
  INVX2TS U559 ( .A(n134), .Y(n157) );
  INVX2TS U560 ( .A(n122), .Y(n1388) );
  INVX2TS U561 ( .A(n1388), .Y(n964) );
  INVX2TS U562 ( .A(n1624), .Y(n139) );
  NOR3XLTS U563 ( .A(n1622), .B(n1617), .C(n125), .Y(n130) );
  INVX2TS U564 ( .A(n130), .Y(n162) );
  INVX2TS U565 ( .A(n162), .Y(n1379) );
  AOI22X1TS U566 ( .A0(n139), .A1(\destinationAddressbuffer[3][8] ), .B0(n1379), .B1(destinationAddressIn_EAST[8]), .Y(n128) );
  OR2X1TS U567 ( .A(n112), .B(n124), .Y(n152) );
  INVX2TS U568 ( .A(n152), .Y(n1801) );
  INVX2TS U569 ( .A(n126), .Y(n143) );
  INVX2TS U570 ( .A(n143), .Y(n1397) );
  CLKBUFX2TS U571 ( .A(n400), .Y(n331) );
  AOI22X1TS U572 ( .A0(n1801), .A1(n333), .B0(n1397), .B1(n331), .Y(n127) );
  OAI211XLTS U573 ( .A0(n157), .A1(n129), .B0(n128), .C0(n127), .Y(n2143) );
  INVX2TS U574 ( .A(n130), .Y(n965) );
  INVX2TS U575 ( .A(n965), .Y(n151) );
  AOI22X1TS U576 ( .A0(n139), .A1(\destinationAddressbuffer[3][9] ), .B0(n151), 
        .B1(destinationAddressIn_EAST[9]), .Y(n132) );
  INVX2TS U577 ( .A(n152), .Y(n1398) );
  INVX2TS U578 ( .A(n967), .Y(n975) );
  CLKBUFX2TS U579 ( .A(n412), .Y(n337) );
  AOI22X1TS U580 ( .A0(n975), .A1(n342), .B0(n1397), .B1(n337), .Y(n131) );
  OAI211XLTS U581 ( .A0(n974), .A1(n133), .B0(n132), .C0(n131), .Y(n2144) );
  INVX2TS U582 ( .A(n134), .Y(n168) );
  INVX2TS U583 ( .A(n162), .Y(n1792) );
  AOI22X1TS U584 ( .A0(n139), .A1(\destinationAddressbuffer[3][11] ), .B0(
        n1792), .B1(destinationAddressIn_EAST[11]), .Y(n137) );
  INVX2TS U585 ( .A(n143), .Y(n135) );
  INVX2TS U586 ( .A(n135), .Y(n957) );
  INVX2TS U587 ( .A(n957), .Y(n147) );
  CLKBUFX2TS U588 ( .A(n391), .Y(n324) );
  AOI22X1TS U589 ( .A0(n1398), .A1(n326), .B0(n147), .B1(n324), .Y(n136) );
  OAI211XLTS U590 ( .A0(n168), .A1(n138), .B0(n137), .C0(n136), .Y(n2146) );
  AOI22X1TS U591 ( .A0(n139), .A1(\destinationAddressbuffer[3][10] ), .B0(
        n1379), .B1(destinationAddressIn_EAST[10]), .Y(n141) );
  INVX2TS U592 ( .A(n152), .Y(n1795) );
  INVX2TS U593 ( .A(n143), .Y(n1787) );
  CLKBUFX2TS U594 ( .A(n406), .Y(n313) );
  AOI22X1TS U595 ( .A0(n1795), .A1(n321), .B0(n1787), .B1(n313), .Y(n140) );
  OAI211XLTS U596 ( .A0(n157), .A1(n142), .B0(n141), .C0(n140), .Y(n2145) );
  INVX2TS U597 ( .A(n1624), .Y(n1805) );
  INVX2TS U598 ( .A(n162), .Y(n1396) );
  AOI22X1TS U599 ( .A0(n1805), .A1(writeOutbuffer[3]), .B0(n1396), .B1(
        writeIn_EAST), .Y(n145) );
  INVX2TS U600 ( .A(n143), .Y(n1809) );
  CLKBUFX2TS U601 ( .A(n420), .Y(n345) );
  AOI22X1TS U602 ( .A0(n1795), .A1(n347), .B0(n1809), .B1(n345), .Y(n144) );
  OAI211XLTS U603 ( .A0(n157), .A1(n146), .B0(n145), .C0(n144), .Y(n2075) );
  INVX2TS U604 ( .A(n1389), .Y(n164) );
  AOI22X1TS U605 ( .A0(n164), .A1(\destinationAddressbuffer[3][5] ), .B0(n1792), .B1(destinationAddressIn_EAST[5]), .Y(n149) );
  CLKBUFX2TS U606 ( .A(destinationAddressIn_WEST[5]), .Y(n678) );
  CLKBUFX2TS U607 ( .A(n678), .Y(n351) );
  AOI22X1TS U608 ( .A0(n975), .A1(n354), .B0(n147), .B1(n351), .Y(n148) );
  OAI211XLTS U609 ( .A0(n168), .A1(n150), .B0(n149), .C0(n148), .Y(n2140) );
  AOI22X1TS U610 ( .A0(n164), .A1(\destinationAddressbuffer[3][6] ), .B0(n151), 
        .B1(destinationAddressIn_EAST[6]), .Y(n155) );
  INVX2TS U611 ( .A(n152), .Y(n153) );
  INVX2TS U612 ( .A(n153), .Y(n967) );
  INVX2TS U613 ( .A(n967), .Y(n158) );
  CLKBUFX2TS U614 ( .A(destinationAddressIn_WEST[6]), .Y(n697) );
  CLKBUFX2TS U615 ( .A(n697), .Y(n363) );
  AOI22X1TS U616 ( .A0(n158), .A1(n367), .B0(n1787), .B1(n363), .Y(n154) );
  OAI211XLTS U617 ( .A0(n157), .A1(n156), .B0(n155), .C0(n154), .Y(n2141) );
  AOI22X1TS U618 ( .A0(n164), .A1(\destinationAddressbuffer[3][7] ), .B0(n1396), .B1(destinationAddressIn_EAST[7]), .Y(n160) );
  CLKBUFX2TS U619 ( .A(destinationAddressIn_WEST[7]), .Y(n712) );
  CLKBUFX2TS U620 ( .A(n712), .Y(n357) );
  AOI22X1TS U621 ( .A0(n158), .A1(n359), .B0(n1809), .B1(n357), .Y(n159) );
  OAI211XLTS U622 ( .A0(n168), .A1(n161), .B0(n160), .C0(n159), .Y(n2142) );
  INVX2TS U623 ( .A(n162), .Y(n163) );
  AOI22X1TS U624 ( .A0(n164), .A1(\destinationAddressbuffer[3][4] ), .B0(n151), 
        .B1(destinationAddressIn_EAST[4]), .Y(n166) );
  CLKBUFX2TS U625 ( .A(destinationAddressIn_WEST[4]), .Y(n665) );
  CLKBUFX2TS U626 ( .A(n665), .Y(n371) );
  AOI22X1TS U627 ( .A0(n1398), .A1(n375), .B0(n135), .B1(n371), .Y(n165) );
  OAI211XLTS U628 ( .A0(n168), .A1(n167), .B0(n166), .C0(n165), .Y(n2139) );
  INVX2TS U629 ( .A(n261), .Y(n307) );
  INVX2TS U630 ( .A(n307), .Y(n380) );
  NOR3XLTS U631 ( .A(n382), .B(n380), .C(n381), .Y(n1631) );
  AOI31XLTS U632 ( .A0(n502), .A1(n385), .A2(n458), .B0(n1628), .Y(n170) );
  AOI21X1TS U633 ( .A0(n173), .A1(n170), .B0(n448), .Y(n172) );
  NAND2X1TS U634 ( .A(n172), .B(n1635), .Y(n174) );
  INVX2TS U635 ( .A(n171), .Y(n1357) );
  INVX2TS U636 ( .A(n1357), .Y(n999) );
  CLKBUFX2TS U637 ( .A(n999), .Y(n182) );
  INVX2TS U638 ( .A(n9), .Y(n989) );
  INVX2TS U639 ( .A(n1356), .Y(n187) );
  OR2X1TS U640 ( .A(n1632), .B(n174), .Y(n185) );
  INVX2TS U641 ( .A(n185), .Y(n1820) );
  AOI22X1TS U642 ( .A0(n187), .A1(\destinationAddressbuffer[2][8] ), .B0(n1820), .B1(n331), .Y(n178) );
  INVX2TS U643 ( .A(n179), .Y(n199) );
  INVX2TS U644 ( .A(n199), .Y(n1821) );
  INVX2TS U645 ( .A(n176), .Y(n190) );
  AOI22X1TS U646 ( .A0(n1821), .A1(n333), .B0(n201), .B1(n332), .Y(n177) );
  OAI211XLTS U647 ( .A0(n204), .A1(n230), .B0(n178), .C0(n177), .Y(n2155) );
  INVX2TS U648 ( .A(n182), .Y(n204) );
  INVX2TS U649 ( .A(n185), .Y(n1814) );
  AOI22X1TS U650 ( .A0(n187), .A1(\destinationAddressbuffer[2][9] ), .B0(n1814), .B1(n337), .Y(n181) );
  INVX2TS U651 ( .A(n179), .Y(n1352) );
  INVX2TS U652 ( .A(n1352), .Y(n994) );
  INVX2TS U653 ( .A(n190), .Y(n1836) );
  INVX2TS U654 ( .A(n190), .Y(n1366) );
  AOI22X1TS U655 ( .A0(n994), .A1(n342), .B0(n1366), .B1(n341), .Y(n180) );
  OAI211XLTS U656 ( .A0(n204), .A1(n226), .B0(n181), .C0(n180), .Y(n2156) );
  INVX2TS U657 ( .A(n182), .Y(n208) );
  INVX2TS U658 ( .A(n185), .Y(n1828) );
  AOI22X1TS U659 ( .A0(n187), .A1(\destinationAddressbuffer[2][10] ), .B0(
        n1828), .B1(n313), .Y(n184) );
  INVX2TS U660 ( .A(n199), .Y(n1830) );
  INVX2TS U661 ( .A(n176), .Y(n993) );
  INVX2TS U662 ( .A(n993), .Y(n201) );
  AOI22X1TS U663 ( .A0(n1830), .A1(n321), .B0(n201), .B1(n319), .Y(n183) );
  OAI211XLTS U664 ( .A0(n208), .A1(n214), .B0(n184), .C0(n183), .Y(n2157) );
  INVX2TS U665 ( .A(n185), .Y(n186) );
  INVX2TS U666 ( .A(n186), .Y(n998) );
  INVX2TS U667 ( .A(n998), .Y(n196) );
  AOI22X1TS U668 ( .A0(n187), .A1(\destinationAddressbuffer[2][11] ), .B0(n196), .B1(n324), .Y(n189) );
  INVX2TS U669 ( .A(n199), .Y(n1361) );
  AOI22X1TS U670 ( .A0(n1361), .A1(n326), .B0(n1836), .B1(n325), .Y(n188) );
  OAI211XLTS U671 ( .A0(n208), .A1(n222), .B0(n189), .C0(n188), .Y(n2158) );
  INVX2TS U672 ( .A(n1636), .Y(n1834) );
  AOI22X1TS U673 ( .A0(n1834), .A1(writeOutbuffer[2]), .B0(n196), .B1(n345), 
        .Y(n192) );
  AOI22X1TS U674 ( .A0(n1830), .A1(n347), .B0(n176), .B1(n346), .Y(n191) );
  OAI211XLTS U675 ( .A0(n204), .A1(n237), .B0(n192), .C0(n191), .Y(n2076) );
  INVX2TS U676 ( .A(n1356), .Y(n205) );
  AOI22X1TS U677 ( .A0(n205), .A1(\destinationAddressbuffer[2][6] ), .B0(n186), 
        .B1(n363), .Y(n195) );
  INVX2TS U678 ( .A(n190), .Y(n193) );
  AOI22X1TS U679 ( .A0(n994), .A1(destinationAddressIn_NORTH[6]), .B0(n193), 
        .B1(n365), .Y(n194) );
  OAI211XLTS U680 ( .A0(n208), .A1(n240), .B0(n195), .C0(n194), .Y(n2153) );
  AOI22X1TS U681 ( .A0(n205), .A1(\destinationAddressbuffer[2][5] ), .B0(n196), 
        .B1(n351), .Y(n198) );
  AOI22X1TS U682 ( .A0(n1361), .A1(destinationAddressIn_NORTH[5]), .B0(n1360), 
        .B1(n353), .Y(n197) );
  OAI211XLTS U683 ( .A0(n1357), .A1(n244), .B0(n198), .C0(n197), .Y(n2152) );
  AOI22X1TS U684 ( .A0(n205), .A1(\destinationAddressbuffer[2][7] ), .B0(n1820), .B1(n357), .Y(n203) );
  INVX2TS U685 ( .A(n199), .Y(n200) );
  AOI22X1TS U686 ( .A0(n200), .A1(destinationAddressIn_NORTH[7]), .B0(n201), 
        .B1(n358), .Y(n202) );
  OAI211XLTS U687 ( .A0(n204), .A1(n255), .B0(n203), .C0(n202), .Y(n2154) );
  AOI22X1TS U688 ( .A0(n205), .A1(\destinationAddressbuffer[2][4] ), .B0(n1828), .B1(n371), .Y(n207) );
  AOI22X1TS U689 ( .A0(n200), .A1(destinationAddressIn_NORTH[4]), .B0(n176), 
        .B1(n374), .Y(n206) );
  OAI211XLTS U690 ( .A0(n208), .A1(n249), .B0(n207), .C0(n206), .Y(n2151) );
  INVX2TS U691 ( .A(n1945), .Y(n387) );
  INVX2TS U692 ( .A(n211), .Y(n267) );
  AOI31XLTS U693 ( .A0(n216), .A1(n1592), .A2(n212), .B0(n267), .Y(n215) );
  INVX2TS U694 ( .A(n1945), .Y(n384) );
  NAND2X1TS U695 ( .A(n215), .B(n1602), .Y(n217) );
  INVX2TS U696 ( .A(n213), .Y(n1440) );
  INVX2TS U697 ( .A(n1440), .Y(n928) );
  CLKBUFX2TS U698 ( .A(n928), .Y(n225) );
  INVX2TS U699 ( .A(n225), .Y(n248) );
  CLKBUFX2TS U700 ( .A(n214), .Y(n411) );
  INVX2TS U701 ( .A(n10), .Y(n920) );
  INVX2TS U702 ( .A(n1451), .Y(n233) );
  OR2X1TS U703 ( .A(n1599), .B(n217), .Y(n231) );
  INVX2TS U704 ( .A(n231), .Y(n1456) );
  AOI22X1TS U705 ( .A0(n233), .A1(\destinationAddressbuffer[5][10] ), .B0(
        n1456), .B1(n755), .Y(n221) );
  INVX2TS U706 ( .A(n227), .Y(n257) );
  INVX2TS U707 ( .A(n257), .Y(n218) );
  OR2X1TS U708 ( .A(n1592), .B(n219), .Y(n245) );
  INVX2TS U709 ( .A(n245), .Y(n1460) );
  AOI22X1TS U710 ( .A0(n218), .A1(n407), .B0(n1460), .B1(n319), .Y(n220) );
  OAI211XLTS U711 ( .A0(n248), .A1(n411), .B0(n221), .C0(n220), .Y(n2121) );
  INVX2TS U712 ( .A(n225), .Y(n254) );
  CLKBUFX2TS U713 ( .A(n222), .Y(n399) );
  INVX2TS U714 ( .A(n231), .Y(n1732) );
  AOI22X1TS U715 ( .A0(n233), .A1(\destinationAddressbuffer[5][11] ), .B0(
        n1732), .B1(n770), .Y(n224) );
  INVX2TS U716 ( .A(n257), .Y(n1447) );
  AOI22X1TS U717 ( .A0(n1447), .A1(n396), .B0(n1460), .B1(n325), .Y(n223) );
  OAI211XLTS U718 ( .A0(n254), .A1(n399), .B0(n224), .C0(n223), .Y(n2122) );
  CLKBUFX2TS U719 ( .A(n226), .Y(n417) );
  INVX2TS U720 ( .A(n231), .Y(n1452) );
  AOI22X1TS U721 ( .A0(n233), .A1(\destinationAddressbuffer[5][9] ), .B0(n1452), .B1(n738), .Y(n229) );
  INVX2TS U722 ( .A(n227), .Y(n1441) );
  INVX2TS U723 ( .A(n1441), .Y(n241) );
  INVX2TS U724 ( .A(n245), .Y(n1744) );
  AOI22X1TS U725 ( .A0(n241), .A1(n414), .B0(n1744), .B1(n341), .Y(n228) );
  OAI211XLTS U726 ( .A0(n248), .A1(n417), .B0(n229), .C0(n228), .Y(n2120) );
  CLKBUFX2TS U727 ( .A(n230), .Y(n404) );
  INVX2TS U728 ( .A(n231), .Y(n232) );
  INVX2TS U729 ( .A(n232), .Y(n927) );
  INVX2TS U730 ( .A(n927), .Y(n250) );
  AOI22X1TS U731 ( .A0(n233), .A1(\destinationAddressbuffer[5][8] ), .B0(n250), 
        .B1(n723), .Y(n236) );
  INVX2TS U732 ( .A(n245), .Y(n234) );
  INVX2TS U733 ( .A(n234), .Y(n916) );
  INVX2TS U734 ( .A(n916), .Y(n251) );
  AOI22X1TS U735 ( .A0(n1447), .A1(n401), .B0(n251), .B1(n332), .Y(n235) );
  OAI211XLTS U736 ( .A0(n248), .A1(n404), .B0(n236), .C0(n235), .Y(n2119) );
  CLKBUFX2TS U737 ( .A(n237), .Y(n424) );
  INVX2TS U738 ( .A(n1603), .Y(n1749) );
  AOI22X1TS U739 ( .A0(n1749), .A1(writeOutbuffer[5]), .B0(n250), .B1(n549), 
        .Y(n239) );
  AOI22X1TS U740 ( .A0(n241), .A1(n421), .B0(n251), .B1(n346), .Y(n238) );
  OAI211XLTS U741 ( .A0(n254), .A1(n424), .B0(n239), .C0(n238), .Y(n2073) );
  CLKBUFX2TS U742 ( .A(n240), .Y(n435) );
  INVX2TS U743 ( .A(n1603), .Y(n256) );
  AOI22X1TS U744 ( .A0(n256), .A1(\destinationAddressbuffer[5][6] ), .B0(n232), 
        .B1(n697), .Y(n243) );
  AOI22X1TS U745 ( .A0(n241), .A1(n432), .B0(n234), .B1(n365), .Y(n242) );
  OAI211XLTS U746 ( .A0(n254), .A1(n435), .B0(n243), .C0(n242), .Y(n2117) );
  CLKBUFX2TS U747 ( .A(n244), .Y(n430) );
  AOI22X1TS U748 ( .A0(n256), .A1(\destinationAddressbuffer[5][5] ), .B0(n1456), .B1(n678), .Y(n247) );
  INVX2TS U749 ( .A(n245), .Y(n1442) );
  AOI22X1TS U750 ( .A0(n218), .A1(n427), .B0(n1442), .B1(n353), .Y(n246) );
  OAI211XLTS U751 ( .A0(n248), .A1(n430), .B0(n247), .C0(n246), .Y(n2116) );
  CLKBUFX2TS U752 ( .A(n249), .Y(n440) );
  AOI22X1TS U753 ( .A0(n256), .A1(\destinationAddressbuffer[5][4] ), .B0(n250), 
        .B1(n665), .Y(n253) );
  INVX2TS U754 ( .A(n257), .Y(n1745) );
  AOI22X1TS U755 ( .A0(n1745), .A1(n437), .B0(n251), .B1(n374), .Y(n252) );
  OAI211XLTS U756 ( .A0(n254), .A1(n440), .B0(n253), .C0(n252), .Y(n2115) );
  CLKBUFX2TS U757 ( .A(n255), .Y(n446) );
  AOI22X1TS U758 ( .A0(n256), .A1(\destinationAddressbuffer[5][7] ), .B0(n1732), .B1(n712), .Y(n259) );
  INVX2TS U759 ( .A(n257), .Y(n1724) );
  AOI22X1TS U760 ( .A0(n1724), .A1(n442), .B0(n1442), .B1(n358), .Y(n258) );
  OAI211XLTS U761 ( .A0(n1440), .A1(n446), .B0(n259), .C0(n258), .Y(n2118) );
  AOI31XLTS U762 ( .A0(n487), .A1(n385), .A2(n387), .B0(n1606), .Y(n264) );
  AOI21X1TS U763 ( .A0(n270), .A1(n264), .B0(n267), .Y(n269) );
  NAND2X1TS U764 ( .A(n269), .B(n1614), .Y(n271) );
  INVX2TS U765 ( .A(n266), .Y(n1407) );
  INVX2TS U766 ( .A(n1407), .Y(n950) );
  CLKBUFX2TS U767 ( .A(n950), .Y(n279) );
  INVX2TS U768 ( .A(n279), .Y(n298) );
  INVX2TS U769 ( .A(n268), .Y(n1419) );
  INVX2TS U770 ( .A(n1419), .Y(n937) );
  INVX2TS U771 ( .A(n1420), .Y(n285) );
  OR2X1TS U772 ( .A(n1610), .B(n271), .Y(n283) );
  INVX2TS U773 ( .A(n283), .Y(n1774) );
  AOI22X1TS U774 ( .A0(n285), .A1(\destinationAddressbuffer[4][11] ), .B0(
        n1774), .B1(n324), .Y(n275) );
  INVX2TS U775 ( .A(n276), .Y(n295) );
  INVX2TS U776 ( .A(n295), .Y(n1422) );
  INVX2TS U777 ( .A(n6), .Y(n273) );
  AOI22X1TS U778 ( .A0(n1422), .A1(n773), .B0(n273), .B1(n396), .Y(n274) );
  OAI211XLTS U779 ( .A0(n298), .A1(n399), .B0(n275), .C0(n274), .Y(n2134) );
  INVX2TS U780 ( .A(n283), .Y(n1764) );
  AOI22X1TS U781 ( .A0(n285), .A1(\destinationAddressbuffer[4][10] ), .B0(
        n1764), .B1(n313), .Y(n278) );
  INVX2TS U782 ( .A(n276), .Y(n1414) );
  INVX2TS U783 ( .A(n1414), .Y(n302) );
  AOI22X1TS U784 ( .A0(n302), .A1(n758), .B0(n273), .B1(n407), .Y(n277) );
  OAI211XLTS U785 ( .A0(n298), .A1(n411), .B0(n278), .C0(n277), .Y(n2133) );
  INVX2TS U786 ( .A(n279), .Y(n305) );
  INVX2TS U787 ( .A(n283), .Y(n1756) );
  INVX2TS U788 ( .A(n1756), .Y(n938) );
  INVX2TS U789 ( .A(n938), .Y(n294) );
  AOI22X1TS U790 ( .A0(n285), .A1(\destinationAddressbuffer[4][9] ), .B0(n294), 
        .B1(n337), .Y(n282) );
  INVX2TS U791 ( .A(n295), .Y(n280) );
  INVX2TS U792 ( .A(n6), .Y(n1757) );
  INVX2TS U793 ( .A(n1757), .Y(n1415) );
  INVX2TS U794 ( .A(n1415), .Y(n940) );
  AOI22X1TS U795 ( .A0(n1766), .A1(n739), .B0(n940), .B1(n414), .Y(n281) );
  OAI211XLTS U796 ( .A0(n305), .A1(n417), .B0(n282), .C0(n281), .Y(n2132) );
  INVX2TS U797 ( .A(n283), .Y(n284) );
  AOI22X1TS U798 ( .A0(n285), .A1(\destinationAddressbuffer[4][8] ), .B0(n284), 
        .B1(n331), .Y(n287) );
  INVX2TS U799 ( .A(n295), .Y(n1781) );
  AOI22X1TS U800 ( .A0(n1781), .A1(n724), .B0(n291), .B1(n401), .Y(n286) );
  OAI211XLTS U801 ( .A0(n298), .A1(n404), .B0(n287), .C0(n286), .Y(n2131) );
  INVX2TS U802 ( .A(n1615), .Y(n1778) );
  INVX2TS U803 ( .A(n938), .Y(n288) );
  AOI22X1TS U804 ( .A0(n1778), .A1(writeOutbuffer[4]), .B0(n288), .B1(n345), 
        .Y(n290) );
  INVX2TS U805 ( .A(n6), .Y(n1765) );
  AOI22X1TS U806 ( .A0(n1781), .A1(n551), .B0(n1765), .B1(n421), .Y(n289) );
  OAI211XLTS U807 ( .A0(n305), .A1(n424), .B0(n290), .C0(n289), .Y(n2074) );
  INVX2TS U808 ( .A(n1615), .Y(n301) );
  AOI22X1TS U809 ( .A0(n301), .A1(\destinationAddressbuffer[4][5] ), .B0(n1764), .B1(n351), .Y(n293) );
  INVX2TS U810 ( .A(n1415), .Y(n291) );
  AOI22X1TS U811 ( .A0(n302), .A1(n679), .B0(n291), .B1(n427), .Y(n292) );
  OAI211XLTS U812 ( .A0(n305), .A1(n430), .B0(n293), .C0(n292), .Y(n2128) );
  AOI22X1TS U813 ( .A0(n301), .A1(\destinationAddressbuffer[4][6] ), .B0(n294), 
        .B1(n363), .Y(n297) );
  INVX2TS U814 ( .A(n295), .Y(n1436) );
  AOI22X1TS U815 ( .A0(n1436), .A1(n699), .B0(n940), .B1(n432), .Y(n296) );
  OAI211XLTS U816 ( .A0(n298), .A1(n435), .B0(n297), .C0(n296), .Y(n2129) );
  AOI22X1TS U817 ( .A0(n301), .A1(\destinationAddressbuffer[4][7] ), .B0(n1774), .B1(n357), .Y(n300) );
  AOI22X1TS U818 ( .A0(n302), .A1(n713), .B0(n1765), .B1(n442), .Y(n299) );
  OAI211XLTS U819 ( .A0(n1407), .A1(n446), .B0(n300), .C0(n299), .Y(n2130) );
  AOI22X1TS U820 ( .A0(n301), .A1(\destinationAddressbuffer[4][4] ), .B0(n284), 
        .B1(n371), .Y(n304) );
  AOI22X1TS U821 ( .A0(n302), .A1(n667), .B0(n940), .B1(n437), .Y(n303) );
  OAI211XLTS U822 ( .A0(n305), .A1(n440), .B0(n304), .C0(n303), .Y(n2127) );
  AOI31XLTS U823 ( .A0(n18), .A1(n384), .A2(n458), .B0(n1640), .Y(n308) );
  AOI21X1TS U824 ( .A0(n314), .A1(n308), .B0(n310), .Y(n312) );
  NAND2X1TS U825 ( .A(n312), .B(n1649), .Y(n315) );
  INVX2TS U826 ( .A(n1), .Y(n1026) );
  CLKBUFX2TS U827 ( .A(n1026), .Y(n329) );
  INVX2TS U828 ( .A(n329), .Y(n362) );
  INVX2TS U829 ( .A(n311), .Y(n1097) );
  INVX2TS U830 ( .A(n1097), .Y(n1010) );
  CLKBUFX2TS U831 ( .A(n350), .Y(n1017) );
  INVX2TS U832 ( .A(n1017), .Y(n338) );
  OR2X1TS U833 ( .A(n1645), .B(n315), .Y(n336) );
  INVX2TS U834 ( .A(n336), .Y(n1854) );
  AOI22X1TS U835 ( .A0(n338), .A1(\destinationAddressbuffer[1][10] ), .B0(
        n1854), .B1(n313), .Y(n323) );
  INVX2TS U836 ( .A(n339), .Y(n352) );
  INVX2TS U837 ( .A(n352), .Y(n316) );
  INVX2TS U838 ( .A(n318), .Y(n340) );
  INVX2TS U839 ( .A(n340), .Y(n1878) );
  INVX2TS U840 ( .A(n340), .Y(n320) );
  AOI22X1TS U841 ( .A0(n316), .A1(n321), .B0(n320), .B1(n319), .Y(n322) );
  OAI211XLTS U842 ( .A0(n362), .A1(n411), .B0(n323), .C0(n322), .Y(n2169) );
  INVX2TS U843 ( .A(n329), .Y(n370) );
  INVX2TS U844 ( .A(n336), .Y(n1866) );
  AOI22X1TS U845 ( .A0(n338), .A1(\destinationAddressbuffer[1][11] ), .B0(
        n1866), .B1(n324), .Y(n328) );
  INVX2TS U846 ( .A(n318), .Y(n1028) );
  INVX2TS U847 ( .A(n1028), .Y(n366) );
  AOI22X1TS U848 ( .A0(n316), .A1(n326), .B0(n366), .B1(n325), .Y(n327) );
  OAI211XLTS U849 ( .A0(n370), .A1(n399), .B0(n328), .C0(n327), .Y(n2170) );
  INVX2TS U850 ( .A(n329), .Y(n378) );
  INVX2TS U851 ( .A(n336), .Y(n330) );
  INVX2TS U852 ( .A(n330), .Y(n1025) );
  INVX2TS U853 ( .A(n1025), .Y(n372) );
  AOI22X1TS U854 ( .A0(n338), .A1(\destinationAddressbuffer[1][8] ), .B0(n372), 
        .B1(n331), .Y(n335) );
  INVX2TS U855 ( .A(n352), .Y(n1846) );
  AOI22X1TS U856 ( .A0(n1846), .A1(n333), .B0(n318), .B1(n332), .Y(n334) );
  OAI211XLTS U857 ( .A0(n378), .A1(n404), .B0(n335), .C0(n334), .Y(n2167) );
  INVX2TS U858 ( .A(n336), .Y(n1843) );
  AOI22X1TS U859 ( .A0(n338), .A1(\destinationAddressbuffer[1][9] ), .B0(n1843), .B1(n337), .Y(n344) );
  INVX2TS U860 ( .A(n339), .Y(n364) );
  INVX2TS U861 ( .A(n364), .Y(n1019) );
  AOI22X1TS U862 ( .A0(n1019), .A1(n342), .B0(n366), .B1(n341), .Y(n343) );
  OAI211XLTS U863 ( .A0(n362), .A1(n417), .B0(n344), .C0(n343), .Y(n2168) );
  INVX2TS U864 ( .A(n350), .Y(n1874) );
  AOI22X1TS U865 ( .A0(n1874), .A1(writeOutbuffer[1]), .B0(n372), .B1(n345), 
        .Y(n349) );
  INVX2TS U866 ( .A(n352), .Y(n1870) );
  AOI22X1TS U867 ( .A0(n1870), .A1(n347), .B0(n318), .B1(n346), .Y(n348) );
  OAI211XLTS U868 ( .A0(n370), .A1(n424), .B0(n349), .C0(n348), .Y(n2077) );
  INVX2TS U869 ( .A(n350), .Y(n373) );
  AOI22X1TS U870 ( .A0(n373), .A1(\destinationAddressbuffer[1][5] ), .B0(n1854), .B1(n351), .Y(n356) );
  INVX2TS U871 ( .A(n352), .Y(n1857) );
  INVX2TS U872 ( .A(n1028), .Y(n1107) );
  AOI22X1TS U873 ( .A0(n1857), .A1(n354), .B0(n1107), .B1(n353), .Y(n355) );
  OAI211XLTS U874 ( .A0(n378), .A1(n430), .B0(n356), .C0(n355), .Y(n2164) );
  AOI22X1TS U875 ( .A0(n373), .A1(\destinationAddressbuffer[1][7] ), .B0(n1866), .B1(n357), .Y(n361) );
  AOI22X1TS U876 ( .A0(n1857), .A1(n359), .B0(n1878), .B1(n358), .Y(n360) );
  OAI211XLTS U877 ( .A0(n362), .A1(n446), .B0(n361), .C0(n360), .Y(n2166) );
  AOI22X1TS U878 ( .A0(n373), .A1(\destinationAddressbuffer[1][6] ), .B0(n330), 
        .B1(n363), .Y(n369) );
  INVX2TS U879 ( .A(n364), .Y(n1880) );
  AOI22X1TS U880 ( .A0(n1880), .A1(n367), .B0(n366), .B1(n365), .Y(n368) );
  OAI211XLTS U881 ( .A0(n370), .A1(n435), .B0(n369), .C0(n368), .Y(n2165) );
  AOI22X1TS U882 ( .A0(n373), .A1(\destinationAddressbuffer[1][4] ), .B0(n372), 
        .B1(n371), .Y(n377) );
  AOI22X1TS U883 ( .A0(n1846), .A1(n375), .B0(n1101), .B1(n374), .Y(n376) );
  OAI211XLTS U884 ( .A0(n378), .A1(n440), .B0(n377), .C0(n376), .Y(n2163) );
  AOI31XLTS U885 ( .A0(n385), .A1(n384), .A2(n449), .B0(n1653), .Y(n386) );
  AOI21X1TS U886 ( .A0(n392), .A1(n386), .B0(n457), .Y(n390) );
  NAND2X1TS U887 ( .A(n390), .B(n1661), .Y(n393) );
  INVX2TS U888 ( .A(n389), .Y(n1068) );
  INVX2TS U889 ( .A(n1068), .Y(n1053) );
  CLKBUFX2TS U890 ( .A(n1053), .Y(n405) );
  INVX2TS U891 ( .A(n405), .Y(n436) );
  INVX2TS U892 ( .A(n11), .Y(n1041) );
  INVX2TS U893 ( .A(n425), .Y(n413) );
  OR2X1TS U894 ( .A(n1658), .B(n393), .Y(n418) );
  INVX2TS U895 ( .A(n418), .Y(n1885) );
  AOI22X1TS U896 ( .A0(n413), .A1(\destinationAddressbuffer[0][11] ), .B0(
        n1885), .B1(n391), .Y(n398) );
  INVX2TS U897 ( .A(n5), .Y(n395) );
  INVX2TS U898 ( .A(n395), .Y(n1036) );
  INVX2TS U899 ( .A(n1036), .Y(n408) );
  AOI22X1TS U900 ( .A0(n431), .A1(n773), .B0(n408), .B1(n396), .Y(n397) );
  OAI211XLTS U901 ( .A0(n436), .A1(n399), .B0(n398), .C0(n397), .Y(n2182) );
  INVX2TS U902 ( .A(n418), .Y(n1894) );
  AOI22X1TS U903 ( .A0(n413), .A1(\destinationAddressbuffer[0][8] ), .B0(n1894), .B1(n400), .Y(n403) );
  INVX2TS U904 ( .A(n5), .Y(n1908) );
  AOI22X1TS U905 ( .A0(n431), .A1(n724), .B0(n1908), .B1(n401), .Y(n402) );
  OAI211XLTS U906 ( .A0(n447), .A1(n404), .B0(n403), .C0(n402), .Y(n2179) );
  INVX2TS U907 ( .A(n405), .Y(n447) );
  INVX2TS U908 ( .A(n418), .Y(n1906) );
  AOI22X1TS U909 ( .A0(n413), .A1(\destinationAddressbuffer[0][10] ), .B0(
        n1906), .B1(n406), .Y(n410) );
  INVX2TS U910 ( .A(n2), .Y(n1070) );
  AOI22X1TS U911 ( .A0(n1070), .A1(n758), .B0(n408), .B1(n407), .Y(n409) );
  OAI211XLTS U912 ( .A0(n447), .A1(n411), .B0(n410), .C0(n409), .Y(n2181) );
  AOI22X1TS U913 ( .A0(n413), .A1(\destinationAddressbuffer[0][9] ), .B0(n419), 
        .B1(n412), .Y(n416) );
  INVX2TS U914 ( .A(n5), .Y(n1896) );
  AOI22X1TS U915 ( .A0(n1070), .A1(n739), .B0(n1896), .B1(n414), .Y(n415) );
  OAI211XLTS U916 ( .A0(n436), .A1(n417), .B0(n416), .C0(n415), .Y(n2180) );
  INVX2TS U917 ( .A(n425), .Y(n1913) );
  INVX2TS U918 ( .A(n418), .Y(n419) );
  INVX2TS U919 ( .A(n419), .Y(n1052) );
  INVX2TS U920 ( .A(n1052), .Y(n426) );
  AOI22X1TS U921 ( .A0(n1913), .A1(writeOutbuffer[0]), .B0(n426), .B1(n420), 
        .Y(n423) );
  INVX2TS U922 ( .A(n2), .Y(n1918) );
  INVX2TS U923 ( .A(n5), .Y(n1059) );
  AOI22X1TS U924 ( .A0(n1918), .A1(n551), .B0(n1059), .B1(n421), .Y(n422) );
  OAI211XLTS U925 ( .A0(n436), .A1(n424), .B0(n423), .C0(n422), .Y(n2078) );
  CLKBUFX2TS U926 ( .A(n425), .Y(n1067) );
  INVX2TS U927 ( .A(n1067), .Y(n441) );
  AOI22X1TS U928 ( .A0(n441), .A1(\destinationAddressbuffer[0][5] ), .B0(n426), 
        .B1(destinationAddressIn_WEST[5]), .Y(n429) );
  AOI22X1TS U929 ( .A0(n431), .A1(n679), .B0(n408), .B1(n427), .Y(n428) );
  OAI211XLTS U930 ( .A0(n447), .A1(n430), .B0(n429), .C0(n428), .Y(n2176) );
  AOI22X1TS U931 ( .A0(n441), .A1(\destinationAddressbuffer[0][6] ), .B0(n426), 
        .B1(destinationAddressIn_WEST[6]), .Y(n434) );
  INVX2TS U932 ( .A(n2), .Y(n431) );
  INVX2TS U933 ( .A(n431), .Y(n1035) );
  INVX2TS U934 ( .A(n1035), .Y(n443) );
  AOI22X1TS U935 ( .A0(n443), .A1(n699), .B0(n395), .B1(n432), .Y(n433) );
  OAI211XLTS U936 ( .A0(n436), .A1(n435), .B0(n434), .C0(n433), .Y(n2177) );
  AOI22X1TS U937 ( .A0(n441), .A1(\destinationAddressbuffer[0][4] ), .B0(n1906), .B1(destinationAddressIn_WEST[4]), .Y(n439) );
  INVX2TS U938 ( .A(n2), .Y(n1898) );
  AOI22X1TS U939 ( .A0(n1898), .A1(n667), .B0(n1908), .B1(n437), .Y(n438) );
  OAI211XLTS U940 ( .A0(n1068), .A1(n440), .B0(n439), .C0(n438), .Y(n2175) );
  AOI22X1TS U941 ( .A0(n441), .A1(\destinationAddressbuffer[0][7] ), .B0(n1894), .B1(destinationAddressIn_WEST[7]), .Y(n445) );
  AOI22X1TS U942 ( .A0(n443), .A1(n713), .B0(n1059), .B1(n442), .Y(n444) );
  OAI211XLTS U943 ( .A0(n447), .A1(n446), .B0(n445), .C0(n444), .Y(n2178) );
  INVX2TS U944 ( .A(n1949), .Y(n534) );
  INVX2TS U945 ( .A(n1949), .Y(n531) );
  INVX2TS U946 ( .A(n1943), .Y(n537) );
  NAND2X1TS U947 ( .A(n531), .B(n537), .Y(n535) );
  OAI21XLTS U948 ( .A0(n534), .A1(n1944), .B0(n535), .Y(n509) );
  INVX2TS U949 ( .A(n1940), .Y(n538) );
  INVX2TS U950 ( .A(n1940), .Y(n533) );
  NOR2XLTS U951 ( .A(n535), .B(n533), .Y(n845) );
  CLKBUFX2TS U952 ( .A(n845), .Y(n803) );
  CLKBUFX2TS U953 ( .A(n803), .Y(n822) );
  AOI21X1TS U954 ( .A0(n535), .A1(n538), .B0(n822), .Y(n506) );
  OAI22X1TS U955 ( .A0(n492), .A1(n509), .B0(n449), .B1(n506), .Y(n450) );
  AOI221XLTS U956 ( .A0(n509), .A1(n463), .B0(n451), .B1(n506), .C0(n450), .Y(
        n455) );
  INVX2TS U957 ( .A(n1937), .Y(n452) );
  NAND2X1TS U958 ( .A(n453), .B(n452), .Y(n468) );
  OAI21XLTS U959 ( .A0(n454), .A1(n1949), .B0(n468), .Y(n472) );
  AOI21X1TS U960 ( .A0(n455), .A1(n472), .B0(n1939), .Y(n456) );
  INVX2TS U961 ( .A(reset), .Y(n499) );
  NAND2X1TS U962 ( .A(n499), .B(n1939), .Y(n510) );
  NOR2XLTS U963 ( .A(reset), .B(n457), .Y(n504) );
  INVX2TS U964 ( .A(n1945), .Y(n469) );
  INVX2TS U965 ( .A(n1948), .Y(n459) );
  INVX2TS U966 ( .A(n1941), .Y(n536) );
  AOI22X1TS U967 ( .A0(n459), .A1(n533), .B0(n536), .B1(n458), .Y(n462) );
  INVX2TS U968 ( .A(n461), .Y(n467) );
  INVX2TS U969 ( .A(n482), .Y(n479) );
  AOI21X1TS U970 ( .A0(n534), .A1(n465), .B0(n464), .Y(n478) );
  ADDHXLTS U971 ( .A(n471), .B(n470), .CO(n482), .S(n484) );
  INVX2TS U972 ( .A(n484), .Y(n473) );
  AOI21X1TS U973 ( .A0(n474), .A1(n473), .B0(n472), .Y(n476) );
  OAI22X1TS U974 ( .A0(n474), .A1(n473), .B0(n480), .B1(n479), .Y(n475) );
  AOI21X1TS U975 ( .A0(n483), .A1(n476), .B0(n475), .Y(n477) );
  AOI211X1TS U976 ( .A0(n480), .A1(n479), .B0(n478), .C0(n477), .Y(n481) );
  INVX2TS U977 ( .A(n481), .Y(n485) );
  NAND2X1TS U978 ( .A(n485), .B(n482), .Y(n489) );
  XNOR2X1TS U979 ( .A(n487), .B(n486), .Y(n488) );
  XOR2X1TS U980 ( .A(n489), .B(n488), .Y(n503) );
  INVX2TS U981 ( .A(n503), .Y(n497) );
  INVX2TS U982 ( .A(n1941), .Y(n532) );
  ADDHXLTS U983 ( .A(n453), .B(n490), .CO(n493), .S(n500) );
  XNOR2X1TS U984 ( .A(n1944), .B(n501), .Y(n494) );
  OAI2BB2XLTS U985 ( .B0(n1951), .B1(n510), .A0N(n504), .A1N(n498), .Y(N2624)
         );
  NAND2X1TS U986 ( .A(n499), .B(n1938), .Y(n508) );
  AOI22X1TS U987 ( .A0(n1937), .A1(n510), .B0(n508), .B1(n452), .Y(n1960) );
  INVX2TS U988 ( .A(n506), .Y(n507) );
  OAI22X1TS U989 ( .A0(n538), .A1(n510), .B0(n507), .B1(n508), .Y(n1965) );
  OAI22X1TS U990 ( .A0(n12), .A1(n510), .B0(n509), .B1(n508), .Y(n1966) );
  CLKBUFX2TS U991 ( .A(readIn_SOUTH), .Y(n1652) );
  CLKBUFX2TS U992 ( .A(n1652), .Y(n1594) );
  CLKBUFX2TS U993 ( .A(n1938), .Y(n851) );
  CLKBUFX2TS U994 ( .A(n550), .Y(n634) );
  CLKBUFX2TS U995 ( .A(n634), .Y(n860) );
  CLKBUFX2TS U996 ( .A(readIn_WEST), .Y(n1612) );
  CLKBUFX2TS U997 ( .A(n1612), .Y(n1647) );
  INVX2TS U998 ( .A(n1938), .Y(n527) );
  NAND2X1TS U999 ( .A(n545), .B(n527), .Y(n515) );
  NOR4XLTS U1000 ( .A(readReady), .B(n518), .C(n461), .D(n515), .Y(n619) );
  CLKBUFX2TS U1001 ( .A(n619), .Y(n635) );
  CLKBUFX2TS U1002 ( .A(n635), .Y(n814) );
  CLKBUFX2TS U1003 ( .A(n814), .Y(n572) );
  AOI22X1TS U1004 ( .A0(n1594), .A1(n860), .B0(n1647), .B1(n572), .Y(n548) );
  CLKBUFX2TS U1005 ( .A(readIn_NORTH), .Y(n1627) );
  CLKBUFX2TS U1006 ( .A(n1627), .Y(n1593) );
  CLKBUFX2TS U1007 ( .A(n698), .Y(n633) );
  CLKBUFX2TS U1008 ( .A(n633), .Y(n571) );
  NOR4XLTS U1009 ( .A(selectBit_WEST), .B(n516), .C(n520), .D(n515), .Y(n653)
         );
  CLKBUFX2TS U1010 ( .A(n653), .Y(n784) );
  CLKBUFX2TS U1011 ( .A(n784), .Y(n676) );
  CLKBUFX2TS U1012 ( .A(n676), .Y(n833) );
  AOI22X1TS U1013 ( .A0(n1593), .A1(n571), .B0(readIn_EAST), .B1(n833), .Y(
        n547) );
  NOR3XLTS U1014 ( .A(n518), .B(n517), .C(n461), .Y(n523) );
  NOR3XLTS U1015 ( .A(selectBit_WEST), .B(n521), .C(n520), .Y(n522) );
  OAI31X1TS U1016 ( .A0(n523), .A1(n544), .A2(n522), .B0(n545), .Y(n526) );
  NAND4XLTS U1017 ( .A(n527), .B(n526), .C(n525), .D(n524), .Y(n681) );
  INVX2TS U1018 ( .A(n681), .Y(n528) );
  INVX2TS U1019 ( .A(n528), .Y(n636) );
  INVX2TS U1020 ( .A(n636), .Y(n529) );
  CLKBUFX2TS U1021 ( .A(n1938), .Y(n607) );
  NOR3XLTS U1022 ( .A(n531), .B(n532), .C(n1943), .Y(n726) );
  CLKBUFX2TS U1023 ( .A(n726), .Y(n637) );
  CLKBUFX2TS U1024 ( .A(n637), .Y(n574) );
  NOR3XLTS U1025 ( .A(n534), .B(n1944), .C(n532), .Y(n700) );
  CLKBUFX2TS U1026 ( .A(n700), .Y(n638) );
  CLKBUFX2TS U1027 ( .A(n638), .Y(n573) );
  AOI22X1TS U1028 ( .A0(readOutbuffer[2]), .A1(n574), .B0(readOutbuffer[0]), 
        .B1(n573), .Y(n542) );
  NOR3XLTS U1029 ( .A(n531), .B(n12), .C(n533), .Y(n727) );
  CLKBUFX2TS U1030 ( .A(n727), .Y(n639) );
  CLKBUFX2TS U1031 ( .A(n639), .Y(n576) );
  NOR3XLTS U1032 ( .A(n534), .B(n537), .C(n538), .Y(n701) );
  CLKBUFX2TS U1033 ( .A(n701), .Y(n640) );
  CLKBUFX2TS U1034 ( .A(n640), .Y(n575) );
  AOI22X1TS U1035 ( .A0(readOutbuffer[6]), .A1(n576), .B0(readOutbuffer[4]), 
        .B1(n575), .Y(n541) );
  NOR2XLTS U1036 ( .A(n536), .B(n535), .Y(n728) );
  CLKBUFX2TS U1037 ( .A(n728), .Y(n641) );
  CLKBUFX2TS U1038 ( .A(n641), .Y(n578) );
  NOR3XLTS U1039 ( .A(n537), .B(n536), .C(n1949), .Y(n702) );
  CLKBUFX2TS U1040 ( .A(n702), .Y(n642) );
  CLKBUFX2TS U1041 ( .A(n642), .Y(n577) );
  AOI22X1TS U1042 ( .A0(readOutbuffer[3]), .A1(n578), .B0(readOutbuffer[1]), 
        .B1(n577), .Y(n540) );
  CLKBUFX2TS U1043 ( .A(n845), .Y(n867) );
  NOR3XLTS U1044 ( .A(n1944), .B(n452), .C(n538), .Y(n868) );
  CLKBUFX2TS U1045 ( .A(n868), .Y(n643) );
  CLKBUFX2TS U1046 ( .A(n643), .Y(n579) );
  AOI22X1TS U1047 ( .A0(readOutbuffer[7]), .A1(n867), .B0(readOutbuffer[5]), 
        .B1(n579), .Y(n539) );
  NAND4XLTS U1048 ( .A(n542), .B(n541), .C(n540), .D(n539), .Y(n543) );
  AOI22X1TS U1049 ( .A0(readOut), .A1(n558), .B0(n607), .B1(n543), .Y(n546) );
  CLKBUFX2TS U1050 ( .A(n676), .Y(n756) );
  AOI22X1TS U1051 ( .A0(writeIn_EAST), .A1(n756), .B0(n549), .B1(n572), .Y(
        n561) );
  CLKBUFX2TS U1052 ( .A(n634), .Y(n772) );
  AOI22X1TS U1053 ( .A0(n552), .A1(n571), .B0(n551), .B1(n772), .Y(n560) );
  AOI22X1TS U1054 ( .A0(writeOutbuffer[2]), .A1(n574), .B0(writeOutbuffer[0]), 
        .B1(n573), .Y(n556) );
  AOI22X1TS U1055 ( .A0(writeOutbuffer[6]), .A1(n576), .B0(writeOutbuffer[4]), 
        .B1(n575), .Y(n555) );
  AOI22X1TS U1056 ( .A0(writeOutbuffer[3]), .A1(n578), .B0(writeOutbuffer[1]), 
        .B1(n577), .Y(n554) );
  AOI22X1TS U1057 ( .A0(writeOutbuffer[7]), .A1(n867), .B0(writeOutbuffer[5]), 
        .B1(n579), .Y(n553) );
  NAND4XLTS U1058 ( .A(n556), .B(n555), .C(n554), .D(n553), .Y(n557) );
  AOI22X1TS U1059 ( .A0(writeOut), .A1(n558), .B0(n607), .B1(n557), .Y(n559)
         );
  CLKBUFX2TS U1060 ( .A(requesterAddressIn_NORTH[0]), .Y(n1005) );
  CLKBUFX2TS U1061 ( .A(requesterAddressIn_EAST[0]), .Y(n1034) );
  CLKBUFX2TS U1062 ( .A(n1034), .Y(n1004) );
  CLKBUFX2TS U1063 ( .A(n676), .Y(n596) );
  AOI22X1TS U1064 ( .A0(n1005), .A1(n571), .B0(n1004), .B1(n596), .Y(n570) );
  CLKBUFX2TS U1065 ( .A(requesterAddressIn_SOUTH[0]), .Y(n1037) );
  CLKBUFX2TS U1066 ( .A(n1037), .Y(n1006) );
  CLKBUFX2TS U1067 ( .A(n550), .Y(n666) );
  CLKBUFX2TS U1068 ( .A(requesterAddressIn_WEST[0]), .Y(n932) );
  CLKBUFX2TS U1069 ( .A(n932), .Y(n958) );
  AOI22X1TS U1070 ( .A0(n1006), .A1(n666), .B0(n958), .B1(n572), .Y(n569) );
  INVX2TS U1071 ( .A(n681), .Y(n708) );
  CLKBUFX2TS U1072 ( .A(n607), .Y(n602) );
  AOI22X1TS U1073 ( .A0(\requesterAddressbuffer[2][0] ), .A1(n574), .B0(
        \requesterAddressbuffer[0][0] ), .B1(n573), .Y(n565) );
  AOI22X1TS U1074 ( .A0(\requesterAddressbuffer[6][0] ), .A1(n576), .B0(
        \requesterAddressbuffer[4][0] ), .B1(n575), .Y(n564) );
  AOI22X1TS U1075 ( .A0(\requesterAddressbuffer[3][0] ), .A1(n578), .B0(
        \requesterAddressbuffer[1][0] ), .B1(n577), .Y(n563) );
  CLKBUFX2TS U1076 ( .A(n803), .Y(n760) );
  CLKBUFX2TS U1077 ( .A(n760), .Y(n608) );
  AOI22X1TS U1078 ( .A0(\requesterAddressbuffer[7][0] ), .A1(n608), .B0(
        \requesterAddressbuffer[5][0] ), .B1(n579), .Y(n562) );
  NAND4XLTS U1079 ( .A(n565), .B(n564), .C(n563), .D(n562), .Y(n566) );
  AOI22X1TS U1080 ( .A0(requesterAddressOut[0]), .A1(n708), .B0(n602), .B1(
        n566), .Y(n568) );
  INVX2TS U1081 ( .A(readRequesterAddress[0]), .Y(n956) );
  INVX2TS U1082 ( .A(n956), .Y(n1003) );
  INVX2TS U1083 ( .A(n567), .Y(n603) );
  NAND2X1TS U1084 ( .A(n1003), .B(n603), .Y(n614) );
  CLKBUFX2TS U1085 ( .A(requesterAddressIn_NORTH[1]), .Y(n1012) );
  CLKBUFX2TS U1086 ( .A(requesterAddressIn_EAST[1]), .Y(n1042) );
  CLKBUFX2TS U1087 ( .A(n1042), .Y(n1011) );
  AOI22X1TS U1088 ( .A0(n1012), .A1(n571), .B0(n1011), .B1(n596), .Y(n587) );
  CLKBUFX2TS U1089 ( .A(requesterAddressIn_SOUTH[1]), .Y(n1043) );
  CLKBUFX2TS U1090 ( .A(n1043), .Y(n1013) );
  CLKBUFX2TS U1091 ( .A(n634), .Y(n815) );
  CLKBUFX2TS U1092 ( .A(requesterAddressIn_WEST[1]), .Y(n939) );
  CLKBUFX2TS U1093 ( .A(n939), .Y(n966) );
  AOI22X1TS U1094 ( .A0(n1013), .A1(n815), .B0(n966), .B1(n572), .Y(n586) );
  AOI22X1TS U1095 ( .A0(\requesterAddressbuffer[2][1] ), .A1(n574), .B0(
        \requesterAddressbuffer[0][1] ), .B1(n573), .Y(n583) );
  AOI22X1TS U1096 ( .A0(\requesterAddressbuffer[6][1] ), .A1(n576), .B0(
        \requesterAddressbuffer[4][1] ), .B1(n575), .Y(n582) );
  AOI22X1TS U1097 ( .A0(\requesterAddressbuffer[3][1] ), .A1(n578), .B0(
        \requesterAddressbuffer[1][1] ), .B1(n577), .Y(n581) );
  AOI22X1TS U1098 ( .A0(\requesterAddressbuffer[7][1] ), .A1(n608), .B0(
        \requesterAddressbuffer[5][1] ), .B1(n579), .Y(n580) );
  NAND4XLTS U1099 ( .A(n583), .B(n582), .C(n581), .D(n580), .Y(n584) );
  AOI22X1TS U1100 ( .A0(requesterAddressOut[1]), .A1(n529), .B0(n602), .B1(
        n584), .Y(n585) );
  INVX2TS U1101 ( .A(readRequesterAddress[1]), .Y(n963) );
  INVX2TS U1102 ( .A(n963), .Y(n1669) );
  NAND2X1TS U1103 ( .A(n1669), .B(n603), .Y(n629) );
  CLKBUFX2TS U1104 ( .A(requesterAddressIn_NORTH[2]), .Y(n1020) );
  CLKBUFX2TS U1105 ( .A(n633), .Y(n618) );
  CLKBUFX2TS U1106 ( .A(requesterAddressIn_EAST[2]), .Y(n1047) );
  CLKBUFX2TS U1107 ( .A(n1047), .Y(n1018) );
  AOI22X1TS U1108 ( .A0(n1020), .A1(n618), .B0(n1018), .B1(n596), .Y(n595) );
  CLKBUFX2TS U1109 ( .A(requesterAddressIn_SOUTH[2]), .Y(n1048) );
  CLKBUFX2TS U1110 ( .A(n1048), .Y(n1021) );
  CLKBUFX2TS U1111 ( .A(requesterAddressIn_WEST[2]), .Y(n945) );
  CLKBUFX2TS U1112 ( .A(n945), .Y(n973) );
  AOI22X1TS U1113 ( .A0(n1021), .A1(n666), .B0(n973), .B1(n635), .Y(n594) );
  INVX2TS U1114 ( .A(n681), .Y(n751) );
  CLKBUFX2TS U1115 ( .A(n637), .Y(n620) );
  AOI22X1TS U1116 ( .A0(\requesterAddressbuffer[2][2] ), .A1(n620), .B0(
        \requesterAddressbuffer[0][2] ), .B1(n700), .Y(n591) );
  CLKBUFX2TS U1117 ( .A(n639), .Y(n621) );
  AOI22X1TS U1118 ( .A0(\requesterAddressbuffer[6][2] ), .A1(n621), .B0(
        \requesterAddressbuffer[4][2] ), .B1(n701), .Y(n590) );
  CLKBUFX2TS U1119 ( .A(n641), .Y(n622) );
  AOI22X1TS U1120 ( .A0(\requesterAddressbuffer[3][2] ), .A1(n622), .B0(
        \requesterAddressbuffer[1][2] ), .B1(n702), .Y(n589) );
  CLKBUFX2TS U1121 ( .A(n643), .Y(n623) );
  AOI22X1TS U1122 ( .A0(\requesterAddressbuffer[7][2] ), .A1(n608), .B0(
        \requesterAddressbuffer[5][2] ), .B1(n623), .Y(n588) );
  NAND4XLTS U1123 ( .A(n591), .B(n590), .C(n589), .D(n588), .Y(n592) );
  AOI22X1TS U1124 ( .A0(requesterAddressOut[2]), .A1(n751), .B0(n602), .B1(
        n592), .Y(n593) );
  INVX2TS U1125 ( .A(readRequesterAddress[2]), .Y(n972) );
  INVX2TS U1126 ( .A(n972), .Y(n1678) );
  NAND2X1TS U1127 ( .A(n1678), .B(n603), .Y(n649) );
  CLKBUFX2TS U1128 ( .A(requesterAddressIn_NORTH[3]), .Y(n1029) );
  CLKBUFX2TS U1129 ( .A(requesterAddressIn_EAST[3]), .Y(n1054) );
  CLKBUFX2TS U1130 ( .A(n1054), .Y(n1027) );
  AOI22X1TS U1131 ( .A0(n1029), .A1(n618), .B0(n1027), .B1(n596), .Y(n606) );
  CLKBUFX2TS U1132 ( .A(requesterAddressIn_SOUTH[3]), .Y(n1055) );
  CLKBUFX2TS U1133 ( .A(n1055), .Y(n1030) );
  CLKBUFX2TS U1134 ( .A(requesterAddressIn_WEST[3]), .Y(n951) );
  CLKBUFX2TS U1135 ( .A(n951), .Y(n981) );
  AOI22X1TS U1136 ( .A0(n1030), .A1(n815), .B0(n981), .B1(n619), .Y(n605) );
  AOI22X1TS U1137 ( .A0(\requesterAddressbuffer[2][3] ), .A1(n620), .B0(
        \requesterAddressbuffer[0][3] ), .B1(n700), .Y(n600) );
  AOI22X1TS U1138 ( .A0(\requesterAddressbuffer[6][3] ), .A1(n621), .B0(
        \requesterAddressbuffer[4][3] ), .B1(n701), .Y(n599) );
  AOI22X1TS U1139 ( .A0(\requesterAddressbuffer[3][3] ), .A1(n622), .B0(
        \requesterAddressbuffer[1][3] ), .B1(n702), .Y(n598) );
  CLKBUFX2TS U1140 ( .A(n760), .Y(n654) );
  AOI22X1TS U1141 ( .A0(\requesterAddressbuffer[7][3] ), .A1(n654), .B0(
        \requesterAddressbuffer[5][3] ), .B1(n623), .Y(n597) );
  NAND4XLTS U1142 ( .A(n600), .B(n599), .C(n598), .D(n597), .Y(n601) );
  AOI22X1TS U1143 ( .A0(requesterAddressOut[3]), .A1(n751), .B0(n602), .B1(
        n601), .Y(n604) );
  INVX2TS U1144 ( .A(readRequesterAddress[3]), .Y(n980) );
  INVX2TS U1145 ( .A(n980), .Y(n1685) );
  NAND2X1TS U1146 ( .A(n1685), .B(n603), .Y(n661) );
  CLKBUFX2TS U1147 ( .A(destinationAddressIn_NORTH[0]), .Y(n1693) );
  CLKBUFX2TS U1148 ( .A(destinationAddressIn_EAST[0]), .Y(n1842) );
  CLKBUFX2TS U1149 ( .A(n1842), .Y(n1722) );
  AOI22X1TS U1150 ( .A0(n1693), .A1(n618), .B0(n1722), .B1(n784), .Y(n617) );
  CLKBUFX2TS U1151 ( .A(destinationAddressIn_WEST[0]), .Y(n1723) );
  CLKBUFX2TS U1152 ( .A(n1723), .Y(n1786) );
  AOI22X1TS U1153 ( .A0(destinationAddressIn_SOUTH[0]), .A1(n666), .B0(n1786), 
        .B1(n619), .Y(n616) );
  CLKBUFX2TS U1154 ( .A(n607), .Y(n660) );
  AOI22X1TS U1155 ( .A0(\destinationAddressbuffer[2][0] ), .A1(n620), .B0(
        \destinationAddressbuffer[0][0] ), .B1(n638), .Y(n612) );
  AOI22X1TS U1156 ( .A0(\destinationAddressbuffer[6][0] ), .A1(n621), .B0(
        \destinationAddressbuffer[4][0] ), .B1(n640), .Y(n611) );
  AOI22X1TS U1157 ( .A0(\destinationAddressbuffer[3][0] ), .A1(n622), .B0(
        \destinationAddressbuffer[1][0] ), .B1(n642), .Y(n610) );
  AOI22X1TS U1158 ( .A0(\destinationAddressbuffer[7][0] ), .A1(n608), .B0(
        \destinationAddressbuffer[5][0] ), .B1(n623), .Y(n609) );
  NAND4XLTS U1159 ( .A(n612), .B(n611), .C(n610), .D(n609), .Y(n613) );
  AOI22X1TS U1160 ( .A0(destinationAddressOut[0]), .A1(n751), .B0(n660), .B1(
        n613), .Y(n615) );
  CLKBUFX2TS U1161 ( .A(destinationAddressIn_NORTH[1]), .Y(n1701) );
  CLKBUFX2TS U1162 ( .A(destinationAddressIn_EAST[1]), .Y(n1852) );
  CLKBUFX2TS U1163 ( .A(n1852), .Y(n1729) );
  AOI22X1TS U1164 ( .A0(n1701), .A1(n618), .B0(n1729), .B1(n653), .Y(n632) );
  CLKBUFX2TS U1165 ( .A(destinationAddressIn_WEST[1]), .Y(n1731) );
  CLKBUFX2TS U1166 ( .A(n1731), .Y(n1793) );
  AOI22X1TS U1167 ( .A0(destinationAddressIn_SOUTH[1]), .A1(n815), .B0(n1793), 
        .B1(n619), .Y(n631) );
  AOI22X1TS U1168 ( .A0(\destinationAddressbuffer[2][1] ), .A1(n620), .B0(
        \destinationAddressbuffer[0][1] ), .B1(n638), .Y(n627) );
  AOI22X1TS U1169 ( .A0(\destinationAddressbuffer[6][1] ), .A1(n621), .B0(
        \destinationAddressbuffer[4][1] ), .B1(n640), .Y(n626) );
  AOI22X1TS U1170 ( .A0(\destinationAddressbuffer[3][1] ), .A1(n622), .B0(
        \destinationAddressbuffer[1][1] ), .B1(n642), .Y(n625) );
  AOI22X1TS U1171 ( .A0(\destinationAddressbuffer[7][1] ), .A1(n654), .B0(
        \destinationAddressbuffer[5][1] ), .B1(n623), .Y(n624) );
  NAND4XLTS U1172 ( .A(n627), .B(n626), .C(n625), .D(n624), .Y(n628) );
  AOI22X1TS U1173 ( .A0(destinationAddressOut[1]), .A1(n708), .B0(n660), .B1(
        n628), .Y(n630) );
  CLKBUFX2TS U1174 ( .A(destinationAddressIn_NORTH[2]), .Y(n1709) );
  CLKBUFX2TS U1175 ( .A(n633), .Y(n680) );
  CLKBUFX2TS U1176 ( .A(destinationAddressIn_EAST[2]), .Y(n1864) );
  CLKBUFX2TS U1177 ( .A(n1864), .Y(n1740) );
  AOI22X1TS U1178 ( .A0(n1709), .A1(n680), .B0(n1740), .B1(n653), .Y(n652) );
  CLKBUFX2TS U1179 ( .A(n634), .Y(n796) );
  CLKBUFX2TS U1180 ( .A(destinationAddressIn_WEST[2]), .Y(n1742) );
  CLKBUFX2TS U1181 ( .A(n1742), .Y(n1800) );
  CLKBUFX2TS U1182 ( .A(n635), .Y(n677) );
  AOI22X1TS U1183 ( .A0(destinationAddressIn_SOUTH[2]), .A1(n796), .B0(n1800), 
        .B1(n677), .Y(n651) );
  INVX2TS U1184 ( .A(n636), .Y(n875) );
  CLKBUFX2TS U1185 ( .A(n637), .Y(n683) );
  CLKBUFX2TS U1186 ( .A(n638), .Y(n682) );
  AOI22X1TS U1187 ( .A0(\destinationAddressbuffer[2][2] ), .A1(n683), .B0(
        \destinationAddressbuffer[0][2] ), .B1(n682), .Y(n647) );
  CLKBUFX2TS U1188 ( .A(n639), .Y(n685) );
  CLKBUFX2TS U1189 ( .A(n640), .Y(n684) );
  AOI22X1TS U1190 ( .A0(\destinationAddressbuffer[6][2] ), .A1(n685), .B0(
        \destinationAddressbuffer[4][2] ), .B1(n684), .Y(n646) );
  CLKBUFX2TS U1191 ( .A(n641), .Y(n687) );
  CLKBUFX2TS U1192 ( .A(n642), .Y(n686) );
  AOI22X1TS U1193 ( .A0(\destinationAddressbuffer[3][2] ), .A1(n687), .B0(
        \destinationAddressbuffer[1][2] ), .B1(n686), .Y(n645) );
  CLKBUFX2TS U1194 ( .A(n643), .Y(n688) );
  AOI22X1TS U1195 ( .A0(\destinationAddressbuffer[7][2] ), .A1(n654), .B0(
        \destinationAddressbuffer[5][2] ), .B1(n688), .Y(n644) );
  NAND4XLTS U1196 ( .A(n647), .B(n646), .C(n645), .D(n644), .Y(n648) );
  AOI22X1TS U1197 ( .A0(destinationAddressOut[2]), .A1(n875), .B0(n660), .B1(
        n648), .Y(n650) );
  CLKBUFX2TS U1198 ( .A(destinationAddressIn_NORTH[3]), .Y(n1717) );
  CLKBUFX2TS U1199 ( .A(destinationAddressIn_EAST[3]), .Y(n1876) );
  CLKBUFX2TS U1200 ( .A(n1876), .Y(n1751) );
  AOI22X1TS U1201 ( .A0(n1717), .A1(n680), .B0(n1751), .B1(n653), .Y(n664) );
  CLKBUFX2TS U1202 ( .A(destinationAddressIn_WEST[3]), .Y(n1752) );
  CLKBUFX2TS U1203 ( .A(n1752), .Y(n1808) );
  AOI22X1TS U1204 ( .A0(destinationAddressIn_SOUTH[3]), .A1(n796), .B0(n1808), 
        .B1(n677), .Y(n663) );
  AOI22X1TS U1205 ( .A0(\destinationAddressbuffer[2][3] ), .A1(n683), .B0(
        \destinationAddressbuffer[0][3] ), .B1(n682), .Y(n658) );
  AOI22X1TS U1206 ( .A0(\destinationAddressbuffer[6][3] ), .A1(n685), .B0(
        \destinationAddressbuffer[4][3] ), .B1(n684), .Y(n657) );
  AOI22X1TS U1207 ( .A0(\destinationAddressbuffer[3][3] ), .A1(n687), .B0(
        \destinationAddressbuffer[1][3] ), .B1(n686), .Y(n656) );
  AOI22X1TS U1208 ( .A0(\destinationAddressbuffer[7][3] ), .A1(n654), .B0(
        \destinationAddressbuffer[5][3] ), .B1(n688), .Y(n655) );
  NAND4XLTS U1209 ( .A(n658), .B(n657), .C(n656), .D(n655), .Y(n659) );
  AOI22X1TS U1210 ( .A0(destinationAddressOut[3]), .A1(n529), .B0(n660), .B1(
        n659), .Y(n662) );
  AOI22X1TS U1211 ( .A0(destinationAddressIn_EAST[4]), .A1(n756), .B0(n665), 
        .B1(n677), .Y(n675) );
  AOI22X1TS U1212 ( .A0(destinationAddressIn_NORTH[4]), .A1(n680), .B0(n667), 
        .B1(n666), .Y(n674) );
  INVX2TS U1213 ( .A(n1939), .Y(n775) );
  CLKBUFX2TS U1214 ( .A(n775), .Y(n874) );
  AOI22X1TS U1215 ( .A0(\destinationAddressbuffer[2][4] ), .A1(n683), .B0(
        \destinationAddressbuffer[0][4] ), .B1(n682), .Y(n671) );
  AOI22X1TS U1216 ( .A0(\destinationAddressbuffer[6][4] ), .A1(n685), .B0(
        \destinationAddressbuffer[4][4] ), .B1(n684), .Y(n670) );
  AOI22X1TS U1217 ( .A0(\destinationAddressbuffer[3][4] ), .A1(n687), .B0(
        \destinationAddressbuffer[1][4] ), .B1(n686), .Y(n669) );
  CLKBUFX2TS U1218 ( .A(n760), .Y(n714) );
  AOI22X1TS U1219 ( .A0(\destinationAddressbuffer[7][4] ), .A1(n714), .B0(
        \destinationAddressbuffer[5][4] ), .B1(n688), .Y(n668) );
  NAND4XLTS U1220 ( .A(n671), .B(n670), .C(n669), .D(n668), .Y(n672) );
  AOI22X1TS U1221 ( .A0(destinationAddressOut[4]), .A1(n708), .B0(n874), .B1(
        n672), .Y(n673) );
  CLKBUFX2TS U1222 ( .A(n676), .Y(n771) );
  AOI22X1TS U1223 ( .A0(destinationAddressIn_EAST[5]), .A1(n771), .B0(n678), 
        .B1(n677), .Y(n696) );
  CLKBUFX2TS U1224 ( .A(n550), .Y(n757) );
  AOI22X1TS U1225 ( .A0(destinationAddressIn_NORTH[5]), .A1(n680), .B0(n679), 
        .B1(n757), .Y(n695) );
  INVX2TS U1226 ( .A(n681), .Y(n840) );
  AOI22X1TS U1227 ( .A0(\destinationAddressbuffer[2][5] ), .A1(n683), .B0(
        \destinationAddressbuffer[0][5] ), .B1(n682), .Y(n692) );
  AOI22X1TS U1228 ( .A0(\destinationAddressbuffer[6][5] ), .A1(n685), .B0(
        \destinationAddressbuffer[4][5] ), .B1(n684), .Y(n691) );
  AOI22X1TS U1229 ( .A0(\destinationAddressbuffer[3][5] ), .A1(n687), .B0(
        \destinationAddressbuffer[1][5] ), .B1(n686), .Y(n690) );
  AOI22X1TS U1230 ( .A0(\destinationAddressbuffer[7][5] ), .A1(n714), .B0(
        \destinationAddressbuffer[5][5] ), .B1(n688), .Y(n689) );
  NAND4XLTS U1231 ( .A(n692), .B(n691), .C(n690), .D(n689), .Y(n693) );
  AOI22X1TS U1232 ( .A0(destinationAddressOut[5]), .A1(n840), .B0(n874), .B1(
        n693), .Y(n694) );
  CLKBUFX2TS U1233 ( .A(n814), .Y(n737) );
  AOI22X1TS U1234 ( .A0(destinationAddressIn_EAST[6]), .A1(n771), .B0(n697), 
        .B1(n737), .Y(n711) );
  CLKBUFX2TS U1235 ( .A(n698), .Y(n740) );
  AOI22X1TS U1236 ( .A0(destinationAddressIn_NORTH[6]), .A1(n740), .B0(n699), 
        .B1(n757), .Y(n710) );
  CLKBUFX2TS U1237 ( .A(n700), .Y(n816) );
  CLKBUFX2TS U1238 ( .A(n816), .Y(n742) );
  AOI22X1TS U1239 ( .A0(\destinationAddressbuffer[2][6] ), .A1(n726), .B0(
        \destinationAddressbuffer[0][6] ), .B1(n742), .Y(n706) );
  CLKBUFX2TS U1240 ( .A(n701), .Y(n818) );
  CLKBUFX2TS U1241 ( .A(n818), .Y(n743) );
  AOI22X1TS U1242 ( .A0(\destinationAddressbuffer[6][6] ), .A1(n727), .B0(
        \destinationAddressbuffer[4][6] ), .B1(n743), .Y(n705) );
  CLKBUFX2TS U1243 ( .A(n702), .Y(n820) );
  CLKBUFX2TS U1244 ( .A(n820), .Y(n744) );
  AOI22X1TS U1245 ( .A0(\destinationAddressbuffer[3][6] ), .A1(n728), .B0(
        \destinationAddressbuffer[1][6] ), .B1(n744), .Y(n704) );
  CLKBUFX2TS U1246 ( .A(n868), .Y(n834) );
  CLKBUFX2TS U1247 ( .A(n834), .Y(n745) );
  AOI22X1TS U1248 ( .A0(\destinationAddressbuffer[7][6] ), .A1(n714), .B0(
        \destinationAddressbuffer[5][6] ), .B1(n745), .Y(n703) );
  NAND4XLTS U1249 ( .A(n706), .B(n705), .C(n704), .D(n703), .Y(n707) );
  AOI22X1TS U1250 ( .A0(destinationAddressOut[6]), .A1(n708), .B0(n874), .B1(
        n707), .Y(n709) );
  AOI22X1TS U1251 ( .A0(destinationAddressIn_EAST[7]), .A1(n833), .B0(n712), 
        .B1(n737), .Y(n722) );
  AOI22X1TS U1252 ( .A0(destinationAddressIn_NORTH[7]), .A1(n740), .B0(n713), 
        .B1(n772), .Y(n721) );
  CLKBUFX2TS U1253 ( .A(n775), .Y(n766) );
  AOI22X1TS U1254 ( .A0(\destinationAddressbuffer[2][7] ), .A1(n726), .B0(
        \destinationAddressbuffer[0][7] ), .B1(n742), .Y(n718) );
  AOI22X1TS U1255 ( .A0(\destinationAddressbuffer[6][7] ), .A1(n727), .B0(
        \destinationAddressbuffer[4][7] ), .B1(n743), .Y(n717) );
  AOI22X1TS U1256 ( .A0(\destinationAddressbuffer[3][7] ), .A1(n728), .B0(
        \destinationAddressbuffer[1][7] ), .B1(n744), .Y(n716) );
  AOI22X1TS U1257 ( .A0(\destinationAddressbuffer[7][7] ), .A1(n714), .B0(
        \destinationAddressbuffer[5][7] ), .B1(n745), .Y(n715) );
  NAND4XLTS U1258 ( .A(n718), .B(n717), .C(n716), .D(n715), .Y(n719) );
  AOI22X1TS U1259 ( .A0(destinationAddressOut[7]), .A1(n528), .B0(n766), .B1(
        n719), .Y(n720) );
  AOI22X1TS U1260 ( .A0(destinationAddressIn_EAST[8]), .A1(n756), .B0(n723), 
        .B1(n737), .Y(n736) );
  AOI22X1TS U1261 ( .A0(n725), .A1(n740), .B0(n724), .B1(n757), .Y(n735) );
  CLKBUFX2TS U1262 ( .A(n726), .Y(n817) );
  AOI22X1TS U1263 ( .A0(\destinationAddressbuffer[2][8] ), .A1(n817), .B0(
        \destinationAddressbuffer[0][8] ), .B1(n742), .Y(n732) );
  CLKBUFX2TS U1264 ( .A(n727), .Y(n819) );
  AOI22X1TS U1265 ( .A0(\destinationAddressbuffer[6][8] ), .A1(n819), .B0(
        \destinationAddressbuffer[4][8] ), .B1(n743), .Y(n731) );
  CLKBUFX2TS U1266 ( .A(n728), .Y(n821) );
  AOI22X1TS U1267 ( .A0(\destinationAddressbuffer[3][8] ), .A1(n821), .B0(
        \destinationAddressbuffer[1][8] ), .B1(n744), .Y(n730) );
  AOI22X1TS U1268 ( .A0(\destinationAddressbuffer[7][8] ), .A1(n822), .B0(
        \destinationAddressbuffer[5][8] ), .B1(n745), .Y(n729) );
  NAND4XLTS U1269 ( .A(n732), .B(n731), .C(n730), .D(n729), .Y(n733) );
  AOI22X1TS U1270 ( .A0(destinationAddressOut[8]), .A1(n875), .B0(n766), .B1(
        n733), .Y(n734) );
  AOI22X1TS U1271 ( .A0(destinationAddressIn_EAST[9]), .A1(n771), .B0(n738), 
        .B1(n737), .Y(n754) );
  AOI22X1TS U1272 ( .A0(n741), .A1(n740), .B0(n739), .B1(n772), .Y(n753) );
  AOI22X1TS U1273 ( .A0(\destinationAddressbuffer[2][9] ), .A1(n817), .B0(
        \destinationAddressbuffer[0][9] ), .B1(n742), .Y(n749) );
  AOI22X1TS U1274 ( .A0(\destinationAddressbuffer[6][9] ), .A1(n819), .B0(
        \destinationAddressbuffer[4][9] ), .B1(n743), .Y(n748) );
  AOI22X1TS U1275 ( .A0(\destinationAddressbuffer[3][9] ), .A1(n821), .B0(
        \destinationAddressbuffer[1][9] ), .B1(n744), .Y(n747) );
  AOI22X1TS U1276 ( .A0(\destinationAddressbuffer[7][9] ), .A1(n822), .B0(
        \destinationAddressbuffer[5][9] ), .B1(n745), .Y(n746) );
  NAND4XLTS U1277 ( .A(n749), .B(n748), .C(n747), .D(n746), .Y(n750) );
  AOI22X1TS U1278 ( .A0(destinationAddressOut[9]), .A1(n751), .B0(n766), .B1(
        n750), .Y(n752) );
  CLKBUFX2TS U1279 ( .A(n814), .Y(n795) );
  AOI22X1TS U1280 ( .A0(destinationAddressIn_EAST[10]), .A1(n756), .B0(n755), 
        .B1(n795), .Y(n769) );
  CLKBUFX2TS U1281 ( .A(n698), .Y(n794) );
  AOI22X1TS U1282 ( .A0(n759), .A1(n794), .B0(n758), .B1(n757), .Y(n768) );
  CLKBUFX2TS U1283 ( .A(n817), .Y(n797) );
  CLKBUFX2TS U1284 ( .A(n816), .Y(n798) );
  AOI22X1TS U1285 ( .A0(\destinationAddressbuffer[2][10] ), .A1(n797), .B0(
        \destinationAddressbuffer[0][10] ), .B1(n798), .Y(n764) );
  CLKBUFX2TS U1286 ( .A(n819), .Y(n799) );
  CLKBUFX2TS U1287 ( .A(n818), .Y(n800) );
  AOI22X1TS U1288 ( .A0(\destinationAddressbuffer[6][10] ), .A1(n799), .B0(
        \destinationAddressbuffer[4][10] ), .B1(n800), .Y(n763) );
  CLKBUFX2TS U1289 ( .A(n821), .Y(n801) );
  CLKBUFX2TS U1290 ( .A(n820), .Y(n802) );
  AOI22X1TS U1291 ( .A0(\destinationAddressbuffer[3][10] ), .A1(n801), .B0(
        \destinationAddressbuffer[1][10] ), .B1(n802), .Y(n762) );
  CLKBUFX2TS U1292 ( .A(n834), .Y(n804) );
  AOI22X1TS U1293 ( .A0(\destinationAddressbuffer[7][10] ), .A1(n760), .B0(
        \destinationAddressbuffer[5][10] ), .B1(n804), .Y(n761) );
  NAND4XLTS U1294 ( .A(n764), .B(n763), .C(n762), .D(n761), .Y(n765) );
  AOI22X1TS U1295 ( .A0(destinationAddressOut[10]), .A1(n875), .B0(n766), .B1(
        n765), .Y(n767) );
  AOI22X1TS U1296 ( .A0(destinationAddressIn_EAST[11]), .A1(n771), .B0(n770), 
        .B1(n795), .Y(n783) );
  AOI22X1TS U1297 ( .A0(n774), .A1(n794), .B0(n773), .B1(n772), .Y(n782) );
  CLKBUFX2TS U1298 ( .A(n775), .Y(n828) );
  AOI22X1TS U1299 ( .A0(\destinationAddressbuffer[2][11] ), .A1(n797), .B0(
        \destinationAddressbuffer[0][11] ), .B1(n798), .Y(n779) );
  AOI22X1TS U1300 ( .A0(\destinationAddressbuffer[6][11] ), .A1(n799), .B0(
        \destinationAddressbuffer[4][11] ), .B1(n800), .Y(n778) );
  AOI22X1TS U1301 ( .A0(\destinationAddressbuffer[3][11] ), .A1(n801), .B0(
        \destinationAddressbuffer[1][11] ), .B1(n802), .Y(n777) );
  AOI22X1TS U1302 ( .A0(\destinationAddressbuffer[7][11] ), .A1(n803), .B0(
        \destinationAddressbuffer[5][11] ), .B1(n804), .Y(n776) );
  NAND4XLTS U1303 ( .A(n779), .B(n778), .C(n777), .D(n776), .Y(n780) );
  AOI22X1TS U1304 ( .A0(destinationAddressOut[11]), .A1(n528), .B0(n828), .B1(
        n780), .Y(n781) );
  CLKBUFX2TS U1305 ( .A(dataIn_NORTH[0]), .Y(n1087) );
  CLKBUFX2TS U1306 ( .A(dataIn_EAST[0]), .Y(n1470) );
  CLKBUFX2TS U1307 ( .A(n1470), .Y(n1346) );
  CLKBUFX2TS U1308 ( .A(n784), .Y(n857) );
  AOI22X1TS U1309 ( .A0(n1087), .A1(n794), .B0(n1346), .B1(n857), .Y(n793) );
  CLKBUFX2TS U1310 ( .A(dataIn_WEST[0]), .Y(n1520) );
  CLKBUFX2TS U1311 ( .A(n1520), .Y(n1408) );
  AOI22X1TS U1312 ( .A0(dataIn_SOUTH[0]), .A1(n796), .B0(n1408), .B1(n795), 
        .Y(n792) );
  AOI22X1TS U1313 ( .A0(\dataoutbuffer[0][0] ), .A1(n798), .B0(
        \dataoutbuffer[2][0] ), .B1(n797), .Y(n788) );
  AOI22X1TS U1314 ( .A0(\dataoutbuffer[4][0] ), .A1(n800), .B0(
        \dataoutbuffer[6][0] ), .B1(n799), .Y(n787) );
  AOI22X1TS U1315 ( .A0(\dataoutbuffer[1][0] ), .A1(n802), .B0(
        \dataoutbuffer[3][0] ), .B1(n801), .Y(n786) );
  AOI22X1TS U1316 ( .A0(\dataoutbuffer[5][0] ), .A1(n804), .B0(
        \dataoutbuffer[7][0] ), .B1(n867), .Y(n785) );
  NAND4XLTS U1317 ( .A(n788), .B(n787), .C(n786), .D(n785), .Y(n789) );
  AOI22X1TS U1318 ( .A0(dataOut[0]), .A1(n529), .B0(n828), .B1(n789), .Y(n791)
         );
  INVX2TS U1319 ( .A(cacheDataOut[0]), .Y(n1086) );
  INVX2TS U1320 ( .A(n567), .Y(n852) );
  NAND2X1TS U1321 ( .A(cacheDataOut[0]), .B(n852), .Y(n790) );
  CLKBUFX2TS U1322 ( .A(dataIn_NORTH[1]), .Y(n1093) );
  CLKBUFX2TS U1323 ( .A(dataIn_EAST[1]), .Y(n1478) );
  CLKBUFX2TS U1324 ( .A(n1478), .Y(n1351) );
  AOI22X1TS U1325 ( .A0(n1093), .A1(n794), .B0(n1351), .B1(n833), .Y(n813) );
  CLKBUFX2TS U1326 ( .A(dataIn_WEST[1]), .Y(n1531) );
  CLKBUFX2TS U1327 ( .A(n1531), .Y(n1413) );
  AOI22X1TS U1328 ( .A0(dataIn_SOUTH[1]), .A1(n796), .B0(n1413), .B1(n795), 
        .Y(n812) );
  AOI22X1TS U1329 ( .A0(\dataoutbuffer[0][1] ), .A1(n798), .B0(
        \dataoutbuffer[2][1] ), .B1(n797), .Y(n808) );
  AOI22X1TS U1330 ( .A0(\dataoutbuffer[4][1] ), .A1(n800), .B0(
        \dataoutbuffer[6][1] ), .B1(n799), .Y(n807) );
  AOI22X1TS U1331 ( .A0(\dataoutbuffer[1][1] ), .A1(n802), .B0(
        \dataoutbuffer[3][1] ), .B1(n801), .Y(n806) );
  AOI22X1TS U1332 ( .A0(\dataoutbuffer[5][1] ), .A1(n804), .B0(
        \dataoutbuffer[7][1] ), .B1(n803), .Y(n805) );
  NAND4XLTS U1333 ( .A(n808), .B(n807), .C(n806), .D(n805), .Y(n809) );
  AOI22X1TS U1334 ( .A0(dataOut[1]), .A1(n840), .B0(n828), .B1(n809), .Y(n811)
         );
  INVX2TS U1335 ( .A(cacheDataOut[1]), .Y(n1091) );
  INVX2TS U1336 ( .A(n567), .Y(n876) );
  NAND2X1TS U1337 ( .A(cacheDataOut[1]), .B(n876), .Y(n810) );
  CLKBUFX2TS U1338 ( .A(dataIn_NORTH[2]), .Y(n1100) );
  CLKBUFX2TS U1339 ( .A(n698), .Y(n858) );
  CLKBUFX2TS U1340 ( .A(dataIn_EAST[2]), .Y(n1487) );
  CLKBUFX2TS U1341 ( .A(n1487), .Y(n1358) );
  AOI22X1TS U1342 ( .A0(n1100), .A1(n858), .B0(n1358), .B1(n857), .Y(n832) );
  CLKBUFX2TS U1343 ( .A(dataIn_WEST[2]), .Y(n1540) );
  CLKBUFX2TS U1344 ( .A(n1540), .Y(n1421) );
  CLKBUFX2TS U1345 ( .A(n814), .Y(n859) );
  AOI22X1TS U1346 ( .A0(dataIn_SOUTH[2]), .A1(n815), .B0(n1421), .B1(n859), 
        .Y(n831) );
  CLKBUFX2TS U1347 ( .A(n816), .Y(n862) );
  CLKBUFX2TS U1348 ( .A(n817), .Y(n861) );
  AOI22X1TS U1349 ( .A0(\dataoutbuffer[0][2] ), .A1(n862), .B0(
        \dataoutbuffer[2][2] ), .B1(n861), .Y(n826) );
  CLKBUFX2TS U1350 ( .A(n818), .Y(n864) );
  CLKBUFX2TS U1351 ( .A(n819), .Y(n863) );
  AOI22X1TS U1352 ( .A0(\dataoutbuffer[4][2] ), .A1(n864), .B0(
        \dataoutbuffer[6][2] ), .B1(n863), .Y(n825) );
  CLKBUFX2TS U1353 ( .A(n820), .Y(n866) );
  CLKBUFX2TS U1354 ( .A(n821), .Y(n865) );
  AOI22X1TS U1355 ( .A0(\dataoutbuffer[1][2] ), .A1(n866), .B0(
        \dataoutbuffer[3][2] ), .B1(n865), .Y(n824) );
  AOI22X1TS U1356 ( .A0(\dataoutbuffer[5][2] ), .A1(n834), .B0(
        \dataoutbuffer[7][2] ), .B1(n822), .Y(n823) );
  NAND4XLTS U1357 ( .A(n826), .B(n825), .C(n824), .D(n823), .Y(n827) );
  AOI22X1TS U1358 ( .A0(dataOut[2]), .A1(n840), .B0(n828), .B1(n827), .Y(n830)
         );
  INVX2TS U1359 ( .A(cacheDataOut[2]), .Y(n1098) );
  NAND2X1TS U1360 ( .A(cacheDataOut[2]), .B(n852), .Y(n829) );
  CLKBUFX2TS U1361 ( .A(dataIn_NORTH[3]), .Y(n1106) );
  CLKBUFX2TS U1362 ( .A(dataIn_EAST[3]), .Y(n1496) );
  CLKBUFX2TS U1363 ( .A(n1496), .Y(n1365) );
  AOI22X1TS U1364 ( .A0(n1106), .A1(n858), .B0(n1365), .B1(n833), .Y(n844) );
  CLKBUFX2TS U1365 ( .A(dataIn_WEST[3]), .Y(n1547) );
  CLKBUFX2TS U1366 ( .A(n1547), .Y(n1426) );
  AOI22X1TS U1367 ( .A0(dataIn_SOUTH[3]), .A1(n860), .B0(n1426), .B1(n859), 
        .Y(n843) );
  AOI22X1TS U1368 ( .A0(\dataoutbuffer[0][3] ), .A1(n862), .B0(
        \dataoutbuffer[2][3] ), .B1(n861), .Y(n838) );
  AOI22X1TS U1369 ( .A0(\dataoutbuffer[4][3] ), .A1(n864), .B0(
        \dataoutbuffer[6][3] ), .B1(n863), .Y(n837) );
  AOI22X1TS U1370 ( .A0(\dataoutbuffer[1][3] ), .A1(n866), .B0(
        \dataoutbuffer[3][3] ), .B1(n865), .Y(n836) );
  AOI22X1TS U1371 ( .A0(\dataoutbuffer[5][3] ), .A1(n834), .B0(
        \dataoutbuffer[7][3] ), .B1(n845), .Y(n835) );
  NAND4XLTS U1372 ( .A(n838), .B(n837), .C(n836), .D(n835), .Y(n839) );
  AOI22X1TS U1373 ( .A0(dataOut[3]), .A1(n840), .B0(n851), .B1(n839), .Y(n842)
         );
  INVX2TS U1374 ( .A(cacheDataOut[3]), .Y(n1105) );
  NAND2X1TS U1375 ( .A(cacheDataOut[3]), .B(n876), .Y(n841) );
  CLKBUFX2TS U1376 ( .A(dataIn_NORTH[4]), .Y(n1112) );
  CLKBUFX2TS U1377 ( .A(dataIn_EAST[4]), .Y(n1504) );
  CLKBUFX2TS U1378 ( .A(n1504), .Y(n1370) );
  AOI22X1TS U1379 ( .A0(n1112), .A1(n858), .B0(n1370), .B1(n857), .Y(n856) );
  CLKBUFX2TS U1380 ( .A(dataIn_WEST[4]), .Y(n1554) );
  CLKBUFX2TS U1381 ( .A(n1554), .Y(n1430) );
  AOI22X1TS U1382 ( .A0(dataIn_SOUTH[4]), .A1(n860), .B0(n1430), .B1(n859), 
        .Y(n855) );
  AOI22X1TS U1383 ( .A0(\dataoutbuffer[0][4] ), .A1(n862), .B0(
        \dataoutbuffer[2][4] ), .B1(n861), .Y(n849) );
  AOI22X1TS U1384 ( .A0(\dataoutbuffer[4][4] ), .A1(n864), .B0(
        \dataoutbuffer[6][4] ), .B1(n863), .Y(n848) );
  AOI22X1TS U1385 ( .A0(\dataoutbuffer[1][4] ), .A1(n866), .B0(
        \dataoutbuffer[3][4] ), .B1(n865), .Y(n847) );
  AOI22X1TS U1386 ( .A0(\dataoutbuffer[5][4] ), .A1(n868), .B0(
        \dataoutbuffer[7][4] ), .B1(n845), .Y(n846) );
  NAND4XLTS U1387 ( .A(n849), .B(n848), .C(n847), .D(n846), .Y(n850) );
  AOI22X1TS U1388 ( .A0(dataOut[4]), .A1(n529), .B0(n851), .B1(n850), .Y(n854)
         );
  INVX2TS U1389 ( .A(cacheDataOut[4]), .Y(n1111) );
  NAND2X1TS U1390 ( .A(cacheDataOut[4]), .B(n852), .Y(n853) );
  CLKBUFX2TS U1391 ( .A(dataIn_NORTH[5]), .Y(n1342) );
  CLKBUFX2TS U1392 ( .A(dataIn_EAST[5]), .Y(n1512) );
  CLKBUFX2TS U1393 ( .A(n1512), .Y(n1375) );
  AOI22X1TS U1394 ( .A0(n1342), .A1(n858), .B0(n1375), .B1(n857), .Y(n880) );
  CLKBUFX2TS U1395 ( .A(dataIn_WEST[5]), .Y(n1563) );
  CLKBUFX2TS U1396 ( .A(n1563), .Y(n1435) );
  AOI22X1TS U1397 ( .A0(dataIn_SOUTH[5]), .A1(n860), .B0(n1435), .B1(n859), 
        .Y(n879) );
  AOI22X1TS U1398 ( .A0(\dataoutbuffer[0][5] ), .A1(n862), .B0(
        \dataoutbuffer[2][5] ), .B1(n861), .Y(n872) );
  AOI22X1TS U1399 ( .A0(\dataoutbuffer[4][5] ), .A1(n864), .B0(
        \dataoutbuffer[6][5] ), .B1(n863), .Y(n871) );
  AOI22X1TS U1400 ( .A0(\dataoutbuffer[1][5] ), .A1(n866), .B0(
        \dataoutbuffer[3][5] ), .B1(n865), .Y(n870) );
  AOI22X1TS U1401 ( .A0(\dataoutbuffer[5][5] ), .A1(n868), .B0(
        \dataoutbuffer[7][5] ), .B1(n867), .Y(n869) );
  NAND4XLTS U1402 ( .A(n872), .B(n871), .C(n870), .D(n869), .Y(n873) );
  AOI22X1TS U1403 ( .A0(dataOut[5]), .A1(n875), .B0(n874), .B1(n873), .Y(n878)
         );
  INVX2TS U1404 ( .A(cacheDataOut[5]), .Y(n1340) );
  NAND2X1TS U1405 ( .A(cacheDataOut[5]), .B(n876), .Y(n877) );
  INVX2TS U1406 ( .A(n956), .Y(n1785) );
  INVX2TS U1407 ( .A(n1579), .Y(n1677) );
  AOI22X1TS U1408 ( .A0(n1785), .A1(n1663), .B0(n1677), .B1(
        \requesterAddressbuffer[7][0] ), .Y(n885) );
  INVX2TS U1409 ( .A(n881), .Y(n1679) );
  INVX2TS U1410 ( .A(n1530), .Y(n1671) );
  AOI22X1TS U1411 ( .A0(n1679), .A1(n958), .B0(n1671), .B1(n1034), .Y(n884) );
  CLKBUFX2TS U1412 ( .A(n1037), .Y(n933) );
  INVX2TS U1413 ( .A(n882), .Y(n1688) );
  CLKBUFX2TS U1414 ( .A(n1005), .Y(n959) );
  AOI22X1TS U1415 ( .A0(n1689), .A1(n933), .B0(n1688), .B1(n959), .Y(n883) );
  INVX2TS U1416 ( .A(n894), .Y(n1670) );
  AOI22X1TS U1417 ( .A0(n1670), .A1(n1669), .B0(n1684), .B1(
        \requesterAddressbuffer[7][1] ), .Y(n888) );
  AOI22X1TS U1418 ( .A0(n1672), .A1(n966), .B0(n889), .B1(n1042), .Y(n887) );
  CLKBUFX2TS U1419 ( .A(n1043), .Y(n941) );
  CLKBUFX2TS U1420 ( .A(n1012), .Y(n968) );
  AOI22X1TS U1421 ( .A0(n1665), .A1(n941), .B0(n1523), .B1(n968), .Y(n886) );
  INVX2TS U1422 ( .A(n1579), .Y(n1528) );
  AOI22X1TS U1423 ( .A0(n32), .A1(n1678), .B0(n1528), .B1(
        \requesterAddressbuffer[7][2] ), .Y(n893) );
  AOI22X1TS U1424 ( .A0(n34), .A1(n973), .B0(n889), .B1(n1047), .Y(n892) );
  INVX2TS U1425 ( .A(n1532), .Y(n1665) );
  CLKBUFX2TS U1426 ( .A(n1048), .Y(n946) );
  CLKBUFX2TS U1427 ( .A(n1020), .Y(n976) );
  AOI22X1TS U1428 ( .A0(n1665), .A1(n946), .B0(n890), .B1(n976), .Y(n891) );
  INVX2TS U1429 ( .A(n894), .Y(n1686) );
  AOI22X1TS U1430 ( .A0(n1686), .A1(n1685), .B0(n1528), .B1(
        \requesterAddressbuffer[7][3] ), .Y(n898) );
  INVX2TS U1431 ( .A(n1530), .Y(n1687) );
  AOI22X1TS U1432 ( .A0(n1521), .A1(n981), .B0(n1687), .B1(n1054), .Y(n897) );
  CLKBUFX2TS U1433 ( .A(n1055), .Y(n952) );
  CLKBUFX2TS U1434 ( .A(n1029), .Y(n982) );
  AOI22X1TS U1435 ( .A0(n895), .A1(n952), .B0(n1556), .B1(n982), .Y(n896) );
  INVX2TS U1436 ( .A(n956), .Y(n1841) );
  INVX2TS U1437 ( .A(n1485), .Y(n1707) );
  AOI22X1TS U1438 ( .A0(n1841), .A1(n902), .B0(n1707), .B1(
        \requesterAddressbuffer[6][0] ), .Y(n901) );
  INVX2TS U1439 ( .A(n1469), .Y(n1699) );
  AOI22X1TS U1440 ( .A0(n932), .A1(n1488), .B0(requesterAddressIn_EAST[0]), 
        .B1(n1699), .Y(n900) );
  AOI22X1TS U1441 ( .A0(n933), .A1(n1718), .B0(n959), .B1(n1703), .Y(n899) );
  INVX2TS U1442 ( .A(n963), .Y(n1762) );
  AOI22X1TS U1443 ( .A0(n1762), .A1(n902), .B0(n1714), .B1(
        \requesterAddressbuffer[6][1] ), .Y(n908) );
  INVX2TS U1444 ( .A(n903), .Y(n1716) );
  INVX2TS U1445 ( .A(n1469), .Y(n1708) );
  AOI22X1TS U1446 ( .A0(n939), .A1(n1716), .B0(requesterAddressIn_EAST[1]), 
        .B1(n1708), .Y(n907) );
  INVX2TS U1447 ( .A(n905), .Y(n1491) );
  AOI22X1TS U1448 ( .A0(n941), .A1(n1498), .B0(n968), .B1(n1491), .Y(n906) );
  INVX2TS U1449 ( .A(n972), .Y(n1772) );
  INVX2TS U1450 ( .A(n1484), .Y(n1698) );
  INVX2TS U1451 ( .A(n1590), .Y(n1476) );
  AOI22X1TS U1452 ( .A0(n1772), .A1(n1698), .B0(n1476), .B1(
        \requesterAddressbuffer[6][2] ), .Y(n911) );
  AOI22X1TS U1453 ( .A0(n945), .A1(n104), .B0(requesterAddressIn_EAST[2]), 
        .B1(n912), .Y(n910) );
  AOI22X1TS U1454 ( .A0(n946), .A1(n1702), .B0(n976), .B1(n100), .Y(n909) );
  INVX2TS U1455 ( .A(n980), .Y(n1779) );
  AOI22X1TS U1456 ( .A0(n1779), .A1(n76), .B0(n1476), .B1(
        \requesterAddressbuffer[6][3] ), .Y(n915) );
  AOI22X1TS U1457 ( .A0(n951), .A1(n94), .B0(requesterAddressIn_EAST[3]), .B1(
        n912), .Y(n914) );
  AOI22X1TS U1458 ( .A0(n952), .A1(n105), .B0(n982), .B1(n1710), .Y(n913) );
  INVX2TS U1459 ( .A(n1451), .Y(n1738) );
  AOI22X1TS U1460 ( .A0(n1003), .A1(n920), .B0(n1738), .B1(
        \requesterAddressbuffer[5][0] ), .Y(n919) );
  INVX2TS U1461 ( .A(n1440), .Y(n1730) );
  AOI22X1TS U1462 ( .A0(n932), .A1(n1452), .B0(requesterAddressIn_EAST[0]), 
        .B1(n1730), .Y(n918) );
  INVX2TS U1463 ( .A(n916), .Y(n1733) );
  AOI22X1TS U1464 ( .A0(n933), .A1(n1733), .B0(requesterAddressIn_NORTH[0]), 
        .B1(n1447), .Y(n917) );
  AOI22X1TS U1465 ( .A0(n1669), .A1(n920), .B0(n1749), .B1(
        \requesterAddressbuffer[5][1] ), .Y(n923) );
  INVX2TS U1466 ( .A(n1440), .Y(n1741) );
  AOI22X1TS U1467 ( .A0(n939), .A1(n1743), .B0(requesterAddressIn_EAST[1]), 
        .B1(n1741), .Y(n922) );
  AOI22X1TS U1468 ( .A0(n941), .A1(n1744), .B0(requesterAddressIn_NORTH[1]), 
        .B1(n1745), .Y(n921) );
  INVX2TS U1469 ( .A(n10), .Y(n1728) );
  INVX2TS U1470 ( .A(n1603), .Y(n1446) );
  AOI22X1TS U1471 ( .A0(n1678), .A1(n1728), .B0(n1446), .B1(
        \requesterAddressbuffer[5][2] ), .Y(n926) );
  AOI22X1TS U1472 ( .A0(n945), .A1(n1456), .B0(requesterAddressIn_EAST[2]), 
        .B1(n928), .Y(n925) );
  AOI22X1TS U1473 ( .A0(n946), .A1(n1442), .B0(requesterAddressIn_NORTH[2]), 
        .B1(n1724), .Y(n924) );
  INVX2TS U1474 ( .A(n10), .Y(n1739) );
  AOI22X1TS U1475 ( .A0(n1685), .A1(n1739), .B0(n1446), .B1(
        \requesterAddressbuffer[5][3] ), .Y(n931) );
  INVX2TS U1476 ( .A(n927), .Y(n1743) );
  AOI22X1TS U1477 ( .A0(n951), .A1(n1743), .B0(requesterAddressIn_EAST[3]), 
        .B1(n928), .Y(n930) );
  AOI22X1TS U1478 ( .A0(n952), .A1(n234), .B0(requesterAddressIn_NORTH[3]), 
        .B1(n1734), .Y(n929) );
  INVX2TS U1479 ( .A(n1420), .Y(n1770) );
  AOI22X1TS U1480 ( .A0(n1003), .A1(n937), .B0(n1770), .B1(
        \requesterAddressbuffer[4][0] ), .Y(n936) );
  INVX2TS U1481 ( .A(n1407), .Y(n1763) );
  AOI22X1TS U1482 ( .A0(n932), .A1(n1756), .B0(requesterAddressIn_EAST[0]), 
        .B1(n1763), .Y(n935) );
  AOI22X1TS U1483 ( .A0(n933), .A1(n280), .B0(requesterAddressIn_NORTH[0]), 
        .B1(n291), .Y(n934) );
  INVX2TS U1484 ( .A(n963), .Y(n1892) );
  AOI22X1TS U1485 ( .A0(n1892), .A1(n937), .B0(n1778), .B1(
        \requesterAddressbuffer[4][1] ), .Y(n944) );
  INVX2TS U1486 ( .A(n1407), .Y(n1773) );
  AOI22X1TS U1487 ( .A0(n939), .A1(n294), .B0(requesterAddressIn_EAST[1]), 
        .B1(n1773), .Y(n943) );
  AOI22X1TS U1488 ( .A0(n941), .A1(n1781), .B0(requesterAddressIn_NORTH[1]), 
        .B1(n940), .Y(n942) );
  INVX2TS U1489 ( .A(n972), .Y(n1904) );
  INVX2TS U1490 ( .A(n1419), .Y(n1761) );
  INVX2TS U1491 ( .A(n1615), .Y(n1412) );
  AOI22X1TS U1492 ( .A0(n1904), .A1(n1761), .B0(n1412), .B1(
        \requesterAddressbuffer[4][2] ), .Y(n949) );
  AOI22X1TS U1493 ( .A0(n945), .A1(n1764), .B0(requesterAddressIn_EAST[2]), 
        .B1(n950), .Y(n948) );
  AOI22X1TS U1494 ( .A0(n946), .A1(n1436), .B0(requesterAddressIn_NORTH[2]), 
        .B1(n1757), .Y(n947) );
  INVX2TS U1495 ( .A(n980), .Y(n1915) );
  INVX2TS U1496 ( .A(n1419), .Y(n1771) );
  AOI22X1TS U1497 ( .A0(n1915), .A1(n1771), .B0(n1412), .B1(
        \requesterAddressbuffer[4][3] ), .Y(n955) );
  AOI22X1TS U1498 ( .A0(n951), .A1(n288), .B0(requesterAddressIn_EAST[3]), 
        .B1(n950), .Y(n954) );
  AOI22X1TS U1499 ( .A0(n952), .A1(n1422), .B0(requesterAddressIn_NORTH[3]), 
        .B1(n1765), .Y(n953) );
  INVX2TS U1500 ( .A(n956), .Y(n1884) );
  INVX2TS U1501 ( .A(n1389), .Y(n1799) );
  AOI22X1TS U1502 ( .A0(n1884), .A1(n964), .B0(n1799), .B1(
        \requesterAddressbuffer[3][0] ), .Y(n962) );
  INVX2TS U1503 ( .A(n957), .Y(n1794) );
  AOI22X1TS U1504 ( .A0(n958), .A1(n1794), .B0(n1004), .B1(n163), .Y(n961) );
  INVX2TS U1505 ( .A(n974), .Y(n1403) );
  AOI22X1TS U1506 ( .A0(n1006), .A1(n1403), .B0(n959), .B1(n1795), .Y(n960) );
  INVX2TS U1507 ( .A(n963), .Y(n1851) );
  AOI22X1TS U1508 ( .A0(n1851), .A1(n964), .B0(n1805), .B1(
        \requesterAddressbuffer[3][1] ), .Y(n971) );
  INVX2TS U1509 ( .A(n965), .Y(n1807) );
  AOI22X1TS U1510 ( .A0(n966), .A1(n126), .B0(n1011), .B1(n1807), .Y(n970) );
  AOI22X1TS U1511 ( .A0(n1013), .A1(n121), .B0(n968), .B1(n975), .Y(n969) );
  INVX2TS U1512 ( .A(n972), .Y(n1863) );
  INVX2TS U1513 ( .A(n1388), .Y(n1791) );
  INVX2TS U1514 ( .A(n1624), .Y(n1383) );
  AOI22X1TS U1515 ( .A0(n1863), .A1(n1791), .B0(n1383), .B1(
        \requesterAddressbuffer[3][2] ), .Y(n979) );
  AOI22X1TS U1516 ( .A0(n973), .A1(n1787), .B0(n1018), .B1(n1379), .Y(n978) );
  INVX2TS U1517 ( .A(n974), .Y(n1810) );
  AOI22X1TS U1518 ( .A0(n1021), .A1(n1810), .B0(n976), .B1(n975), .Y(n977) );
  INVX2TS U1519 ( .A(n980), .Y(n1875) );
  AOI22X1TS U1520 ( .A0(n1875), .A1(n122), .B0(n1383), .B1(
        \requesterAddressbuffer[3][3] ), .Y(n985) );
  AOI22X1TS U1521 ( .A0(n981), .A1(n1794), .B0(n1027), .B1(n1396), .Y(n984) );
  AOI22X1TS U1522 ( .A0(n1030), .A1(n1403), .B0(n982), .B1(n1801), .Y(n983) );
  INVX2TS U1523 ( .A(n1636), .Y(n1825) );
  AOI22X1TS U1524 ( .A0(n1785), .A1(n989), .B0(n1825), .B1(
        \requesterAddressbuffer[2][0] ), .Y(n988) );
  INVX2TS U1525 ( .A(n1357), .Y(n1819) );
  AOI22X1TS U1526 ( .A0(requesterAddressIn_WEST[0]), .A1(n1814), .B0(n1004), 
        .B1(n1819), .Y(n987) );
  AOI22X1TS U1527 ( .A0(n1006), .A1(n1836), .B0(n1005), .B1(n1830), .Y(n986)
         );
  AOI22X1TS U1528 ( .A0(n1892), .A1(n989), .B0(n1834), .B1(
        \requesterAddressbuffer[2][1] ), .Y(n992) );
  INVX2TS U1529 ( .A(n1357), .Y(n1827) );
  AOI22X1TS U1530 ( .A0(requesterAddressIn_WEST[1]), .A1(n1359), .B0(n1011), 
        .B1(n1827), .Y(n991) );
  INVX2TS U1531 ( .A(n993), .Y(n1829) );
  AOI22X1TS U1532 ( .A0(n1013), .A1(n1829), .B0(n1012), .B1(n1837), .Y(n990)
         );
  INVX2TS U1533 ( .A(n9), .Y(n1818) );
  INVX2TS U1534 ( .A(n1636), .Y(n1350) );
  AOI22X1TS U1535 ( .A0(n1904), .A1(n1818), .B0(n1350), .B1(
        \requesterAddressbuffer[2][2] ), .Y(n997) );
  AOI22X1TS U1536 ( .A0(requesterAddressIn_WEST[2]), .A1(n1820), .B0(n1018), 
        .B1(n999), .Y(n996) );
  INVX2TS U1537 ( .A(n993), .Y(n1360) );
  AOI22X1TS U1538 ( .A0(n1021), .A1(n1360), .B0(n1020), .B1(n994), .Y(n995) );
  INVX2TS U1539 ( .A(n9), .Y(n1826) );
  AOI22X1TS U1540 ( .A0(n1915), .A1(n1826), .B0(n1350), .B1(
        \requesterAddressbuffer[2][3] ), .Y(n1002) );
  INVX2TS U1541 ( .A(n998), .Y(n1359) );
  AOI22X1TS U1542 ( .A0(requesterAddressIn_WEST[3]), .A1(n1359), .B0(n1027), 
        .B1(n999), .Y(n1001) );
  AOI22X1TS U1543 ( .A0(n1030), .A1(n193), .B0(n1029), .B1(n1821), .Y(n1000)
         );
  INVX2TS U1544 ( .A(n1017), .Y(n1861) );
  AOI22X1TS U1545 ( .A0(n1003), .A1(n1010), .B0(n1861), .B1(
        \requesterAddressbuffer[1][0] ), .Y(n1009) );
  INVX2TS U1546 ( .A(n1), .Y(n1853) );
  AOI22X1TS U1547 ( .A0(requesterAddressIn_WEST[0]), .A1(n1843), .B0(n1004), 
        .B1(n1853), .Y(n1008) );
  AOI22X1TS U1548 ( .A0(n1006), .A1(n1878), .B0(n1005), .B1(n1857), .Y(n1007)
         );
  AOI22X1TS U1549 ( .A0(n1762), .A1(n1010), .B0(n1874), .B1(
        \requesterAddressbuffer[1][1] ), .Y(n1016) );
  INVX2TS U1550 ( .A(n1), .Y(n1865) );
  AOI22X1TS U1551 ( .A0(requesterAddressIn_WEST[1]), .A1(n1099), .B0(n1011), 
        .B1(n1865), .Y(n1015) );
  INVX2TS U1552 ( .A(n340), .Y(n1868) );
  AOI22X1TS U1553 ( .A0(n1013), .A1(n1868), .B0(n1012), .B1(n1019), .Y(n1014)
         );
  INVX2TS U1554 ( .A(n1097), .Y(n1850) );
  INVX2TS U1555 ( .A(n1017), .Y(n1092) );
  AOI22X1TS U1556 ( .A0(n1772), .A1(n1850), .B0(n1092), .B1(
        \requesterAddressbuffer[1][2] ), .Y(n1024) );
  AOI22X1TS U1557 ( .A0(requesterAddressIn_WEST[2]), .A1(n1854), .B0(n1018), 
        .B1(n1026), .Y(n1023) );
  AOI22X1TS U1558 ( .A0(n1021), .A1(n320), .B0(n1020), .B1(n1019), .Y(n1022)
         );
  INVX2TS U1559 ( .A(n1097), .Y(n1862) );
  AOI22X1TS U1560 ( .A0(n1779), .A1(n1862), .B0(n1092), .B1(
        \requesterAddressbuffer[1][3] ), .Y(n1033) );
  INVX2TS U1561 ( .A(n1025), .Y(n1099) );
  AOI22X1TS U1562 ( .A0(requesterAddressIn_WEST[3]), .A1(n1099), .B0(n1027), 
        .B1(n1026), .Y(n1032) );
  INVX2TS U1563 ( .A(n1028), .Y(n1101) );
  AOI22X1TS U1564 ( .A0(n1030), .A1(n1101), .B0(n1029), .B1(n1870), .Y(n1031)
         );
  INVX2TS U1565 ( .A(n1067), .Y(n1902) );
  AOI22X1TS U1566 ( .A0(readRequesterAddress[0]), .A1(n1041), .B0(n1902), .B1(
        \requesterAddressbuffer[0][0] ), .Y(n1040) );
  INVX2TS U1567 ( .A(n1068), .Y(n1893) );
  AOI22X1TS U1568 ( .A0(requesterAddressIn_WEST[0]), .A1(n1885), .B0(n1034), 
        .B1(n1893), .Y(n1039) );
  INVX2TS U1569 ( .A(n1035), .Y(n1082) );
  INVX2TS U1570 ( .A(n1036), .Y(n1077) );
  AOI22X1TS U1571 ( .A0(n1037), .A1(n1082), .B0(requesterAddressIn_NORTH[0]), 
        .B1(n1077), .Y(n1038) );
  AOI22X1TS U1572 ( .A0(n1851), .A1(n1041), .B0(n1913), .B1(
        \requesterAddressbuffer[0][1] ), .Y(n1046) );
  INVX2TS U1573 ( .A(n1068), .Y(n1905) );
  AOI22X1TS U1574 ( .A0(requesterAddressIn_WEST[1]), .A1(n1069), .B0(n1042), 
        .B1(n1905), .Y(n1045) );
  AOI22X1TS U1575 ( .A0(n1043), .A1(n1070), .B0(requesterAddressIn_NORTH[1]), 
        .B1(n1077), .Y(n1044) );
  INVX2TS U1576 ( .A(n11), .Y(n1891) );
  INVX2TS U1577 ( .A(n1067), .Y(n1063) );
  AOI22X1TS U1578 ( .A0(n1863), .A1(n1891), .B0(n1063), .B1(
        \requesterAddressbuffer[0][2] ), .Y(n1051) );
  AOI22X1TS U1579 ( .A0(requesterAddressIn_WEST[2]), .A1(n1894), .B0(n1047), 
        .B1(n1053), .Y(n1050) );
  AOI22X1TS U1580 ( .A0(n1048), .A1(n1918), .B0(requesterAddressIn_NORTH[2]), 
        .B1(n1896), .Y(n1049) );
  INVX2TS U1581 ( .A(n11), .Y(n1903) );
  AOI22X1TS U1582 ( .A0(n1875), .A1(n1903), .B0(n1063), .B1(
        \requesterAddressbuffer[0][3] ), .Y(n1058) );
  INVX2TS U1583 ( .A(n1052), .Y(n1069) );
  AOI22X1TS U1584 ( .A0(requesterAddressIn_WEST[3]), .A1(n1069), .B0(n1054), 
        .B1(n1053), .Y(n1057) );
  AOI22X1TS U1585 ( .A0(n1055), .A1(n1898), .B0(requesterAddressIn_NORTH[3]), 
        .B1(n1059), .Y(n1056) );
  INVX2TS U1586 ( .A(n1086), .Y(n1468) );
  AOI22X1TS U1587 ( .A0(n1891), .A1(n1468), .B0(n1063), .B1(
        \dataoutbuffer[0][0] ), .Y(n1062) );
  AOI22X1TS U1588 ( .A0(n1069), .A1(n1408), .B0(n1893), .B1(n1346), .Y(n1061)
         );
  CLKBUFX2TS U1589 ( .A(n1087), .Y(n1472) );
  AOI22X1TS U1590 ( .A0(n1918), .A1(dataIn_SOUTH[0]), .B0(n1059), .B1(n1472), 
        .Y(n1060) );
  INVX2TS U1591 ( .A(n1091), .Y(n1477) );
  AOI22X1TS U1592 ( .A0(n1903), .A1(n1477), .B0(n1063), .B1(
        \dataoutbuffer[0][1] ), .Y(n1066) );
  AOI22X1TS U1593 ( .A0(n419), .A1(n1413), .B0(n1905), .B1(n1351), .Y(n1065)
         );
  CLKBUFX2TS U1594 ( .A(n1093), .Y(n1480) );
  AOI22X1TS U1595 ( .A0(n1082), .A1(dataIn_SOUTH[1]), .B0(n395), .B1(n1480), 
        .Y(n1064) );
  INVX2TS U1596 ( .A(n11), .Y(n1914) );
  INVX2TS U1597 ( .A(n1098), .Y(n1486) );
  INVX2TS U1598 ( .A(n1067), .Y(n1081) );
  AOI22X1TS U1599 ( .A0(n1914), .A1(n1486), .B0(n1081), .B1(
        \dataoutbuffer[0][2] ), .Y(n1073) );
  AOI22X1TS U1600 ( .A0(n1069), .A1(n1421), .B0(n389), .B1(n1358), .Y(n1072)
         );
  CLKBUFX2TS U1601 ( .A(n1100), .Y(n1490) );
  AOI22X1TS U1602 ( .A0(n1070), .A1(dataIn_SOUTH[2]), .B0(n1077), .B1(n1490), 
        .Y(n1071) );
  INVX2TS U1603 ( .A(n1105), .Y(n1495) );
  AOI22X1TS U1604 ( .A0(n1891), .A1(n1495), .B0(n1081), .B1(
        \dataoutbuffer[0][3] ), .Y(n1076) );
  AOI22X1TS U1605 ( .A0(n1906), .A1(n1426), .B0(n1893), .B1(n1365), .Y(n1075)
         );
  CLKBUFX2TS U1606 ( .A(n1106), .Y(n1499) );
  AOI22X1TS U1607 ( .A0(n1082), .A1(dataIn_SOUTH[3]), .B0(n1908), .B1(n1499), 
        .Y(n1074) );
  INVX2TS U1608 ( .A(n1111), .Y(n1503) );
  AOI22X1TS U1609 ( .A0(n1903), .A1(n1503), .B0(n1081), .B1(
        \dataoutbuffer[0][4] ), .Y(n1080) );
  AOI22X1TS U1610 ( .A0(n1885), .A1(n1430), .B0(n1905), .B1(n1370), .Y(n1079)
         );
  CLKBUFX2TS U1611 ( .A(n1112), .Y(n1506) );
  AOI22X1TS U1612 ( .A0(n443), .A1(dataIn_SOUTH[4]), .B0(n1077), .B1(n1506), 
        .Y(n1078) );
  INVX2TS U1613 ( .A(n1340), .Y(n1511) );
  AOI22X1TS U1614 ( .A0(n1914), .A1(n1511), .B0(n1081), .B1(
        \dataoutbuffer[0][5] ), .Y(n1085) );
  AOI22X1TS U1615 ( .A0(n419), .A1(n1435), .B0(n389), .B1(n1375), .Y(n1084) );
  CLKBUFX2TS U1616 ( .A(n1342), .Y(n1515) );
  AOI22X1TS U1617 ( .A0(n1082), .A1(dataIn_SOUTH[5]), .B0(n395), .B1(n1515), 
        .Y(n1083) );
  INVX2TS U1618 ( .A(n1086), .Y(n1519) );
  AOI22X1TS U1619 ( .A0(n1850), .A1(n1519), .B0(n1092), .B1(
        \dataoutbuffer[1][0] ), .Y(n1090) );
  AOI22X1TS U1620 ( .A0(n1099), .A1(dataIn_WEST[0]), .B0(n1853), .B1(n1346), 
        .Y(n1089) );
  CLKBUFX2TS U1621 ( .A(n1087), .Y(n1522) );
  CLKBUFX2TS U1622 ( .A(dataIn_SOUTH[0]), .Y(n1524) );
  CLKBUFX2TS U1623 ( .A(n1524), .Y(n1471) );
  AOI22X1TS U1624 ( .A0(n1019), .A1(n1522), .B0(n1107), .B1(n1471), .Y(n1088)
         );
  INVX2TS U1625 ( .A(n1091), .Y(n1529) );
  AOI22X1TS U1626 ( .A0(n1862), .A1(n1529), .B0(n1092), .B1(
        \dataoutbuffer[1][1] ), .Y(n1096) );
  AOI22X1TS U1627 ( .A0(n330), .A1(dataIn_WEST[1]), .B0(n1865), .B1(n1351), 
        .Y(n1095) );
  CLKBUFX2TS U1628 ( .A(n1093), .Y(n1533) );
  CLKBUFX2TS U1629 ( .A(dataIn_SOUTH[1]), .Y(n1534) );
  CLKBUFX2TS U1630 ( .A(n1534), .Y(n1479) );
  AOI22X1TS U1631 ( .A0(n1880), .A1(n1533), .B0(n1101), .B1(n1479), .Y(n1094)
         );
  INVX2TS U1632 ( .A(n1098), .Y(n1539) );
  INVX2TS U1633 ( .A(n1017), .Y(n1341) );
  AOI22X1TS U1634 ( .A0(n311), .A1(n1539), .B0(n1341), .B1(
        \dataoutbuffer[1][2] ), .Y(n1104) );
  AOI22X1TS U1635 ( .A0(n1099), .A1(dataIn_WEST[2]), .B0(n309), .B1(n1358), 
        .Y(n1103) );
  CLKBUFX2TS U1636 ( .A(n1100), .Y(n1541) );
  CLKBUFX2TS U1637 ( .A(dataIn_SOUTH[2]), .Y(n1542) );
  CLKBUFX2TS U1638 ( .A(n1542), .Y(n1489) );
  AOI22X1TS U1639 ( .A0(n316), .A1(n1541), .B0(n1101), .B1(n1489), .Y(n1102)
         );
  INVX2TS U1640 ( .A(n1105), .Y(n1546) );
  AOI22X1TS U1641 ( .A0(n1850), .A1(n1546), .B0(n1341), .B1(
        \dataoutbuffer[1][3] ), .Y(n1110) );
  AOI22X1TS U1642 ( .A0(n1866), .A1(dataIn_WEST[3]), .B0(n1853), .B1(n1365), 
        .Y(n1109) );
  CLKBUFX2TS U1643 ( .A(n1106), .Y(n1548) );
  CLKBUFX2TS U1644 ( .A(dataIn_SOUTH[3]), .Y(n1549) );
  CLKBUFX2TS U1645 ( .A(n1549), .Y(n1497) );
  AOI22X1TS U1646 ( .A0(n1870), .A1(n1548), .B0(n1107), .B1(n1497), .Y(n1108)
         );
  INVX2TS U1647 ( .A(n1111), .Y(n1553) );
  AOI22X1TS U1648 ( .A0(n1862), .A1(n1553), .B0(n1341), .B1(
        \dataoutbuffer[1][4] ), .Y(n1339) );
  AOI22X1TS U1649 ( .A0(n1843), .A1(dataIn_WEST[4]), .B0(n1865), .B1(n1370), 
        .Y(n1338) );
  CLKBUFX2TS U1650 ( .A(n1112), .Y(n1555) );
  CLKBUFX2TS U1651 ( .A(dataIn_SOUTH[4]), .Y(n1557) );
  CLKBUFX2TS U1652 ( .A(n1557), .Y(n1505) );
  AOI22X1TS U1653 ( .A0(n1846), .A1(n1555), .B0(n1868), .B1(n1505), .Y(n1337)
         );
  INVX2TS U1654 ( .A(n1340), .Y(n1562) );
  AOI22X1TS U1655 ( .A0(n1010), .A1(n1562), .B0(n1341), .B1(
        \dataoutbuffer[1][5] ), .Y(n1345) );
  AOI22X1TS U1656 ( .A0(n330), .A1(dataIn_WEST[5]), .B0(n309), .B1(n1375), .Y(
        n1344) );
  CLKBUFX2TS U1657 ( .A(n1342), .Y(n1564) );
  CLKBUFX2TS U1658 ( .A(dataIn_SOUTH[5]), .Y(n1565) );
  CLKBUFX2TS U1659 ( .A(n1565), .Y(n1513) );
  AOI22X1TS U1660 ( .A0(n1880), .A1(n1564), .B0(n366), .B1(n1513), .Y(n1343)
         );
  AOI22X1TS U1661 ( .A0(n1818), .A1(n1468), .B0(n1350), .B1(
        \dataoutbuffer[2][0] ), .Y(n1349) );
  AOI22X1TS U1662 ( .A0(n1359), .A1(dataIn_WEST[0]), .B0(n1819), .B1(n1346), 
        .Y(n1348) );
  AOI22X1TS U1663 ( .A0(n1361), .A1(n1522), .B0(n1366), .B1(dataIn_SOUTH[0]), 
        .Y(n1347) );
  AOI22X1TS U1664 ( .A0(n1826), .A1(n1477), .B0(n1350), .B1(
        \dataoutbuffer[2][1] ), .Y(n1355) );
  AOI22X1TS U1665 ( .A0(n186), .A1(dataIn_WEST[1]), .B0(n1827), .B1(n1351), 
        .Y(n1354) );
  INVX2TS U1666 ( .A(n1352), .Y(n1837) );
  AOI22X1TS U1667 ( .A0(n1837), .A1(n1533), .B0(n1360), .B1(dataIn_SOUTH[1]), 
        .Y(n1353) );
  INVX2TS U1668 ( .A(n9), .Y(n1835) );
  INVX2TS U1669 ( .A(n1356), .Y(n1374) );
  AOI22X1TS U1670 ( .A0(n1835), .A1(n1486), .B0(n1374), .B1(
        \dataoutbuffer[2][2] ), .Y(n1364) );
  AOI22X1TS U1671 ( .A0(n1359), .A1(dataIn_WEST[2]), .B0(n171), .B1(n1358), 
        .Y(n1363) );
  AOI22X1TS U1672 ( .A0(n1361), .A1(n1541), .B0(n1360), .B1(dataIn_SOUTH[2]), 
        .Y(n1362) );
  AOI22X1TS U1673 ( .A0(n1818), .A1(n1495), .B0(n1374), .B1(
        \dataoutbuffer[2][3] ), .Y(n1369) );
  AOI22X1TS U1674 ( .A0(n1828), .A1(dataIn_WEST[3]), .B0(n1819), .B1(n1365), 
        .Y(n1368) );
  AOI22X1TS U1675 ( .A0(n994), .A1(n1548), .B0(n1366), .B1(dataIn_SOUTH[3]), 
        .Y(n1367) );
  AOI22X1TS U1676 ( .A0(n1826), .A1(n1503), .B0(n1374), .B1(
        \dataoutbuffer[2][4] ), .Y(n1373) );
  AOI22X1TS U1677 ( .A0(n1814), .A1(dataIn_WEST[4]), .B0(n1827), .B1(n1370), 
        .Y(n1372) );
  AOI22X1TS U1678 ( .A0(n1821), .A1(n1555), .B0(n193), .B1(dataIn_SOUTH[4]), 
        .Y(n1371) );
  AOI22X1TS U1679 ( .A0(n1835), .A1(n1511), .B0(n1374), .B1(
        \dataoutbuffer[2][5] ), .Y(n1378) );
  AOI22X1TS U1680 ( .A0(n186), .A1(dataIn_WEST[5]), .B0(n171), .B1(n1375), .Y(
        n1377) );
  AOI22X1TS U1681 ( .A0(n1837), .A1(n1564), .B0(n201), .B1(dataIn_SOUTH[5]), 
        .Y(n1376) );
  AOI22X1TS U1682 ( .A0(n1791), .A1(n1468), .B0(n1383), .B1(
        \dataoutbuffer[3][0] ), .Y(n1382) );
  AOI22X1TS U1683 ( .A0(n1397), .A1(dataIn_WEST[0]), .B0(n1379), .B1(
        dataIn_EAST[0]), .Y(n1381) );
  AOI22X1TS U1684 ( .A0(n153), .A1(n1472), .B0(n1384), .B1(n1471), .Y(n1380)
         );
  AOI22X1TS U1685 ( .A0(n122), .A1(n1477), .B0(n1383), .B1(
        \dataoutbuffer[3][1] ), .Y(n1387) );
  AOI22X1TS U1686 ( .A0(n1809), .A1(dataIn_WEST[1]), .B0(n1807), .B1(
        dataIn_EAST[1]), .Y(n1386) );
  AOI22X1TS U1687 ( .A0(n1398), .A1(n1480), .B0(n1384), .B1(n1479), .Y(n1385)
         );
  INVX2TS U1688 ( .A(n1388), .Y(n1806) );
  INVX2TS U1689 ( .A(n1389), .Y(n1402) );
  AOI22X1TS U1690 ( .A0(n1806), .A1(n1486), .B0(n1402), .B1(
        \dataoutbuffer[3][2] ), .Y(n1392) );
  AOI22X1TS U1691 ( .A0(n147), .A1(dataIn_WEST[2]), .B0(n163), .B1(
        dataIn_EAST[2]), .Y(n1391) );
  AOI22X1TS U1692 ( .A0(n153), .A1(n1490), .B0(n1403), .B1(n1489), .Y(n1390)
         );
  AOI22X1TS U1693 ( .A0(n1791), .A1(n1495), .B0(n1402), .B1(
        \dataoutbuffer[3][3] ), .Y(n1395) );
  AOI22X1TS U1694 ( .A0(n1794), .A1(dataIn_WEST[3]), .B0(n151), .B1(
        dataIn_EAST[3]), .Y(n1394) );
  AOI22X1TS U1695 ( .A0(n1801), .A1(n1499), .B0(n134), .B1(n1497), .Y(n1393)
         );
  AOI22X1TS U1696 ( .A0(n964), .A1(n1503), .B0(n1402), .B1(
        \dataoutbuffer[3][4] ), .Y(n1401) );
  AOI22X1TS U1697 ( .A0(n1397), .A1(dataIn_WEST[4]), .B0(n1396), .B1(
        dataIn_EAST[4]), .Y(n1400) );
  AOI22X1TS U1698 ( .A0(n1398), .A1(n1506), .B0(n1810), .B1(n1505), .Y(n1399)
         );
  AOI22X1TS U1699 ( .A0(n1806), .A1(n1511), .B0(n1402), .B1(
        \dataoutbuffer[3][5] ), .Y(n1406) );
  AOI22X1TS U1700 ( .A0(n135), .A1(dataIn_WEST[5]), .B0(n1807), .B1(
        dataIn_EAST[5]), .Y(n1405) );
  AOI22X1TS U1701 ( .A0(n153), .A1(n1515), .B0(n1403), .B1(n1513), .Y(n1404)
         );
  AOI22X1TS U1702 ( .A0(n1761), .A1(n1519), .B0(n1412), .B1(
        \dataoutbuffer[4][0] ), .Y(n1411) );
  AOI22X1TS U1703 ( .A0(n284), .A1(n1408), .B0(n950), .B1(dataIn_EAST[0]), .Y(
        n1410) );
  AOI22X1TS U1704 ( .A0(n1422), .A1(n1524), .B0(n273), .B1(n1522), .Y(n1409)
         );
  AOI22X1TS U1705 ( .A0(n1771), .A1(n1529), .B0(n1412), .B1(
        \dataoutbuffer[4][1] ), .Y(n1418) );
  AOI22X1TS U1706 ( .A0(n288), .A1(n1413), .B0(n1763), .B1(dataIn_EAST[1]), 
        .Y(n1417) );
  INVX2TS U1707 ( .A(n1414), .Y(n1766) );
  INVX2TS U1708 ( .A(n1415), .Y(n1780) );
  AOI22X1TS U1709 ( .A0(n1766), .A1(n1534), .B0(n1780), .B1(n1533), .Y(n1416)
         );
  INVX2TS U1710 ( .A(n1420), .Y(n1434) );
  AOI22X1TS U1711 ( .A0(n268), .A1(n1539), .B0(n1434), .B1(
        \dataoutbuffer[4][2] ), .Y(n1425) );
  AOI22X1TS U1712 ( .A0(n284), .A1(n1421), .B0(n1773), .B1(dataIn_EAST[2]), 
        .Y(n1424) );
  AOI22X1TS U1713 ( .A0(n1422), .A1(n1542), .B0(n273), .B1(n1541), .Y(n1423)
         );
  AOI22X1TS U1714 ( .A0(n1761), .A1(n1546), .B0(n1434), .B1(
        \dataoutbuffer[4][3] ), .Y(n1429) );
  AOI22X1TS U1715 ( .A0(n1774), .A1(n1426), .B0(n266), .B1(dataIn_EAST[3]), 
        .Y(n1428) );
  AOI22X1TS U1716 ( .A0(n1436), .A1(n1549), .B0(n1780), .B1(n1548), .Y(n1427)
         );
  AOI22X1TS U1717 ( .A0(n1771), .A1(n1553), .B0(n1434), .B1(
        \dataoutbuffer[4][4] ), .Y(n1433) );
  AOI22X1TS U1718 ( .A0(n1756), .A1(n1430), .B0(n1763), .B1(dataIn_EAST[4]), 
        .Y(n1432) );
  AOI22X1TS U1719 ( .A0(n1766), .A1(n1557), .B0(n1757), .B1(n1555), .Y(n1431)
         );
  AOI22X1TS U1720 ( .A0(n937), .A1(n1562), .B0(n1434), .B1(
        \dataoutbuffer[4][5] ), .Y(n1439) );
  AOI22X1TS U1721 ( .A0(n294), .A1(n1435), .B0(n1773), .B1(dataIn_EAST[5]), 
        .Y(n1438) );
  AOI22X1TS U1722 ( .A0(n1436), .A1(n1565), .B0(n1780), .B1(n1564), .Y(n1437)
         );
  AOI22X1TS U1723 ( .A0(n1728), .A1(n1519), .B0(n1446), .B1(
        \dataoutbuffer[5][0] ), .Y(n1445) );
  AOI22X1TS U1724 ( .A0(n1452), .A1(n1520), .B0(n928), .B1(n1470), .Y(n1444)
         );
  INVX2TS U1725 ( .A(n1441), .Y(n1734) );
  AOI22X1TS U1726 ( .A0(n1734), .A1(n1472), .B0(n1442), .B1(n1471), .Y(n1443)
         );
  AOI22X1TS U1727 ( .A0(n1739), .A1(n1529), .B0(n1446), .B1(
        \dataoutbuffer[5][1] ), .Y(n1450) );
  AOI22X1TS U1728 ( .A0(n250), .A1(n1531), .B0(n1730), .B1(n1478), .Y(n1449)
         );
  AOI22X1TS U1729 ( .A0(n1447), .A1(n1480), .B0(n251), .B1(n1479), .Y(n1448)
         );
  INVX2TS U1730 ( .A(n10), .Y(n1750) );
  INVX2TS U1731 ( .A(n1451), .Y(n1464) );
  AOI22X1TS U1732 ( .A0(n1750), .A1(n1539), .B0(n1464), .B1(
        \dataoutbuffer[5][2] ), .Y(n1455) );
  AOI22X1TS U1733 ( .A0(n1452), .A1(n1540), .B0(n1741), .B1(n1487), .Y(n1454)
         );
  AOI22X1TS U1734 ( .A0(n218), .A1(n1490), .B0(n1460), .B1(n1489), .Y(n1453)
         );
  AOI22X1TS U1735 ( .A0(n1728), .A1(n1546), .B0(n1464), .B1(
        \dataoutbuffer[5][3] ), .Y(n1459) );
  AOI22X1TS U1736 ( .A0(n1456), .A1(n1547), .B0(n213), .B1(n1496), .Y(n1458)
         );
  AOI22X1TS U1737 ( .A0(n1734), .A1(n1499), .B0(n1744), .B1(n1497), .Y(n1457)
         );
  AOI22X1TS U1738 ( .A0(n1739), .A1(n1553), .B0(n1464), .B1(
        \dataoutbuffer[5][4] ), .Y(n1463) );
  AOI22X1TS U1739 ( .A0(n1732), .A1(n1554), .B0(n1730), .B1(n1504), .Y(n1462)
         );
  AOI22X1TS U1740 ( .A0(n1745), .A1(n1506), .B0(n1460), .B1(n1505), .Y(n1461)
         );
  AOI22X1TS U1741 ( .A0(n1750), .A1(n1562), .B0(n1464), .B1(
        \dataoutbuffer[5][5] ), .Y(n1467) );
  AOI22X1TS U1742 ( .A0(n232), .A1(n1563), .B0(n1741), .B1(n1512), .Y(n1466)
         );
  AOI22X1TS U1743 ( .A0(n1724), .A1(n1515), .B0(n234), .B1(n1513), .Y(n1465)
         );
  AOI22X1TS U1744 ( .A0(n1698), .A1(n1468), .B0(n1476), .B1(
        \dataoutbuffer[6][0] ), .Y(n1475) );
  AOI22X1TS U1745 ( .A0(n1488), .A1(n1520), .B0(n912), .B1(n1470), .Y(n1474)
         );
  AOI22X1TS U1746 ( .A0(n1491), .A1(n1472), .B0(n1498), .B1(n1471), .Y(n1473)
         );
  AOI22X1TS U1747 ( .A0(n76), .A1(n1477), .B0(n1476), .B1(
        \dataoutbuffer[6][1] ), .Y(n1483) );
  AOI22X1TS U1748 ( .A0(n1716), .A1(n1531), .B0(n1699), .B1(n1478), .Y(n1482)
         );
  AOI22X1TS U1749 ( .A0(n97), .A1(n1480), .B0(n83), .B1(n1479), .Y(n1481) );
  INVX2TS U1750 ( .A(n1484), .Y(n1715) );
  INVX2TS U1751 ( .A(n1485), .Y(n1510) );
  AOI22X1TS U1752 ( .A0(n1715), .A1(n1486), .B0(n1510), .B1(
        \dataoutbuffer[6][2] ), .Y(n1494) );
  AOI22X1TS U1753 ( .A0(n1488), .A1(n1540), .B0(n1708), .B1(n1487), .Y(n1493)
         );
  AOI22X1TS U1754 ( .A0(n1491), .A1(n1490), .B0(n83), .B1(n1489), .Y(n1492) );
  AOI22X1TS U1755 ( .A0(n1698), .A1(n1495), .B0(n1510), .B1(
        \dataoutbuffer[6][3] ), .Y(n1502) );
  AOI22X1TS U1756 ( .A0(n94), .A1(n1547), .B0(n74), .B1(n1496), .Y(n1501) );
  AOI22X1TS U1757 ( .A0(n1710), .A1(n1499), .B0(n1498), .B1(n1497), .Y(n1500)
         );
  AOI22X1TS U1758 ( .A0(n902), .A1(n1503), .B0(n1510), .B1(
        \dataoutbuffer[6][4] ), .Y(n1509) );
  AOI22X1TS U1759 ( .A0(n1700), .A1(n1554), .B0(n1699), .B1(n1504), .Y(n1508)
         );
  AOI22X1TS U1760 ( .A0(n1694), .A1(n1506), .B0(n1514), .B1(n1505), .Y(n1507)
         );
  AOI22X1TS U1761 ( .A0(n1715), .A1(n1511), .B0(n1510), .B1(
        \dataoutbuffer[6][5] ), .Y(n1518) );
  AOI22X1TS U1762 ( .A0(n1716), .A1(n1563), .B0(n1708), .B1(n1512), .Y(n1517)
         );
  AOI22X1TS U1763 ( .A0(n1491), .A1(n1515), .B0(n1514), .B1(n1513), .Y(n1516)
         );
  AOI22X1TS U1764 ( .A0(n1670), .A1(n1519), .B0(n1528), .B1(
        \dataoutbuffer[7][0] ), .Y(n1527) );
  AOI22X1TS U1765 ( .A0(n1521), .A1(n1520), .B0(n1671), .B1(dataIn_EAST[0]), 
        .Y(n1526) );
  AOI22X1TS U1766 ( .A0(n65), .A1(n1524), .B0(n1523), .B1(n1522), .Y(n1525) );
  AOI22X1TS U1767 ( .A0(n32), .A1(n1529), .B0(n1528), .B1(
        \dataoutbuffer[7][1] ), .Y(n1537) );
  AOI22X1TS U1768 ( .A0(n1679), .A1(n1531), .B0(n889), .B1(dataIn_EAST[1]), 
        .Y(n1536) );
  INVX2TS U1769 ( .A(n1532), .Y(n1689) );
  AOI22X1TS U1770 ( .A0(n1689), .A1(n1534), .B0(n1688), .B1(n1533), .Y(n1535)
         );
  INVX2TS U1771 ( .A(n1538), .Y(n1561) );
  AOI22X1TS U1772 ( .A0(n1686), .A1(n1539), .B0(n1561), .B1(
        \dataoutbuffer[7][2] ), .Y(n1545) );
  AOI22X1TS U1773 ( .A0(n1672), .A1(n1540), .B0(n1687), .B1(dataIn_EAST[2]), 
        .Y(n1544) );
  AOI22X1TS U1774 ( .A0(n49), .A1(n1542), .B0(n38), .B1(n1541), .Y(n1543) );
  AOI22X1TS U1775 ( .A0(n1670), .A1(n1546), .B0(n1561), .B1(
        \dataoutbuffer[7][3] ), .Y(n1552) );
  AOI22X1TS U1776 ( .A0(n1679), .A1(n1547), .B0(n1671), .B1(dataIn_EAST[3]), 
        .Y(n1551) );
  AOI22X1TS U1777 ( .A0(n1680), .A1(n1549), .B0(n38), .B1(n1548), .Y(n1550) );
  AOI22X1TS U1778 ( .A0(n32), .A1(n1553), .B0(n1561), .B1(
        \dataoutbuffer[7][4] ), .Y(n1560) );
  AOI22X1TS U1779 ( .A0(n1664), .A1(n1554), .B0(n31), .B1(dataIn_EAST[4]), .Y(
        n1559) );
  AOI22X1TS U1780 ( .A0(n1689), .A1(n1557), .B0(n1556), .B1(n1555), .Y(n1558)
         );
  AOI22X1TS U1781 ( .A0(n1686), .A1(n1562), .B0(n1561), .B1(
        \dataoutbuffer[7][5] ), .Y(n1568) );
  AOI22X1TS U1782 ( .A0(n63), .A1(n1563), .B0(n1687), .B1(dataIn_EAST[5]), .Y(
        n1567) );
  AOI22X1TS U1783 ( .A0(n1665), .A1(n1565), .B0(n1688), .B1(n1564), .Y(n1566)
         );
  INVX2TS U1784 ( .A(n1569), .Y(n1643) );
  AOI22X1TS U1785 ( .A0(n1571), .A1(n1594), .B0(n1593), .B1(n1570), .Y(n1573)
         );
  AOI22X1TS U1786 ( .A0(n1574), .A1(n1643), .B0(n1573), .B1(n1572), .Y(n1576)
         );
  AOI22X1TS U1787 ( .A0(n1577), .A1(n1647), .B0(n1576), .B1(n1575), .Y(n1580)
         );
  AOI32X1TS U1788 ( .A0(n1580), .A1(n1579), .A2(n1578), .B0(n1684), .B1(n1952), 
        .Y(n2079) );
  INVX2TS U1789 ( .A(n1569), .Y(n1656) );
  AOI22X1TS U1790 ( .A0(n1582), .A1(n1594), .B0(n1593), .B1(n1581), .Y(n1584)
         );
  AOI22X1TS U1791 ( .A0(n1585), .A1(n1656), .B0(n1584), .B1(n1583), .Y(n1587)
         );
  AOI22X1TS U1792 ( .A0(n1588), .A1(n1612), .B0(n1587), .B1(n1586), .Y(n1591)
         );
  AOI32X1TS U1793 ( .A0(n1591), .A1(n1590), .A2(n1589), .B0(n1714), .B1(n1953), 
        .Y(n2080) );
  AOI22X1TS U1794 ( .A0(n1595), .A1(n1594), .B0(n1593), .B1(n1592), .Y(n1597)
         );
  AOI22X1TS U1795 ( .A0(n1598), .A1(n1656), .B0(n1597), .B1(n1596), .Y(n1600)
         );
  AOI22X1TS U1796 ( .A0(n1601), .A1(n1612), .B0(n1600), .B1(n1599), .Y(n1604)
         );
  AOI32X1TS U1797 ( .A0(n1604), .A1(n1603), .A2(n1602), .B0(n1749), .B1(n1954), 
        .Y(n2081) );
  CLKBUFX2TS U1798 ( .A(n1652), .Y(n1639) );
  AOI22X1TS U1799 ( .A0(n1606), .A1(n1639), .B0(n1627), .B1(n1605), .Y(n1608)
         );
  AOI22X1TS U1800 ( .A0(n1609), .A1(n1643), .B0(n1608), .B1(n1607), .Y(n1611)
         );
  AOI22X1TS U1801 ( .A0(n1613), .A1(n1612), .B0(n1611), .B1(n1610), .Y(n1616)
         );
  AOI32X1TS U1802 ( .A0(n1616), .A1(n1615), .A2(n1614), .B0(n1778), .B1(n1955), 
        .Y(n2082) );
  AOI22X1TS U1803 ( .A0(n112), .A1(n1639), .B0(readIn_NORTH), .B1(n25), .Y(
        n1618) );
  AOI22X1TS U1804 ( .A0(n1619), .A1(n1643), .B0(n1618), .B1(n1617), .Y(n1621)
         );
  AOI22X1TS U1805 ( .A0(n1622), .A1(readIn_WEST), .B0(n1621), .B1(n1620), .Y(
        n1625) );
  AOI32X1TS U1806 ( .A0(n1625), .A1(n1624), .A2(n1623), .B0(n1805), .B1(n1956), 
        .Y(n2083) );
  AOI22X1TS U1807 ( .A0(n1628), .A1(n1639), .B0(n1627), .B1(n1626), .Y(n1630)
         );
  AOI22X1TS U1808 ( .A0(n1631), .A1(n1656), .B0(n1630), .B1(n1629), .Y(n1633)
         );
  AOI22X1TS U1809 ( .A0(n1634), .A1(readIn_WEST), .B0(n1633), .B1(n1632), .Y(
        n1637) );
  AOI32X1TS U1810 ( .A0(n1637), .A1(n1636), .A2(n1635), .B0(n1834), .B1(n1957), 
        .Y(n2084) );
  AOI22X1TS U1811 ( .A0(n1640), .A1(n1639), .B0(readIn_NORTH), .B1(n1638), .Y(
        n1642) );
  AOI22X1TS U1812 ( .A0(n1644), .A1(n1643), .B0(n1642), .B1(n1641), .Y(n1646)
         );
  AOI22X1TS U1813 ( .A0(n1648), .A1(n1647), .B0(n1646), .B1(n1645), .Y(n1650)
         );
  AOI32X1TS U1814 ( .A0(n1650), .A1(n350), .A2(n1649), .B0(n1874), .B1(n1958), 
        .Y(n2085) );
  AOI22X1TS U1815 ( .A0(n1653), .A1(n1652), .B0(readIn_NORTH), .B1(n1651), .Y(
        n1655) );
  AOI22X1TS U1816 ( .A0(n1657), .A1(n1656), .B0(n1655), .B1(n1654), .Y(n1659)
         );
  AOI22X1TS U1817 ( .A0(n1660), .A1(readIn_WEST), .B0(n1659), .B1(n1658), .Y(
        n1662) );
  AOI32X1TS U1818 ( .A0(n1662), .A1(n425), .A2(n1661), .B0(n1913), .B1(n1959), 
        .Y(n2086) );
  AOI22X1TS U1819 ( .A0(n1841), .A1(n1663), .B0(n1677), .B1(
        \destinationAddressbuffer[7][0] ), .Y(n1668) );
  AOI22X1TS U1820 ( .A0(n1664), .A1(n1723), .B0(n31), .B1(n1722), .Y(n1667) );
  CLKBUFX2TS U1821 ( .A(n1693), .Y(n1845) );
  AOI22X1TS U1822 ( .A0(n1665), .A1(destinationAddressIn_SOUTH[0]), .B0(n1673), 
        .B1(n1845), .Y(n1666) );
  AOI22X1TS U1823 ( .A0(n1670), .A1(n1669), .B0(n1677), .B1(
        \destinationAddressbuffer[7][1] ), .Y(n1676) );
  AOI22X1TS U1824 ( .A0(n1672), .A1(n1731), .B0(n1671), .B1(n1729), .Y(n1675)
         );
  CLKBUFX2TS U1825 ( .A(n1701), .Y(n1856) );
  AOI22X1TS U1826 ( .A0(n65), .A1(destinationAddressIn_SOUTH[1]), .B0(n1673), 
        .B1(n1856), .Y(n1674) );
  AOI22X1TS U1827 ( .A0(n1663), .A1(n1678), .B0(n1677), .B1(
        \destinationAddressbuffer[7][2] ), .Y(n1683) );
  AOI22X1TS U1828 ( .A0(n1679), .A1(n1742), .B0(n31), .B1(n1740), .Y(n1682) );
  CLKBUFX2TS U1829 ( .A(n1709), .Y(n1869) );
  AOI22X1TS U1830 ( .A0(n1680), .A1(destinationAddressIn_SOUTH[2]), .B0(n890), 
        .B1(n1869), .Y(n1681) );
  AOI22X1TS U1831 ( .A0(n1686), .A1(n1685), .B0(n1684), .B1(
        \destinationAddressbuffer[7][3] ), .Y(n1692) );
  AOI22X1TS U1832 ( .A0(n34), .A1(n1752), .B0(n1687), .B1(n1751), .Y(n1691) );
  CLKBUFX2TS U1833 ( .A(n1717), .Y(n1879) );
  AOI22X1TS U1834 ( .A0(n1689), .A1(destinationAddressIn_SOUTH[3]), .B0(n1688), 
        .B1(n1879), .Y(n1690) );
  AOI22X1TS U1835 ( .A0(n1884), .A1(n1715), .B0(n1707), .B1(
        \destinationAddressbuffer[6][0] ), .Y(n1697) );
  AOI22X1TS U1836 ( .A0(n90), .A1(n1723), .B0(n74), .B1(n1722), .Y(n1696) );
  CLKBUFX2TS U1837 ( .A(n1693), .Y(n1886) );
  CLKBUFX2TS U1838 ( .A(destinationAddressIn_SOUTH[0]), .Y(n1887) );
  CLKBUFX2TS U1839 ( .A(n1887), .Y(n1844) );
  AOI22X1TS U1840 ( .A0(n1694), .A1(n1886), .B0(n105), .B1(n1844), .Y(n1695)
         );
  AOI22X1TS U1841 ( .A0(n1762), .A1(n1698), .B0(n1707), .B1(
        \destinationAddressbuffer[6][1] ), .Y(n1706) );
  AOI22X1TS U1842 ( .A0(n1700), .A1(n1731), .B0(n1699), .B1(n1729), .Y(n1705)
         );
  CLKBUFX2TS U1843 ( .A(n1701), .Y(n1895) );
  CLKBUFX2TS U1844 ( .A(destinationAddressIn_SOUTH[1]), .Y(n1897) );
  CLKBUFX2TS U1845 ( .A(n1897), .Y(n1855) );
  AOI22X1TS U1846 ( .A0(n1703), .A1(n1895), .B0(n1702), .B1(n1855), .Y(n1704)
         );
  AOI22X1TS U1847 ( .A0(n1772), .A1(n76), .B0(n1707), .B1(
        \destinationAddressbuffer[6][2] ), .Y(n1713) );
  AOI22X1TS U1848 ( .A0(n90), .A1(n1742), .B0(n1708), .B1(n1740), .Y(n1712) );
  CLKBUFX2TS U1849 ( .A(n1709), .Y(n1907) );
  CLKBUFX2TS U1850 ( .A(destinationAddressIn_SOUTH[2]), .Y(n1909) );
  CLKBUFX2TS U1851 ( .A(n1909), .Y(n1867) );
  AOI22X1TS U1852 ( .A0(n1710), .A1(n1907), .B0(n105), .B1(n1867), .Y(n1711)
         );
  AOI22X1TS U1853 ( .A0(n1779), .A1(n1715), .B0(n1714), .B1(
        \destinationAddressbuffer[6][3] ), .Y(n1721) );
  AOI22X1TS U1854 ( .A0(n1716), .A1(n1752), .B0(n74), .B1(n1751), .Y(n1720) );
  CLKBUFX2TS U1855 ( .A(n1717), .Y(n1916) );
  CLKBUFX2TS U1856 ( .A(destinationAddressIn_SOUTH[3]), .Y(n1917) );
  CLKBUFX2TS U1857 ( .A(n1917), .Y(n1877) );
  AOI22X1TS U1858 ( .A0(n100), .A1(n1916), .B0(n1718), .B1(n1877), .Y(n1719)
         );
  AOI22X1TS U1859 ( .A0(n1884), .A1(n1750), .B0(n1738), .B1(
        \destinationAddressbuffer[5][0] ), .Y(n1727) );
  AOI22X1TS U1860 ( .A0(n1743), .A1(n1723), .B0(n213), .B1(n1722), .Y(n1726)
         );
  AOI22X1TS U1861 ( .A0(n1724), .A1(n1886), .B0(n1733), .B1(
        destinationAddressIn_SOUTH[0]), .Y(n1725) );
  AOI22X1TS U1862 ( .A0(readRequesterAddress[1]), .A1(n1728), .B0(n1738), .B1(
        \destinationAddressbuffer[5][1] ), .Y(n1737) );
  AOI22X1TS U1863 ( .A0(n1732), .A1(n1731), .B0(n1730), .B1(n1729), .Y(n1736)
         );
  AOI22X1TS U1864 ( .A0(n1734), .A1(n1895), .B0(n1733), .B1(
        destinationAddressIn_SOUTH[1]), .Y(n1735) );
  AOI22X1TS U1865 ( .A0(readRequesterAddress[2]), .A1(n1739), .B0(n1738), .B1(
        \destinationAddressbuffer[5][2] ), .Y(n1748) );
  AOI22X1TS U1866 ( .A0(n1743), .A1(n1742), .B0(n1741), .B1(n1740), .Y(n1747)
         );
  AOI22X1TS U1867 ( .A0(n1745), .A1(n1907), .B0(n1744), .B1(
        destinationAddressIn_SOUTH[2]), .Y(n1746) );
  AOI22X1TS U1868 ( .A0(readRequesterAddress[3]), .A1(n1750), .B0(n1749), .B1(
        \destinationAddressbuffer[5][3] ), .Y(n1755) );
  AOI22X1TS U1869 ( .A0(n232), .A1(n1752), .B0(n213), .B1(n1751), .Y(n1754) );
  AOI22X1TS U1870 ( .A0(n241), .A1(n1916), .B0(n1733), .B1(
        destinationAddressIn_SOUTH[3]), .Y(n1753) );
  AOI22X1TS U1871 ( .A0(n1785), .A1(n268), .B0(n1770), .B1(
        \destinationAddressbuffer[4][0] ), .Y(n1760) );
  AOI22X1TS U1872 ( .A0(n1756), .A1(n1786), .B0(n266), .B1(
        destinationAddressIn_EAST[0]), .Y(n1759) );
  AOI22X1TS U1873 ( .A0(n280), .A1(n1887), .B0(n1757), .B1(n1886), .Y(n1758)
         );
  AOI22X1TS U1874 ( .A0(n1762), .A1(n1761), .B0(n1770), .B1(
        \destinationAddressbuffer[4][1] ), .Y(n1769) );
  AOI22X1TS U1875 ( .A0(n1764), .A1(n1793), .B0(n1763), .B1(
        destinationAddressIn_EAST[1]), .Y(n1768) );
  AOI22X1TS U1876 ( .A0(n1766), .A1(n1897), .B0(n1765), .B1(n1895), .Y(n1767)
         );
  AOI22X1TS U1877 ( .A0(n1772), .A1(n1771), .B0(n1770), .B1(
        \destinationAddressbuffer[4][2] ), .Y(n1777) );
  AOI22X1TS U1878 ( .A0(n1774), .A1(n1800), .B0(n1773), .B1(
        destinationAddressIn_EAST[2]), .Y(n1776) );
  AOI22X1TS U1879 ( .A0(n280), .A1(n1909), .B0(n291), .B1(n1907), .Y(n1775) );
  AOI22X1TS U1880 ( .A0(n1779), .A1(n268), .B0(n1778), .B1(
        \destinationAddressbuffer[4][3] ), .Y(n1784) );
  AOI22X1TS U1881 ( .A0(n288), .A1(n1808), .B0(n266), .B1(
        destinationAddressIn_EAST[3]), .Y(n1783) );
  AOI22X1TS U1882 ( .A0(n1781), .A1(n1917), .B0(n1780), .B1(n1916), .Y(n1782)
         );
  AOI22X1TS U1883 ( .A0(n1785), .A1(n1806), .B0(n1799), .B1(
        \destinationAddressbuffer[3][0] ), .Y(n1790) );
  AOI22X1TS U1884 ( .A0(n1787), .A1(n1786), .B0(n1792), .B1(
        destinationAddressIn_EAST[0]), .Y(n1789) );
  AOI22X1TS U1885 ( .A0(n158), .A1(n1845), .B0(n1384), .B1(n1844), .Y(n1788)
         );
  AOI22X1TS U1886 ( .A0(n1851), .A1(n1791), .B0(n1799), .B1(
        \destinationAddressbuffer[3][1] ), .Y(n1798) );
  AOI22X1TS U1887 ( .A0(n1794), .A1(n1793), .B0(n1792), .B1(
        destinationAddressIn_EAST[1]), .Y(n1797) );
  AOI22X1TS U1888 ( .A0(n1795), .A1(n1856), .B0(n1810), .B1(n1855), .Y(n1796)
         );
  AOI22X1TS U1889 ( .A0(n1863), .A1(n122), .B0(n1799), .B1(
        \destinationAddressbuffer[3][2] ), .Y(n1804) );
  AOI22X1TS U1890 ( .A0(n135), .A1(n1800), .B0(n163), .B1(
        destinationAddressIn_EAST[2]), .Y(n1803) );
  AOI22X1TS U1891 ( .A0(n1801), .A1(n1869), .B0(n121), .B1(n1867), .Y(n1802)
         );
  AOI22X1TS U1892 ( .A0(n1875), .A1(n1806), .B0(n1805), .B1(
        \destinationAddressbuffer[3][3] ), .Y(n1813) );
  AOI22X1TS U1893 ( .A0(n1809), .A1(n1808), .B0(n1807), .B1(
        destinationAddressIn_EAST[3]), .Y(n1812) );
  AOI22X1TS U1894 ( .A0(n158), .A1(n1879), .B0(n1810), .B1(n1877), .Y(n1811)
         );
  AOI22X1TS U1895 ( .A0(n1841), .A1(n1835), .B0(n1825), .B1(
        \destinationAddressbuffer[2][0] ), .Y(n1817) );
  AOI22X1TS U1896 ( .A0(n1814), .A1(destinationAddressIn_WEST[0]), .B0(n999), 
        .B1(n1842), .Y(n1816) );
  AOI22X1TS U1897 ( .A0(n200), .A1(n1845), .B0(n1829), .B1(n1844), .Y(n1815)
         );
  AOI22X1TS U1898 ( .A0(n1892), .A1(n1818), .B0(n1825), .B1(
        \destinationAddressbuffer[2][1] ), .Y(n1824) );
  AOI22X1TS U1899 ( .A0(n1820), .A1(destinationAddressIn_WEST[1]), .B0(n1819), 
        .B1(n1852), .Y(n1823) );
  AOI22X1TS U1900 ( .A0(n1821), .A1(n1856), .B0(n193), .B1(n1855), .Y(n1822)
         );
  AOI22X1TS U1901 ( .A0(n1904), .A1(n1826), .B0(n1825), .B1(
        \destinationAddressbuffer[2][2] ), .Y(n1833) );
  AOI22X1TS U1902 ( .A0(n1828), .A1(destinationAddressIn_WEST[2]), .B0(n1827), 
        .B1(n1864), .Y(n1832) );
  AOI22X1TS U1903 ( .A0(n1830), .A1(n1869), .B0(n1829), .B1(n1867), .Y(n1831)
         );
  AOI22X1TS U1904 ( .A0(n1915), .A1(n1835), .B0(n1834), .B1(
        \destinationAddressbuffer[2][3] ), .Y(n1840) );
  AOI22X1TS U1905 ( .A0(n196), .A1(destinationAddressIn_WEST[3]), .B0(n171), 
        .B1(n1876), .Y(n1839) );
  AOI22X1TS U1906 ( .A0(n1837), .A1(n1879), .B0(n1836), .B1(n1877), .Y(n1838)
         );
  AOI22X1TS U1907 ( .A0(n1841), .A1(n311), .B0(n1861), .B1(
        \destinationAddressbuffer[1][0] ), .Y(n1849) );
  AOI22X1TS U1908 ( .A0(n1843), .A1(destinationAddressIn_WEST[0]), .B0(n1026), 
        .B1(n1842), .Y(n1848) );
  AOI22X1TS U1909 ( .A0(n1846), .A1(n1845), .B0(n1868), .B1(n1844), .Y(n1847)
         );
  AOI22X1TS U1910 ( .A0(n1851), .A1(n1850), .B0(n1861), .B1(
        \destinationAddressbuffer[1][1] ), .Y(n1860) );
  AOI22X1TS U1911 ( .A0(n1854), .A1(destinationAddressIn_WEST[1]), .B0(n1853), 
        .B1(n1852), .Y(n1859) );
  AOI22X1TS U1912 ( .A0(n1857), .A1(n1856), .B0(n320), .B1(n1855), .Y(n1858)
         );
  AOI22X1TS U1913 ( .A0(n1863), .A1(n1862), .B0(n1861), .B1(
        \destinationAddressbuffer[1][2] ), .Y(n1873) );
  AOI22X1TS U1914 ( .A0(n1866), .A1(destinationAddressIn_WEST[2]), .B0(n1865), 
        .B1(n1864), .Y(n1872) );
  AOI22X1TS U1915 ( .A0(n1870), .A1(n1869), .B0(n1868), .B1(n1867), .Y(n1871)
         );
  AOI22X1TS U1916 ( .A0(n1875), .A1(n311), .B0(n1874), .B1(
        \destinationAddressbuffer[1][3] ), .Y(n1883) );
  AOI22X1TS U1917 ( .A0(n372), .A1(destinationAddressIn_WEST[3]), .B0(n309), 
        .B1(n1876), .Y(n1882) );
  AOI22X1TS U1918 ( .A0(n1880), .A1(n1879), .B0(n1878), .B1(n1877), .Y(n1881)
         );
  AOI22X1TS U1919 ( .A0(n1884), .A1(n1914), .B0(n1902), .B1(
        \destinationAddressbuffer[0][0] ), .Y(n1890) );
  AOI22X1TS U1920 ( .A0(n1885), .A1(destinationAddressIn_WEST[0]), .B0(n405), 
        .B1(destinationAddressIn_EAST[0]), .Y(n1889) );
  AOI22X1TS U1921 ( .A0(n1898), .A1(n1887), .B0(n1896), .B1(n1886), .Y(n1888)
         );
  AOI22X1TS U1922 ( .A0(n1892), .A1(n1891), .B0(n1902), .B1(
        \destinationAddressbuffer[0][1] ), .Y(n1901) );
  AOI22X1TS U1923 ( .A0(n1894), .A1(destinationAddressIn_WEST[1]), .B0(n1893), 
        .B1(destinationAddressIn_EAST[1]), .Y(n1900) );
  AOI22X1TS U1924 ( .A0(n1898), .A1(n1897), .B0(n1896), .B1(n1895), .Y(n1899)
         );
  AOI22X1TS U1925 ( .A0(n1904), .A1(n1903), .B0(n1902), .B1(
        \destinationAddressbuffer[0][2] ), .Y(n1912) );
  AOI22X1TS U1926 ( .A0(n1906), .A1(destinationAddressIn_WEST[2]), .B0(n1905), 
        .B1(destinationAddressIn_EAST[2]), .Y(n1911) );
  AOI22X1TS U1927 ( .A0(n443), .A1(n1909), .B0(n1908), .B1(n1907), .Y(n1910)
         );
  AOI22X1TS U1928 ( .A0(n1915), .A1(n1914), .B0(n1913), .B1(
        \destinationAddressbuffer[0][3] ), .Y(n1921) );
  AOI22X1TS U1929 ( .A0(n426), .A1(destinationAddressIn_WEST[3]), .B0(n1053), 
        .B1(destinationAddressIn_EAST[3]), .Y(n1920) );
  AOI22X1TS U1930 ( .A0(n1918), .A1(n1917), .B0(n408), .B1(n1916), .Y(n1919)
         );
endmodule


module router ( clk, reset, localRouterAddress, destinationAddressIn_NORTH, 
        requesterAddressIn_NORTH, readIn_NORTH, writeIn_NORTH, dataIn_NORTH, 
        destinationAddressOut_NORTH, requesterAddressOut_NORTH, readOut_NORTH, 
        writeOut_NORTH, dataOut_NORTH, destinationAddressIn_SOUTH, 
        requesterAddressIn_SOUTH, readIn_SOUTH, writeIn_SOUTH, dataIn_SOUTH, 
        destinationAddressOut_SOUTH, requesterAddressOut_SOUTH, readOut_SOUTH, 
        writeOut_SOUTH, dataOut_SOUTH, destinationAddressIn_EAST, 
        requesterAddressIn_EAST, readIn_EAST, writeIn_EAST, dataIn_EAST, 
        destinationAddressOut_EAST, requesterAddressOut_EAST, readOut_EAST, 
        writeOut_EAST, dataOut_EAST, destinationAddressIn_WEST, 
        requesterAddressIn_WEST, readIn_WEST, writeIn_WEST, dataIn_WEST, 
        destinationAddressOut_WEST, requesterAddressOut_WEST, readOut_WEST, 
        writeOut_WEST, dataOut_WEST, cacheDataIn_A, cacheAddressIn_A, 
        cacheDataOut_A, memWrite_A, cacheDataIn_B, cacheAddressIn_B, 
        cacheDataOut_B, memWrite_B );
  input [3:0] localRouterAddress;
  input [11:0] destinationAddressIn_NORTH;
  input [3:0] requesterAddressIn_NORTH;
  input [5:0] dataIn_NORTH;
  output [11:0] destinationAddressOut_NORTH;
  output [3:0] requesterAddressOut_NORTH;
  output [5:0] dataOut_NORTH;
  input [11:0] destinationAddressIn_SOUTH;
  input [3:0] requesterAddressIn_SOUTH;
  input [5:0] dataIn_SOUTH;
  output [11:0] destinationAddressOut_SOUTH;
  output [3:0] requesterAddressOut_SOUTH;
  output [5:0] dataOut_SOUTH;
  input [11:0] destinationAddressIn_EAST;
  input [3:0] requesterAddressIn_EAST;
  input [5:0] dataIn_EAST;
  output [11:0] destinationAddressOut_EAST;
  output [3:0] requesterAddressOut_EAST;
  output [5:0] dataOut_EAST;
  input [11:0] destinationAddressIn_WEST;
  input [3:0] requesterAddressIn_WEST;
  input [5:0] dataIn_WEST;
  output [11:0] destinationAddressOut_WEST;
  output [3:0] requesterAddressOut_WEST;
  output [5:0] dataOut_WEST;
  output [5:0] cacheDataIn_A;
  output [7:0] cacheAddressIn_A;
  input [5:0] cacheDataOut_A;
  output [5:0] cacheDataIn_B;
  output [7:0] cacheAddressIn_B;
  input [5:0] cacheDataOut_B;
  input clk, reset, readIn_NORTH, writeIn_NORTH, readIn_SOUTH, writeIn_SOUTH,
         readIn_EAST, writeIn_EAST, readIn_WEST, writeIn_WEST;
  output readOut_NORTH, writeOut_NORTH, readOut_SOUTH, writeOut_SOUTH,
         readOut_EAST, writeOut_EAST, readOut_WEST, writeOut_WEST, memWrite_A,
         memWrite_B;
  wire   readInBuffer_NORTH, writeInBuffer_NORTH, memRead_NORTH,
         memWrite_NORTH, readInBuffer_SOUTH, writeInBuffer_SOUTH,
         memRead_SOUTH, memWrite_SOUTH, readInBuffer_EAST, writeInBuffer_EAST,
         memRead_EAST, memWrite_EAST, readInBuffer_WEST, writeInBuffer_WEST,
         memRead_WEST, memWrite_WEST, readReady_NORTH, readReady_SOUTH,
         readReady_EAST, readReady_WEST, N4, N5, N6, N7, N8, N9, N10, N11, N12,
         N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26,
         N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40,
         N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54,
         N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68,
         N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82,
         N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96,
         N97, N98, N99, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670;
  wire   [3:0] outputPortSelect_NORTH;
  wire   [3:0] outputPortSelect_SOUTH;
  wire   [3:0] outputPortSelect_EAST;
  wire   [3:0] outputPortSelect_WEST;
  wire   [11:0] destinationAddressInBuffer_NORTH;
  wire   [3:0] requesterAddressInBuffer_NORTH;
  wire   [5:0] dataInBuffer_NORTH;
  wire   [3:0] cacheRequesterAddress_NORTH;
  wire   [5:0] cacheDataOut_NORTH;
  wire   [11:0] destinationAddressInBuffer_SOUTH;
  wire   [3:0] requesterAddressInBuffer_SOUTH;
  wire   [5:0] dataInBuffer_SOUTH;
  wire   [3:0] cacheRequesterAddress_SOUTH;
  wire   [5:0] cacheDataOut_SOUTH;
  wire   [11:0] destinationAddressInBuffer_EAST;
  wire   [3:0] requesterAddressInBuffer_EAST;
  wire   [5:0] dataInBuffer_EAST;
  wire   [3:0] cacheRequesterAddress_EAST;
  wire   [5:0] cacheDataOut_EAST;
  wire   [11:0] destinationAddressInBuffer_WEST;
  wire   [3:0] requesterAddressInBuffer_WEST;
  wire   [5:0] dataInBuffer_WEST;
  wire   [3:0] cacheRequesterAddress_WEST;
  wire   [5:0] cacheDataOut_WEST;

  cacheAccessArbiter cacheController ( .clk(clk), .reset(n670), 
        .cacheAddressIn_NORTH({n431, n430, n429, n428, n427, n425, n423, n421}), .requesterAddressIn_NORTH({n641, n637, n633, n629}), .memRead_NORTH(
        memRead_NORTH), .memWrite_NORTH(memWrite_NORTH), .dataIn_NORTH({n419, 
        n417, n415, n413, n411, n409}), .readReady_NORTH(readReady_NORTH), 
        .requesterAddressOut_NORTH(cacheRequesterAddress_NORTH), 
        .cacheDataOut_NORTH(cacheDataOut_NORTH), .cacheAddressIn_SOUTH({n625, 
        n623, n621, n619, n617, n612, n607, n602}), .requesterAddressIn_SOUTH(
        {n407, n405, n403, n401}), .memRead_SOUTH(memRead_SOUTH), 
        .memWrite_SOUTH(memWrite_SOUTH), .dataIn_SOUTH({n597, n592, n587, n582, 
        n577, n572}), .readReady_SOUTH(readReady_SOUTH), 
        .requesterAddressOut_SOUTH(cacheRequesterAddress_SOUTH), 
        .cacheDataOut_SOUTH(cacheDataOut_SOUTH), .cacheAddressIn_EAST({n381, 
        n379, n377, n375, n567, n562, n557, n552}), .requesterAddressIn_EAST({
        n547, n546, n545, n544}), .memRead_EAST(memRead_EAST), .memWrite_EAST(
        n291), .dataIn_EAST({n543, n538, n533, n528, n523, n518}), 
        .readReady_EAST(readReady_EAST), .requesterAddressOut_EAST(
        cacheRequesterAddress_EAST), .cacheDataOut_EAST(cacheDataOut_EAST), 
        .cacheAddressIn_WEST({n513, n509, n505, n501, n497, n493, n489, n485}), 
        .requesterAddressIn_WEST({n481, n476, n471, n466}), .memRead_WEST(
        memRead_WEST), .memWrite_WEST(n328), .dataIn_WEST({n461, n457, n453, 
        n449, n445, n441}), .readReady_WEST(readReady_WEST), 
        .requesterAddressOut_WEST(cacheRequesterAddress_WEST), 
        .cacheDataOut_WEST(cacheDataOut_WEST), .cacheDataIn_A(cacheDataIn_A), 
        .cacheAddressIn_A(cacheAddressIn_A), .cacheDataOut_A(cacheDataOut_A), 
        .memWrite_A(memWrite_A), .cacheDataIn_B(cacheDataIn_B), 
        .cacheAddressIn_B(cacheAddressIn_B), .cacheDataOut_B(cacheDataOut_B), 
        .memWrite_B(memWrite_B) );
  outputPortArbiter_0 outNorth ( .clk(clk), .reset(n668), .selectBit_NORTH(
        n350), .destinationAddressIn_NORTH({
        destinationAddressInBuffer_NORTH[11:8], n657, n653, n649, n645, 
        destinationAddressInBuffer_NORTH[3:0]}), .requesterAddressIn_NORTH({
        n641, n637, n633, n629}), .readIn_NORTH(n434), .writeIn_NORTH(n663), 
        .dataIn_NORTH(dataInBuffer_NORTH), .selectBit_SOUTH(n362), 
        .destinationAddressIn_SOUTH({destinationAddressInBuffer_SOUTH[11:8], 
        n624, n622, n620, n618, n616, n611, n606, n601}), 
        .requesterAddressIn_SOUTH(requesterAddressInBuffer_SOUTH), 
        .readIn_SOUTH(n435), .writeIn_SOUTH(n662), .dataIn_SOUTH({n596, n591, 
        n586, n581, n576, n571}), .selectBit_EAST(n387), 
        .destinationAddressIn_EAST({n374, n371, n368, n365, n357, n355, n353, 
        n351, n566, n561, n556, n551}), .requesterAddressIn_EAST({n399, n397, 
        n395, n393}), .readIn_EAST(n390), .writeIn_EAST(n386), .dataIn_EAST({
        n542, n537, n532, n527, n522, n517}), .selectBit_WEST(
        outputPortSelect_WEST[0]), .destinationAddressIn_WEST({
        destinationAddressInBuffer_WEST[11:8], n513, n509, n505, n501, n497, 
        n493, n489, n485}), .requesterAddressIn_WEST({n480, n475, n470, n465}), 
        .readIn_WEST(n437), .writeIn_WEST(n658), .dataIn_WEST({n461, n457, 
        n453, n449, n445, n441}), .readReady(readReady_NORTH), 
        .readRequesterAddress(cacheRequesterAddress_NORTH), .cacheDataOut(
        cacheDataOut_NORTH), .destinationAddressOut(
        destinationAddressOut_NORTH), .requesterAddressOut(
        requesterAddressOut_NORTH), .readOut(readOut_NORTH), .writeOut(
        writeOut_NORTH), .dataOut(dataOut_NORTH) );
  outputPortArbiter_3 outSouth ( .clk(clk), .reset(n669), .selectBit_NORTH(
        n349), .destinationAddressIn_NORTH({
        destinationAddressInBuffer_NORTH[11:8], n654, n650, n646, n642, n426, 
        n424, n422, n420}), .requesterAddressIn_NORTH({n638, n634, n630, n626}), .readIn_NORTH(n665), .writeIn_NORTH(n433), .dataIn_NORTH({n418, n416, n414, 
        n412, n410, n408}), .selectBit_SOUTH(n360), 
        .destinationAddressIn_SOUTH({destinationAddressInBuffer_SOUTH[11:8], 
        n624, n622, n620, n618, n613, n608, n603, n598}), 
        .requesterAddressIn_SOUTH({n406, n404, n402, n400}), .readIn_SOUTH(
        n432), .writeIn_SOUTH(n662), .dataIn_SOUTH({n593, n588, n583, n578, 
        n573, n568}), .selectBit_EAST(n388), .destinationAddressIn_EAST({
        destinationAddressInBuffer_EAST[11:4], n563, n558, n553, n548}), 
        .requesterAddressIn_EAST({n398, n396, n394, n392}), .readIn_EAST(n389), 
        .writeIn_EAST(n384), .dataIn_EAST({n539, n534, n529, n524, n519, n514}), .selectBit_WEST(outputPortSelect_WEST[1]), .destinationAddressIn_WEST({
        destinationAddressInBuffer_WEST[11:8], n510, n506, n502, n498, n494, 
        n490, n486, n482}), .requesterAddressIn_WEST({n477, n472, n467, n462}), 
        .readIn_WEST(n660), .writeIn_WEST(n436), .dataIn_WEST({n458, n454, 
        n450, n446, n442, n438}), .readReady(readReady_SOUTH), 
        .readRequesterAddress(cacheRequesterAddress_SOUTH), .cacheDataOut(
        cacheDataOut_SOUTH), .destinationAddressOut(
        destinationAddressOut_SOUTH), .requesterAddressOut(
        requesterAddressOut_SOUTH), .readOut(readOut_SOUTH), .writeOut(
        writeOut_SOUTH), .dataOut(dataOut_SOUTH) );
  outputPortArbiter_2 outEast ( .clk(clk), .reset(n670), .selectBit_NORTH(n348), .destinationAddressIn_NORTH({destinationAddressInBuffer_NORTH[11:8], n655, 
        n651, n647, n643, n426, n424, n422, n420}), .requesterAddressIn_NORTH(
        {n639, n635, n631, n627}), .readIn_NORTH(n666), .writeIn_NORTH(n433), 
        .dataIn_NORTH({n418, n416, n414, n412, n410, n408}), .selectBit_SOUTH(
        n359), .destinationAddressIn_SOUTH({
        destinationAddressInBuffer_SOUTH[11:8], n624, n622, n620, n618, n614, 
        n609, n604, n599}), .requesterAddressIn_SOUTH({n406, n404, n402, n400}), .readIn_SOUTH(n432), .writeIn_SOUTH(n662), .dataIn_SOUTH({n594, n589, n584, 
        n579, n574, n569}), .selectBit_EAST(n308), .destinationAddressIn_EAST(
        {n372, n369, n366, n363, n358, n356, n354, n352, n564, n559, n554, 
        n549}), .requesterAddressIn_EAST(requesterAddressInBuffer_EAST), 
        .readIn_EAST(n391), .writeIn_EAST(n383), .dataIn_EAST({n540, n535, 
        n530, n525, n520, n515}), .selectBit_WEST(outputPortSelect_WEST[2]), 
        .destinationAddressIn_WEST({destinationAddressInBuffer_WEST[11:8], 
        n511, n507, n503, n499, n495, n491, n487, n483}), 
        .requesterAddressIn_WEST({n478, n473, n468, n463}), .readIn_WEST(n661), 
        .writeIn_WEST(n436), .dataIn_WEST({n459, n455, n451, n447, n443, n439}), .readReady(readReady_EAST), .readRequesterAddress(cacheRequesterAddress_EAST), .cacheDataOut(cacheDataOut_EAST), .destinationAddressOut(
        destinationAddressOut_EAST), .requesterAddressOut(
        requesterAddressOut_EAST), .readOut(readOut_EAST), .writeOut(
        writeOut_EAST), .dataOut(dataOut_EAST) );
  outputPortArbiter_1 outWest ( .clk(clk), .reset(n667), .selectBit_NORTH(n255), .destinationAddressIn_NORTH({destinationAddressInBuffer_NORTH[11:8], n656, 
        n652, n648, n644, destinationAddressInBuffer_NORTH[3:0]}), 
        .requesterAddressIn_NORTH({n640, n636, n632, n628}), .readIn_NORTH(
        n434), .writeIn_NORTH(n664), .dataIn_NORTH(dataInBuffer_NORTH), 
        .selectBit_SOUTH(n361), .destinationAddressIn_SOUTH({
        destinationAddressInBuffer_SOUTH[11:8], n624, n622, n620, n618, n615, 
        n610, n605, n600}), .requesterAddressIn_SOUTH(
        requesterAddressInBuffer_SOUTH), .readIn_SOUTH(n435), .writeIn_SOUTH(
        n662), .dataIn_SOUTH({n595, n590, n585, n580, n575, n570}), 
        .selectBit_EAST(n310), .destinationAddressIn_EAST({n373, n370, n367, 
        n364, n382, n380, n378, n376, n565, n560, n555, n550}), 
        .requesterAddressIn_EAST(requesterAddressInBuffer_EAST), .readIn_EAST(
        n389), .writeIn_EAST(n385), .dataIn_EAST({n541, n536, n531, n526, n521, 
        n516}), .selectBit_WEST(outputPortSelect_WEST[3]), 
        .destinationAddressIn_WEST({destinationAddressInBuffer_WEST[11:8], 
        n512, n508, n504, n500, n496, n492, n488, n484}), 
        .requesterAddressIn_WEST({n479, n474, n469, n464}), .readIn_WEST(n437), 
        .writeIn_WEST(n659), .dataIn_WEST({n460, n456, n452, n448, n444, n440}), .readReady(readReady_WEST), .readRequesterAddress(cacheRequesterAddress_WEST), .cacheDataOut(cacheDataOut_WEST), .destinationAddressOut(
        destinationAddressOut_WEST), .requesterAddressOut(
        requesterAddressOut_WEST), .readOut(readOut_WEST), .writeOut(
        writeOut_WEST), .dataOut(dataOut_WEST) );
  DFFQX1TS writeInBuffer_SOUTH_reg ( .D(N45), .CK(clk), .Q(writeInBuffer_SOUTH) );
  DFFQX1TS \requesterAddressInBuffer_WEST_reg[3]  ( .D(N91), .CK(clk), .Q(
        requesterAddressInBuffer_WEST[3]) );
  DFFQX1TS \requesterAddressInBuffer_WEST_reg[2]  ( .D(N90), .CK(clk), .Q(
        requesterAddressInBuffer_WEST[2]) );
  DFFQX1TS \requesterAddressInBuffer_WEST_reg[1]  ( .D(N89), .CK(clk), .Q(
        requesterAddressInBuffer_WEST[1]) );
  DFFQX1TS \requesterAddressInBuffer_WEST_reg[0]  ( .D(N88), .CK(clk), .Q(
        requesterAddressInBuffer_WEST[0]) );
  DFFQX1TS \destinationAddressInBuffer_SOUTH_reg[3]  ( .D(N31), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[3]) );
  DFFQX1TS \destinationAddressInBuffer_EAST_reg[3]  ( .D(N55), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[3]) );
  DFFQX1TS \destinationAddressInBuffer_SOUTH_reg[2]  ( .D(N30), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[2]) );
  DFFQX1TS \destinationAddressInBuffer_EAST_reg[2]  ( .D(N54), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[2]) );
  DFFQX1TS \destinationAddressInBuffer_SOUTH_reg[1]  ( .D(N29), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[1]) );
  DFFQX1TS \destinationAddressInBuffer_EAST_reg[1]  ( .D(N53), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[1]) );
  DFFQX1TS \destinationAddressInBuffer_SOUTH_reg[0]  ( .D(N28), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[0]) );
  DFFQX1TS \destinationAddressInBuffer_EAST_reg[0]  ( .D(N52), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[0]) );
  DFFQX1TS \dataInBuffer_SOUTH_reg[5]  ( .D(N51), .CK(clk), .Q(
        dataInBuffer_SOUTH[5]) );
  DFFQX1TS \dataInBuffer_EAST_reg[5]  ( .D(N75), .CK(clk), .Q(
        dataInBuffer_EAST[5]) );
  DFFQX1TS \dataInBuffer_SOUTH_reg[4]  ( .D(N50), .CK(clk), .Q(
        dataInBuffer_SOUTH[4]) );
  DFFQX1TS \dataInBuffer_EAST_reg[4]  ( .D(N74), .CK(clk), .Q(
        dataInBuffer_EAST[4]) );
  DFFQX1TS \dataInBuffer_SOUTH_reg[3]  ( .D(N49), .CK(clk), .Q(
        dataInBuffer_SOUTH[3]) );
  DFFQX1TS \dataInBuffer_EAST_reg[3]  ( .D(N73), .CK(clk), .Q(
        dataInBuffer_EAST[3]) );
  DFFQX1TS \dataInBuffer_SOUTH_reg[2]  ( .D(N48), .CK(clk), .Q(
        dataInBuffer_SOUTH[2]) );
  DFFQX1TS \dataInBuffer_EAST_reg[2]  ( .D(N72), .CK(clk), .Q(
        dataInBuffer_EAST[2]) );
  DFFQX1TS \dataInBuffer_SOUTH_reg[1]  ( .D(N47), .CK(clk), .Q(
        dataInBuffer_SOUTH[1]) );
  DFFQX1TS \dataInBuffer_EAST_reg[1]  ( .D(N71), .CK(clk), .Q(
        dataInBuffer_EAST[1]) );
  DFFQX1TS \dataInBuffer_SOUTH_reg[0]  ( .D(N46), .CK(clk), .Q(
        dataInBuffer_SOUTH[0]) );
  DFFQX1TS \dataInBuffer_EAST_reg[0]  ( .D(N70), .CK(clk), .Q(
        dataInBuffer_EAST[0]) );
  DFFQX1TS \destinationAddressInBuffer_NORTH_reg[7]  ( .D(N11), .CK(clk), .Q(
        destinationAddressInBuffer_NORTH[7]) );
  DFFQX1TS \destinationAddressInBuffer_NORTH_reg[6]  ( .D(N10), .CK(clk), .Q(
        destinationAddressInBuffer_NORTH[6]) );
  DFFQX1TS \destinationAddressInBuffer_NORTH_reg[5]  ( .D(N9), .CK(clk), .Q(
        destinationAddressInBuffer_NORTH[5]) );
  DFFQX1TS \destinationAddressInBuffer_NORTH_reg[4]  ( .D(N8), .CK(clk), .Q(
        destinationAddressInBuffer_NORTH[4]) );
  DFFQX1TS writeInBuffer_NORTH_reg ( .D(N21), .CK(clk), .Q(writeInBuffer_NORTH) );
  DFFQX1TS writeInBuffer_WEST_reg ( .D(N93), .CK(clk), .Q(writeInBuffer_WEST)
         );
  DFFQX1TS readInBuffer_WEST_reg ( .D(N92), .CK(clk), .Q(readInBuffer_WEST) );
  DFFQX1TS readInBuffer_NORTH_reg ( .D(N20), .CK(clk), .Q(readInBuffer_NORTH)
         );
  DFFQX1TS \destinationAddressInBuffer_WEST_reg[11]  ( .D(N87), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[11]) );
  DFFQX1TS \destinationAddressInBuffer_WEST_reg[10]  ( .D(N86), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[10]) );
  DFFQX1TS \destinationAddressInBuffer_WEST_reg[9]  ( .D(N85), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[9]) );
  DFFQX1TS \destinationAddressInBuffer_WEST_reg[8]  ( .D(N84), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[8]) );
  DFFQX1TS readInBuffer_EAST_reg ( .D(N68), .CK(clk), .Q(readInBuffer_EAST) );
  DFFQX1TS \destinationAddressInBuffer_EAST_reg[11]  ( .D(N63), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[11]) );
  DFFQX1TS \destinationAddressInBuffer_EAST_reg[10]  ( .D(N62), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[10]) );
  DFFQX1TS \destinationAddressInBuffer_EAST_reg[9]  ( .D(N61), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[9]) );
  DFFQX1TS \destinationAddressInBuffer_EAST_reg[8]  ( .D(N60), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[8]) );
  DFFQX1TS \destinationAddressInBuffer_SOUTH_reg[7]  ( .D(N35), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[7]) );
  DFFQX1TS \destinationAddressInBuffer_SOUTH_reg[6]  ( .D(N34), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[6]) );
  DFFQX1TS \destinationAddressInBuffer_SOUTH_reg[5]  ( .D(N33), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[5]) );
  DFFQX1TS \destinationAddressInBuffer_SOUTH_reg[4]  ( .D(N32), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[4]) );
  DFFQX1TS writeInBuffer_EAST_reg ( .D(N69), .CK(clk), .Q(writeInBuffer_EAST)
         );
  DFFQX1TS \destinationAddressInBuffer_EAST_reg[7]  ( .D(N59), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[7]) );
  DFFQX1TS \destinationAddressInBuffer_EAST_reg[6]  ( .D(N58), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[6]) );
  DFFQX1TS \destinationAddressInBuffer_EAST_reg[5]  ( .D(N57), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[5]) );
  DFFQX1TS \destinationAddressInBuffer_EAST_reg[4]  ( .D(N56), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[4]) );
  DFFQX1TS \destinationAddressInBuffer_SOUTH_reg[11]  ( .D(N39), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[11]) );
  DFFQX1TS \destinationAddressInBuffer_SOUTH_reg[10]  ( .D(N38), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[10]) );
  DFFQX1TS \destinationAddressInBuffer_SOUTH_reg[9]  ( .D(N37), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[9]) );
  DFFQX1TS \destinationAddressInBuffer_SOUTH_reg[8]  ( .D(N36), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[8]) );
  DFFQX1TS \destinationAddressInBuffer_NORTH_reg[11]  ( .D(N15), .CK(clk), .Q(
        destinationAddressInBuffer_NORTH[11]) );
  DFFQX1TS \destinationAddressInBuffer_NORTH_reg[10]  ( .D(N14), .CK(clk), .Q(
        destinationAddressInBuffer_NORTH[10]) );
  DFFQX1TS \destinationAddressInBuffer_NORTH_reg[9]  ( .D(N13), .CK(clk), .Q(
        destinationAddressInBuffer_NORTH[9]) );
  DFFQX1TS \destinationAddressInBuffer_NORTH_reg[8]  ( .D(N12), .CK(clk), .Q(
        destinationAddressInBuffer_NORTH[8]) );
  DFFQX1TS \destinationAddressInBuffer_NORTH_reg[3]  ( .D(N7), .CK(clk), .Q(
        destinationAddressInBuffer_NORTH[3]) );
  DFFQX1TS \destinationAddressInBuffer_NORTH_reg[2]  ( .D(N6), .CK(clk), .Q(
        destinationAddressInBuffer_NORTH[2]) );
  DFFQX1TS \destinationAddressInBuffer_NORTH_reg[1]  ( .D(N5), .CK(clk), .Q(
        destinationAddressInBuffer_NORTH[1]) );
  DFFQX1TS \destinationAddressInBuffer_NORTH_reg[0]  ( .D(N4), .CK(clk), .Q(
        destinationAddressInBuffer_NORTH[0]) );
  DFFQX1TS \dataInBuffer_NORTH_reg[5]  ( .D(N27), .CK(clk), .Q(
        dataInBuffer_NORTH[5]) );
  DFFQX1TS \dataInBuffer_NORTH_reg[4]  ( .D(N26), .CK(clk), .Q(
        dataInBuffer_NORTH[4]) );
  DFFQX1TS \dataInBuffer_NORTH_reg[3]  ( .D(N25), .CK(clk), .Q(
        dataInBuffer_NORTH[3]) );
  DFFQX1TS \dataInBuffer_NORTH_reg[2]  ( .D(N24), .CK(clk), .Q(
        dataInBuffer_NORTH[2]) );
  DFFQX1TS \dataInBuffer_NORTH_reg[1]  ( .D(N23), .CK(clk), .Q(
        dataInBuffer_NORTH[1]) );
  DFFQX1TS \dataInBuffer_NORTH_reg[0]  ( .D(N22), .CK(clk), .Q(
        dataInBuffer_NORTH[0]) );
  DFFQX1TS \requesterAddressInBuffer_SOUTH_reg[3]  ( .D(N43), .CK(clk), .Q(
        requesterAddressInBuffer_SOUTH[3]) );
  DFFQX1TS \requesterAddressInBuffer_SOUTH_reg[2]  ( .D(N42), .CK(clk), .Q(
        requesterAddressInBuffer_SOUTH[2]) );
  DFFQX1TS \requesterAddressInBuffer_SOUTH_reg[1]  ( .D(N41), .CK(clk), .Q(
        requesterAddressInBuffer_SOUTH[1]) );
  DFFQX1TS \requesterAddressInBuffer_SOUTH_reg[0]  ( .D(N40), .CK(clk), .Q(
        requesterAddressInBuffer_SOUTH[0]) );
  DFFQX1TS \requesterAddressInBuffer_EAST_reg[3]  ( .D(N67), .CK(clk), .Q(
        requesterAddressInBuffer_EAST[3]) );
  DFFQX1TS \requesterAddressInBuffer_EAST_reg[2]  ( .D(N66), .CK(clk), .Q(
        requesterAddressInBuffer_EAST[2]) );
  DFFQX1TS \requesterAddressInBuffer_EAST_reg[1]  ( .D(N65), .CK(clk), .Q(
        requesterAddressInBuffer_EAST[1]) );
  DFFQX1TS \requesterAddressInBuffer_EAST_reg[0]  ( .D(N64), .CK(clk), .Q(
        requesterAddressInBuffer_EAST[0]) );
  DFFQX1TS readInBuffer_SOUTH_reg ( .D(N44), .CK(clk), .Q(readInBuffer_SOUTH)
         );
  DFFQX1TS \dataInBuffer_WEST_reg[5]  ( .D(N99), .CK(clk), .Q(
        dataInBuffer_WEST[5]) );
  DFFQX1TS \dataInBuffer_WEST_reg[4]  ( .D(N98), .CK(clk), .Q(
        dataInBuffer_WEST[4]) );
  DFFQX1TS \dataInBuffer_WEST_reg[3]  ( .D(N97), .CK(clk), .Q(
        dataInBuffer_WEST[3]) );
  DFFQX1TS \dataInBuffer_WEST_reg[2]  ( .D(N96), .CK(clk), .Q(
        dataInBuffer_WEST[2]) );
  DFFQX1TS \dataInBuffer_WEST_reg[1]  ( .D(N95), .CK(clk), .Q(
        dataInBuffer_WEST[1]) );
  DFFQX1TS \dataInBuffer_WEST_reg[0]  ( .D(N94), .CK(clk), .Q(
        dataInBuffer_WEST[0]) );
  DFFQX1TS \requesterAddressInBuffer_NORTH_reg[3]  ( .D(N19), .CK(clk), .Q(
        requesterAddressInBuffer_NORTH[3]) );
  DFFQX1TS \requesterAddressInBuffer_NORTH_reg[2]  ( .D(N18), .CK(clk), .Q(
        requesterAddressInBuffer_NORTH[2]) );
  DFFQX1TS \requesterAddressInBuffer_NORTH_reg[1]  ( .D(N17), .CK(clk), .Q(
        requesterAddressInBuffer_NORTH[1]) );
  DFFQX1TS \requesterAddressInBuffer_NORTH_reg[0]  ( .D(N16), .CK(clk), .Q(
        requesterAddressInBuffer_NORTH[0]) );
  DFFQX1TS \destinationAddressInBuffer_WEST_reg[7]  ( .D(N83), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[7]) );
  DFFQX1TS \destinationAddressInBuffer_WEST_reg[6]  ( .D(N82), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[6]) );
  DFFQX1TS \destinationAddressInBuffer_WEST_reg[5]  ( .D(N81), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[5]) );
  DFFQX1TS \destinationAddressInBuffer_WEST_reg[4]  ( .D(N80), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[4]) );
  DFFQX1TS \destinationAddressInBuffer_WEST_reg[3]  ( .D(N79), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[3]) );
  DFFQX1TS \destinationAddressInBuffer_WEST_reg[2]  ( .D(N78), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[2]) );
  DFFQX1TS \destinationAddressInBuffer_WEST_reg[1]  ( .D(N77), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[1]) );
  DFFQX1TS \destinationAddressInBuffer_WEST_reg[0]  ( .D(N76), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[0]) );
  DFFQX1TS \inWest/memRead_reg  ( .D(n73), .CK(clk), .Q(memRead_WEST) );
  DFFQX1TS \inWest/memWrite_reg  ( .D(n78), .CK(clk), .Q(memWrite_WEST) );
  DFFQX1TS \inEast/memRead_reg  ( .D(n79), .CK(clk), .Q(memRead_EAST) );
  DFFQX1TS \inEast/memWrite_reg  ( .D(n84), .CK(clk), .Q(memWrite_EAST) );
  DFFHQX1TS \inNorth/outputPortSelect_reg[0]  ( .D(n95), .CK(clk), .Q(
        outputPortSelect_NORTH[0]) );
  DFFHQX1TS \inNorth/outputPortSelect_reg[3]  ( .D(n92), .CK(clk), .Q(
        outputPortSelect_NORTH[3]) );
  DFFHQX1TS \inNorth/outputPortSelect_reg[1]  ( .D(n94), .CK(clk), .Q(
        outputPortSelect_NORTH[1]) );
  DFFHQX1TS \inNorth/outputPortSelect_reg[2]  ( .D(n93), .CK(clk), .Q(
        outputPortSelect_NORTH[2]) );
  DFFHQX1TS \inSouth/outputPortSelect_reg[0]  ( .D(n89), .CK(clk), .Q(
        outputPortSelect_SOUTH[0]) );
  DFFHQX1TS \inSouth/outputPortSelect_reg[3]  ( .D(n86), .CK(clk), .Q(
        outputPortSelect_SOUTH[3]) );
  DFFHQX1TS \inSouth/outputPortSelect_reg[1]  ( .D(n88), .CK(clk), .Q(
        outputPortSelect_SOUTH[1]) );
  DFFHQX1TS \inSouth/outputPortSelect_reg[2]  ( .D(n87), .CK(clk), .Q(
        outputPortSelect_SOUTH[2]) );
  DFFHQX1TS \inEast/outputPortSelect_reg[0]  ( .D(n83), .CK(clk), .Q(
        outputPortSelect_EAST[0]) );
  DFFHQX1TS \inEast/outputPortSelect_reg[3]  ( .D(n80), .CK(clk), .Q(
        outputPortSelect_EAST[3]) );
  DFFHQX1TS \inEast/outputPortSelect_reg[1]  ( .D(n82), .CK(clk), .Q(
        outputPortSelect_EAST[1]) );
  DFFQX1TS \inSouth/memWrite_reg  ( .D(n90), .CK(clk), .Q(memWrite_SOUTH) );
  DFFQX1TS \inSouth/memRead_reg  ( .D(n85), .CK(clk), .Q(memRead_SOUTH) );
  DFFQX1TS \inWest/outputPortSelect_reg[2]  ( .D(n75), .CK(clk), .Q(
        outputPortSelect_WEST[2]) );
  DFFQX1TS \inWest/outputPortSelect_reg[3]  ( .D(n74), .CK(clk), .Q(
        outputPortSelect_WEST[3]) );
  DFFQX1TS \inWest/outputPortSelect_reg[0]  ( .D(n77), .CK(clk), .Q(
        outputPortSelect_WEST[0]) );
  DFFQX1TS \inWest/outputPortSelect_reg[1]  ( .D(n76), .CK(clk), .Q(
        outputPortSelect_WEST[1]) );
  DFFHQX1TS \inEast/outputPortSelect_reg[2]  ( .D(n81), .CK(clk), .Q(
        outputPortSelect_EAST[2]) );
  DFFQX1TS \inNorth/memRead_reg  ( .D(n91), .CK(clk), .Q(memRead_NORTH) );
  DFFQX1TS \inNorth/memWrite_reg  ( .D(n96), .CK(clk), .Q(memWrite_NORTH) );
  CLKBUFX2TS U258 ( .A(memWrite_WEST), .Y(n328) );
  CLKBUFX2TS U259 ( .A(memWrite_EAST), .Y(n291) );
  CLKBUFX2TS U260 ( .A(outputPortSelect_EAST[2]), .Y(n308) );
  CLKBUFX2TS U261 ( .A(outputPortSelect_EAST[3]), .Y(n310) );
  INVX2TS U262 ( .A(n236), .Y(n326) );
  INVX2TS U263 ( .A(n236), .Y(n289) );
  INVX2TS U264 ( .A(n236), .Y(n668) );
  CLKBUFX2TS U265 ( .A(n237), .Y(n241) );
  CLKBUFX2TS U266 ( .A(n327), .Y(n330) );
  CLKBUFX2TS U267 ( .A(n290), .Y(n294) );
  BUFX3TS U268 ( .A(outputPortSelect_NORTH[3]), .Y(n255) );
  CLKBUFX2TS U269 ( .A(n201), .Y(n286) );
  CLKBUFX2TS U270 ( .A(n224), .Y(n230) );
  CLKBUFX2TS U271 ( .A(n190), .Y(n315) );
  CLKBUFX2TS U272 ( .A(n212), .Y(n260) );
  INVX2TS U273 ( .A(n158), .Y(n194) );
  AO22XLTS U274 ( .A0(n345), .A1(n344), .B0(n327), .B1(
        outputPortSelect_WEST[2]), .Y(n75) );
  AO22XLTS U275 ( .A0(readInBuffer_SOUTH), .A1(n285), .B0(n284), .B1(
        memRead_SOUTH), .Y(n85) );
  AO22XLTS U276 ( .A0(writeInBuffer_SOUTH), .A1(n285), .B0(n284), .B1(
        memWrite_SOUTH), .Y(n90) );
  AO22XLTS U277 ( .A0(readInBuffer_NORTH), .A1(n258), .B0(n237), .B1(
        memRead_NORTH), .Y(n91) );
  AO22XLTS U278 ( .A0(writeInBuffer_NORTH), .A1(n258), .B0(n241), .B1(
        memWrite_NORTH), .Y(n96) );
  AO22XLTS U279 ( .A0(n384), .A1(n313), .B0(n294), .B1(memWrite_EAST), .Y(n84)
         );
  AO22XLTS U280 ( .A0(n390), .A1(n313), .B0(n294), .B1(memRead_EAST), .Y(n79)
         );
  INVX2TS U281 ( .A(n231), .Y(n232) );
  INVX2TS U282 ( .A(n187), .Y(n188) );
  INVX2TS U283 ( .A(outputPortSelect_NORTH[2]), .Y(n253) );
  INVX2TS U284 ( .A(n253), .Y(n348) );
  INVX2TS U285 ( .A(outputPortSelect_NORTH[1]), .Y(n245) );
  INVX2TS U286 ( .A(n245), .Y(n349) );
  INVX2TS U287 ( .A(outputPortSelect_NORTH[0]), .Y(n240) );
  INVX2TS U288 ( .A(n240), .Y(n350) );
  INVX2TS U289 ( .A(destinationAddressInBuffer_EAST[4]), .Y(n152) );
  INVX2TS U290 ( .A(n152), .Y(n351) );
  INVX2TS U291 ( .A(n152), .Y(n352) );
  INVX2TS U292 ( .A(destinationAddressInBuffer_EAST[5]), .Y(n153) );
  INVX2TS U293 ( .A(n153), .Y(n353) );
  INVX2TS U294 ( .A(n153), .Y(n354) );
  INVX2TS U295 ( .A(destinationAddressInBuffer_EAST[6]), .Y(n154) );
  INVX2TS U296 ( .A(n154), .Y(n355) );
  INVX2TS U297 ( .A(n154), .Y(n356) );
  INVX2TS U298 ( .A(destinationAddressInBuffer_EAST[7]), .Y(n155) );
  INVX2TS U299 ( .A(n155), .Y(n357) );
  INVX2TS U300 ( .A(n155), .Y(n358) );
  INVX2TS U301 ( .A(outputPortSelect_SOUTH[2]), .Y(n278) );
  INVX2TS U302 ( .A(n278), .Y(n359) );
  INVX2TS U303 ( .A(outputPortSelect_SOUTH[1]), .Y(n270) );
  INVX2TS U304 ( .A(n270), .Y(n360) );
  INVX2TS U305 ( .A(outputPortSelect_SOUTH[3]), .Y(n281) );
  INVX2TS U306 ( .A(n281), .Y(n361) );
  INVX2TS U307 ( .A(outputPortSelect_SOUTH[0]), .Y(n265) );
  INVX2TS U308 ( .A(n265), .Y(n362) );
  INVX2TS U309 ( .A(destinationAddressInBuffer_EAST[8]), .Y(n148) );
  INVX2TS U310 ( .A(n148), .Y(n363) );
  INVX2TS U311 ( .A(n148), .Y(n364) );
  INVX2TS U312 ( .A(n148), .Y(n365) );
  INVX2TS U313 ( .A(destinationAddressInBuffer_EAST[9]), .Y(n149) );
  INVX2TS U314 ( .A(n149), .Y(n366) );
  INVX2TS U315 ( .A(n149), .Y(n367) );
  INVX2TS U316 ( .A(n149), .Y(n368) );
  INVX2TS U317 ( .A(destinationAddressInBuffer_EAST[10]), .Y(n150) );
  INVX2TS U318 ( .A(n150), .Y(n369) );
  INVX2TS U319 ( .A(n150), .Y(n370) );
  INVX2TS U320 ( .A(n150), .Y(n371) );
  INVX2TS U321 ( .A(destinationAddressInBuffer_EAST[11]), .Y(n151) );
  INVX2TS U322 ( .A(n151), .Y(n372) );
  INVX2TS U323 ( .A(n151), .Y(n373) );
  INVX2TS U324 ( .A(n151), .Y(n374) );
  INVX2TS U325 ( .A(n152), .Y(n375) );
  INVX2TS U326 ( .A(n152), .Y(n376) );
  INVX2TS U327 ( .A(n153), .Y(n377) );
  INVX2TS U328 ( .A(n153), .Y(n378) );
  INVX2TS U329 ( .A(n154), .Y(n379) );
  INVX2TS U330 ( .A(n154), .Y(n380) );
  INVX2TS U331 ( .A(n155), .Y(n381) );
  INVX2TS U332 ( .A(n155), .Y(n382) );
  INVX2TS U333 ( .A(writeInBuffer_EAST), .Y(n156) );
  INVX2TS U334 ( .A(n156), .Y(n383) );
  INVX2TS U335 ( .A(n156), .Y(n384) );
  INVX2TS U336 ( .A(n156), .Y(n385) );
  INVX2TS U337 ( .A(n156), .Y(n386) );
  CLKBUFX2TS U338 ( .A(outputPortSelect_EAST[0]), .Y(n387) );
  INVX2TS U339 ( .A(outputPortSelect_EAST[1]), .Y(n299) );
  INVX2TS U340 ( .A(n299), .Y(n388) );
  INVX2TS U341 ( .A(readInBuffer_EAST), .Y(n157) );
  INVX2TS U342 ( .A(n157), .Y(n389) );
  INVX2TS U343 ( .A(n157), .Y(n390) );
  INVX2TS U344 ( .A(n157), .Y(n391) );
  CLKBUFX2TS U345 ( .A(reset), .Y(n158) );
  CLKBUFX2TS U346 ( .A(n194), .Y(n220) );
  CLKBUFX2TS U347 ( .A(n220), .Y(n236) );
  INVX2TS U348 ( .A(n236), .Y(n670) );
  CLKBUFX2TS U349 ( .A(writeInBuffer_SOUTH), .Y(n662) );
  CLKBUFX2TS U350 ( .A(destinationAddressInBuffer_SOUTH[7]), .Y(n624) );
  CLKBUFX2TS U351 ( .A(destinationAddressInBuffer_SOUTH[4]), .Y(n618) );
  CLKBUFX2TS U352 ( .A(destinationAddressInBuffer_SOUTH[6]), .Y(n622) );
  CLKBUFX2TS U353 ( .A(destinationAddressInBuffer_SOUTH[5]), .Y(n620) );
  CLKBUFX2TS U354 ( .A(readInBuffer_SOUTH), .Y(n435) );
  CLKBUFX2TS U355 ( .A(requesterAddressInBuffer_WEST[1]), .Y(n170) );
  CLKBUFX2TS U356 ( .A(n170), .Y(n469) );
  CLKBUFX2TS U357 ( .A(destinationAddressInBuffer_SOUTH[3]), .Y(n179) );
  CLKBUFX2TS U358 ( .A(n179), .Y(n615) );
  CLKBUFX2TS U359 ( .A(destinationAddressInBuffer_EAST[3]), .Y(n165) );
  CLKBUFX2TS U360 ( .A(n165), .Y(n565) );
  CLKBUFX2TS U361 ( .A(n170), .Y(n470) );
  CLKBUFX2TS U362 ( .A(n179), .Y(n616) );
  CLKBUFX2TS U363 ( .A(n165), .Y(n566) );
  CLKBUFX2TS U364 ( .A(destinationAddressInBuffer_SOUTH[2]), .Y(n180) );
  CLKBUFX2TS U365 ( .A(n180), .Y(n610) );
  CLKBUFX2TS U366 ( .A(destinationAddressInBuffer_EAST[2]), .Y(n166) );
  CLKBUFX2TS U367 ( .A(n166), .Y(n560) );
  CLKBUFX2TS U368 ( .A(destinationAddressInBuffer_SOUTH[1]), .Y(n178) );
  CLKBUFX2TS U369 ( .A(n178), .Y(n605) );
  CLKBUFX2TS U370 ( .A(destinationAddressInBuffer_EAST[1]), .Y(n164) );
  CLKBUFX2TS U371 ( .A(n164), .Y(n555) );
  CLKBUFX2TS U372 ( .A(requesterAddressInBuffer_WEST[0]), .Y(n169) );
  CLKBUFX2TS U373 ( .A(n169), .Y(n464) );
  CLKBUFX2TS U374 ( .A(destinationAddressInBuffer_SOUTH[0]), .Y(n173) );
  CLKBUFX2TS U375 ( .A(n173), .Y(n600) );
  CLKBUFX2TS U376 ( .A(destinationAddressInBuffer_EAST[0]), .Y(n159) );
  CLKBUFX2TS U377 ( .A(n159), .Y(n550) );
  CLKBUFX2TS U378 ( .A(n178), .Y(n606) );
  CLKBUFX2TS U379 ( .A(n164), .Y(n556) );
  CLKBUFX2TS U380 ( .A(n180), .Y(n611) );
  CLKBUFX2TS U381 ( .A(n166), .Y(n561) );
  CLKBUFX2TS U382 ( .A(n173), .Y(n601) );
  CLKBUFX2TS U383 ( .A(n159), .Y(n551) );
  CLKBUFX2TS U384 ( .A(n169), .Y(n465) );
  CLKBUFX2TS U385 ( .A(n170), .Y(n467) );
  CLKBUFX2TS U386 ( .A(n179), .Y(n613) );
  CLKBUFX2TS U387 ( .A(n165), .Y(n563) );
  CLKBUFX2TS U388 ( .A(requesterAddressInBuffer_WEST[3]), .Y(n171) );
  CLKBUFX2TS U389 ( .A(n171), .Y(n479) );
  CLKBUFX2TS U390 ( .A(requesterAddressInBuffer_WEST[2]), .Y(n172) );
  CLKBUFX2TS U391 ( .A(n172), .Y(n474) );
  CLKBUFX2TS U392 ( .A(n172), .Y(n475) );
  CLKBUFX2TS U393 ( .A(n171), .Y(n480) );
  CLKBUFX2TS U394 ( .A(n180), .Y(n608) );
  CLKBUFX2TS U395 ( .A(n166), .Y(n558) );
  CLKBUFX2TS U396 ( .A(n178), .Y(n603) );
  CLKBUFX2TS U397 ( .A(n164), .Y(n553) );
  CLKBUFX2TS U398 ( .A(n169), .Y(n462) );
  CLKBUFX2TS U399 ( .A(n173), .Y(n598) );
  CLKBUFX2TS U400 ( .A(n159), .Y(n548) );
  CLKBUFX2TS U401 ( .A(dataInBuffer_SOUTH[0]), .Y(n182) );
  CLKBUFX2TS U402 ( .A(n182), .Y(n570) );
  CLKBUFX2TS U403 ( .A(dataInBuffer_EAST[0]), .Y(n168) );
  CLKBUFX2TS U404 ( .A(n168), .Y(n516) );
  CLKBUFX2TS U405 ( .A(dataInBuffer_SOUTH[5]), .Y(n175) );
  CLKBUFX2TS U406 ( .A(n175), .Y(n595) );
  CLKBUFX2TS U407 ( .A(dataInBuffer_EAST[5]), .Y(n161) );
  CLKBUFX2TS U408 ( .A(n161), .Y(n541) );
  CLKBUFX2TS U409 ( .A(n182), .Y(n571) );
  CLKBUFX2TS U410 ( .A(n168), .Y(n517) );
  CLKBUFX2TS U411 ( .A(dataInBuffer_SOUTH[1]), .Y(n181) );
  CLKBUFX2TS U412 ( .A(n181), .Y(n576) );
  CLKBUFX2TS U413 ( .A(dataInBuffer_EAST[1]), .Y(n167) );
  CLKBUFX2TS U414 ( .A(n167), .Y(n522) );
  CLKBUFX2TS U415 ( .A(dataInBuffer_SOUTH[3]), .Y(n176) );
  CLKBUFX2TS U416 ( .A(n176), .Y(n586) );
  CLKBUFX2TS U417 ( .A(dataInBuffer_EAST[3]), .Y(n162) );
  CLKBUFX2TS U418 ( .A(n162), .Y(n532) );
  CLKBUFX2TS U419 ( .A(dataInBuffer_SOUTH[4]), .Y(n177) );
  CLKBUFX2TS U420 ( .A(n177), .Y(n590) );
  CLKBUFX2TS U421 ( .A(dataInBuffer_EAST[4]), .Y(n163) );
  CLKBUFX2TS U422 ( .A(n163), .Y(n536) );
  CLKBUFX2TS U423 ( .A(n181), .Y(n575) );
  CLKBUFX2TS U424 ( .A(n167), .Y(n521) );
  CLKBUFX2TS U425 ( .A(dataInBuffer_SOUTH[2]), .Y(n174) );
  CLKBUFX2TS U426 ( .A(n174), .Y(n580) );
  CLKBUFX2TS U427 ( .A(dataInBuffer_EAST[2]), .Y(n160) );
  CLKBUFX2TS U428 ( .A(n160), .Y(n526) );
  CLKBUFX2TS U429 ( .A(n175), .Y(n596) );
  CLKBUFX2TS U430 ( .A(n161), .Y(n542) );
  CLKBUFX2TS U431 ( .A(n177), .Y(n591) );
  CLKBUFX2TS U432 ( .A(n163), .Y(n537) );
  CLKBUFX2TS U433 ( .A(n174), .Y(n581) );
  CLKBUFX2TS U434 ( .A(n160), .Y(n527) );
  CLKBUFX2TS U435 ( .A(n176), .Y(n585) );
  CLKBUFX2TS U436 ( .A(n162), .Y(n531) );
  CLKBUFX2TS U437 ( .A(n171), .Y(n477) );
  CLKBUFX2TS U438 ( .A(n172), .Y(n472) );
  CLKBUFX2TS U439 ( .A(n175), .Y(n593) );
  CLKBUFX2TS U440 ( .A(n161), .Y(n539) );
  CLKBUFX2TS U441 ( .A(n174), .Y(n578) );
  CLKBUFX2TS U442 ( .A(n160), .Y(n524) );
  CLKBUFX2TS U443 ( .A(n181), .Y(n573) );
  CLKBUFX2TS U444 ( .A(n167), .Y(n519) );
  CLKBUFX2TS U445 ( .A(n182), .Y(n568) );
  CLKBUFX2TS U446 ( .A(n168), .Y(n514) );
  CLKBUFX2TS U447 ( .A(n177), .Y(n588) );
  CLKBUFX2TS U448 ( .A(n163), .Y(n534) );
  CLKBUFX2TS U449 ( .A(n176), .Y(n583) );
  CLKBUFX2TS U450 ( .A(n162), .Y(n529) );
  CLKBUFX2TS U451 ( .A(readInBuffer_NORTH), .Y(n434) );
  CLKBUFX2TS U452 ( .A(writeInBuffer_NORTH), .Y(n433) );
  CLKBUFX2TS U453 ( .A(readInBuffer_WEST), .Y(n437) );
  CLKBUFX2TS U454 ( .A(writeInBuffer_WEST), .Y(n436) );
  CLKBUFX2TS U455 ( .A(n220), .Y(n223) );
  INVX2TS U456 ( .A(n223), .Y(n667) );
  INVX2TS U457 ( .A(n223), .Y(n669) );
  CLKBUFX2TS U458 ( .A(readInBuffer_WEST), .Y(n660) );
  CLKBUFX2TS U459 ( .A(writeInBuffer_NORTH), .Y(n663) );
  CLKBUFX2TS U460 ( .A(writeInBuffer_WEST), .Y(n658) );
  CLKBUFX2TS U461 ( .A(destinationAddressInBuffer_WEST[5]), .Y(n505) );
  CLKBUFX2TS U462 ( .A(destinationAddressInBuffer_WEST[7]), .Y(n513) );
  CLKBUFX2TS U463 ( .A(destinationAddressInBuffer_WEST[4]), .Y(n501) );
  CLKBUFX2TS U464 ( .A(destinationAddressInBuffer_WEST[6]), .Y(n509) );
  CLKBUFX2TS U465 ( .A(destinationAddressInBuffer_NORTH[4]), .Y(n428) );
  CLKBUFX2TS U466 ( .A(destinationAddressInBuffer_WEST[4]), .Y(n500) );
  CLKBUFX2TS U467 ( .A(destinationAddressInBuffer_NORTH[5]), .Y(n429) );
  CLKBUFX2TS U468 ( .A(destinationAddressInBuffer_WEST[5]), .Y(n504) );
  CLKBUFX2TS U469 ( .A(destinationAddressInBuffer_NORTH[6]), .Y(n430) );
  CLKBUFX2TS U470 ( .A(destinationAddressInBuffer_WEST[6]), .Y(n508) );
  CLKBUFX2TS U471 ( .A(destinationAddressInBuffer_NORTH[7]), .Y(n431) );
  CLKBUFX2TS U472 ( .A(destinationAddressInBuffer_WEST[7]), .Y(n512) );
  CLKBUFX2TS U473 ( .A(destinationAddressInBuffer_NORTH[7]), .Y(n654) );
  CLKBUFX2TS U474 ( .A(destinationAddressInBuffer_WEST[7]), .Y(n510) );
  CLKBUFX2TS U475 ( .A(destinationAddressInBuffer_NORTH[7]), .Y(n655) );
  CLKBUFX2TS U476 ( .A(destinationAddressInBuffer_WEST[7]), .Y(n511) );
  CLKBUFX2TS U477 ( .A(destinationAddressInBuffer_NORTH[4]), .Y(n642) );
  CLKBUFX2TS U478 ( .A(destinationAddressInBuffer_WEST[4]), .Y(n498) );
  CLKBUFX2TS U479 ( .A(destinationAddressInBuffer_NORTH[6]), .Y(n650) );
  CLKBUFX2TS U480 ( .A(destinationAddressInBuffer_WEST[6]), .Y(n506) );
  CLKBUFX2TS U481 ( .A(destinationAddressInBuffer_NORTH[4]), .Y(n643) );
  CLKBUFX2TS U482 ( .A(destinationAddressInBuffer_WEST[4]), .Y(n499) );
  CLKBUFX2TS U483 ( .A(destinationAddressInBuffer_NORTH[6]), .Y(n651) );
  CLKBUFX2TS U484 ( .A(destinationAddressInBuffer_WEST[6]), .Y(n507) );
  CLKBUFX2TS U485 ( .A(destinationAddressInBuffer_NORTH[5]), .Y(n647) );
  CLKBUFX2TS U486 ( .A(destinationAddressInBuffer_WEST[5]), .Y(n503) );
  CLKBUFX2TS U487 ( .A(destinationAddressInBuffer_NORTH[5]), .Y(n646) );
  CLKBUFX2TS U488 ( .A(destinationAddressInBuffer_WEST[5]), .Y(n502) );
  CLKBUFX2TS U489 ( .A(requesterAddressInBuffer_NORTH[1]), .Y(n632) );
  CLKBUFX2TS U490 ( .A(destinationAddressInBuffer_WEST[3]), .Y(n496) );
  CLKBUFX2TS U491 ( .A(requesterAddressInBuffer_NORTH[1]), .Y(n633) );
  CLKBUFX2TS U492 ( .A(requesterAddressInBuffer_EAST[1]), .Y(n395) );
  CLKBUFX2TS U493 ( .A(destinationAddressInBuffer_WEST[3]), .Y(n497) );
  CLKBUFX2TS U494 ( .A(destinationAddressInBuffer_WEST[2]), .Y(n492) );
  CLKBUFX2TS U495 ( .A(destinationAddressInBuffer_WEST[1]), .Y(n488) );
  CLKBUFX2TS U496 ( .A(requesterAddressInBuffer_NORTH[0]), .Y(n628) );
  CLKBUFX2TS U497 ( .A(destinationAddressInBuffer_WEST[0]), .Y(n484) );
  CLKBUFX2TS U498 ( .A(destinationAddressInBuffer_WEST[1]), .Y(n489) );
  CLKBUFX2TS U499 ( .A(destinationAddressInBuffer_WEST[2]), .Y(n493) );
  CLKBUFX2TS U500 ( .A(destinationAddressInBuffer_WEST[0]), .Y(n485) );
  CLKBUFX2TS U501 ( .A(requesterAddressInBuffer_NORTH[0]), .Y(n629) );
  CLKBUFX2TS U502 ( .A(requesterAddressInBuffer_EAST[0]), .Y(n393) );
  CLKBUFX2TS U503 ( .A(requesterAddressInBuffer_NORTH[1]), .Y(n630) );
  CLKBUFX2TS U504 ( .A(requesterAddressInBuffer_EAST[1]), .Y(n394) );
  CLKBUFX2TS U505 ( .A(destinationAddressInBuffer_WEST[3]), .Y(n494) );
  CLKBUFX2TS U506 ( .A(requesterAddressInBuffer_NORTH[1]), .Y(n631) );
  CLKBUFX2TS U507 ( .A(requesterAddressInBuffer_SOUTH[1]), .Y(n402) );
  CLKBUFX2TS U508 ( .A(requesterAddressInBuffer_WEST[1]), .Y(n468) );
  CLKBUFX2TS U509 ( .A(destinationAddressInBuffer_SOUTH[3]), .Y(n614) );
  CLKBUFX2TS U510 ( .A(destinationAddressInBuffer_NORTH[3]), .Y(n426) );
  CLKBUFX2TS U511 ( .A(destinationAddressInBuffer_EAST[3]), .Y(n564) );
  CLKBUFX2TS U512 ( .A(destinationAddressInBuffer_WEST[3]), .Y(n495) );
  CLKBUFX2TS U513 ( .A(requesterAddressInBuffer_NORTH[3]), .Y(n640) );
  CLKBUFX2TS U514 ( .A(requesterAddressInBuffer_NORTH[2]), .Y(n636) );
  CLKBUFX2TS U515 ( .A(requesterAddressInBuffer_NORTH[2]), .Y(n637) );
  CLKBUFX2TS U516 ( .A(requesterAddressInBuffer_EAST[2]), .Y(n397) );
  CLKBUFX2TS U517 ( .A(requesterAddressInBuffer_NORTH[3]), .Y(n641) );
  CLKBUFX2TS U518 ( .A(requesterAddressInBuffer_EAST[3]), .Y(n399) );
  CLKBUFX2TS U519 ( .A(destinationAddressInBuffer_WEST[2]), .Y(n490) );
  CLKBUFX2TS U520 ( .A(destinationAddressInBuffer_WEST[1]), .Y(n486) );
  CLKBUFX2TS U521 ( .A(destinationAddressInBuffer_SOUTH[1]), .Y(n604) );
  CLKBUFX2TS U522 ( .A(destinationAddressInBuffer_NORTH[1]), .Y(n422) );
  CLKBUFX2TS U523 ( .A(destinationAddressInBuffer_EAST[1]), .Y(n554) );
  CLKBUFX2TS U524 ( .A(destinationAddressInBuffer_WEST[1]), .Y(n487) );
  CLKBUFX2TS U525 ( .A(destinationAddressInBuffer_SOUTH[2]), .Y(n609) );
  CLKBUFX2TS U526 ( .A(destinationAddressInBuffer_NORTH[2]), .Y(n424) );
  CLKBUFX2TS U527 ( .A(destinationAddressInBuffer_EAST[2]), .Y(n559) );
  CLKBUFX2TS U528 ( .A(destinationAddressInBuffer_WEST[2]), .Y(n491) );
  CLKBUFX2TS U529 ( .A(requesterAddressInBuffer_NORTH[0]), .Y(n626) );
  CLKBUFX2TS U530 ( .A(requesterAddressInBuffer_EAST[0]), .Y(n392) );
  CLKBUFX2TS U531 ( .A(destinationAddressInBuffer_SOUTH[0]), .Y(n599) );
  CLKBUFX2TS U532 ( .A(destinationAddressInBuffer_EAST[0]), .Y(n549) );
  CLKBUFX2TS U533 ( .A(destinationAddressInBuffer_WEST[0]), .Y(n483) );
  CLKBUFX2TS U534 ( .A(destinationAddressInBuffer_NORTH[0]), .Y(n420) );
  CLKBUFX2TS U535 ( .A(destinationAddressInBuffer_WEST[0]), .Y(n482) );
  CLKBUFX2TS U536 ( .A(requesterAddressInBuffer_NORTH[0]), .Y(n627) );
  CLKBUFX2TS U537 ( .A(requesterAddressInBuffer_SOUTH[0]), .Y(n400) );
  CLKBUFX2TS U538 ( .A(requesterAddressInBuffer_WEST[0]), .Y(n463) );
  CLKBUFX2TS U539 ( .A(dataInBuffer_WEST[0]), .Y(n440) );
  CLKBUFX2TS U540 ( .A(dataInBuffer_WEST[5]), .Y(n460) );
  CLKBUFX2TS U541 ( .A(dataInBuffer_WEST[0]), .Y(n441) );
  CLKBUFX2TS U542 ( .A(dataInBuffer_WEST[1]), .Y(n445) );
  CLKBUFX2TS U543 ( .A(dataInBuffer_WEST[3]), .Y(n453) );
  CLKBUFX2TS U544 ( .A(dataInBuffer_WEST[4]), .Y(n456) );
  CLKBUFX2TS U545 ( .A(dataInBuffer_WEST[1]), .Y(n444) );
  CLKBUFX2TS U546 ( .A(dataInBuffer_WEST[2]), .Y(n448) );
  CLKBUFX2TS U547 ( .A(dataInBuffer_WEST[5]), .Y(n461) );
  CLKBUFX2TS U548 ( .A(dataInBuffer_WEST[4]), .Y(n457) );
  CLKBUFX2TS U549 ( .A(dataInBuffer_WEST[2]), .Y(n449) );
  CLKBUFX2TS U550 ( .A(dataInBuffer_WEST[3]), .Y(n452) );
  CLKBUFX2TS U551 ( .A(requesterAddressInBuffer_NORTH[3]), .Y(n638) );
  CLKBUFX2TS U552 ( .A(requesterAddressInBuffer_EAST[3]), .Y(n398) );
  CLKBUFX2TS U553 ( .A(requesterAddressInBuffer_NORTH[3]), .Y(n639) );
  CLKBUFX2TS U554 ( .A(requesterAddressInBuffer_SOUTH[3]), .Y(n406) );
  CLKBUFX2TS U555 ( .A(requesterAddressInBuffer_WEST[3]), .Y(n478) );
  CLKBUFX2TS U556 ( .A(requesterAddressInBuffer_NORTH[2]), .Y(n634) );
  CLKBUFX2TS U557 ( .A(requesterAddressInBuffer_EAST[2]), .Y(n396) );
  CLKBUFX2TS U558 ( .A(requesterAddressInBuffer_NORTH[2]), .Y(n635) );
  CLKBUFX2TS U559 ( .A(requesterAddressInBuffer_SOUTH[2]), .Y(n404) );
  CLKBUFX2TS U560 ( .A(requesterAddressInBuffer_WEST[2]), .Y(n473) );
  CLKBUFX2TS U561 ( .A(dataInBuffer_SOUTH[4]), .Y(n589) );
  CLKBUFX2TS U562 ( .A(dataInBuffer_EAST[4]), .Y(n535) );
  CLKBUFX2TS U563 ( .A(dataInBuffer_WEST[4]), .Y(n455) );
  CLKBUFX2TS U564 ( .A(dataInBuffer_SOUTH[3]), .Y(n584) );
  CLKBUFX2TS U565 ( .A(dataInBuffer_EAST[3]), .Y(n530) );
  CLKBUFX2TS U566 ( .A(dataInBuffer_WEST[3]), .Y(n451) );
  CLKBUFX2TS U567 ( .A(dataInBuffer_SOUTH[2]), .Y(n579) );
  CLKBUFX2TS U568 ( .A(dataInBuffer_EAST[2]), .Y(n525) );
  CLKBUFX2TS U569 ( .A(dataInBuffer_WEST[2]), .Y(n447) );
  CLKBUFX2TS U570 ( .A(dataInBuffer_WEST[5]), .Y(n458) );
  CLKBUFX2TS U571 ( .A(dataInBuffer_NORTH[2]), .Y(n412) );
  CLKBUFX2TS U572 ( .A(dataInBuffer_WEST[2]), .Y(n446) );
  CLKBUFX2TS U573 ( .A(dataInBuffer_WEST[1]), .Y(n442) );
  CLKBUFX2TS U574 ( .A(dataInBuffer_NORTH[5]), .Y(n418) );
  CLKBUFX2TS U575 ( .A(dataInBuffer_SOUTH[5]), .Y(n594) );
  CLKBUFX2TS U576 ( .A(dataInBuffer_EAST[5]), .Y(n540) );
  CLKBUFX2TS U577 ( .A(dataInBuffer_WEST[5]), .Y(n459) );
  CLKBUFX2TS U578 ( .A(dataInBuffer_WEST[0]), .Y(n438) );
  CLKBUFX2TS U579 ( .A(dataInBuffer_NORTH[4]), .Y(n416) );
  CLKBUFX2TS U580 ( .A(dataInBuffer_WEST[4]), .Y(n454) );
  CLKBUFX2TS U581 ( .A(dataInBuffer_NORTH[3]), .Y(n414) );
  CLKBUFX2TS U582 ( .A(dataInBuffer_WEST[3]), .Y(n450) );
  CLKBUFX2TS U583 ( .A(dataInBuffer_NORTH[0]), .Y(n408) );
  CLKBUFX2TS U584 ( .A(dataInBuffer_SOUTH[0]), .Y(n569) );
  CLKBUFX2TS U585 ( .A(dataInBuffer_EAST[0]), .Y(n515) );
  CLKBUFX2TS U586 ( .A(dataInBuffer_WEST[0]), .Y(n439) );
  CLKBUFX2TS U587 ( .A(dataInBuffer_NORTH[1]), .Y(n410) );
  CLKBUFX2TS U588 ( .A(dataInBuffer_SOUTH[1]), .Y(n574) );
  CLKBUFX2TS U589 ( .A(dataInBuffer_EAST[1]), .Y(n520) );
  CLKBUFX2TS U590 ( .A(dataInBuffer_WEST[1]), .Y(n443) );
  CLKBUFX2TS U591 ( .A(n159), .Y(n552) );
  CLKBUFX2TS U592 ( .A(n160), .Y(n528) );
  CLKBUFX2TS U593 ( .A(n161), .Y(n543) );
  CLKBUFX2TS U594 ( .A(n162), .Y(n533) );
  CLKBUFX2TS U595 ( .A(n163), .Y(n538) );
  CLKBUFX2TS U596 ( .A(n164), .Y(n557) );
  CLKBUFX2TS U597 ( .A(n165), .Y(n567) );
  CLKBUFX2TS U598 ( .A(n166), .Y(n562) );
  CLKBUFX2TS U599 ( .A(n167), .Y(n523) );
  CLKBUFX2TS U600 ( .A(n168), .Y(n518) );
  CLKBUFX2TS U601 ( .A(n169), .Y(n466) );
  CLKBUFX2TS U602 ( .A(n393), .Y(n544) );
  CLKBUFX2TS U603 ( .A(n395), .Y(n545) );
  CLKBUFX2TS U604 ( .A(n170), .Y(n471) );
  CLKBUFX2TS U605 ( .A(n399), .Y(n547) );
  CLKBUFX2TS U606 ( .A(n171), .Y(n481) );
  CLKBUFX2TS U607 ( .A(n397), .Y(n546) );
  CLKBUFX2TS U608 ( .A(n172), .Y(n476) );
  CLKBUFX2TS U609 ( .A(readInBuffer_NORTH), .Y(n665) );
  CLKBUFX2TS U610 ( .A(n434), .Y(n666) );
  CLKBUFX2TS U611 ( .A(n437), .Y(n661) );
  CLKBUFX2TS U612 ( .A(n173), .Y(n602) );
  CLKBUFX2TS U613 ( .A(destinationAddressInBuffer_SOUTH[7]), .Y(n625) );
  CLKBUFX2TS U614 ( .A(destinationAddressInBuffer_SOUTH[4]), .Y(n619) );
  CLKBUFX2TS U615 ( .A(destinationAddressInBuffer_SOUTH[6]), .Y(n623) );
  CLKBUFX2TS U616 ( .A(destinationAddressInBuffer_SOUTH[5]), .Y(n621) );
  CLKBUFX2TS U617 ( .A(n174), .Y(n582) );
  CLKBUFX2TS U618 ( .A(n175), .Y(n597) );
  CLKBUFX2TS U619 ( .A(n176), .Y(n587) );
  CLKBUFX2TS U620 ( .A(n177), .Y(n592) );
  CLKBUFX2TS U621 ( .A(n178), .Y(n607) );
  CLKBUFX2TS U622 ( .A(n179), .Y(n617) );
  CLKBUFX2TS U623 ( .A(n180), .Y(n612) );
  CLKBUFX2TS U624 ( .A(n181), .Y(n577) );
  CLKBUFX2TS U625 ( .A(n182), .Y(n572) );
  CLKBUFX2TS U626 ( .A(n433), .Y(n664) );
  CLKBUFX2TS U627 ( .A(n436), .Y(n659) );
  CLKBUFX2TS U628 ( .A(n429), .Y(n649) );
  CLKBUFX2TS U629 ( .A(n431), .Y(n657) );
  CLKBUFX2TS U630 ( .A(n428), .Y(n645) );
  CLKBUFX2TS U631 ( .A(n430), .Y(n653) );
  CLKBUFX2TS U632 ( .A(n428), .Y(n644) );
  CLKBUFX2TS U633 ( .A(n429), .Y(n648) );
  CLKBUFX2TS U634 ( .A(n430), .Y(n652) );
  CLKBUFX2TS U635 ( .A(n431), .Y(n656) );
  CLKBUFX2TS U636 ( .A(readInBuffer_SOUTH), .Y(n432) );
  CLKBUFX2TS U637 ( .A(requesterAddressInBuffer_SOUTH[0]), .Y(n401) );
  CLKBUFX2TS U638 ( .A(requesterAddressInBuffer_SOUTH[1]), .Y(n403) );
  CLKBUFX2TS U639 ( .A(requesterAddressInBuffer_SOUTH[2]), .Y(n405) );
  CLKBUFX2TS U640 ( .A(requesterAddressInBuffer_SOUTH[3]), .Y(n407) );
  CLKBUFX2TS U641 ( .A(destinationAddressInBuffer_NORTH[0]), .Y(n421) );
  CLKBUFX2TS U642 ( .A(dataInBuffer_NORTH[0]), .Y(n409) );
  CLKBUFX2TS U643 ( .A(dataInBuffer_NORTH[1]), .Y(n411) );
  CLKBUFX2TS U644 ( .A(dataInBuffer_NORTH[2]), .Y(n413) );
  CLKBUFX2TS U645 ( .A(dataInBuffer_NORTH[3]), .Y(n415) );
  CLKBUFX2TS U646 ( .A(dataInBuffer_NORTH[4]), .Y(n417) );
  CLKBUFX2TS U647 ( .A(dataInBuffer_NORTH[5]), .Y(n419) );
  CLKBUFX2TS U648 ( .A(destinationAddressInBuffer_NORTH[3]), .Y(n427) );
  CLKBUFX2TS U649 ( .A(destinationAddressInBuffer_NORTH[2]), .Y(n425) );
  CLKBUFX2TS U650 ( .A(destinationAddressInBuffer_NORTH[1]), .Y(n423) );
  NOR2BX1TS U651 ( .AN(dataIn_WEST[0]), .B(n289), .Y(N94) );
  CLKBUFX2TS U652 ( .A(n194), .Y(n206) );
  CLKBUFX2TS U653 ( .A(n206), .Y(n238) );
  INVX2TS U654 ( .A(n238), .Y(n183) );
  NOR2BX1TS U655 ( .AN(dataIn_WEST[1]), .B(n183), .Y(N95) );
  NOR2BX1TS U656 ( .AN(dataIn_WEST[2]), .B(n183), .Y(N96) );
  NOR2BX1TS U657 ( .AN(dataIn_WEST[3]), .B(n183), .Y(N97) );
  NOR2BX1TS U658 ( .AN(dataIn_WEST[4]), .B(n183), .Y(N98) );
  INVX2TS U659 ( .A(n238), .Y(n184) );
  NOR2BX1TS U660 ( .AN(dataIn_WEST[5]), .B(n184), .Y(N99) );
  NOR2BX1TS U661 ( .AN(writeIn_WEST), .B(n184), .Y(N93) );
  NOR2BX1TS U662 ( .AN(readIn_WEST), .B(n184), .Y(N92) );
  NOR2BX1TS U663 ( .AN(requesterAddressIn_WEST[0]), .B(n184), .Y(N88) );
  INVX2TS U664 ( .A(n238), .Y(n185) );
  NOR2BX1TS U665 ( .AN(requesterAddressIn_WEST[1]), .B(n185), .Y(N89) );
  NOR2BX1TS U666 ( .AN(requesterAddressIn_WEST[2]), .B(n185), .Y(N90) );
  NOR2BX1TS U667 ( .AN(requesterAddressIn_WEST[3]), .B(n185), .Y(N91) );
  NOR2BX1TS U668 ( .AN(destinationAddressIn_WEST[0]), .B(n185), .Y(N76) );
  CLKBUFX2TS U669 ( .A(n194), .Y(n218) );
  CLKBUFX2TS U670 ( .A(n218), .Y(n263) );
  INVX2TS U671 ( .A(n263), .Y(n186) );
  NOR2BX1TS U672 ( .AN(destinationAddressIn_WEST[1]), .B(n186), .Y(N77) );
  NOR2BX1TS U673 ( .AN(destinationAddressIn_WEST[2]), .B(n186), .Y(N78) );
  NOR2BX1TS U674 ( .AN(destinationAddressIn_WEST[3]), .B(n186), .Y(N79) );
  NOR2BX1TS U675 ( .AN(destinationAddressIn_WEST[4]), .B(n186), .Y(N80) );
  INVX2TS U676 ( .A(n263), .Y(n189) );
  NOR2BX1TS U677 ( .AN(destinationAddressIn_WEST[5]), .B(n189), .Y(N81) );
  NOR2BX1TS U678 ( .AN(destinationAddressIn_WEST[6]), .B(n189), .Y(N82) );
  NOR2BX1TS U679 ( .AN(destinationAddressIn_WEST[7]), .B(n189), .Y(N83) );
  CLKBUFX2TS U680 ( .A(destinationAddressIn_WEST[8]), .Y(n187) );
  NOR2BX1TS U681 ( .AN(n187), .B(n189), .Y(N84) );
  CLKBUFX2TS U682 ( .A(destinationAddressIn_WEST[9]), .Y(n190) );
  INVX2TS U683 ( .A(n263), .Y(n193) );
  NOR2BX1TS U684 ( .AN(n190), .B(n193), .Y(N85) );
  CLKBUFX2TS U685 ( .A(destinationAddressIn_WEST[10]), .Y(n191) );
  NOR2BX1TS U686 ( .AN(n191), .B(n193), .Y(N86) );
  CLKBUFX2TS U687 ( .A(destinationAddressIn_WEST[11]), .Y(n192) );
  NOR2BX1TS U688 ( .AN(n192), .B(n193), .Y(N87) );
  NOR2BX1TS U689 ( .AN(dataIn_EAST[0]), .B(n193), .Y(N70) );
  CLKBUFX2TS U690 ( .A(n194), .Y(n211) );
  CLKBUFX2TS U691 ( .A(n211), .Y(n292) );
  INVX2TS U692 ( .A(n292), .Y(n195) );
  NOR2BX1TS U693 ( .AN(dataIn_EAST[1]), .B(n195), .Y(N71) );
  NOR2BX1TS U694 ( .AN(dataIn_EAST[2]), .B(n195), .Y(N72) );
  NOR2BX1TS U695 ( .AN(dataIn_EAST[3]), .B(n195), .Y(N73) );
  NOR2BX1TS U696 ( .AN(dataIn_EAST[4]), .B(n195), .Y(N74) );
  INVX2TS U697 ( .A(n292), .Y(n196) );
  NOR2BX1TS U698 ( .AN(dataIn_EAST[5]), .B(n196), .Y(N75) );
  NOR2BX1TS U699 ( .AN(writeIn_EAST), .B(n196), .Y(N69) );
  NOR2BX1TS U700 ( .AN(readIn_EAST), .B(n196), .Y(N68) );
  NOR2BX1TS U701 ( .AN(requesterAddressIn_EAST[0]), .B(n196), .Y(N64) );
  INVX2TS U702 ( .A(n292), .Y(n197) );
  NOR2BX1TS U703 ( .AN(requesterAddressIn_EAST[1]), .B(n197), .Y(N65) );
  NOR2BX1TS U704 ( .AN(requesterAddressIn_EAST[2]), .B(n197), .Y(N66) );
  NOR2BX1TS U705 ( .AN(requesterAddressIn_EAST[3]), .B(n197), .Y(N67) );
  NOR2BX1TS U706 ( .AN(destinationAddressIn_EAST[0]), .B(n197), .Y(N52) );
  CLKBUFX2TS U707 ( .A(n220), .Y(n329) );
  INVX2TS U708 ( .A(n329), .Y(n198) );
  NOR2BX1TS U709 ( .AN(destinationAddressIn_EAST[1]), .B(n198), .Y(N53) );
  NOR2BX1TS U710 ( .AN(destinationAddressIn_EAST[2]), .B(n198), .Y(N54) );
  NOR2BX1TS U711 ( .AN(destinationAddressIn_EAST[3]), .B(n198), .Y(N55) );
  NOR2BX1TS U712 ( .AN(destinationAddressIn_EAST[4]), .B(n198), .Y(N56) );
  INVX2TS U713 ( .A(n329), .Y(n200) );
  NOR2BX1TS U714 ( .AN(destinationAddressIn_EAST[5]), .B(n200), .Y(N57) );
  NOR2BX1TS U715 ( .AN(destinationAddressIn_EAST[6]), .B(n200), .Y(N58) );
  NOR2BX1TS U716 ( .AN(destinationAddressIn_EAST[7]), .B(n200), .Y(N59) );
  CLKBUFX2TS U717 ( .A(destinationAddressIn_EAST[8]), .Y(n199) );
  NOR2BX1TS U718 ( .AN(n199), .B(n200), .Y(N60) );
  CLKBUFX2TS U719 ( .A(destinationAddressIn_EAST[9]), .Y(n201) );
  INVX2TS U720 ( .A(n329), .Y(n204) );
  NOR2BX1TS U721 ( .AN(n201), .B(n204), .Y(N61) );
  CLKBUFX2TS U722 ( .A(destinationAddressIn_EAST[10]), .Y(n202) );
  NOR2BX1TS U723 ( .AN(n202), .B(n204), .Y(N62) );
  CLKBUFX2TS U724 ( .A(destinationAddressIn_EAST[11]), .Y(n203) );
  NOR2BX1TS U725 ( .AN(n203), .B(n204), .Y(N63) );
  NOR2BX1TS U726 ( .AN(dataIn_SOUTH[0]), .B(n204), .Y(N46) );
  INVX2TS U727 ( .A(n206), .Y(n217) );
  NOR2BX1TS U728 ( .AN(dataIn_SOUTH[1]), .B(n217), .Y(N47) );
  NOR2BX1TS U729 ( .AN(dataIn_SOUTH[2]), .B(n217), .Y(N48) );
  NOR2BX1TS U730 ( .AN(dataIn_SOUTH[3]), .B(n217), .Y(N49) );
  INVX2TS U731 ( .A(n206), .Y(n205) );
  NOR2BX1TS U732 ( .AN(dataIn_SOUTH[4]), .B(n205), .Y(N50) );
  NOR2BX1TS U733 ( .AN(dataIn_SOUTH[5]), .B(n205), .Y(N51) );
  NOR2BX1TS U734 ( .AN(writeIn_SOUTH), .B(n205), .Y(N45) );
  NOR2BX1TS U735 ( .AN(readIn_SOUTH), .B(n205), .Y(N44) );
  INVX2TS U736 ( .A(n206), .Y(n207) );
  NOR2BX1TS U737 ( .AN(requesterAddressIn_SOUTH[0]), .B(n207), .Y(N40) );
  NOR2BX1TS U738 ( .AN(requesterAddressIn_SOUTH[1]), .B(n207), .Y(N41) );
  NOR2BX1TS U739 ( .AN(requesterAddressIn_SOUTH[2]), .B(n207), .Y(N42) );
  NOR2BX1TS U740 ( .AN(requesterAddressIn_SOUTH[3]), .B(n207), .Y(N43) );
  INVX2TS U741 ( .A(n211), .Y(n208) );
  NOR2BX1TS U742 ( .AN(destinationAddressIn_SOUTH[0]), .B(n208), .Y(N28) );
  NOR2BX1TS U743 ( .AN(destinationAddressIn_SOUTH[1]), .B(n208), .Y(N29) );
  NOR2BX1TS U744 ( .AN(destinationAddressIn_SOUTH[2]), .B(n208), .Y(N30) );
  NOR2BX1TS U745 ( .AN(destinationAddressIn_SOUTH[3]), .B(n208), .Y(N31) );
  INVX2TS U746 ( .A(n211), .Y(n209) );
  NOR2BX1TS U747 ( .AN(destinationAddressIn_SOUTH[4]), .B(n209), .Y(N32) );
  NOR2BX1TS U748 ( .AN(destinationAddressIn_SOUTH[5]), .B(n209), .Y(N33) );
  NOR2BX1TS U749 ( .AN(destinationAddressIn_SOUTH[6]), .B(n209), .Y(N34) );
  NOR2BX1TS U750 ( .AN(destinationAddressIn_SOUTH[7]), .B(n209), .Y(N35) );
  CLKBUFX2TS U751 ( .A(destinationAddressIn_SOUTH[8]), .Y(n210) );
  INVX2TS U752 ( .A(n211), .Y(n215) );
  NOR2BX1TS U753 ( .AN(n210), .B(n215), .Y(N36) );
  CLKBUFX2TS U754 ( .A(destinationAddressIn_SOUTH[9]), .Y(n212) );
  NOR2BX1TS U755 ( .AN(n212), .B(n215), .Y(N37) );
  CLKBUFX2TS U756 ( .A(destinationAddressIn_SOUTH[10]), .Y(n213) );
  NOR2BX1TS U757 ( .AN(n213), .B(n215), .Y(N38) );
  CLKBUFX2TS U758 ( .A(destinationAddressIn_SOUTH[11]), .Y(n214) );
  NOR2BX1TS U759 ( .AN(n214), .B(n215), .Y(N39) );
  INVX2TS U760 ( .A(n218), .Y(n216) );
  NOR2BX1TS U761 ( .AN(dataIn_NORTH[0]), .B(n216), .Y(N22) );
  NOR2BX1TS U762 ( .AN(dataIn_NORTH[1]), .B(n216), .Y(N23) );
  NOR2BX1TS U763 ( .AN(dataIn_NORTH[2]), .B(n216), .Y(N24) );
  NOR2BX1TS U764 ( .AN(dataIn_NORTH[3]), .B(n216), .Y(N25) );
  INVX2TS U765 ( .A(n218), .Y(n325) );
  NOR2BX1TS U766 ( .AN(dataIn_NORTH[4]), .B(n325), .Y(N26) );
  NOR2BX1TS U767 ( .AN(dataIn_NORTH[5]), .B(n217), .Y(N27) );
  NOR2BX1TS U768 ( .AN(writeIn_NORTH), .B(n325), .Y(N21) );
  NOR2BX1TS U769 ( .AN(readIn_NORTH), .B(n325), .Y(N20) );
  INVX2TS U770 ( .A(n218), .Y(n219) );
  NOR2BX1TS U771 ( .AN(requesterAddressIn_NORTH[0]), .B(n219), .Y(N16) );
  NOR2BX1TS U772 ( .AN(requesterAddressIn_NORTH[1]), .B(n219), .Y(N17) );
  NOR2BX1TS U773 ( .AN(requesterAddressIn_NORTH[2]), .B(n219), .Y(N18) );
  NOR2BX1TS U774 ( .AN(requesterAddressIn_NORTH[3]), .B(n219), .Y(N19) );
  NOR2BX1TS U775 ( .AN(destinationAddressIn_NORTH[0]), .B(n668), .Y(N4) );
  NOR2BX1TS U776 ( .AN(destinationAddressIn_NORTH[1]), .B(n667), .Y(N5) );
  NOR2BX1TS U777 ( .AN(destinationAddressIn_NORTH[2]), .B(n669), .Y(N6) );
  NOR2BX1TS U778 ( .AN(destinationAddressIn_NORTH[3]), .B(n158), .Y(N7) );
  INVX2TS U779 ( .A(n223), .Y(n221) );
  NOR2BX1TS U780 ( .AN(destinationAddressIn_NORTH[4]), .B(n221), .Y(N8) );
  NOR2BX1TS U781 ( .AN(destinationAddressIn_NORTH[5]), .B(n221), .Y(N9) );
  NOR2BX1TS U782 ( .AN(destinationAddressIn_NORTH[6]), .B(n221), .Y(N10) );
  NOR2BX1TS U783 ( .AN(destinationAddressIn_NORTH[7]), .B(n221), .Y(N11) );
  CLKBUFX2TS U784 ( .A(destinationAddressIn_NORTH[8]), .Y(n222) );
  INVX2TS U785 ( .A(n223), .Y(n227) );
  NOR2BX1TS U786 ( .AN(n222), .B(n227), .Y(N12) );
  CLKBUFX2TS U787 ( .A(destinationAddressIn_NORTH[9]), .Y(n224) );
  NOR2BX1TS U788 ( .AN(n224), .B(n227), .Y(N13) );
  CLKBUFX2TS U789 ( .A(destinationAddressIn_NORTH[10]), .Y(n225) );
  NOR2BX1TS U790 ( .AN(n225), .B(n227), .Y(N14) );
  CLKBUFX2TS U791 ( .A(destinationAddressIn_NORTH[11]), .Y(n226) );
  NOR2BX1TS U792 ( .AN(n226), .B(n227), .Y(N15) );
  CLKBUFX2TS U793 ( .A(localRouterAddress[2]), .Y(n259) );
  INVX2TS U794 ( .A(n259), .Y(n298) );
  CLKBUFX2TS U795 ( .A(localRouterAddress[3]), .Y(n228) );
  INVX2TS U796 ( .A(n228), .Y(n229) );
  INVX2TS U797 ( .A(n229), .Y(n317) );
  CLKAND2X2TS U798 ( .A(n226), .B(n229), .Y(n243) );
  INVX2TS U799 ( .A(n259), .Y(n314) );
  INVX2TS U800 ( .A(n317), .Y(n267) );
  OAI22X1TS U801 ( .A0(n225), .A1(n314), .B0(n226), .B1(n267), .Y(n239) );
  AOI211XLTS U802 ( .A0(n225), .A1(n298), .B0(n243), .C0(n239), .Y(n252) );
  CLKBUFX2TS U803 ( .A(localRouterAddress[1]), .Y(n231) );
  INVX2TS U804 ( .A(n232), .Y(n302) );
  INVX2TS U805 ( .A(n231), .Y(n335) );
  OR2X1TS U806 ( .A(n230), .B(n335), .Y(n235) );
  CLKBUFX2TS U807 ( .A(localRouterAddress[0]), .Y(n233) );
  INVX2TS U808 ( .A(n233), .Y(n324) );
  INVX2TS U809 ( .A(n302), .Y(n336) );
  AOI22X1TS U810 ( .A0(n222), .A1(n324), .B0(n230), .B1(n336), .Y(n234) );
  INVX2TS U811 ( .A(n233), .Y(n322) );
  OR2X1TS U812 ( .A(n222), .B(n322), .Y(n248) );
  NAND4XLTS U813 ( .A(n252), .B(n235), .C(n234), .D(n248), .Y(n250) );
  NOR2XLTS U814 ( .A(n289), .B(n250), .Y(n258) );
  NOR3XLTS U815 ( .A(n326), .B(n434), .C(n433), .Y(n237) );
  OAI21XLTS U816 ( .A0(readInBuffer_NORTH), .A1(writeInBuffer_NORTH), .B0(n238), .Y(n246) );
  INVX2TS U817 ( .A(n246), .Y(n251) );
  NAND2X1TS U818 ( .A(n251), .B(n239), .Y(n242) );
  OAI2BB2XLTS U819 ( .B0(n243), .B1(n242), .A0N(outputPortSelect_NORTH[0]), 
        .A1N(n241), .Y(n95) );
  OR2X1TS U820 ( .A(n226), .B(n267), .Y(n244) );
  AOI31XLTS U821 ( .A0(n225), .A1(n314), .A2(n244), .B0(n243), .Y(n247) );
  OAI2BB2XLTS U822 ( .B0(n247), .B1(n246), .A0N(n237), .A1N(
        outputPortSelect_NORTH[1]), .Y(n94) );
  INVX2TS U823 ( .A(n302), .Y(n316) );
  CLKAND2X2TS U824 ( .A(n224), .B(n316), .Y(n249) );
  OAI22X1TS U825 ( .A0(n224), .A1(n232), .B0(n249), .B1(n248), .Y(n254) );
  NAND3XLTS U826 ( .A(n252), .B(n251), .C(n250), .Y(n257) );
  OAI2BB2XLTS U827 ( .B0(n254), .B1(n257), .A0N(n241), .A1N(
        outputPortSelect_NORTH[2]), .Y(n93) );
  INVX2TS U828 ( .A(n254), .Y(n256) );
  OAI2BB2XLTS U829 ( .B0(n257), .B1(n256), .A0N(outputPortSelect_NORTH[3]), 
        .A1N(n241), .Y(n92) );
  INVX2TS U830 ( .A(n259), .Y(n318) );
  NOR2BX1TS U831 ( .AN(n214), .B(n228), .Y(n268) );
  OAI22X1TS U832 ( .A0(n213), .A1(n298), .B0(n214), .B1(n267), .Y(n264) );
  AOI211XLTS U833 ( .A0(n213), .A1(n318), .B0(n268), .C0(n264), .Y(n277) );
  AOI22X1TS U834 ( .A0(n210), .A1(n324), .B0(n260), .B1(n335), .Y(n262) );
  OR2X1TS U835 ( .A(n260), .B(n335), .Y(n261) );
  OR2X1TS U836 ( .A(n210), .B(n322), .Y(n273) );
  NAND4XLTS U837 ( .A(n277), .B(n262), .C(n261), .D(n273), .Y(n275) );
  NOR2XLTS U838 ( .A(n289), .B(n275), .Y(n285) );
  NOR3XLTS U839 ( .A(n326), .B(n435), .C(writeInBuffer_SOUTH), .Y(n279) );
  CLKBUFX2TS U840 ( .A(n279), .Y(n284) );
  OAI21XLTS U841 ( .A0(readInBuffer_SOUTH), .A1(writeInBuffer_SOUTH), .B0(n263), .Y(n271) );
  INVX2TS U842 ( .A(n271), .Y(n276) );
  NAND2X1TS U843 ( .A(n276), .B(n264), .Y(n266) );
  OAI2BB2XLTS U844 ( .B0(n268), .B1(n266), .A0N(outputPortSelect_SOUTH[0]), 
        .A1N(n279), .Y(n89) );
  OR2X1TS U845 ( .A(n214), .B(n267), .Y(n269) );
  AOI31XLTS U846 ( .A0(n213), .A1(n318), .A2(n269), .B0(n268), .Y(n272) );
  OAI2BB2XLTS U847 ( .B0(n272), .B1(n271), .A0N(n279), .A1N(
        outputPortSelect_SOUTH[1]), .Y(n88) );
  NOR2BX1TS U848 ( .AN(n212), .B(n302), .Y(n274) );
  OAI22X1TS U849 ( .A0(n212), .A1(n316), .B0(n274), .B1(n273), .Y(n280) );
  NAND3XLTS U850 ( .A(n277), .B(n276), .C(n275), .Y(n283) );
  OAI2BB2XLTS U851 ( .B0(n280), .B1(n283), .A0N(n279), .A1N(
        outputPortSelect_SOUTH[2]), .Y(n87) );
  INVX2TS U852 ( .A(n280), .Y(n282) );
  OAI2BB2XLTS U853 ( .B0(n283), .B1(n282), .A0N(outputPortSelect_SOUTH[3]), 
        .A1N(n284), .Y(n86) );
  NOR2BX1TS U854 ( .AN(n203), .B(n228), .Y(n296) );
  OAI22X1TS U855 ( .A0(n202), .A1(n318), .B0(n203), .B1(n229), .Y(n293) );
  AOI211XLTS U856 ( .A0(n202), .A1(n314), .B0(n296), .C0(n293), .Y(n307) );
  AOI22X1TS U857 ( .A0(n199), .A1(n324), .B0(n286), .B1(n232), .Y(n288) );
  OR2X1TS U858 ( .A(n286), .B(n316), .Y(n287) );
  OR2X1TS U859 ( .A(n199), .B(n322), .Y(n303) );
  NAND4XLTS U860 ( .A(n307), .B(n288), .C(n287), .D(n303), .Y(n305) );
  NOR2XLTS U861 ( .A(n289), .B(n305), .Y(n313) );
  NOR3XLTS U862 ( .A(n326), .B(n391), .C(n386), .Y(n290) );
  OAI21XLTS U863 ( .A0(n390), .A1(n385), .B0(n292), .Y(n300) );
  INVX2TS U864 ( .A(n300), .Y(n306) );
  NAND2X1TS U865 ( .A(n306), .B(n293), .Y(n295) );
  OAI2BB2XLTS U866 ( .B0(n296), .B1(n295), .A0N(outputPortSelect_EAST[0]), 
        .A1N(n290), .Y(n83) );
  OR2X1TS U867 ( .A(n203), .B(n229), .Y(n297) );
  AOI31XLTS U868 ( .A0(n202), .A1(n298), .A2(n297), .B0(n296), .Y(n301) );
  OAI2BB2XLTS U869 ( .B0(n301), .B1(n300), .A0N(n294), .A1N(
        outputPortSelect_EAST[1]), .Y(n82) );
  NOR2BX1TS U870 ( .AN(n201), .B(n302), .Y(n304) );
  OAI22X1TS U871 ( .A0(n201), .A1(n336), .B0(n304), .B1(n303), .Y(n309) );
  NAND3XLTS U872 ( .A(n307), .B(n306), .C(n305), .Y(n312) );
  OAI2BB2XLTS U873 ( .B0(n309), .B1(n312), .A0N(n290), .A1N(
        outputPortSelect_EAST[2]), .Y(n81) );
  INVX2TS U874 ( .A(n309), .Y(n311) );
  OAI2BB2XLTS U875 ( .B0(n312), .B1(n311), .A0N(outputPortSelect_EAST[3]), 
        .A1N(n294), .Y(n80) );
  NAND2X1TS U876 ( .A(n191), .B(n314), .Y(n338) );
  INVX2TS U877 ( .A(n338), .Y(n333) );
  NOR2XLTS U878 ( .A(n315), .B(n316), .Y(n319) );
  INVX2TS U879 ( .A(n317), .Y(n320) );
  OAI22X1TS U880 ( .A0(n191), .A1(n318), .B0(n192), .B1(n320), .Y(n342) );
  AOI211XLTS U881 ( .A0(n315), .A1(n336), .B0(n319), .C0(n342), .Y(n321) );
  NAND2X1TS U882 ( .A(n192), .B(n320), .Y(n339) );
  OAI211XLTS U883 ( .A0(n187), .A1(n322), .B0(n321), .C0(n339), .Y(n323) );
  AOI211XLTS U884 ( .A0(n187), .A1(n324), .B0(n333), .C0(n323), .Y(n343) );
  NOR2BX1TS U885 ( .AN(n343), .B(n325), .Y(n347) );
  NOR3XLTS U886 ( .A(n326), .B(n437), .C(n436), .Y(n327) );
  AO22XLTS U887 ( .A0(writeInBuffer_WEST), .A1(n347), .B0(n330), .B1(
        memWrite_WEST), .Y(n78) );
  OAI21XLTS U888 ( .A0(readInBuffer_WEST), .A1(writeInBuffer_WEST), .B0(n329), 
        .Y(n341) );
  NAND2X1TS U889 ( .A(n342), .B(n339), .Y(n331) );
  OAI2BB2XLTS U890 ( .B0(n341), .B1(n331), .A0N(n330), .A1N(
        outputPortSelect_WEST[0]), .Y(n77) );
  INVX2TS U891 ( .A(n339), .Y(n332) );
  OAI22X1TS U892 ( .A0(n333), .A1(n332), .B0(n192), .B1(n320), .Y(n334) );
  OAI2BB2XLTS U893 ( .B0(n334), .B1(n341), .A0N(n330), .A1N(
        outputPortSelect_WEST[1]), .Y(n76) );
  NAND2X1TS U894 ( .A(n315), .B(n335), .Y(n337) );
  AOI2BB2XLTS U895 ( .B0(n188), .B1(n337), .A0N(n315), .A1N(n336), .Y(n345) );
  NAND2X1TS U896 ( .A(n339), .B(n338), .Y(n340) );
  NOR4XLTS U897 ( .A(n343), .B(n342), .C(n341), .D(n340), .Y(n344) );
  INVX2TS U898 ( .A(n344), .Y(n346) );
  OAI2BB2XLTS U899 ( .B0(n346), .B1(n345), .A0N(outputPortSelect_WEST[3]), 
        .A1N(n330), .Y(n74) );
  AO22XLTS U900 ( .A0(readInBuffer_WEST), .A1(n347), .B0(n327), .B1(
        memRead_WEST), .Y(n73) );
endmodule

