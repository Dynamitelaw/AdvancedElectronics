

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO router 
  PIN localRouterAddress[5] 
    ANTENNAPARTIALMETALAREA 2.04 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.696 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.94 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.878 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 48.8 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 162.096 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.72 LAYER MQ ; 
    ANTENNAMAXAREACAR 239.936 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 867.291 LAYER MQ ;
    ANTENNAMAXCUTCAR 2.6732 LAYER VQ ;
  END localRouterAddress[5]
  PIN localRouterAddress[4] 
    ANTENNAPARTIALMETALAREA 0.24 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.62 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.694 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 75.52 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 250.8 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0368 LAYER MQ ; 
    ANTENNAMAXAREACAR 131.732 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 460.725 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAMAXCUTCAR 2.61728 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 120.48 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 398.112 LAYER MG ;
    ANTENNAGATEAREA 1.3824 LAYER MG ; 
    ANTENNAMAXAREACAR 218.884 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 748.711 LAYER MG ;
    ANTENNAMAXCUTCAR 2.61728 LAYER FY ;
  END localRouterAddress[4]
  PIN localRouterAddress[3] 
    ANTENNAPARTIALMETALAREA 0.32 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.184 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.98 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.326 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 88.8 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 295.152 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9072 LAYER MQ ; 
    ANTENNAMAXAREACAR 174.972 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 612.528 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAMAXCUTCAR 4.34303 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 119.84 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 396 LAYER MG ;
    ANTENNAGATEAREA 1.2096 LAYER MG ; 
    ANTENNAMAXAREACAR 274.046 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 939.909 LAYER MG ;
    ANTENNAMAXCUTCAR 4.34303 LAYER FY ;
  END localRouterAddress[3]
  PIN localRouterAddress[2] 
    ANTENNAPARTIALMETALAREA 10.44 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 38.776 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 194.324 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3984 LAYER M3 ; 
    ANTENNAMAXAREACAR 194.853 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 727.44 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER VL ;
    ANTENNAMAXCUTCAR 2.02273 LAYER VL ;
    ANTENNAPARTIALMETALAREA 53.12 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 176.352 LAYER MQ ;
    ANTENNAGATEAREA 0.7968 LAYER MQ ; 
    ANTENNAMAXAREACAR 261.52 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 948.765 LAYER MQ ;
    ANTENNAMAXCUTCAR 2.02273 LAYER VQ ;
  END localRouterAddress[2]
  PIN localRouterAddress[1] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.78 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.286 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 77.6 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 260.304 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8064 LAYER MQ ; 
    ANTENNAMAXAREACAR 181.067 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 639.391 LAYER MQ ;
    ANTENNAMAXCUTCAR 2.38095 LAYER VQ ;
  END localRouterAddress[1]
  PIN localRouterAddress[0] 
    ANTENNAPARTIALMETALAREA 27.64 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 102.416 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0696 LAYER M3 ; 
    ANTENNAMAXAREACAR 8.75862 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 33.8161 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.14943 LAYER VL ;
  END localRouterAddress[0]
  PIN destinationAddressIn_NORTH[13] 
    ANTENNAPARTIALMETALAREA 8.76 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 32.412 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.98 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.326 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 59.68 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 198 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 0.96 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 4.224 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 LAYER MG ; 
    ANTENNAMAXAREACAR 26.5194 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 112.041 LAYER MG ;
    ANTENNAMAXCUTCAR 6.94444 LAYER FY ;
  END destinationAddressIn_NORTH[13]
  PIN destinationAddressIn_NORTH[12] 
    ANTENNAPARTIALMETALAREA 9.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 33.67 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.78 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.886 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 33.12 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 109.824 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 2.88 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 12.672 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 LAYER MG ; 
    ANTENNAMAXAREACAR 84.3221 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 320.921 LAYER MG ;
    ANTENNAMAXCUTCAR 9.72222 LAYER FY ;
  END destinationAddressIn_NORTH[12]
  PIN destinationAddressIn_NORTH[11] 
    ANTENNAPARTIALMETALAREA 39.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 147.186 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.504 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3744 LAYER M3 ; 
    ANTENNAMAXAREACAR 21.8886 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 81.0612 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END destinationAddressIn_NORTH[11]
  PIN destinationAddressIn_NORTH[10] 
    ANTENNAPARTIALMETALAREA 10.66 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 39.442 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.46 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.702 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 25.12 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 83.424 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 3.36 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 14.784 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 LAYER MG ; 
    ANTENNAMAXAREACAR 95.0401 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 363.219 LAYER MG ;
    ANTENNAMAXCUTCAR 9.72222 LAYER FY ;
  END destinationAddressIn_NORTH[10]
  PIN destinationAddressIn_NORTH[9] 
    ANTENNAPARTIALMETALAREA 9.4 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 34.78 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.1 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.07 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 34.72 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 115.104 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 2.88 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 12.672 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 LAYER MG ; 
    ANTENNAMAXAREACAR 86.0582 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 325.123 LAYER MG ;
    ANTENNAMAXCUTCAR 9.72222 LAYER FY ;
  END destinationAddressIn_NORTH[9]
  PIN destinationAddressIn_NORTH[8] 
    ANTENNAPARTIALMETALAREA 6.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.57 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.02 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.874 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 67.68 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 224.4 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.32 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 4.64 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 16.896 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2304 LAYER MG ; 
    ANTENNAMAXAREACAR 45.7356 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 175.453 LAYER MG ;
    ANTENNAMAXCUTCAR 6.94444 LAYER FY ;
  END destinationAddressIn_NORTH[8]
  PIN destinationAddressIn_NORTH[7] 
    ANTENNAPARTIALMETALAREA 7.04 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 26.196 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.184 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 40.5 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 155.222 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END destinationAddressIn_NORTH[7]
  PIN destinationAddressIn_NORTH[6] 
    ANTENNAPARTIALMETALAREA 7.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 26.418 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 8.38 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 31.006 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 34.24 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 114.048 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 0.96 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 4.224 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER MG ; 
    ANTENNAMAXAREACAR 95.0139 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 370.743 LAYER MG ;
    ANTENNAMAXCUTCAR 6.94444 LAYER FY ;
  END destinationAddressIn_NORTH[6]
  PIN destinationAddressIn_NORTH[5] 
    ANTENNAPARTIALMETALAREA 4.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.688 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 75.9167 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 283.694 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END destinationAddressIn_NORTH[5]
  PIN destinationAddressIn_NORTH[4] 
    ANTENNAPARTIALMETALAREA 3.42 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.802 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 62.375 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 233.59 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END destinationAddressIn_NORTH[4]
  PIN destinationAddressIn_NORTH[3] 
    ANTENNAPARTIALMETALAREA 6.24 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.236 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 111.333 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 414.736 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END destinationAddressIn_NORTH[3]
  PIN destinationAddressIn_NORTH[2] 
    ANTENNAPARTIALMETALAREA 5.98 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.274 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 106.819 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 398.035 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END destinationAddressIn_NORTH[2]
  PIN destinationAddressIn_NORTH[1] 
    ANTENNAPARTIALMETALAREA 5.58 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.794 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 99.875 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 372.34 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END destinationAddressIn_NORTH[1]
  PIN destinationAddressIn_NORTH[0] 
    ANTENNAPARTIALMETALAREA 6.46 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 24.05 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.48 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 21.0556 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 83.2778 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END destinationAddressIn_NORTH[0]
  PIN requesterAddressIn_NORTH[5] 
    ANTENNAPARTIALMETALAREA 6.96 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 25.9 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 123.833 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 460.986 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END requesterAddressIn_NORTH[5]
  PIN requesterAddressIn_NORTH[4] 
    ANTENNAPARTIALMETALAREA 7.66 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 28.49 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 135.986 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 505.951 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END requesterAddressIn_NORTH[4]
  PIN requesterAddressIn_NORTH[3] 
    ANTENNAPARTIALMETALAREA 6.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.162 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 110.986 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 413.451 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END requesterAddressIn_NORTH[3]
  PIN requesterAddressIn_NORTH[2] 
    ANTENNAPARTIALMETALAREA 6.42 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.902 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 114.458 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 426.299 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END requesterAddressIn_NORTH[2]
  PIN requesterAddressIn_NORTH[1] 
    ANTENNAPARTIALMETALAREA 8.04 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 29.896 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 142.583 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 530.361 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END requesterAddressIn_NORTH[1]
  PIN requesterAddressIn_NORTH[0] 
    ANTENNAPARTIALMETALAREA 6.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.754 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 113.764 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 423.729 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END requesterAddressIn_NORTH[0]
  PIN dataIn_NORTH[31] 
    ANTENNAPARTIALMETALAREA 5.7 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 21.09 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.98 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.774 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 29.0417 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 112.826 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_NORTH[31]
  PIN dataIn_NORTH[30] 
    ANTENNAPARTIALMETALAREA 5.9 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 21.83 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.032 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 57.1667 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 216.889 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_NORTH[30]
  PIN dataIn_NORTH[29] 
    ANTENNAPARTIALMETALAREA 4.84 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.908 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.216 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 43.2778 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 165.5 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_NORTH[29]
  PIN dataIn_NORTH[28] 
    ANTENNAPARTIALMETALAREA 5.7 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 21.09 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.368 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 34.9444 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 134.667 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_NORTH[28]
  PIN dataIn_NORTH[27] 
    ANTENNAPARTIALMETALAREA 6.26 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.162 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.26 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.11 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 59.5972 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 225.882 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_NORTH[27]
  PIN dataIn_NORTH[26] 
    ANTENNAPARTIALMETALAREA 6.58 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 24.346 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.22 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 18.9722 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 75.5694 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_NORTH[26]
  PIN dataIn_NORTH[25] 
    ANTENNAPARTIALMETALAREA 5.96 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.052 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.552 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 48.8333 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 186.056 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_NORTH[25]
  PIN dataIn_NORTH[24] 
    ANTENNAPARTIALMETALAREA 2.58 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.546 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.216 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 52.3056 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 201.472 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_NORTH[24]
  PIN dataIn_NORTH[23] 
    ANTENNAPARTIALMETALAREA 7.64 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 28.268 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 135.639 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 502.097 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END dataIn_NORTH[23]
  PIN dataIn_NORTH[22] 
    ANTENNAPARTIALMETALAREA 5.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.498 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 98.4861 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 367.201 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END dataIn_NORTH[22]
  PIN dataIn_NORTH[21] 
    ANTENNAPARTIALMETALAREA 5.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.498 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 98.4861 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 367.201 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END dataIn_NORTH[21]
  PIN dataIn_NORTH[20] 
    ANTENNAPARTIALMETALAREA 8.7 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 32.338 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 154.042 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 572.757 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END dataIn_NORTH[20]
  PIN dataIn_NORTH[19] 
    ANTENNAPARTIALMETALAREA 7.8 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 28.86 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.848 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 30.7778 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 119.25 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_NORTH[19]
  PIN dataIn_NORTH[18] 
    ANTENNAPARTIALMETALAREA 6.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.162 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 110.986 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 413.451 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END dataIn_NORTH[18]
  PIN dataIn_NORTH[17] 
    ANTENNAPARTIALMETALAREA 5.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.498 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 98.4861 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 367.201 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END dataIn_NORTH[17]
  PIN dataIn_NORTH[16] 
    ANTENNAPARTIALMETALAREA 5.7 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 21.09 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.368 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 22.4444 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 88.4167 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_NORTH[16]
  PIN dataIn_NORTH[15] 
    ANTENNAPARTIALMETALAREA 4.78 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.834 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 85.9861 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 320.951 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END dataIn_NORTH[15]
  PIN dataIn_NORTH[14] 
    ANTENNAPARTIALMETALAREA 6.42 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.754 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.516 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 50.9167 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 193.764 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_NORTH[14]
  PIN dataIn_NORTH[13] 
    ANTENNAPARTIALMETALAREA 7.44 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 27.528 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 132.167 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 489.25 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END dataIn_NORTH[13]
  PIN dataIn_NORTH[12] 
    ANTENNAPARTIALMETALAREA 7.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 26.122 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 125.569 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 464.84 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END dataIn_NORTH[12]
  PIN dataIn_NORTH[11] 
    ANTENNAPARTIALMETALAREA 6.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.976 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.184 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 9.94444 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 42.1667 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_NORTH[11]
  PIN dataIn_NORTH[10] 
    ANTENNAPARTIALMETALAREA 4.54 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.798 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.48 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 32.1667 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 124.389 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_NORTH[10]
  PIN dataIn_NORTH[9] 
    ANTENNAPARTIALMETALAREA 4.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.576 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 80.7778 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 299.111 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END dataIn_NORTH[9]
  PIN dataIn_NORTH[8] 
    ANTENNAPARTIALMETALAREA 3.34 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.506 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 60.9861 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 228.451 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END dataIn_NORTH[8]
  PIN dataIn_NORTH[7] 
    ANTENNAPARTIALMETALAREA 6.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.754 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 113.764 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 423.729 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END dataIn_NORTH[7]
  PIN dataIn_NORTH[6] 
    ANTENNAPARTIALMETALAREA 5.78 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 21.386 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 103.347 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 382.618 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END dataIn_NORTH[6]
  PIN dataIn_NORTH[5] 
    ANTENNAPARTIALMETALAREA 6.68 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 24.716 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 28 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 108.972 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_NORTH[5]
  PIN dataIn_NORTH[4] 
    ANTENNAPARTIALMETALAREA 6.82 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 25.234 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.184 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 9.94444 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 42.1667 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_NORTH[4]
  PIN dataIn_NORTH[3] 
    ANTENNAPARTIALMETALAREA 6.68 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 24.716 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.256 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 34.9444 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 134.667 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_NORTH[3]
  PIN dataIn_NORTH[2] 
    ANTENNAPARTIALMETALAREA 3.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.47 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.256 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 87.7222 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 329.944 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_NORTH[2]
  PIN dataIn_NORTH[1] 
    ANTENNAPARTIALMETALAREA 6.78 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 25.234 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 120.708 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 449.424 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END dataIn_NORTH[1]
  PIN dataIn_NORTH[0] 
    ANTENNAPARTIALMETALAREA 5.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 19.018 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.48 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 14.1111 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 57.5833 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_NORTH[0]
  PIN destinationAddressOut_NORTH[13] 
    ANTENNAPARTIALMETALAREA 0.26 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.962 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.48 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 2.112 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 41.12 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 136.224 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5588 LAYER MG ; 
    ANTENNAMAXAREACAR 28.6573 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 98.3986 LAYER MG ;
    ANTENNAMAXCUTCAR 0.552881 LAYER FY ;
  END destinationAddressOut_NORTH[13]
  PIN destinationAddressOut_NORTH[12] 
    ANTENNAPARTIALMETALAREA 5.26 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 19.61 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 24.42 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 90.502 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 32 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 106.128 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5588 LAYER MQ ; 
    ANTENNAMAXAREACAR 15.6713 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 57.1251 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.970885 LAYER VQ ;
  END destinationAddressOut_NORTH[12]
  PIN destinationAddressOut_NORTH[11] 
    ANTENNAPARTIALMETALAREA 3.44 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.728 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 22.94 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 84.878 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 29.12 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 96.624 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5588 LAYER MQ ; 
    ANTENNAMAXAREACAR 62.4281 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 230.611 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.739403 LAYER VQ ;
  END destinationAddressOut_NORTH[11]
  PIN destinationAddressOut_NORTH[10] 
    ANTENNAPARTIALMETALAREA 4.34 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.058 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 13.94 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 51.726 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 4.32 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 14.784 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5588 LAYER MQ ; 
    ANTENNAMAXAREACAR 15.2543 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 59.3044 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.28768 LAYER VQ ;
  END destinationAddressOut_NORTH[10]
  PIN destinationAddressOut_NORTH[9] 
    ANTENNAPARTIALMETALAREA 4.46 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.65 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 10.54 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 38.998 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 2.72 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 9.504 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 22.56 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 74.976 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5588 LAYER MG ; 
    ANTENNAMAXAREACAR 21.1475 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 74.3534 LAYER MG ;
    ANTENNAMAXCUTCAR 0.552881 LAYER FY ;
  END destinationAddressOut_NORTH[9]
  PIN destinationAddressOut_NORTH[8] 
    ANTENNAPARTIALMETALAREA 0.7 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.738 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 53.28 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 176.352 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5588 LAYER MQ ; 
    ANTENNAMAXAREACAR 17.6493 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 58.7753 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.28768 LAYER VQ ;
  END destinationAddressOut_NORTH[8]
  PIN destinationAddressOut_NORTH[7] 
    ANTENNAPARTIALMETALAREA 0.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.85 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.664 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 13.12 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 43.824 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 43.36 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 143.616 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5588 LAYER MG ; 
    ANTENNAMAXAREACAR 22.546 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 77.3766 LAYER MG ;
    ANTENNAMAXCUTCAR 0.552881 LAYER FY ;
  END destinationAddressOut_NORTH[7]
  PIN destinationAddressOut_NORTH[6] 
    ANTENNAPARTIALMETALAREA 2.34 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.658 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 20.7 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 76.59 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 47.04 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 155.76 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5588 LAYER MQ ; 
    ANTENNAMAXAREACAR 25.1055 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 89.4126 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.507922 LAYER VQ ;
  END destinationAddressOut_NORTH[6]
  PIN destinationAddressOut_NORTH[5] 
    ANTENNAPARTIALMETALAREA 3.68 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.616 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 14.7 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 54.39 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.8 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 3.168 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 57.76 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 191.136 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 31.7713 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 105.986 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END destinationAddressOut_NORTH[5]
  PIN destinationAddressOut_NORTH[4] 
    ANTENNAPARTIALMETALAREA 2.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.954 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 31.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 104.016 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 10.2769 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 34.4098 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END destinationAddressOut_NORTH[4]
  PIN destinationAddressOut_NORTH[3] 
    ANTENNAPARTIALMETALAREA 2.4 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.028 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 40.16 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 133.056 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 18.4 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 61.248 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 6.20724 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 20.9822 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END destinationAddressOut_NORTH[3]
  PIN destinationAddressOut_NORTH[2] 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 45.1 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 166.87 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 28.96 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 96.096 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 11.0507 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 37.5563 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END destinationAddressOut_NORTH[2]
  PIN destinationAddressOut_NORTH[1] 
    ANTENNAPARTIALMETALAREA 2.28 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.584 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 35.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 117.216 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 11.0507 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 36.8002 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END destinationAddressOut_NORTH[1]
  PIN destinationAddressOut_NORTH[0] 
    ANTENNAPARTIALMETALAREA 2.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.066 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 52.42 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 193.954 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 33.6 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 111.408 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 10.7436 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 35.8717 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END destinationAddressOut_NORTH[0]
  PIN requesterAddressOut_NORTH[5] 
    ANTENNAPARTIALMETALAREA 6.4 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.828 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M2 ; 
    ANTENNAMAXAREACAR 2.04303 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 7.49309 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0118133 LAYER V2 ;
  END requesterAddressOut_NORTH[5]
  PIN requesterAddressOut_NORTH[4] 
    ANTENNAPARTIALMETALAREA 6.7 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 24.938 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M2 ; 
    ANTENNAMAXAREACAR 2.13163 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 7.82091 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0118133 LAYER V2 ;
  END requesterAddressOut_NORTH[4]
  PIN requesterAddressOut_NORTH[3] 
    ANTENNAPARTIALMETALAREA 0.4 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.48 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 44.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 164.576 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 14.7542 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 54.5681 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END requesterAddressOut_NORTH[3]
  PIN requesterAddressOut_NORTH[2] 
    ANTENNAPARTIALMETALAREA 0.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.518 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 42.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 158.656 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 14.8251 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 54.8304 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END requesterAddressOut_NORTH[2]
  PIN requesterAddressOut_NORTH[1] 
    ANTENNAPARTIALMETALAREA 0.52 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.924 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 12.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 47.064 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 5.62247 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 20.8245 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END requesterAddressOut_NORTH[1]
  PIN requesterAddressOut_NORTH[0] 
    ANTENNAPARTIALMETALAREA 5.66 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 21.09 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M2 ; 
    ANTENNAMAXAREACAR 1.82448 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 6.68447 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0118133 LAYER V2 ;
  END requesterAddressOut_NORTH[0]
  PIN dataOut_NORTH[31] 
    ANTENNAPARTIALMETALAREA 3.84 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.208 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 32.3 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 119.51 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 54.4 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 180.048 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 17.0283 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 56.6679 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END dataOut_NORTH[31]
  PIN dataOut_NORTH[30] 
    ANTENNAPARTIALMETALAREA 3.46 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.802 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.18 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.48 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 2.112 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 57.12 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 189.024 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 49.4441 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 163.834 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_NORTH[30]
  PIN dataOut_NORTH[29] 
    ANTENNAPARTIALMETALAREA 2.34 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.658 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.48 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 2.112 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 67.36 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 222.816 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 42.0489 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 139.496 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_NORTH[29]
  PIN dataOut_NORTH[28] 
    ANTENNAPARTIALMETALAREA 5.42 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.202 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.024 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.48 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 2.112 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 37.6 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 124.608 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 33.7796 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 112.453 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_NORTH[28]
  PIN dataOut_NORTH[27] 
    ANTENNAPARTIALMETALAREA 0.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.85 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.036 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 3.2 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 11.088 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 97.12 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 321.024 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 46.2072 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 153.483 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_NORTH[27]
  PIN dataOut_NORTH[26] 
    ANTENNAPARTIALMETALAREA 3.78 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.986 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.26 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.962 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.48 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 2.112 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 67.04 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 221.76 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 39.072 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 129.445 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_NORTH[26]
  PIN dataOut_NORTH[25] 
    ANTENNAPARTIALMETALAREA 2.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.954 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 81.76 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 270.336 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 29.92 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 99.264 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 10.3183 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 34.7943 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_NORTH[25]
  PIN dataOut_NORTH[24] 
    ANTENNAPARTIALMETALAREA 2.66 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.842 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 32.3 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 119.51 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 5.92 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 20.064 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 47.2 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 157.344 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 32.1494 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 107.338 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_NORTH[24]
  PIN dataOut_NORTH[23] 
    ANTENNAPARTIALMETALAREA 0.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.85 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 1.6 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 5.808 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 95.2 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 314.688 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 49.7985 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 165.07 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_NORTH[23]
  PIN dataOut_NORTH[22] 
    ANTENNAPARTIALMETALAREA 2.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.066 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.5 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.85 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 10.72 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 35.904 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 114.08 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 376.992 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 56.0832 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 185.639 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_NORTH[22]
  PIN dataOut_NORTH[21] 
    ANTENNAPARTIALMETALAREA 4.66 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.242 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.64 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 2.64 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 107.52 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 355.872 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 47.4358 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 157.656 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_NORTH[21]
  PIN dataOut_NORTH[20] 
    ANTENNAPARTIALMETALAREA 3.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.618 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.48 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 2.112 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 115.84 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 383.328 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 45.9237 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 152.212 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_NORTH[20]
  PIN dataOut_NORTH[19] 
    ANTENNAPARTIALMETALAREA 5.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 18.722 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.036 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.48 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 2.112 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 95.84 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 316.8 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 57.2409 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 190.735 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_NORTH[19]
  PIN dataOut_NORTH[18] 
    ANTENNAPARTIALMETALAREA 0.12 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 48.8 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 161.568 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 14.8074 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 49.1121 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END dataOut_NORTH[18]
  PIN dataOut_NORTH[17] 
    ANTENNAPARTIALMETALAREA 2.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.362 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 67.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 222.816 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 20.5959 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 68.3372 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END dataOut_NORTH[17]
  PIN dataOut_NORTH[16] 
    ANTENNAPARTIALMETALAREA 2.78 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.434 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 29.34 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 108.558 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 41.12 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 136.224 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 30.72 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 102.432 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 10.0111 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 33.7193 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_NORTH[16]
  PIN dataOut_NORTH[15] 
    ANTENNAPARTIALMETALAREA 5.28 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 19.536 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.26 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.662 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 4 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 13.728 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 105.76 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 350.592 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 39.5209 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 131.305 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_NORTH[15]
  PIN dataOut_NORTH[14] 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.37 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.18 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.48 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 2.112 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 121.76 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 402.336 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 56.9338 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 188.616 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_NORTH[14]
  PIN dataOut_NORTH[13] 
    ANTENNAPARTIALMETALAREA 5.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.276 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.74 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.438 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.96 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 3.696 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 123.68 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 408.672 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 60.7849 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 201.599 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_NORTH[13]
  PIN dataOut_NORTH[12] 
    ANTENNAPARTIALMETALAREA 2.58 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.842 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 76.96 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 254.496 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 24.5534 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 81.8894 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END dataOut_NORTH[12]
  PIN dataOut_NORTH[11] 
    ANTENNAPARTIALMETALAREA 6 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.2 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.22 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.614 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 22.4 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 74.448 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 73.44 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 242.88 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 46.6892 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 154.995 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_NORTH[11]
  PIN dataOut_NORTH[10] 
    ANTENNAPARTIALMETALAREA 3.9 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.43 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.62 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.694 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.96 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 3.696 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 67.2 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 222.816 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 30.59 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 101.847 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_NORTH[10]
  PIN dataOut_NORTH[9] 
    ANTENNAPARTIALMETALAREA 3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.1 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 38.02 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 140.822 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 89.76 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 296.736 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 27.359 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 90.7146 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END dataOut_NORTH[9]
  PIN dataOut_NORTH[8] 
    ANTENNAPARTIALMETALAREA 0.08 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.296 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.18 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.766 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 2.08 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 7.392 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 73.76 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 243.936 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 45.8292 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 151.971 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_NORTH[8]
  PIN dataOut_NORTH[7] 
    ANTENNAPARTIALMETALAREA 0.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.85 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.48 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 2.112 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 70.88 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 234.432 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 48.0737 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 159.898 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_NORTH[7]
  PIN dataOut_NORTH[6] 
    ANTENNAPARTIALMETALAREA 5.82 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 21.534 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 41.82 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 154.734 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 87.04 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 287.76 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 26.5144 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 87.9544 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END dataOut_NORTH[6]
  PIN dataOut_NORTH[5] 
    ANTENNAPARTIALMETALAREA 4.44 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.428 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 32.86 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 121.582 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.48 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 2.112 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 1.76 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 6.336 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 29.2905 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 97.9603 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_NORTH[5]
  PIN dataOut_NORTH[4] 
    ANTENNAPARTIALMETALAREA 6.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.57 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.78 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 17.686 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 47.68 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 157.872 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 61.44 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 203.808 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 30.6845 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 102.65 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_NORTH[4]
  PIN dataOut_NORTH[3] 
    ANTENNAPARTIALMETALAREA 4.72 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.464 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.7 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 17.39 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.48 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 2.112 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 85.6 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 283.008 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 54.1458 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 179.586 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_NORTH[3]
  PIN dataOut_NORTH[2] 
    ANTENNAPARTIALMETALAREA 0.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.85 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.26 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.962 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 2.56 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 8.976 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 92.96 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 307.296 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 59.7217 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 197.684 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_NORTH[2]
  PIN dataOut_NORTH[1] 
    ANTENNAPARTIALMETALAREA 3.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.876 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 7.9 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 29.23 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 1.76 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 6.336 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 77.28 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 255.552 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 55.6815 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 184.096 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_NORTH[1]
  PIN dataOut_NORTH[0] 
    ANTENNAPARTIALMETALAREA 6.26 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.162 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.5 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.35 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 51.84 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 171.6 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 64.8 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 214.368 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 26.8806 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 89.4594 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_NORTH[0]
  PIN destinationAddressIn_SOUTH[13] 
    ANTENNAPARTIALMETALAREA 6.76 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 25.012 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.032 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 LAYER M3 ; 
    ANTENNAMAXAREACAR 16.4684 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 64.8701 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END destinationAddressIn_SOUTH[13]
  PIN destinationAddressIn_SOUTH[12] 
    ANTENNAPARTIALMETALAREA 17.8 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 65.86 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 9.76 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 32.736 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 LAYER MQ ; 
    ANTENNAMAXAREACAR 110.377 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 389.31 LAYER MQ ;
    ANTENNAMAXCUTCAR 2.64675 LAYER VQ ;
  END destinationAddressIn_SOUTH[12]
  PIN destinationAddressIn_SOUTH[11] 
    ANTENNAPARTIALMETALAREA 35.08 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 129.796 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.512 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3744 LAYER M3 ; 
    ANTENNAMAXAREACAR 28.8286 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 108.442 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.14943 LAYER VL ;
  END destinationAddressIn_SOUTH[11]
  PIN destinationAddressIn_SOUTH[10] 
    ANTENNAPARTIALMETALAREA 3.7 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.69 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.46 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.702 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 45.28 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 149.952 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 3.04 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 12.672 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 LAYER MG ; 
    ANTENNAMAXAREACAR 153.34 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 578.392 LAYER MG ;
    ANTENNAMAXCUTCAR 4.23986 LAYER FY ;
  END destinationAddressIn_SOUTH[10]
  PIN destinationAddressIn_SOUTH[9] 
    ANTENNAPARTIALMETALAREA 37.88 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 140.156 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.184 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 LAYER M3 ; 
    ANTENNAMAXAREACAR 8.92128 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 34.6185 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END destinationAddressIn_SOUTH[9]
  PIN destinationAddressIn_SOUTH[8] 
    ANTENNAPARTIALMETALAREA 12.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 45.658 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.8 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 3.168 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2304 LAYER MQ ; 
    ANTENNAMAXAREACAR 94.0272 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 353.185 LAYER MQ ;
    ANTENNAMAXCUTCAR 3.36111 LAYER VQ ;
  END destinationAddressIn_SOUTH[8]
  PIN destinationAddressIn_SOUTH[7] 
    ANTENNAPARTIALMETALAREA 8.76 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 32.412 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.88 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 59.9444 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 227.167 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END destinationAddressIn_SOUTH[7]
  PIN destinationAddressIn_SOUTH[6] 
    ANTENNAPARTIALMETALAREA 9.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 34.114 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 16.8889 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 67.8611 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END destinationAddressIn_SOUTH[6]
  PIN destinationAddressIn_SOUTH[5] 
    ANTENNAPARTIALMETALAREA 3.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.322 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 55.4306 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 207.896 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END destinationAddressIn_SOUTH[5]
  PIN destinationAddressIn_SOUTH[4] 
    ANTENNAPARTIALMETALAREA 4.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 18.278 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.208 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 86.3333 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 324.806 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END destinationAddressIn_SOUTH[4]
  PIN destinationAddressIn_SOUTH[3] 
    ANTENNAPARTIALMETALAREA 4.54 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.946 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 81.8194 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 305.535 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END destinationAddressIn_SOUTH[3]
  PIN destinationAddressIn_SOUTH[2] 
    ANTENNAPARTIALMETALAREA 3.78 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.986 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.88 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 68.2778 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 258 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END destinationAddressIn_SOUTH[2]
  PIN destinationAddressIn_SOUTH[1] 
    ANTENNAPARTIALMETALAREA 3.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.986 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 67.9306 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 254.146 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END destinationAddressIn_SOUTH[1]
  PIN destinationAddressIn_SOUTH[0] 
    ANTENNAPARTIALMETALAREA 6.62 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 24.642 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 117.931 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 439.146 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END destinationAddressIn_SOUTH[0]
  PIN requesterAddressIn_SOUTH[5] 
    ANTENNAPARTIALMETALAREA 24.84 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 91.908 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.184 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 36.3333 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 139.806 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END requesterAddressIn_SOUTH[5]
  PIN requesterAddressIn_SOUTH[4] 
    ANTENNAPARTIALMETALAREA 6.82 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 25.234 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.94 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.478 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 30.4 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 100.848 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 0.96 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 4.224 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER MG ; 
    ANTENNAMAXAREACAR 92.2361 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 354.91 LAYER MG ;
    ANTENNAMAXCUTCAR 6.94444 LAYER FY ;
  END requesterAddressIn_SOUTH[4]
  PIN requesterAddressIn_SOUTH[3] 
    ANTENNAPARTIALMETALAREA 23.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 85.914 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 1.44 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 5.28 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER MQ ; 
    ANTENNAMAXAREACAR 80.0833 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 298.278 LAYER MQ ;
    ANTENNAMAXCUTCAR 4.16667 LAYER VQ ;
  END requesterAddressIn_SOUTH[3]
  PIN requesterAddressIn_SOUTH[2] 
    ANTENNAPARTIALMETALAREA 17.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 64.898 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.736 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 25.2222 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 103.833 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END requesterAddressIn_SOUTH[2]
  PIN requesterAddressIn_SOUTH[1] 
    ANTENNAPARTIALMETALAREA 24.56 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 90.872 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 34.9444 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 134.667 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END requesterAddressIn_SOUTH[1]
  PIN requesterAddressIn_SOUTH[0] 
    ANTENNAPARTIALMETALAREA 3.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.578 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.62 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.694 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 30.72 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 101.904 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 0.96 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 4.224 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER MG ; 
    ANTENNAMAXAREACAR 111.681 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 429.076 LAYER MG ;
    ANTENNAMAXCUTCAR 6.94444 LAYER FY ;
  END requesterAddressIn_SOUTH[0]
  PIN dataIn_SOUTH[31] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 38.24 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 127.248 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 0.48 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 2.112 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER MG ; 
    ANTENNAMAXAREACAR 243.625 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 888.104 LAYER MG ;
    ANTENNAMAXCUTCAR 6.94444 LAYER FY ;
  END dataIn_SOUTH[31]
  PIN dataIn_SOUTH[30] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.18 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 43.52 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 144.672 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 0.48 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 2.112 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER MG ; 
    ANTENNAMAXAREACAR 192.931 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 687.549 LAYER MG ;
    ANTENNAMAXCUTCAR 6.94444 LAYER FY ;
  END dataIn_SOUTH[30]
  PIN dataIn_SOUTH[29] 
    ANTENNAPARTIALMETALAREA 2.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.658 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 42.9306 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 161.646 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END dataIn_SOUTH[29]
  PIN dataIn_SOUTH[28] 
    ANTENNAPARTIALMETALAREA 2.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.658 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 42.9306 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 161.646 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END dataIn_SOUTH[28]
  PIN dataIn_SOUTH[27] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 14.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 55.204 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 1.44 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 6.336 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 0.48 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 2.112 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER MG ; 
    ANTENNAMAXAREACAR 45.0139 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 181.021 LAYER MG ;
    ANTENNAMAXCUTCAR 6.94444 LAYER FY ;
  END dataIn_SOUTH[27]
  PIN dataIn_SOUTH[26] 
    ANTENNAPARTIALMETALAREA 3.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.95 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 15.06 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 55.87 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.48 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 2.112 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 1.28 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 5.28 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER MG ; 
    ANTENNAMAXAREACAR 64.4583 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 256.576 LAYER MG ;
    ANTENNAMAXCUTCAR 6.94444 LAYER FY ;
  END dataIn_SOUTH[26]
  PIN dataIn_SOUTH[25] 
    ANTENNAPARTIALMETALAREA 3.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.322 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 55.4306 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 207.896 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END dataIn_SOUTH[25]
  PIN dataIn_SOUTH[24] 
    ANTENNAPARTIALMETALAREA 4.7 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.538 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 84.5972 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 315.812 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END dataIn_SOUTH[24]
  PIN dataIn_SOUTH[23] 
    ANTENNAPARTIALMETALAREA 3.82 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.282 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 69.3194 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 259.285 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END dataIn_SOUTH[23]
  PIN dataIn_SOUTH[22] 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 12.7 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 47.138 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 1.92 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 8.448 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER MQ ; 
    ANTENNAMAXAREACAR 90.1528 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 362.271 LAYER MQ ;
    ANTENNAMAXCUTCAR 4.16667 LAYER VQ ;
  END dataIn_SOUTH[22]
  PIN dataIn_SOUTH[21] 
    ANTENNAPARTIALMETALAREA 3.04 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.396 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 55.7778 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 209.181 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END dataIn_SOUTH[21]
  PIN dataIn_SOUTH[20] 
    ANTENNAPARTIALMETALAREA 3.42 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.802 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 62.375 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 233.59 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END dataIn_SOUTH[20]
  PIN dataIn_SOUTH[19] 
    ANTENNAPARTIALMETALAREA 2.46 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.25 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 45.7083 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 171.924 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END dataIn_SOUTH[19]
  PIN dataIn_SOUTH[18] 
    ANTENNAPARTIALMETALAREA 4.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.022 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 72.7917 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 272.132 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END dataIn_SOUTH[18]
  PIN dataIn_SOUTH[17] 
    ANTENNAPARTIALMETALAREA 2.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.954 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 44.3194 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 166.785 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END dataIn_SOUTH[17]
  PIN dataIn_SOUTH[16] 
    ANTENNAPARTIALMETALAREA 3.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.914 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 58.2083 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 218.174 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END dataIn_SOUTH[16]
  PIN dataIn_SOUTH[15] 
    ANTENNAPARTIALMETALAREA 4.8 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.76 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 11.1 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 41.366 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 1.44 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 6.336 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 0.48 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 2.112 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER MG ; 
    ANTENNAMAXAREACAR 176.264 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 669.215 LAYER MG ;
    ANTENNAMAXCUTCAR 6.94444 LAYER FY ;
  END dataIn_SOUTH[15]
  PIN dataIn_SOUTH[14] 
    ANTENNAPARTIALMETALAREA 3.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.766 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 8.78 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 32.486 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.48 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 2.112 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 4.32 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 14.784 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER MG ; 
    ANTENNAMAXAREACAR 107.514 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 385.604 LAYER MG ;
    ANTENNAMAXCUTCAR 6.94444 LAYER FY ;
  END dataIn_SOUTH[14]
  PIN dataIn_SOUTH[13] 
    ANTENNAPARTIALMETALAREA 2.62 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.842 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 48.4861 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 182.201 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END dataIn_SOUTH[13]
  PIN dataIn_SOUTH[12] 
    ANTENNAPARTIALMETALAREA 4.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.318 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 74.875 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 277.271 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END dataIn_SOUTH[12]
  PIN dataIn_SOUTH[11] 
    ANTENNAPARTIALMETALAREA 2.36 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.88 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 43.9722 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 165.5 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END dataIn_SOUTH[11]
  PIN dataIn_SOUTH[10] 
    ANTENNAPARTIALMETALAREA 2.78 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.286 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.34 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.958 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.48 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 2.112 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 2.4 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 8.448 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER MG ; 
    ANTENNAMAXAREACAR 195.014 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 722.687 LAYER MG ;
    ANTENNAMAXCUTCAR 6.94444 LAYER FY ;
  END dataIn_SOUTH[10]
  PIN dataIn_SOUTH[9] 
    ANTENNAPARTIALMETALAREA 2.6 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.768 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 48.1389 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 180.917 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END dataIn_SOUTH[9]
  PIN dataIn_SOUTH[8] 
    ANTENNAPARTIALMETALAREA 2.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.138 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.48 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 39.1111 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 150.083 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_SOUTH[8]
  PIN dataIn_SOUTH[7] 
    ANTENNAPARTIALMETALAREA 3.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.322 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 55.4306 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 207.896 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END dataIn_SOUTH[7]
  PIN dataIn_SOUTH[6] 
    ANTENNAPARTIALMETALAREA 2.46 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.25 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 45.7083 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 171.924 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END dataIn_SOUTH[6]
  PIN dataIn_SOUTH[5] 
    ANTENNAPARTIALMETALAREA 3.84 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.208 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 69.6667 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 258 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END dataIn_SOUTH[5]
  PIN dataIn_SOUTH[4] 
    ANTENNAPARTIALMETALAREA 6.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.57 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 108.208 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 403.174 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END dataIn_SOUTH[4]
  PIN dataIn_SOUTH[3] 
    ANTENNAPARTIALMETALAREA 5.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.276 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 98.1389 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 363.347 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END dataIn_SOUTH[3]
  PIN dataIn_SOUTH[2] 
    ANTENNAPARTIALMETALAREA 2.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.51 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 42.9306 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 159.076 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END dataIn_SOUTH[2]
  PIN dataIn_SOUTH[1] 
    ANTENNAPARTIALMETALAREA 6.8 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 25.16 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 121.056 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 448.139 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END dataIn_SOUTH[1]
  PIN dataIn_SOUTH[0] 
    ANTENNAPARTIALMETALAREA 6.98 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 25.826 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.48 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 30.7778 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 119.25 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_SOUTH[0]
  PIN destinationAddressOut_SOUTH[13] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.292 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 67.2 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 222.288 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5588 LAYER MQ ; 
    ANTENNAMAXAREACAR 22.6543 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 76.0817 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.28768 LAYER VQ ;
  END destinationAddressOut_SOUTH[13]
  PIN destinationAddressOut_SOUTH[12] 
    ANTENNAPARTIALMETALAREA 2.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.214 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.02 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.174 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 82.88 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 274.032 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5588 LAYER MQ ; 
    ANTENNAMAXAREACAR 26.5938 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 89.3991 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.507922 LAYER VQ ;
  END destinationAddressOut_SOUTH[12]
  PIN destinationAddressOut_SOUTH[11] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 81.76 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 270.336 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 7.84 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 26.4 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5588 LAYER MG ; 
    ANTENNAMAXAREACAR 8.39035 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 32.1391 LAYER MG ;
    ANTENNAMAXCUTCAR 0.552881 LAYER FY ;
  END destinationAddressOut_SOUTH[11]
  PIN destinationAddressOut_SOUTH[10] 
    ANTENNAPARTIALMETALAREA 5.86 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 21.682 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.46 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.702 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 71.2 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 235.488 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5588 LAYER MQ ; 
    ANTENNAMAXAREACAR 22.578 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 74.997 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.28768 LAYER VQ ;
  END destinationAddressOut_SOUTH[10]
  PIN destinationAddressOut_SOUTH[9] 
    ANTENNAPARTIALMETALAREA 4.82 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.834 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.288 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 74.4 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 246.048 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5588 LAYER MQ ; 
    ANTENNAMAXAREACAR 30.6271 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 105.196 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.507922 LAYER VQ ;
  END destinationAddressOut_SOUTH[9]
  PIN destinationAddressOut_SOUTH[8] 
    ANTENNAPARTIALMETALAREA 2.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.77 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.3 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.81 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 67.84 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 224.4 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5588 LAYER MQ ; 
    ANTENNAMAXAREACAR 24.8314 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 85.1143 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.28768 LAYER VQ ;
  END destinationAddressOut_SOUTH[8]
  PIN destinationAddressOut_SOUTH[7] 
    ANTENNAPARTIALMETALAREA 2.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.138 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 66.4 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 219.648 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5588 LAYER MQ ; 
    ANTENNAMAXAREACAR 25.6242 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 88.9937 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.507922 LAYER VQ ;
  END destinationAddressOut_SOUTH[7]
  PIN destinationAddressOut_SOUTH[6] 
    ANTENNAPARTIALMETALAREA 2.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.77 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.1 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.47 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 64.96 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 214.896 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5588 LAYER MQ ; 
    ANTENNAMAXAREACAR 21.1168 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 70.2921 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.28768 LAYER VQ ;
  END destinationAddressOut_SOUTH[6]
  PIN destinationAddressOut_SOUTH[5] 
    ANTENNAPARTIALMETALAREA 3.58 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.394 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M2 ; 
    ANTENNAMAXAREACAR 1.21019 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 4.41158 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0118133 LAYER V2 ;
  END destinationAddressOut_SOUTH[5]
  PIN destinationAddressOut_SOUTH[4] 
    ANTENNAPARTIALMETALAREA 3.66 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.69 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M2 ; 
    ANTENNAMAXAREACAR 1.23382 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 4.499 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0118133 LAYER V2 ;
  END destinationAddressOut_SOUTH[4]
  PIN destinationAddressOut_SOUTH[3] 
    ANTENNAPARTIALMETALAREA 3.96 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.652 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 24.864 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.30292 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 8.49841 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END destinationAddressOut_SOUTH[3]
  PIN destinationAddressOut_SOUTH[2] 
    ANTENNAPARTIALMETALAREA 3.7 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.69 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.984 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.73588 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 6.40035 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END destinationAddressOut_SOUTH[2]
  PIN destinationAddressOut_SOUTH[1] 
    ANTENNAPARTIALMETALAREA 5.24 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 19.388 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M2 ; 
    ANTENNAMAXAREACAR 1.70044 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 6.18181 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0118133 LAYER V2 ;
  END destinationAddressOut_SOUTH[1]
  PIN destinationAddressOut_SOUTH[0] 
    ANTENNAPARTIALMETALAREA 5.26 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 19.61 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M2 ; 
    ANTENNAMAXAREACAR 1.70635 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 6.24737 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0118133 LAYER V2 ;
  END destinationAddressOut_SOUTH[0]
  PIN requesterAddressOut_SOUTH[5] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.036 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 47.04 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 155.76 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 14.3112 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 47.4842 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END requesterAddressOut_SOUTH[5]
  PIN requesterAddressOut_SOUTH[4] 
    ANTENNAPARTIALMETALAREA 4.42 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.354 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.62 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 24.494 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 39.52 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 130.944 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 12.0962 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 40.1771 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END requesterAddressOut_SOUTH[4]
  PIN requesterAddressOut_SOUTH[3] 
    ANTENNAPARTIALMETALAREA 3.08 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.396 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.06 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 22.422 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 35.84 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 118.8 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 11.7418 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 39.3005 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END requesterAddressOut_SOUTH[3]
  PIN requesterAddressOut_SOUTH[2] 
    ANTENNAPARTIALMETALAREA 2.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.622 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.14 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.918 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 42.72 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 141.504 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 13.1771 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 43.7985 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END requesterAddressOut_SOUTH[2]
  PIN requesterAddressOut_SOUTH[1] 
    ANTENNAPARTIALMETALAREA 1.88 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.956 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.5 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.55 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 43.68 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 144.672 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 13.2716 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 44.0347 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END requesterAddressOut_SOUTH[1]
  PIN requesterAddressOut_SOUTH[0] 
    ANTENNAPARTIALMETALAREA 2.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.25 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.62 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.694 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 43.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 143.616 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 13.2952 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 44.16 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END requesterAddressOut_SOUTH[0]
  PIN dataOut_SOUTH[31] 
    ANTENNAPARTIALMETALAREA 3.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.84 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 10.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 40.552 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.63783 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 13.5687 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END dataOut_SOUTH[31]
  PIN dataOut_SOUTH[30] 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.18 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.64 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 2.64 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 13.28 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 44.352 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 25.3685 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 84.4506 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_SOUTH[30]
  PIN dataOut_SOUTH[29] 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.772 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 78.24 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 258.72 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 23.5965 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 78.154 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END dataOut_SOUTH[29]
  PIN dataOut_SOUTH[28] 
    ANTENNAPARTIALMETALAREA 1.86 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.882 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.1 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.07 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 60.48 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 200.112 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 15.2 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 50.688 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 7.30588 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 25.0908 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_SOUTH[28]
  PIN dataOut_SOUTH[27] 
    ANTENNAPARTIALMETALAREA 6.54 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 24.346 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 11.78 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 43.734 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 27.84 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 92.4 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 12.4211 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 42.7589 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END dataOut_SOUTH[27]
  PIN dataOut_SOUTH[26] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.18 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 54.88 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 181.632 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 18.08 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 60.192 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 10.4837 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 35.3874 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_SOUTH[26]
  PIN dataOut_SOUTH[25] 
    ANTENNAPARTIALMETALAREA 2.8 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.36 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 9.14 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 33.966 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 55.04 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 182.16 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 17.6071 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 58.7778 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END dataOut_SOUTH[25]
  PIN dataOut_SOUTH[24] 
    ANTENNAPARTIALMETALAREA 3.78 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.986 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.7 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 17.39 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 66.56 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 220.176 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 20.147 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 66.7707 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END dataOut_SOUTH[24]
  PIN dataOut_SOUTH[23] 
    ANTENNAPARTIALMETALAREA 2.24 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.288 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 10.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 39.368 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 9.60357 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 35.5108 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END dataOut_SOUTH[23]
  PIN dataOut_SOUTH[22] 
    ANTENNAPARTIALMETALAREA 2.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.214 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.3 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.11 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 39.84 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 132 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 12.7436 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 42.5467 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END dataOut_SOUTH[22]
  PIN dataOut_SOUTH[21] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.8 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 3.168 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 14.88 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 49.632 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 19.7099 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 68.7175 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_SOUTH[21]
  PIN dataOut_SOUTH[20] 
    ANTENNAPARTIALMETALAREA 2.66 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.842 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.94 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 25.678 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 70.08 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 231.792 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 21.7772 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 72.3868 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END dataOut_SOUTH[20]
  PIN dataOut_SOUTH[19] 
    ANTENNAPARTIALMETALAREA 2.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.14 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.94 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.478 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 43.04 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 142.56 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 13.5079 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 44.9845 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END dataOut_SOUTH[19]
  PIN dataOut_SOUTH[18] 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.9 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.33 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 52.8 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 174.768 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 25.76 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 85.536 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 10.8853 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 36.3442 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_SOUTH[18]
  PIN dataOut_SOUTH[17] 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.37 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 39.2 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 129.888 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 13.5315 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 45.5256 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END dataOut_SOUTH[17]
  PIN dataOut_SOUTH[16] 
    ANTENNAPARTIALMETALAREA 19.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 70.818 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 2.56 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 8.976 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 1.88355 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 6.75653 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END dataOut_SOUTH[16]
  PIN dataOut_SOUTH[15] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 6.88 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 23.232 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 15.84 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 52.8 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 17.4535 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 59.1015 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_SOUTH[15]
  PIN dataOut_SOUTH[14] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.18 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 2.08 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 7.392 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 26.08 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 86.592 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 21.5504 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 72.3961 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_SOUTH[14]
  PIN dataOut_SOUTH[13] 
    ANTENNAPARTIALMETALAREA 2.24 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.436 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M2 ; 
    ANTENNAMAXAREACAR 0.814442 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 2.94731 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0118133 LAYER V2 ;
  END dataOut_SOUTH[13]
  PIN dataOut_SOUTH[12] 
    ANTENNAPARTIALMETALAREA 2.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.066 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M2 ; 
    ANTENNAMAXAREACAR 0.784908 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 2.83804 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0118133 LAYER V2 ;
  END dataOut_SOUTH[12]
  PIN dataOut_SOUTH[11] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.036 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 11.68 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 39.072 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 28 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 92.928 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 17.9379 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 59.6473 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_SOUTH[11]
  PIN dataOut_SOUTH[10] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.26 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.962 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.48 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 2.112 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 34.08 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 112.992 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 22.4801 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 74.8091 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_SOUTH[10]
  PIN dataOut_SOUTH[9] 
    ANTENNAPARTIALMETALAREA 2.04 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.548 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 21 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 77.848 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 6.39034 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 23.6219 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END dataOut_SOUTH[9]
  PIN dataOut_SOUTH[8] 
    ANTENNAPARTIALMETALAREA 2.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.954 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M2 ; 
    ANTENNAMAXAREACAR 0.855789 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 3.1003 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0118133 LAYER V2 ;
  END dataOut_SOUTH[8]
  PIN dataOut_SOUTH[7] 
    ANTENNAPARTIALMETALAREA 2.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.362 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M2 ; 
    ANTENNAMAXAREACAR 0.808535 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 2.92546 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0118133 LAYER V2 ;
  END dataOut_SOUTH[7]
  PIN dataOut_SOUTH[6] 
    ANTENNAPARTIALMETALAREA 2.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.288 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M2 ; 
    ANTENNAMAXAREACAR 0.835706 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 3.03816 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0118133 LAYER V2 ;
  END dataOut_SOUTH[6]
  PIN dataOut_SOUTH[5] 
    ANTENNAPARTIALMETALAREA 2.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.658 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M2 ; 
    ANTENNAMAXAREACAR 0.832162 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 3.01288 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0118133 LAYER V2 ;
  END dataOut_SOUTH[5]
  PIN dataOut_SOUTH[4] 
    ANTENNAPARTIALMETALAREA 4.54 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.946 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M2 ; 
    ANTENNAMAXAREACAR 1.49371 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 5.4606 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0118133 LAYER V2 ;
  END dataOut_SOUTH[4]
  PIN dataOut_SOUTH[3] 
    ANTENNAPARTIALMETALAREA 2.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.14 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M2 ; 
    ANTENNAMAXAREACAR 0.790815 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 2.85989 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0118133 LAYER V2 ;
  END dataOut_SOUTH[3]
  PIN dataOut_SOUTH[2] 
    ANTENNAPARTIALMETALAREA 3.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.914 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M2 ; 
    ANTENNAMAXAREACAR 1.09206 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 3.97448 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0118133 LAYER V2 ;
  END dataOut_SOUTH[2]
  PIN dataOut_SOUTH[1] 
    ANTENNAPARTIALMETALAREA 3.64 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.616 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M2 ; 
    ANTENNAMAXAREACAR 1.22791 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 4.47714 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0118133 LAYER V2 ;
  END dataOut_SOUTH[1]
  PIN dataOut_SOUTH[0] 
    ANTENNAPARTIALMETALAREA 3.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.618 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M2 ; 
    ANTENNAMAXAREACAR 1.06843 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 3.88706 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0118133 LAYER V2 ;
  END dataOut_SOUTH[0]
  PIN destinationAddressIn_EAST[13] 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.37 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 12.3 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 45.51 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 47.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 159.456 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 2.4 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 10.56 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 LAYER MG ; 
    ANTENNAMAXAREACAR 112.604 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 432.426 LAYER MG ;
    ANTENNAMAXCUTCAR 4.59906 LAYER FY ;
  END destinationAddressIn_EAST[13]
  PIN destinationAddressIn_EAST[12] 
    ANTENNAPARTIALMETALAREA 6.32 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.532 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 34.58 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 128.39 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 1.28 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 4.752 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 1.92 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 8.448 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 LAYER MG ; 
    ANTENNAMAXAREACAR 156.236 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 595.248 LAYER MG ;
    ANTENNAMAXCUTCAR 4.59906 LAYER FY ;
  END destinationAddressIn_EAST[12]
  PIN destinationAddressIn_EAST[11] 
    ANTENNAPARTIALMETALAREA 6.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.754 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 7.62 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 28.342 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 120.912 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3744 LAYER MQ ; 
    ANTENNAMAXAREACAR 164.45 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 576.083 LAYER MQ ;
    ANTENNAMAXCUTCAR 1.81624 LAYER VQ ;
  END destinationAddressIn_EAST[11]
  PIN destinationAddressIn_EAST[10] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 19.9 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 73.926 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 16.8 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 55.968 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 1.92 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 8.448 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 LAYER MG ; 
    ANTENNAMAXAREACAR 153.121 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 580.466 LAYER MG ;
    ANTENNAMAXCUTCAR 3.90461 LAYER FY ;
  END destinationAddressIn_EAST[10]
  PIN destinationAddressIn_EAST[9] 
    ANTENNAPARTIALMETALAREA 12.34 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 45.806 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 27.62 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 102.342 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 25.92 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 87.12 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 1.92 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 8.448 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 LAYER MG ; 
    ANTENNAMAXAREACAR 82.5185 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 316.731 LAYER MG ;
    ANTENNAMAXCUTCAR 3.90461 LAYER FY ;
  END destinationAddressIn_EAST[9]
  PIN destinationAddressIn_EAST[8] 
    ANTENNAPARTIALMETALAREA 0.12 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.444 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 48.3 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 179.006 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 34.08 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 112.992 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 2.88 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 12.672 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2304 LAYER MG ; 
    ANTENNAMAXAREACAR 113.614 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 431.924 LAYER MG ;
    ANTENNAMAXCUTCAR 2.77778 LAYER FY ;
  END destinationAddressIn_EAST[8]
  PIN destinationAddressIn_EAST[7] 
    ANTENNAPARTIALMETALAREA 8.46 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 31.45 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.664 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 19.6667 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 78.1389 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END destinationAddressIn_EAST[7]
  PIN destinationAddressIn_EAST[6] 
    ANTENNAPARTIALMETALAREA 5.72 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 21.312 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 102.306 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 381.333 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END destinationAddressIn_EAST[6]
  PIN destinationAddressIn_EAST[5] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 7.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 26.64 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 148.833 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 556.056 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END destinationAddressIn_EAST[5]
  PIN destinationAddressIn_EAST[4] 
    ANTENNAPARTIALMETALAREA 0.12 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.444 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 7.7 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 28.638 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 138.764 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 518.799 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END destinationAddressIn_EAST[4]
  PIN destinationAddressIn_EAST[3] 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.37 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 15.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 58.756 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.48 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 2.112 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 4 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 13.728 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER MG ; 
    ANTENNAMAXAREACAR 120.014 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 434.076 LAYER MG ;
    ANTENNAMAXCUTCAR 6.94444 LAYER FY ;
  END destinationAddressIn_EAST[3]
  PIN destinationAddressIn_EAST[2] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 13.42 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 49.654 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.96 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 4.224 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 1.28 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 5.28 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER MG ; 
    ANTENNAMAXAREACAR 61.6806 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 246.299 LAYER MG ;
    ANTENNAMAXCUTCAR 6.94444 LAYER FY ;
  END destinationAddressIn_EAST[2]
  PIN destinationAddressIn_EAST[1] 
    ANTENNAPARTIALMETALAREA 0.34 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.406 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.184 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 11.3333 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 47.3056 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END destinationAddressIn_EAST[1]
  PIN destinationAddressIn_EAST[0] 
    ANTENNAPARTIALMETALAREA 4.8 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.908 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 86.3333 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 322.236 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END destinationAddressIn_EAST[0]
  PIN requesterAddressIn_EAST[5] 
    ANTENNAPARTIALMETALAREA 16.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 59.866 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 7.16667 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 31.8889 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END requesterAddressIn_EAST[5]
  PIN requesterAddressIn_EAST[4] 
    ANTENNAPARTIALMETALAREA 15.88 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 58.904 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.312 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 125.222 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 468.694 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END requesterAddressIn_EAST[4]
  PIN requesterAddressIn_EAST[3] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.984 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 97.4444 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 371.056 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END requesterAddressIn_EAST[3]
  PIN requesterAddressIn_EAST[2] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.54 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.798 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 1.92 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 6.864 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER MQ ; 
    ANTENNAMAXAREACAR 57.5139 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 216.576 LAYER MQ ;
    ANTENNAMAXCUTCAR 4.16667 LAYER VQ ;
  END requesterAddressIn_EAST[2]
  PIN requesterAddressIn_EAST[1] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 8.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 30.488 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 160.639 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 602.306 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END requesterAddressIn_EAST[1]
  PIN requesterAddressIn_EAST[0] 
    ANTENNAPARTIALMETALAREA 17.96 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 66.6 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.136 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 65.5 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 247.722 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END requesterAddressIn_EAST[0]
  PIN dataIn_EAST[31] 
    ANTENNAPARTIALMETALAREA 2.96 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.952 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.584 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 44.6667 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 170.639 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_EAST[31]
  PIN dataIn_EAST[30] 
    ANTENNAPARTIALMETALAREA 1.28 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.884 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 25.2222 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 96.125 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END dataIn_EAST[30]
  PIN dataIn_EAST[29] 
    ANTENNAPARTIALMETALAREA 1.66 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.29 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 31.8194 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 120.535 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END dataIn_EAST[29]
  PIN dataIn_EAST[28] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.24 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 94.6667 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 355.639 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_EAST[28]
  PIN dataIn_EAST[27] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.728 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 68.2778 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 258 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_EAST[27]
  PIN dataIn_EAST[26] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.46 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.102 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 4.64 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 15.84 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER MQ ; 
    ANTENNAMAXAREACAR 96.75 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 337.722 LAYER MQ ;
    ANTENNAMAXCUTCAR 4.16667 LAYER VQ ;
  END dataIn_EAST[26]
  PIN dataIn_EAST[25] 
    ANTENNAPARTIALMETALAREA 0.12 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.444 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 9.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 33.744 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 168.278 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 628 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_EAST[25]
  PIN dataIn_EAST[24] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.28 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 93.2778 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 350.5 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_EAST[24]
  PIN dataIn_EAST[23] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.064 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 51.6111 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 196.333 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_EAST[23]
  PIN dataIn_EAST[22] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.904 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 114.111 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 427.583 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_EAST[22]
  PIN dataIn_EAST[21] 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.37 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.688 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 78 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 293.972 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_EAST[21]
  PIN dataIn_EAST[20] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 22.2 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 112.722 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 422.444 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_EAST[20]
  PIN dataIn_EAST[19] 
    ANTENNAPARTIALMETALAREA 0.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.518 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.472 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 48.8333 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 186.056 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_EAST[19]
  PIN dataIn_EAST[18] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 18.056 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 90.5 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 340.222 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_EAST[18]
  PIN dataIn_EAST[17] 
    ANTENNAPARTIALMETALAREA 0.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.518 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 22.496 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 109.944 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 412.167 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_EAST[17]
  PIN dataIn_EAST[16] 
    ANTENNAPARTIALMETALAREA 0.08 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.296 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.096 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 82.1667 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 309.389 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_EAST[16]
  PIN dataIn_EAST[15] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.976 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 116.889 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 437.861 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_EAST[15]
  PIN dataIn_EAST[14] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.88 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 53 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 201.472 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_EAST[14]
  PIN dataIn_EAST[13] 
    ANTENNAPARTIALMETALAREA 0.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.518 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 17.464 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 87.7222 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 329.944 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_EAST[13]
  PIN dataIn_EAST[12] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 22.2 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 115.5 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 432.722 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_EAST[12]
  PIN dataIn_EAST[11] 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.37 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 17.464 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 103 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 386.472 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_EAST[11]
  PIN dataIn_EAST[10] 
    ANTENNAPARTIALMETALAREA 0.88 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.404 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 18.2778 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 70.4306 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END dataIn_EAST[10]
  PIN dataIn_EAST[9] 
    ANTENNAPARTIALMETALAREA 0.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.518 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.064 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 84.25 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 319.667 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_EAST[9]
  PIN dataIn_EAST[8] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.976 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 116.889 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 437.861 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_EAST[8]
  PIN dataIn_EAST[7] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.088 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 121.75 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 458.417 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_EAST[7]
  PIN dataIn_EAST[6] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 17.464 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 86.3333 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 324.806 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_EAST[6]
  PIN dataIn_EAST[5] 
    ANTENNAPARTIALMETALAREA 0.9 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.478 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 18.625 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 71.7153 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END dataIn_EAST[5]
  PIN dataIn_EAST[4] 
    ANTENNAPARTIALMETALAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.738 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.28 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 101.611 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 381.333 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_EAST[4]
  PIN dataIn_EAST[3] 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.37 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.54 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.798 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 3.52 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 12.144 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER MQ ; 
    ANTENNAMAXAREACAR 92.5833 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 330.083 LAYER MQ ;
    ANTENNAMAXCUTCAR 4.16667 LAYER VQ ;
  END dataIn_EAST[3]
  PIN dataIn_EAST[2] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 24.272 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 162.722 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 607.444 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_EAST[2]
  PIN dataIn_EAST[1] 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.37 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 18.648 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 122.444 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 458.417 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_EAST[1]
  PIN dataIn_EAST[0] 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.088 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 112.722 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 422.444 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_EAST[0]
  PIN destinationAddressOut_EAST[13] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.38 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.406 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 25.12 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 83.952 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 71.2 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 235.488 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5588 LAYER MG ; 
    ANTENNAMAXAREACAR 32.9864 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 119.21 LAYER MG ;
    ANTENNAMAXCUTCAR 0.332639 LAYER FY ;
  END destinationAddressOut_EAST[13]
  PIN destinationAddressOut_EAST[12] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.86 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.182 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 103.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 341.616 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 62.24 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 205.92 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5588 LAYER MG ; 
    ANTENNAMAXAREACAR 25.0148 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 87.4451 LAYER MG ;
    ANTENNAMAXCUTCAR 0.332639 LAYER FY ;
  END destinationAddressOut_EAST[12]
  PIN destinationAddressOut_EAST[11] 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.37 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.66 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.142 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 99.68 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 329.472 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 75.36 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 249.216 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5588 LAYER MG ; 
    ANTENNAMAXAREACAR 27.8675 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 94.9562 LAYER MG ;
    ANTENNAMAXCUTCAR 0.552881 LAYER FY ;
  END destinationAddressOut_EAST[11]
  PIN destinationAddressOut_EAST[10] 
    ANTENNAPARTIALMETALAREA 13.64 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 50.616 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.02 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.774 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 63.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 209.616 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 53.92 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 178.464 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5588 LAYER MG ; 
    ANTENNAMAXAREACAR 25.7788 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 90.6974 LAYER MG ;
    ANTENNAMAXCUTCAR 0.552881 LAYER FY ;
  END destinationAddressOut_EAST[10]
  PIN destinationAddressOut_EAST[9] 
    ANTENNAPARTIALMETALAREA 8.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 30.118 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.3 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.11 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 13.6 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 45.936 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 56.48 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 186.912 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5588 LAYER MG ; 
    ANTENNAMAXAREACAR 20.8462 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 71.9438 LAYER MG ;
    ANTENNAMAXCUTCAR 0.552881 LAYER FY ;
  END destinationAddressOut_EAST[9]
  PIN destinationAddressOut_EAST[8] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.3 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.51 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 99.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 328.416 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 74.08 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 244.992 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5588 LAYER MG ; 
    ANTENNAMAXAREACAR 23.1343 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 76.8263 LAYER MG ;
    ANTENNAMAXCUTCAR 0.332639 LAYER FY ;
  END destinationAddressOut_EAST[8]
  PIN destinationAddressOut_EAST[7] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.1 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.47 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 102.56 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 338.976 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 44.64 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 147.84 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5588 LAYER MG ; 
    ANTENNAMAXAREACAR 20.6109 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 71.6136 LAYER MG ;
    ANTENNAMAXCUTCAR 0.552881 LAYER FY ;
  END destinationAddressOut_EAST[7]
  PIN destinationAddressOut_EAST[6] 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.22 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.614 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 100.96 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 333.696 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 42.72 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 141.504 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5588 LAYER MG ; 
    ANTENNAMAXAREACAR 17.9369 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 62.0735 LAYER MG ;
    ANTENNAMAXCUTCAR 0.332639 LAYER FY ;
  END destinationAddressOut_EAST[6]
  PIN destinationAddressOut_EAST[5] 
    ANTENNAPARTIALMETALAREA 35.26 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 130.758 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M2 ; 
    ANTENNAMAXAREACAR 10.5664 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 39.0731 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0118133 LAYER V2 ;
  END destinationAddressOut_EAST[5]
  PIN destinationAddressOut_EAST[4] 
    ANTENNAPARTIALMETALAREA 0.12 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.444 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 8.74 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 32.486 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 19.52 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 64.944 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 14.24 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 47.52 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 14.512 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 49.1641 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END destinationAddressOut_EAST[4]
  PIN destinationAddressOut_EAST[3] 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.37 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.34 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.958 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 65.12 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 215.424 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 28.64 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 95.04 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 9.11332 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 30.525 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END destinationAddressOut_EAST[3]
  PIN destinationAddressOut_EAST[2] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.22 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 62.4 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 206.448 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 50.4 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 166.848 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 15.782 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 52.4582 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END destinationAddressOut_EAST[2]
  PIN destinationAddressOut_EAST[1] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.14 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 22.718 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 61.92 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 204.864 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 20 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 66.528 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 6.75065 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 22.8038 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END destinationAddressOut_EAST[1]
  PIN destinationAddressOut_EAST[0] 
    ANTENNAPARTIALMETALAREA 9.84 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 36.556 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.22 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 9.6 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 32.208 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 7.5067 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 26.818 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END destinationAddressOut_EAST[0]
  PIN requesterAddressOut_EAST[5] 
    ANTENNAPARTIALMETALAREA 12.7 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 47.138 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.208 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 6.69749 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 24.7583 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END requesterAddressOut_EAST[5]
  PIN requesterAddressOut_EAST[4] 
    ANTENNAPARTIALMETALAREA 20.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 75.258 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.4 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.91308 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 7.0997 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END requesterAddressOut_EAST[4]
  PIN requesterAddressOut_EAST[3] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.9 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.43 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 7.84 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 26.4 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 3.56105 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 12.4269 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END requesterAddressOut_EAST[3]
  PIN requesterAddressOut_EAST[2] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.02 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.774 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 51.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 170.016 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 42.72 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 141.504 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 13.4606 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 44.9467 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END requesterAddressOut_EAST[2]
  PIN requesterAddressOut_EAST[1] 
    ANTENNAPARTIALMETALAREA 10.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 38.554 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 3.52 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 13.2 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 25.12 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 83.424 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 8.121 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 27.2692 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END requesterAddressOut_EAST[1]
  PIN requesterAddressOut_EAST[0] 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.128 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.48 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 2.112 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 0.8 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 3.168 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 3.17711 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 11.4588 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END requesterAddressOut_EAST[0]
  PIN dataOut_EAST[31] 
    ANTENNAPARTIALMETALAREA 0.86 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.182 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.5 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.35 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 17.28 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 57.552 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 23.2 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 77.088 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 13.8741 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 46.7093 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_EAST[31]
  PIN dataOut_EAST[30] 
    ANTENNAPARTIALMETALAREA 0.12 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.444 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.78 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 17.686 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 18.56 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 61.776 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 27.36 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 90.816 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 13.756 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 45.8753 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_EAST[30]
  PIN dataOut_EAST[29] 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.37 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 8.06 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 29.822 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 13.28 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 44.352 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 20 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 66.528 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 18.3041 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 60.7884 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_EAST[29]
  PIN dataOut_EAST[28] 
    ANTENNAPARTIALMETALAREA 19 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 70.448 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.98 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.774 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 5.28 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 17.952 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 24.8 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 82.368 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 8.62897 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 29.2302 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_EAST[28]
  PIN dataOut_EAST[27] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.14 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.918 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 78.56 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 259.776 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 54.56 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 180.576 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 16.8156 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 55.9615 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_EAST[27]
  PIN dataOut_EAST[26] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.34 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.758 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 12 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 40.128 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 41.44 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 137.28 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 29.5268 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 98.5321 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_EAST[26]
  PIN dataOut_EAST[25] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.46 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.102 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 60.16 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 199.584 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 55.84 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 184.8 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 19.5091 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 65.0767 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_EAST[25]
  PIN dataOut_EAST[24] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.54 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.998 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 3.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 11.616 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 55.52 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 183.744 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 37.5599 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 124.72 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_EAST[24]
  PIN dataOut_EAST[23] 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.37 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.74 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.838 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 73.28 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 242.352 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 47.84 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 158.4 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 16.8156 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 56.2261 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_EAST[23]
  PIN dataOut_EAST[22] 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.42 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.554 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 3.52 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 12.144 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 60.32 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 199.584 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 35.6934 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 118.267 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_EAST[22]
  PIN dataOut_EAST[21] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.62 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.694 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 48 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 158.928 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 57.76 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 191.136 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 20.0761 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 66.929 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_EAST[21]
  PIN dataOut_EAST[20] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.7 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.59 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 34.24 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 113.52 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 56.8 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 187.968 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 23.4311 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 77.9249 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_EAST[20]
  PIN dataOut_EAST[19] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.94 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.878 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 14.88 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 49.632 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 57.44 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 190.08 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 25.9355 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 86.4541 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_EAST[19]
  PIN dataOut_EAST[18] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.02 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.774 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 13.92 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 46.464 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 58.24 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 193.248 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 18.8239 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 62.8298 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_EAST[18]
  PIN dataOut_EAST[17] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.544 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 12.616 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 46.7004 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END dataOut_EAST[17]
  PIN dataOut_EAST[16] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.5 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.55 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 51.04 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 168.96 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 18.7766 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 63.5338 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END dataOut_EAST[16]
  PIN dataOut_EAST[15] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.54 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.798 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 17.28 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 57.552 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 42.4 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 140.448 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 34.9137 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 116.328 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_EAST[15]
  PIN dataOut_EAST[14] 
    ANTENNAPARTIALMETALAREA 29.36 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 108.78 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.184 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.52324 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 5.61359 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END dataOut_EAST[14]
  PIN dataOut_EAST[13] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.38 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.206 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 77.12 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 255.024 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 53.92 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 178.464 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 16.916 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 56.3141 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_EAST[13]
  PIN dataOut_EAST[12] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.984 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.35431 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 12.4323 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END dataOut_EAST[12]
  PIN dataOut_EAST[11] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.06 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.022 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 22.24 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 73.92 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 9.04244 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 30.9196 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END dataOut_EAST[11]
  PIN dataOut_EAST[10] 
    ANTENNAPARTIALMETALAREA 0.12 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.444 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 7.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 27.232 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.30706 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 12.2574 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END dataOut_EAST[10]
  PIN dataOut_EAST[9] 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.37 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.088 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.00759 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 7.44938 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END dataOut_EAST[9]
  PIN dataOut_EAST[8] 
    ANTENNAPARTIALMETALAREA 11.4 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 42.328 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.48 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.14522 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 4.21488 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END dataOut_EAST[8]
  PIN dataOut_EAST[7] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 10.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 40.848 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.54333 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 13.1316 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END dataOut_EAST[7]
  PIN dataOut_EAST[6] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.22 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 23.68 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 78.672 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 27.36 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 90.816 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 11.665 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 39.7205 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_EAST[6]
  PIN dataOut_EAST[5] 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.37 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.74 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.838 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 6.56 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 22.176 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 36 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 119.328 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 19.5091 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 64.831 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_EAST[5]
  PIN dataOut_EAST[4] 
    ANTENNAPARTIALMETALAREA 0.66 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.442 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.46 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.902 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 6.56 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 22.176 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 33.76 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 111.936 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 17.8552 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 59.5244 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_EAST[4]
  PIN dataOut_EAST[3] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.22 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.214 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 31.68 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 105.072 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 50.4 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 166.848 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 15.9237 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 52.8882 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_EAST[3]
  PIN dataOut_EAST[2] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.26 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.062 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 24.8 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 82.368 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 59.04 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 195.36 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 20.2474 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 67.4305 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_EAST[2]
  PIN dataOut_EAST[1] 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.37 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.74 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.238 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 33.12 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 109.824 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 41.76 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 138.336 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 14.4648 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 48.6868 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_EAST[1]
  PIN dataOut_EAST[0] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.46 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.902 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 11.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 38.016 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 46.24 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 153.12 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 21.4228 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 71.3826 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_EAST[0]
  PIN destinationAddressIn_WEST[13] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.98 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.326 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 38.08 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 126.192 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 1.92 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 8.448 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 LAYER MG ; 
    ANTENNAMAXAREACAR 130.612 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 493.669 LAYER MG ;
    ANTENNAMAXCUTCAR 4.23986 LAYER FY ;
  END destinationAddressIn_WEST[13]
  PIN destinationAddressIn_WEST[12] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.3 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.51 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 40 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 132.528 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 2.56 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 10.56 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 LAYER MG ; 
    ANTENNAMAXAREACAR 71.5053 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 267.544 LAYER MG ;
    ANTENNAMAXCUTCAR 3.52463 LAYER FY ;
  END destinationAddressIn_WEST[12]
  PIN destinationAddressIn_WEST[11] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 25.6 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 85.008 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3744 LAYER MQ ; 
    ANTENNAMAXAREACAR 183.506 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 657.032 LAYER MQ ;
    ANTENNAMAXCUTCAR 1.81624 LAYER VQ ;
  END destinationAddressIn_WEST[11]
  PIN destinationAddressIn_WEST[10] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.768 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 LAYER M3 ; 
    ANTENNAMAXAREACAR 34.6169 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 134.376 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END destinationAddressIn_WEST[10]
  PIN destinationAddressIn_WEST[9] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 32.16 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 106.656 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 4.64 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 15.84 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 LAYER MG ; 
    ANTENNAMAXAREACAR 194.754 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 695.282 LAYER MG ;
    ANTENNAMAXCUTCAR 4.23986 LAYER FY ;
  END destinationAddressIn_WEST[9]
  PIN destinationAddressIn_WEST[8] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.924 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 30.08 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 100.32 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2304 LAYER MQ ; 
    ANTENNAMAXAREACAR 243.995 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 854.568 LAYER MQ ;
    ANTENNAMAXCUTCAR 4.16667 LAYER VQ ;
  END destinationAddressIn_WEST[8]
  PIN destinationAddressIn_WEST[7] 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.37 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.38 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.054 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 134.597 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 503.382 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END destinationAddressIn_WEST[7]
  PIN destinationAddressIn_WEST[6] 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 7.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 27.232 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 159.944 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 597.167 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END destinationAddressIn_WEST[6]
  PIN destinationAddressIn_WEST[5] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 9.54 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 35.446 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.64 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 2.64 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER MQ ; 
    ANTENNAMAXAREACAR 18.9722 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 77.7222 LAYER MQ ;
    ANTENNAMAXCUTCAR 4.16667 LAYER VQ ;
  END destinationAddressIn_WEST[5]
  PIN destinationAddressIn_WEST[4] 
    ANTENNAPARTIALMETALAREA 0.12 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.444 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.78 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.534 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 108.208 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 405.743 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END destinationAddressIn_WEST[4]
  PIN destinationAddressIn_WEST[3] 
    ANTENNAPARTIALMETALAREA 0.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.518 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 7.8 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 29.008 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 148.833 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 556.056 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END destinationAddressIn_WEST[3]
  PIN destinationAddressIn_WEST[2] 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 7.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 29.6 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 143.278 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 535.5 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END destinationAddressIn_WEST[2]
  PIN destinationAddressIn_WEST[1] 
    ANTENNAPARTIALMETALAREA 1.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.07 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 21.4028 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 81.9931 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END destinationAddressIn_WEST[1]
  PIN destinationAddressIn_WEST[0] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.432 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 71.75 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 273.417 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END destinationAddressIn_WEST[0]
  PIN requesterAddressIn_WEST[5] 
    ANTENNAPARTIALMETALAREA 3.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.098 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.46 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.702 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 7.2 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 24.288 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 0.96 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 4.224 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER MG ; 
    ANTENNAMAXAREACAR 61.6806 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 237.41 LAYER MG ;
    ANTENNAMAXCUTCAR 6.94444 LAYER FY ;
  END requesterAddressIn_WEST[5]
  PIN requesterAddressIn_WEST[4] 
    ANTENNAPARTIALMETALAREA 12.32 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 45.88 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 21.0556 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 83.2778 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END requesterAddressIn_WEST[4]
  PIN requesterAddressIn_WEST[3] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.8 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 73.1389 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 278.556 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END requesterAddressIn_WEST[3]
  PIN requesterAddressIn_WEST[2] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 7.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 27.824 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 155.778 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 581.75 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END requesterAddressIn_WEST[2]
  PIN requesterAddressIn_WEST[1] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.544 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 58.5556 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 222.028 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END requesterAddressIn_WEST[1]
  PIN requesterAddressIn_WEST[0] 
    ANTENNAPARTIALMETALAREA 0.9 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.33 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 7.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 26.344 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 128 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 478.972 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END requesterAddressIn_WEST[0]
  PIN dataIn_WEST[31] 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.42 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.102 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 169.319 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 631.854 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_WEST[31]
  PIN dataIn_WEST[30] 
    ANTENNAPARTIALMETALAREA 6.8 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 25.308 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.136 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 61.3333 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 232.306 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_WEST[30]
  PIN dataIn_WEST[29] 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.984 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 190.5 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 710.222 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_WEST[29]
  PIN dataIn_WEST[28] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 17.168 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 132.861 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 499.528 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_WEST[28]
  PIN dataIn_WEST[27] 
    ANTENNAPARTIALMETALAREA 2.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.878 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.584 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 78 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 293.972 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_WEST[27]
  PIN dataIn_WEST[26] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.88 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 53 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 201.472 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_WEST[26]
  PIN dataIn_WEST[25] 
    ANTENNAPARTIALMETALAREA 6.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 25.826 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 123.486 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 459.701 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END dataIn_WEST[25]
  PIN dataIn_WEST[24] 
    ANTENNAPARTIALMETALAREA 6.04 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.496 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 34.9444 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 134.667 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_WEST[24]
  PIN dataIn_WEST[23] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.984 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 100.222 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 376.194 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_WEST[23]
  PIN dataIn_WEST[22] 
    ANTENNAPARTIALMETALAREA 0.12 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.444 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.872 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 110.639 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 417.306 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_WEST[22]
  PIN dataIn_WEST[21] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.912 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 78.6944 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 299.111 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_WEST[21]
  PIN dataIn_WEST[20] 
    ANTENNAPARTIALMETALAREA 4.6 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.168 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 12.7222 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 52.4444 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_WEST[20]
  PIN dataIn_WEST[19] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.584 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 51.6111 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 196.333 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_WEST[19]
  PIN dataIn_WEST[18] 
    ANTENNAPARTIALMETALAREA 0.12 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.444 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.36 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.88 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 46.0556 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 175.778 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_WEST[18]
  PIN dataIn_WEST[17] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.8 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 101.611 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 381.333 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_WEST[17]
  PIN dataIn_WEST[16] 
    ANTENNAPARTIALMETALAREA 0.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.85 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.872 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 100.222 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 376.194 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_WEST[16]
  PIN dataIn_WEST[15] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.392 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 76.6111 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 288.833 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_WEST[15]
  PIN dataIn_WEST[14] 
    ANTENNAPARTIALMETALAREA 0.64 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.516 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2 ; 
    ANTENNAMAXAREACAR 14.1111 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 55.0139 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2 ;
  END dataIn_WEST[14]
  PIN dataIn_WEST[13] 
    ANTENNAPARTIALMETALAREA 0.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.518 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.096 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 79.3889 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 299.111 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_WEST[13]
  PIN dataIn_WEST[12] 
    ANTENNAPARTIALMETALAREA 0.34 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.258 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.584 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 44.6667 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 170.639 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_WEST[12]
  PIN dataIn_WEST[11] 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.22 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.162 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 113.069 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 423.729 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_WEST[11]
  PIN dataIn_WEST[10] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.688 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 79.3889 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 299.111 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_WEST[10]
  PIN dataIn_WEST[9] 
    ANTENNAPARTIALMETALAREA 0.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.518 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.176 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 47.4444 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 180.917 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_WEST[9]
  PIN dataIn_WEST[8] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.68 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 114.806 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 432.722 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_WEST[8]
  PIN dataIn_WEST[7] 
    ANTENNAPARTIALMETALAREA 0.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.258 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.96 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 28 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 108.972 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_WEST[7]
  PIN dataIn_WEST[6] 
    ANTENNAPARTIALMETALAREA 0.12 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.444 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.872 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 83.5556 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 314.528 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_WEST[6]
  PIN dataIn_WEST[5] 
    ANTENNAPARTIALMETALAREA 0.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.518 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.84 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 101.611 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 381.333 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_WEST[5]
  PIN dataIn_WEST[4] 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.064 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 51.6111 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 196.333 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_WEST[4]
  PIN dataIn_WEST[3] 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.37 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.76 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.36 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 57.1667 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 216.889 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_WEST[3]
  PIN dataIn_WEST[2] 
    ANTENNAPARTIALMETALAREA 0.12 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.444 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 24.864 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 121.056 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 453.278 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_WEST[2]
  PIN dataIn_WEST[1] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 18.352 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 94.6667 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 355.639 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_WEST[1]
  PIN dataIn_WEST[0] 
    ANTENNAPARTIALMETALAREA 0.08 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.296 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.64 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.016 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 116.889 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 437.861 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END dataIn_WEST[0]
  PIN destinationAddressOut_WEST[13] 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.37 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.14 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.766 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 125.12 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 413.424 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5588 LAYER MQ ; 
    ANTENNAMAXAREACAR 44.6372 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 154.051 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.519162 LAYER VQ ;
  END destinationAddressOut_WEST[13]
  PIN destinationAddressOut_WEST[12] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.22 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 129.76 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 429.264 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5588 LAYER MQ ; 
    ANTENNAMAXAREACAR 39.6768 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 132.686 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.507922 LAYER VQ ;
  END destinationAddressOut_WEST[12]
  PIN destinationAddressOut_WEST[11] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.66 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.942 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 105.76 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 349.536 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 5.92 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 20.064 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5588 LAYER MG ; 
    ANTENNAMAXAREACAR 11.659 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 41.9377 LAYER MG ;
    ANTENNAMAXCUTCAR 0.552881 LAYER FY ;
  END destinationAddressOut_WEST[11]
  PIN destinationAddressOut_WEST[10] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.9 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.43 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 138.72 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 458.304 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5588 LAYER MQ ; 
    ANTENNAMAXAREACAR 52.2041 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 178.589 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.507922 LAYER VQ ;
  END destinationAddressOut_WEST[10]
  PIN destinationAddressOut_WEST[9] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.3 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.31 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 121.12 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 400.224 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5588 LAYER MQ ; 
    ANTENNAMAXAREACAR 54.9447 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 190.514 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.739403 LAYER VQ ;
  END destinationAddressOut_WEST[9]
  PIN destinationAddressOut_WEST[8] 
    ANTENNAPARTIALMETALAREA 0.08 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.296 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.98 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.326 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 122.08 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 403.392 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5588 LAYER MQ ; 
    ANTENNAMAXAREACAR 38.1233 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 127.79 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.507922 LAYER VQ ;
  END destinationAddressOut_WEST[8]
  PIN destinationAddressOut_WEST[7] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.3 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.51 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 5.12 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 17.424 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 20.48 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 68.64 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5588 LAYER MG ; 
    ANTENNAMAXAREACAR 28.8443 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 98.3889 LAYER MG ;
    ANTENNAMAXCUTCAR 0.552881 LAYER FY ;
  END destinationAddressOut_WEST[7]
  PIN destinationAddressOut_WEST[6] 
    ANTENNAPARTIALMETALAREA 0.12 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.444 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.54 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.798 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 74.72 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 247.104 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.5588 LAYER MQ ; 
    ANTENNAMAXAREACAR 29.4654 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 102.139 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.507922 LAYER VQ ;
  END destinationAddressOut_WEST[6]
  PIN destinationAddressOut_WEST[5] 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.256 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 9.6 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 32.208 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 58.88 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 195.36 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 28.1564 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 93.5232 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END destinationAddressOut_WEST[5]
  PIN destinationAddressOut_WEST[4] 
    ANTENNAPARTIALMETALAREA 0.08 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.296 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.54 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.998 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.8 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 3.168 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 57.44 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 190.08 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 53.7146 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 177.845 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END destinationAddressOut_WEST[4]
  PIN destinationAddressOut_WEST[3] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.38 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.406 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 15.52 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 51.744 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 50.08 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 165.792 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 50.0584 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 165.672 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END destinationAddressOut_WEST[3]
  PIN destinationAddressOut_WEST[2] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.7 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.59 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 7.84 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 26.4 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 52.96 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 175.296 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 53.0448 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 175.43 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END destinationAddressOut_WEST[2]
  PIN destinationAddressOut_WEST[1] 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.37 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.34 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.958 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 6.08 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 20.592 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 46.4 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 154.176 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 15.0554 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 50.5179 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END destinationAddressOut_WEST[1]
  PIN destinationAddressOut_WEST[0] 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.18 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.166 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.48 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 2.112 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 29.28 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 97.152 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 51.1452 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 169.731 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END destinationAddressOut_WEST[0]
  PIN requesterAddressOut_WEST[5] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.962 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 7.1 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 26.27 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 116.96 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 387.024 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 28.64 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 95.04 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 9.98751 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 33.6083 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END requesterAddressOut_WEST[5]
  PIN requesterAddressOut_WEST[4] 
    ANTENNAPARTIALMETALAREA 0.12 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.444 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.78 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.286 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 4.16 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 14.256 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 26.88 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 89.76 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 44.6006 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 148.488 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END requesterAddressOut_WEST[4]
  PIN requesterAddressOut_WEST[3] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.7 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.59 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.8 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 3.168 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 53.92 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 178.464 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 54.0159 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 178.927 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END requesterAddressOut_WEST[3]
  PIN requesterAddressOut_WEST[2] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.54 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.998 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.8 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 3.168 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 40.8 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 135.168 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 50.7908 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 168.817 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END requesterAddressOut_WEST[2]
  PIN requesterAddressOut_WEST[1] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 24.272 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 30.08 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 99.792 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 20.32 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 67.584 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 36.7566 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 122.315 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END requesterAddressOut_WEST[1]
  PIN requesterAddressOut_WEST[0] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.7 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 17.39 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 45.28 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 150.48 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 25.76 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 85.536 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 15.2563 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 51.6284 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END requesterAddressOut_WEST[0]
  PIN dataOut_WEST[31] 
    ANTENNAPARTIALMETALAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.738 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.02 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.774 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 84.64 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 279.84 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 59.04 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 195.36 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 18.5876 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 61.9887 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_WEST[31]
  PIN dataOut_WEST[30] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.82 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.734 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 2.88 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 10.032 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 70.4 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 233.376 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 22.675 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 75.6236 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_WEST[30]
  PIN dataOut_WEST[29] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.54 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.998 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.48 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 2.112 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 58.4 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 193.248 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 25.6638 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 85.5492 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_WEST[29]
  PIN dataOut_WEST[28] 
    ANTENNAPARTIALMETALAREA 7.36 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 27.38 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.66 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.59 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.48 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 2.112 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 37.6 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 124.608 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 12.2557 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 41.0932 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_WEST[28]
  PIN dataOut_WEST[27] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.58 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.294 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 82.4 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 272.448 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 65.44 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 216.48 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 20.9975 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 69.7146 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_WEST[27]
  PIN dataOut_WEST[26] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.54 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.998 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.48 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 2.112 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 63.52 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 210.144 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 47.2232 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 156.41 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_WEST[26]
  PIN dataOut_WEST[25] 
    ANTENNAPARTIALMETALAREA 0.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.518 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.54 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.998 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.48 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 2.112 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 79.68 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 264 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 25.5339 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 85.0483 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_WEST[25]
  PIN dataOut_WEST[24] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.02 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.174 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 27.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 90.816 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 61.6 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 203.808 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 23.3366 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 77.8776 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_WEST[24]
  PIN dataOut_WEST[23] 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.37 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 8.86 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 32.782 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 20.96 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 69.696 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 35.68 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 118.272 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 16.792 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 55.8552 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_WEST[23]
  PIN dataOut_WEST[22] 
    ANTENNAPARTIALMETALAREA 0.08 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.296 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.54 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.998 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.8 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 3.168 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 67.84 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 224.928 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 28.688 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 96.0253 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_WEST[22]
  PIN dataOut_WEST[21] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.78 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 25.086 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 7.52 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 25.344 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 58.56 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 194.304 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 20.0348 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 66.6106 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_WEST[21]
  PIN dataOut_WEST[20] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.02 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.774 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 1.44 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 5.28 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 69.44 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 230.208 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 25.1417 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 83.8361 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_WEST[20]
  PIN dataOut_WEST[19] 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.37 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 5.1 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 18.87 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 22.56 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 74.976 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 56 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 185.856 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 18.7235 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 62.8233 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_WEST[19]
  PIN dataOut_WEST[18] 
    ANTENNAPARTIALMETALAREA 0.08 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.296 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.54 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.998 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.64 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 2.64 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 65.92 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 218.592 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 47.359 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 157.226 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_WEST[18]
  PIN dataOut_WEST[17] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.94 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.726 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 22.24 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 73.92 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 55.2 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 182.688 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 22.297 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 74.258 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_WEST[17]
  PIN dataOut_WEST[16] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.34 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.958 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 6.4 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 21.648 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 52.48 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 174.24 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 18.8003 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 63.1204 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_WEST[16]
  PIN dataOut_WEST[15] 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.37 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.34 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.958 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.48 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 2.112 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 65.28 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 216.48 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 39.1901 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 130.189 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_WEST[15]
  PIN dataOut_WEST[14] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.86 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.182 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 14.08 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 46.992 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 34.4 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 114.048 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 22.1789 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 73.6886 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_WEST[14]
  PIN dataOut_WEST[13] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.74 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.838 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 68.48 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 226.512 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 23.9627 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 80.7057 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END dataOut_WEST[13]
  PIN dataOut_WEST[12] 
    ANTENNAPARTIALMETALAREA 0.12 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.444 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.26 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.062 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 81.76 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 270.336 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 26.7955 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 89.5869 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END dataOut_WEST[12]
  PIN dataOut_WEST[11] 
    ANTENNAPARTIALMETALAREA 3.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.098 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.86 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 25.382 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 18.88 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 62.832 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 36 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 119.328 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 17.7843 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 59.5646 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_WEST[11]
  PIN dataOut_WEST[10] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.54 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.998 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.48 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 2.112 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 54.88 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 181.632 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 30.2509 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 100.449 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_WEST[10]
  PIN dataOut_WEST[9] 
    ANTENNAPARTIALMETALAREA 1.36 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.032 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.7 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.59 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.48 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 2.112 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 44.32 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 146.784 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 28.3218 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 94.0737 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END dataOut_WEST[9]
  PIN dataOut_WEST[8] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.14 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.918 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 88.32 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 291.984 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 26.5734 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 87.978 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END dataOut_WEST[8]
  PIN dataOut_WEST[7] 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.37 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.58 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.246 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 24 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 79.728 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 16.7447 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 59.2102 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END dataOut_WEST[7]
  PIN dataOut_WEST[6] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.18 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.366 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 79.36 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 262.416 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 24.5274 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 81.4782 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END dataOut_WEST[6]
  PIN dataOut_WEST[5] 
    ANTENNAPARTIALMETALAREA 0.9 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.478 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 55.68 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 184.272 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 17.5221 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 58.3996 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END dataOut_WEST[5]
  PIN dataOut_WEST[4] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.7 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.59 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 57.12 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 189.024 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 18.753 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 62.7282 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END dataOut_WEST[4]
  PIN dataOut_WEST[3] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.66 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.142 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 52.48 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 173.712 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 17.7465 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 59.5644 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END dataOut_WEST[3]
  PIN dataOut_WEST[2] 
    ANTENNAPARTIALMETALAREA 0.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.06 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.022 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 16.8 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 55.968 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 8.07374 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 28.0654 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END dataOut_WEST[2]
  PIN dataOut_WEST[1] 
    ANTENNAPARTIALMETALAREA 0.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.46 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.102 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 52.16 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 172.656 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 17.2409 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 57.7193 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END dataOut_WEST[1]
  PIN dataOut_WEST[0] 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 7.82 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 28.934 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 58.88 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 194.832 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 18.6821 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 62.258 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END dataOut_WEST[0]
  PIN cacheDataIn_A[31] 
    ANTENNAPARTIALMETALAREA 1.88 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.956 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.02 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.174 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 56.64 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 187.44 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 34.08 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 112.992 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 10.5309 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 35.1275 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END cacheDataIn_A[31]
  PIN cacheDataIn_A[30] 
    ANTENNAPARTIALMETALAREA 5.78 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 21.386 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.9 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.03 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 49.12 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 162.624 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 40.8 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 135.168 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 12.4919 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 41.5894 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END cacheDataIn_A[30]
  PIN cacheDataIn_A[29] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.18 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.48 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 2.112 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 35.52 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 118.272 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 12.7755 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 43.2669 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END cacheDataIn_A[29]
  PIN cacheDataIn_A[28] 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.86 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.882 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 52.16 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 172.656 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 45.92 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 152.064 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 15.0436 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 50.4258 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END cacheDataIn_A[28]
  PIN cacheDataIn_A[27] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.48 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 54.24 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 179.52 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 43.36 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 143.616 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 13.2303 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 44.0188 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END cacheDataIn_A[27]
  PIN cacheDataIn_A[26] 
    ANTENNAPARTIALMETALAREA 3.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.506 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 14.34 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 53.206 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 21.76 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 72.336 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 8.07374 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 27.3921 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END cacheDataIn_A[26]
  PIN cacheDataIn_A[25] 
    ANTENNAPARTIALMETALAREA 2.56 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.472 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.98 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.726 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 51.52 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 170.544 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 33.76 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 111.936 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 10.8617 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 36.2568 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END cacheDataIn_A[25]
  PIN cacheDataIn_A[24] 
    ANTENNAPARTIALMETALAREA 2.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.878 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 10.06 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 37.222 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 50.08 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 165.792 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 1.12 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 4.224 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 4.48249 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 16.623 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END cacheDataIn_A[24]
  PIN cacheDataIn_A[23] 
    ANTENNAPARTIALMETALAREA 3.32 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.284 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 1.6 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 5.808 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 46.4 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 154.176 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 15.3035 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 51.1842 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END cacheDataIn_A[23]
  PIN cacheDataIn_A[22] 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.46 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.702 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.96 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 3.696 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 41.76 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 138.336 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 27.3531 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 90.9243 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END cacheDataIn_A[22]
  PIN cacheDataIn_A[21] 
    ANTENNAPARTIALMETALAREA 1.92 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.104 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.54 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.998 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 33.6 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 111.408 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 53.28 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 176.352 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 18.186 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 61.183 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END cacheDataIn_A[21]
  PIN cacheDataIn_A[20] 
    ANTENNAPARTIALMETALAREA 7.26 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 27.01 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.46 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.902 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 34.4 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 114.048 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 29.28 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 97.152 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 9.86937 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 33.2468 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END cacheDataIn_A[20]
  PIN cacheDataIn_A[19] 
    ANTENNAPARTIALMETALAREA 4.44 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.576 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.22 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 26.72 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 88.704 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 9.57404 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 32.4009 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END cacheDataIn_A[19]
  PIN cacheDataIn_A[18] 
    ANTENNAPARTIALMETALAREA 17.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 64.01 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 8.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 29.896 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.56282 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 9.46001 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END cacheDataIn_A[18]
  PIN cacheDataIn_A[17] 
    ANTENNAPARTIALMETALAREA 2.8 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.36 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 24.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 90.28 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 7.58349 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 28.0802 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END cacheDataIn_A[17]
  PIN cacheDataIn_A[16] 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.37 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.06 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.322 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 13.76 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 45.936 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 41.76 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 138.336 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 20.2887 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 67.9237 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END cacheDataIn_A[16]
  PIN cacheDataIn_A[15] 
    ANTENNAPARTIALMETALAREA 6.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 25.826 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.848 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 0.814442 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 3.07844 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END cacheDataIn_A[15]
  PIN cacheDataIn_A[14] 
    ANTENNAPARTIALMETALAREA 3.86 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.282 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.22 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 29.76 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 98.736 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 16.1304 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 56.2568 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END cacheDataIn_A[14]
  PIN cacheDataIn_A[13] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.036 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 7.52 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 25.344 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 50.72 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 167.904 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 18.1151 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 61.1286 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END cacheDataIn_A[13]
  PIN cacheDataIn_A[12] 
    ANTENNAPARTIALMETALAREA 5.82 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 21.682 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 11 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 40.848 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 4.67504 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 17.2874 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END cacheDataIn_A[12]
  PIN cacheDataIn_A[11] 
    ANTENNAPARTIALMETALAREA 10.88 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 40.256 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.3 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.11 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 5.12 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 17.424 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 10.6963 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 39.0613 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END cacheDataIn_A[11]
  PIN cacheDataIn_A[10] 
    ANTENNAPARTIALMETALAREA 4.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.466 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 22.54 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 83.398 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 24 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 79.728 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 7.7666 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 25.991 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END cacheDataIn_A[10]
  PIN cacheDataIn_A[9] 
    ANTENNAPARTIALMETALAREA 2.28 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.584 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M2 ; 
    ANTENNAMAXAREACAR 0.826255 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 2.99102 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0118133 LAYER V2 ;
  END cacheDataIn_A[9]
  PIN cacheDataIn_A[8] 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.86 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.282 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.64 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 2.64 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 60 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 198.528 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 19.1369 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 63.5108 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END cacheDataIn_A[8]
  PIN cacheDataIn_A[7] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 1.12 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 4.224 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 63.2 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 209.088 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 19.7217 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 65.4476 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END cacheDataIn_A[7]
  PIN cacheDataIn_A[6] 
    ANTENNAPARTIALMETALAREA 4.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.874 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 30.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 113.368 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 9.22555 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 34.1121 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END cacheDataIn_A[6]
  PIN cacheDataIn_A[5] 
    ANTENNAPARTIALMETALAREA 2.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.658 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M2 ; 
    ANTENNAMAXAREACAR 0.832162 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 3.01288 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0118133 LAYER V2 ;
  END cacheDataIn_A[5]
  PIN cacheDataIn_A[4] 
    ANTENNAPARTIALMETALAREA 3.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.914 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M2 ; 
    ANTENNAMAXAREACAR 1.09206 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 3.97448 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0118133 LAYER V2 ;
  END cacheDataIn_A[4]
  PIN cacheDataIn_A[3] 
    ANTENNAPARTIALMETALAREA 3.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.986 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M2 ; 
    ANTENNAMAXAREACAR 1.25744 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 4.58641 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0118133 LAYER V2 ;
  END cacheDataIn_A[3]
  PIN cacheDataIn_A[2] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.22 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 2.72 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 9.504 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 76.96 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 254.496 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 23.2952 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 77.2332 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END cacheDataIn_A[2]
  PIN cacheDataIn_A[1] 
    ANTENNAPARTIALMETALAREA 3.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.618 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M2 ; 
    ANTENNAMAXAREACAR 1.06843 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 3.88706 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0118133 LAYER V2 ;
  END cacheDataIn_A[1]
  PIN cacheDataIn_A[0] 
    ANTENNAPARTIALMETALAREA 4.7 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.538 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M2 ; 
    ANTENNAMAXAREACAR 1.54096 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 5.63544 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0118133 LAYER V2 ;
  END cacheDataIn_A[0]
  PIN cacheAddressIn_A[7] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.656 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 29.6 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 98.208 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 12.74 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 43.7748 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END cacheAddressIn_A[7]
  PIN cacheAddressIn_A[6] 
    ANTENNAPARTIALMETALAREA 6.98 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 25.826 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 19.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 71.04 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 6.85106 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 25.3702 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END cacheAddressIn_A[6]
  PIN cacheAddressIn_A[5] 
    ANTENNAPARTIALMETALAREA 6.24 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.088 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 24.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 89.392 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 7.91426 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 29.3041 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END cacheAddressIn_A[5]
  PIN cacheAddressIn_A[4] 
    ANTENNAPARTIALMETALAREA 7.66 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 28.342 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 16.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 61.568 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 5.51615 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 20.3874 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END cacheAddressIn_A[4]
  PIN cacheAddressIn_A[3] 
    ANTENNAPARTIALMETALAREA 11.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 42.476 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 16.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 60.088 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 5.39802 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 19.9503 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END cacheAddressIn_A[3]
  PIN cacheAddressIn_A[2] 
    ANTENNAPARTIALMETALAREA 2.74 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.138 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 16.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 62.16 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 5.12631 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 18.9887 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END cacheAddressIn_A[2]
  PIN cacheAddressIn_A[1] 
    ANTENNAPARTIALMETALAREA 10.28 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 38.036 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 20.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 77.552 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 6.4376 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 23.7967 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END cacheAddressIn_A[1]
  PIN cacheAddressIn_A[0] 
    ANTENNAPARTIALMETALAREA 4.78 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.834 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 21.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 79.624 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 7.08733 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 26.2444 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END cacheAddressIn_A[0]
  PIN cacheDataOut_A[31] 
    ANTENNAPARTIALMETALAREA 2.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.102 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1152 LAYER M2 ; 
    ANTENNAMAXAREACAR 22.0937 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 84.1458 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.347222 LAYER V2 ;
  END cacheDataOut_A[31]
  PIN cacheDataOut_A[30] 
    ANTENNAPARTIALMETALAREA 2.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.658 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1152 LAYER M2 ; 
    ANTENNAMAXAREACAR 21.3993 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 80.2917 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.347222 LAYER V2 ;
  END cacheDataOut_A[30]
  PIN cacheDataOut_A[29] 
    ANTENNAPARTIALMETALAREA 4.08 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.244 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1152 LAYER M2 ; 
    ANTENNAMAXAREACAR 36.8507 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 137.462 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.347222 LAYER V2 ;
  END cacheDataOut_A[29]
  PIN cacheDataOut_A[28] 
    ANTENNAPARTIALMETALAREA 3.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.322 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1152 LAYER M2 ; 
    ANTENNAMAXAREACAR 27.6493 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 103.417 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.347222 LAYER V2 ;
  END cacheDataOut_A[28]
  PIN cacheDataOut_A[27] 
    ANTENNAPARTIALMETALAREA 5.66 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 21.09 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 65.2838 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 243.856 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END cacheDataOut_A[27]
  PIN cacheDataOut_A[26] 
    ANTENNAPARTIALMETALAREA 3.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.21 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.664 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1656 LAYER M3 ; 
    ANTENNAMAXAREACAR 8.38164 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 32.1715 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.483092 LAYER VL ;
  END cacheDataOut_A[26]
  PIN cacheDataOut_A[25] 
    ANTENNAPARTIALMETALAREA 4.92 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 18.204 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1152 LAYER M2 ; 
    ANTENNAMAXAREACAR 44.1424 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 163.156 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.347222 LAYER V2 ;
  END cacheDataOut_A[25]
  PIN cacheDataOut_A[24] 
    ANTENNAPARTIALMETALAREA 2.54 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.546 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 30.1486 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 113.856 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END cacheDataOut_A[24]
  PIN cacheDataOut_A[23] 
    ANTENNAPARTIALMETALAREA 4.52 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.724 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 52.4459 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 194.689 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END cacheDataOut_A[23]
  PIN cacheDataOut_A[22] 
    ANTENNAPARTIALMETALAREA 4.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.91 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1152 LAYER M2 ; 
    ANTENNAMAXAREACAR 38.7604 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 143.243 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.347222 LAYER V2 ;
  END cacheDataOut_A[22]
  PIN cacheDataOut_A[21] 
    ANTENNAPARTIALMETALAREA 3.34 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.506 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 39.1577 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 147.189 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END cacheDataOut_A[21]
  PIN cacheDataOut_A[20] 
    ANTENNAPARTIALMETALAREA 2.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.026 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 34.6532 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 130.523 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END cacheDataOut_A[20]
  PIN cacheDataOut_A[19] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 13.12 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 43.824 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER MQ ; 
    ANTENNAMAXAREACAR 160.329 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 542.369 LAYER MQ ;
    ANTENNAMAXCUTCAR 2.7027 LAYER VQ ;
  END cacheDataOut_A[19]
  PIN cacheDataOut_A[18] 
    ANTENNAPARTIALMETALAREA 3.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.578 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1152 LAYER M2 ; 
    ANTENNAMAXAREACAR 35.6354 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 131.681 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.347222 LAYER V2 ;
  END cacheDataOut_A[18]
  PIN cacheDataOut_A[17] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 5.76 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 19.536 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER MQ ; 
    ANTENNAMAXAREACAR 82.8514 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 288.856 LAYER MQ ;
    ANTENNAMAXCUTCAR 2.7027 LAYER VQ ;
  END cacheDataOut_A[17]
  PIN cacheDataOut_A[16] 
    ANTENNAPARTIALMETALAREA 2.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.25 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 29.6982 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 110.523 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END cacheDataOut_A[16]
  PIN cacheDataOut_A[15] 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.184 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 8.48 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 28.512 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1152 LAYER MQ ; 
    ANTENNAMAXAREACAR 78.8646 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 268.052 LAYER MQ ;
    ANTENNAMAXCUTCAR 2.08333 LAYER VQ ;
  END cacheDataOut_A[15]
  PIN cacheDataOut_A[14] 
    ANTENNAPARTIALMETALAREA 2.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.77 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.664 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1152 LAYER M3 ; 
    ANTENNAMAXAREACAR 36.8507 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 138.747 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END cacheDataOut_A[14]
  PIN cacheDataOut_A[13] 
    ANTENNAPARTIALMETALAREA 2.16 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.992 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1608 LAYER M3 ; 
    ANTENNAMAXAREACAR 12.4876 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 49.0647 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.497512 LAYER VL ;
  END cacheDataOut_A[13]
  PIN cacheDataOut_A[12] 
    ANTENNAPARTIALMETALAREA 4.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 47.2658 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 177.189 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END cacheDataOut_A[12]
  PIN cacheDataOut_A[11] 
    ANTENNAPARTIALMETALAREA 2.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.954 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 28.3468 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 107.189 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END cacheDataOut_A[11]
  PIN cacheDataOut_A[10] 
    ANTENNAPARTIALMETALAREA 2.98 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.026 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 35.1036 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 130.523 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END cacheDataOut_A[10]
  PIN cacheDataOut_A[9] 
    ANTENNAPARTIALMETALAREA 2.96 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.952 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 34.8784 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 129.689 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END cacheDataOut_A[9]
  PIN cacheDataOut_A[8] 
    ANTENNAPARTIALMETALAREA 3.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.174 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.664 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 18.6622 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 73.0225 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END cacheDataOut_A[8]
  PIN cacheDataOut_A[7] 
    ANTENNAPARTIALMETALAREA 3.96 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.652 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 46.1396 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 171.356 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END cacheDataOut_A[7]
  PIN cacheDataOut_A[6] 
    ANTENNAPARTIALMETALAREA 2.58 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.546 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.552 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 15.9595 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 63.0225 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END cacheDataOut_A[6]
  PIN cacheDataOut_A[5] 
    ANTENNAPARTIALMETALAREA 3.52 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.024 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 41.1847 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 153.023 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END cacheDataOut_A[5]
  PIN cacheDataOut_A[4] 
    ANTENNAPARTIALMETALAREA 2.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.214 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 9.96 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 37 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0696 LAYER M3 ; 
    ANTENNAMAXAREACAR 151.471 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 562.195 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.14943 LAYER VL ;
  END cacheDataOut_A[4]
  PIN cacheDataOut_A[3] 
    ANTENNAPARTIALMETALAREA 2.52 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.324 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 29.9234 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 111.356 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END cacheDataOut_A[3]
  PIN cacheDataOut_A[2] 
    ANTENNAPARTIALMETALAREA 2.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.77 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.504 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 47.5563 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 181.439 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END cacheDataOut_A[2]
  PIN cacheDataOut_A[1] 
    ANTENNAPARTIALMETALAREA 3.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.914 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 36.9054 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 140.523 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END cacheDataOut_A[1]
  PIN cacheDataOut_A[0] 
    ANTENNAPARTIALMETALAREA 2.54 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.546 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 30.1486 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 113.856 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END cacheDataOut_A[0]
  PIN cacheDataIn_B[31] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.036 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.8 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 3.168 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 27.36 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 90.816 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 17.6898 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 58.7424 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END cacheDataIn_B[31]
  PIN cacheDataIn_B[30] 
    ANTENNAPARTIALMETALAREA 6.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.718 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 11.22 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 41.662 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 14.08 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 46.992 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 5.43937 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 18.5959 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END cacheDataIn_B[30]
  PIN cacheDataIn_B[29] 
    ANTENNAPARTIALMETALAREA 18.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 67.858 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M2 ; 
    ANTENNAMAXAREACAR 5.5575 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 20.4966 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0118133 LAYER V2 ;
  END cacheDataIn_B[29]
  PIN cacheDataIn_B[28] 
    ANTENNAPARTIALMETALAREA 5.64 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 21.016 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.664 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 4.59471 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 16.978 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END cacheDataIn_B[28]
  PIN cacheDataIn_B[27] 
    ANTENNAPARTIALMETALAREA 2.32 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.584 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.22 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.214 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 35.04 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 116.16 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 14.8782 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 50.9999 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END cacheDataIn_B[27]
  PIN cacheDataIn_B[26] 
    ANTENNAPARTIALMETALAREA 2.7 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.99 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 12.22 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 45.214 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 5.44 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 18.48 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 3.76187 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 13.4098 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END cacheDataIn_B[26]
  PIN cacheDataIn_B[25] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.036 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 41.44 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 137.28 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 34.88 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 116.16 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 10.8853 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 36.5002 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END cacheDataIn_B[25]
  PIN cacheDataIn_B[24] 
    ANTENNAPARTIALMETALAREA 2.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.77 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.06 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 22.422 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 2.08 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 7.392 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 24.16 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 80.256 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 19.2492 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 64.0773 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END cacheDataIn_B[24]
  PIN cacheDataIn_B[23] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 4 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 13.728 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 43.36 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 143.616 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 21.73 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 73.4452 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END cacheDataIn_B[23]
  PIN cacheDataIn_B[22] 
    ANTENNAPARTIALMETALAREA 4.86 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.982 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 18.3 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 67.71 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 33.6 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 111.408 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 10.7554 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 35.9591 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END cacheDataIn_B[22]
  PIN cacheDataIn_B[21] 
    ANTENNAPARTIALMETALAREA 8.36 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 30.932 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 17.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 66.008 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 6.42342 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 23.8438 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END cacheDataIn_B[21]
  PIN cacheDataIn_B[20] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.38 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.406 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 3.04 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 10.56 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 42.08 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 139.392 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 19.867 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 66.1734 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END cacheDataIn_B[20]
  PIN cacheDataIn_B[19] 
    ANTENNAPARTIALMETALAREA 16.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 59.57 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M2 ; 
    ANTENNAMAXAREACAR 4.92903 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 18.1835 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0118133 LAYER V2 ;
  END cacheDataIn_B[19]
  PIN cacheDataIn_B[18] 
    ANTENNAPARTIALMETALAREA 4.86 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.982 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 16.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 62.752 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 6.40216 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 23.7093 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END cacheDataIn_B[18]
  PIN cacheDataIn_B[17] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 3.68 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 12.672 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 41.12 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 136.224 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 21.9284 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 72.793 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END cacheDataIn_B[17]
  PIN cacheDataIn_B[16] 
    ANTENNAPARTIALMETALAREA 18.58 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 69.042 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M2 ; 
    ANTENNAMAXAREACAR 5.64019 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 20.8463 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0118133 LAYER V2 ;
  END cacheDataIn_B[16]
  PIN cacheDataIn_B[15] 
    ANTENNAPARTIALMETALAREA 4.46 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.65 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 15.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 57.424 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 4.90186 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 18.1145 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END cacheDataIn_B[15]
  PIN cacheDataIn_B[14] 
    ANTENNAPARTIALMETALAREA 6.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.606 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 22.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 84.656 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 9.46181 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 34.9863 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END cacheDataIn_B[14]
  PIN cacheDataIn_B[13] 
    ANTENNAPARTIALMETALAREA 3.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.876 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 16.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 59.496 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 4.99637 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 18.4641 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END cacheDataIn_B[13]
  PIN cacheDataIn_B[12] 
    ANTENNAPARTIALMETALAREA 9.62 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 35.89 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M2 ; 
    ANTENNAMAXAREACAR 2.994 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 11.0554 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0118133 LAYER V2 ;
  END cacheDataIn_B[12]
  PIN cacheDataIn_B[11] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 4.64 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 15.84 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 46.24 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 153.12 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 17.6898 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 59.6118 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END cacheDataIn_B[11]
  PIN cacheDataIn_B[10] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.18 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.48 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 2.112 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 43.68 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 144.672 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 21.3756 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 70.9432 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END cacheDataIn_B[10]
  PIN cacheDataIn_B[9] 
    ANTENNAPARTIALMETALAREA 3.96 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.652 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 22.92 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 84.952 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 7.02826 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 25.9822 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END cacheDataIn_B[9]
  PIN cacheDataIn_B[8] 
    ANTENNAPARTIALMETALAREA 2.06 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.77 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M2 ; 
    ANTENNAMAXAREACAR 0.761282 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 2.75062 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0118133 LAYER V2 ;
  END cacheDataIn_B[8]
  PIN cacheDataIn_B[7] 
    ANTENNAPARTIALMETALAREA 3.28 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.136 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 27.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 100.64 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 8.2096 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 30.3531 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END cacheDataIn_B[7]
  PIN cacheDataIn_B[6] 
    ANTENNAPARTIALMETALAREA 2.54 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.398 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 25.88 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 95.904 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 7.97333 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 29.4789 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END cacheDataIn_B[6]
  PIN cacheDataIn_B[5] 
    ANTENNAPARTIALMETALAREA 2.52 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.472 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M2 ; 
    ANTENNAMAXAREACAR 0.897135 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 3.25328 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0118133 LAYER V2 ;
  END cacheDataIn_B[5]
  PIN cacheDataIn_B[4] 
    ANTENNAPARTIALMETALAREA 6.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.866 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 25.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 94.128 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 7.68981 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 28.4299 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END cacheDataIn_B[4]
  PIN cacheDataIn_B[3] 
    ANTENNAPARTIALMETALAREA 3.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.618 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M2 ; 
    ANTENNAMAXAREACAR 1.06843 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 3.88706 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0118133 LAYER V2 ;
  END cacheDataIn_B[3]
  PIN cacheDataIn_B[2] 
    ANTENNAPARTIALMETALAREA 2.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.658 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M2 ; 
    ANTENNAMAXAREACAR 0.832162 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 3.01288 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0118133 LAYER V2 ;
  END cacheDataIn_B[2]
  PIN cacheDataIn_B[1] 
    ANTENNAPARTIALMETALAREA 6.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 23.458 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M2 ; 
    ANTENNAMAXAREACAR 2.0135 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 7.38382 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0118133 LAYER V2 ;
  END cacheDataIn_B[1]
  PIN cacheDataIn_B[0] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 1.44 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 5.28 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 49.44 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 163.68 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 15.5457 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 51.6597 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END cacheDataIn_B[0]
  PIN cacheAddressIn_B[7] 
    ANTENNAPARTIALMETALAREA 4.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.576 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 10.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 37.592 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.30706 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 12.2574 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END cacheAddressIn_B[7]
  PIN cacheAddressIn_B[6] 
    ANTENNAPARTIALMETALAREA 7.26 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 26.862 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 10.08 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 37.592 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.63783 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 13.4813 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END cacheAddressIn_B[6]
  PIN cacheAddressIn_B[5] 
    ANTENNAPARTIALMETALAREA 12.7 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 47.138 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M2 ; 
    ANTENNAMAXAREACAR 3.90363 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 14.3773 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0118133 LAYER V2 ;
  END cacheAddressIn_B[5]
  PIN cacheAddressIn_B[4] 
    ANTENNAPARTIALMETALAREA 2.14 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.066 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M2 ; 
    ANTENNAMAXAREACAR 0.784908 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 2.83804 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0118133 LAYER V2 ;
  END cacheAddressIn_B[4]
  PIN cacheAddressIn_B[3] 
    ANTENNAPARTIALMETALAREA 3.4 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.728 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M2 ; 
    ANTENNAMAXAREACAR 1.15703 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 4.21488 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0118133 LAYER V2 ;
  END cacheAddressIn_B[3]
  PIN cacheAddressIn_B[2] 
    ANTENNAPARTIALMETALAREA 6.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 24.198 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M2 ; 
    ANTENNAMAXAREACAR 2.07256 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 7.60236 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0118133 LAYER V2 ;
  END cacheAddressIn_B[2]
  PIN cacheAddressIn_B[1] 
    ANTENNAPARTIALMETALAREA 5.64 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 20.868 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 10 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 37.296 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.14167 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 11.6455 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END cacheAddressIn_B[1]
  PIN cacheAddressIn_B[0] 
    ANTENNAPARTIALMETALAREA 3.7 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.69 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 8.44 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 31.376 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 4.52383 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 16.7158 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END cacheAddressIn_B[0]
  PIN cacheDataOut_B[31] 
    ANTENNAPARTIALMETALAREA 2.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.176 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 3 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.248 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1152 LAYER M3 ; 
    ANTENNAMAXAREACAR 31.9896 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 120.76 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END cacheDataOut_B[31]
  PIN cacheDataOut_B[30] 
    ANTENNAPARTIALMETALAREA 4.7 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.39 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1152 LAYER M2 ; 
    ANTENNAMAXAREACAR 42.2326 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 156.09 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.347222 LAYER V2 ;
  END cacheDataOut_B[30]
  PIN cacheDataOut_B[29] 
    ANTENNAPARTIALMETALAREA 3.98 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.874 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1152 LAYER M2 ; 
    ANTENNAMAXAREACAR 35.9826 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 134.25 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.347222 LAYER V2 ;
  END cacheDataOut_B[29]
  PIN cacheDataOut_B[28] 
    ANTENNAPARTIALMETALAREA 4.7 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.39 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1152 LAYER M2 ; 
    ANTENNAMAXAREACAR 42.2326 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 156.09 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.347222 LAYER V2 ;
  END cacheDataOut_B[28]
  PIN cacheDataOut_B[27] 
    ANTENNAPARTIALMETALAREA 4.04 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.096 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 47.0405 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 176.356 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END cacheDataOut_B[27]
  PIN cacheDataOut_B[26] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.72 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.212 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1152 LAYER M3 ; 
    ANTENNAMAXAREACAR 62.8924 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 235.049 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END cacheDataOut_B[26]
  PIN cacheDataOut_B[25] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.16 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.592 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 8.32 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 27.984 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1152 LAYER MQ ; 
    ANTENNAMAXAREACAR 78.691 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 267.965 LAYER MQ ;
    ANTENNAMAXCUTCAR 2.08333 LAYER VQ ;
  END cacheDataOut_B[25]
  PIN cacheDataOut_B[24] 
    ANTENNAPARTIALMETALAREA 3.22 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.914 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.84 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.256 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 18.6622 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 73.0225 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END cacheDataOut_B[24]
  PIN cacheDataOut_B[23] 
    ANTENNAPARTIALMETALAREA 3.88 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.356 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 45.2387 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 168.023 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END cacheDataOut_B[23]
  PIN cacheDataOut_B[22] 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.26 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.962 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 8 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 26.928 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1152 LAYER MQ ; 
    ANTENNAMAXAREACAR 75.8958 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 258.656 LAYER MQ ;
    ANTENNAMAXCUTCAR 2.08333 LAYER VQ ;
  END cacheDataOut_B[22]
  PIN cacheDataOut_B[21] 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.4 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.18 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 7.68 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 25.872 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER MQ ; 
    ANTENNAMAXAREACAR 94.5631 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 323.541 LAYER MQ ;
    ANTENNAMAXCUTCAR 2.7027 LAYER VQ ;
  END cacheDataOut_B[21]
  PIN cacheDataOut_B[20] 
    ANTENNAPARTIALMETALAREA 4.72 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.464 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.3 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.258 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1584 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.82071 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 15.8434 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.505051 LAYER VL ;
  END cacheDataOut_B[20]
  PIN cacheDataOut_B[19] 
    ANTENNAPARTIALMETALAREA 3.76 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.912 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 15.0586 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 59.6892 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END cacheDataOut_B[19]
  PIN cacheDataOut_B[18] 
    ANTENNAPARTIALMETALAREA 3.9 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.578 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1152 LAYER M2 ; 
    ANTENNAMAXAREACAR 35.2882 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 131.681 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.347222 LAYER V2 ;
  END cacheDataOut_B[18]
  PIN cacheDataOut_B[17] 
    ANTENNAPARTIALMETALAREA 2.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.026 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 34.6532 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 130.523 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END cacheDataOut_B[17]
  PIN cacheDataOut_B[16] 
    ANTENNAPARTIALMETALAREA 5.38 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 19.906 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 62.1306 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 230.523 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END cacheDataOut_B[16]
  PIN cacheDataOut_B[15] 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.48 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.776 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 7.84 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 26.4 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER MQ ; 
    ANTENNAMAXAREACAR 104.473 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 359.486 LAYER MQ ;
    ANTENNAMAXCUTCAR 2.7027 LAYER VQ ;
  END cacheDataOut_B[15]
  PIN cacheDataOut_B[14] 
    ANTENNAPARTIALMETALAREA 4.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.798 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.184 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1152 LAYER M3 ; 
    ANTENNAMAXAREACAR 4.90625 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 20.5521 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END cacheDataOut_B[14]
  PIN cacheDataOut_B[13] 
    ANTENNAPARTIALMETALAREA 4.48 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.576 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 51.9955 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 193.023 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END cacheDataOut_B[13]
  PIN cacheDataOut_B[12] 
    ANTENNAPARTIALMETALAREA 2.98 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.026 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.184 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 6.04955 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 26.3559 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END cacheDataOut_B[12]
  PIN cacheDataOut_B[11] 
    ANTENNAPARTIALMETALAREA 3.02 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.322 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1152 LAYER M2 ; 
    ANTENNAMAXAREACAR 27.6493 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 103.417 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.347222 LAYER V2 ;
  END cacheDataOut_B[11]
  PIN cacheDataOut_B[10] 
    ANTENNAPARTIALMETALAREA 2.998 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.0926 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1152 LAYER M2 ; 
    ANTENNAMAXAREACAR 27.6319 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 102.016 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.347222 LAYER V2 ;
  END cacheDataOut_B[10]
  PIN cacheDataOut_B[9] 
    ANTENNAPARTIALMETALAREA 5.08 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 18.796 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.68 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.664 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1152 LAYER M3 ; 
    ANTENNAMAXAREACAR 10.4618 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 41.1076 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.694444 LAYER VL ;
  END cacheDataOut_B[9]
  PIN cacheDataOut_B[8] 
    ANTENNAPARTIALMETALAREA 4.58 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.946 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 53.1216 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 197.189 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END cacheDataOut_B[8]
  PIN cacheDataOut_B[7] 
    ANTENNAPARTIALMETALAREA 4.52 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.724 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 52.4459 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 194.689 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END cacheDataOut_B[7]
  PIN cacheDataOut_B[6] 
    ANTENNAPARTIALMETALAREA 3.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.618 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1584 LAYER M2 ; 
    ANTENNAMAXAREACAR 20.6136 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 77.0808 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.252525 LAYER V2 ;
  END cacheDataOut_B[6]
  PIN cacheDataOut_B[5] 
    ANTENNAPARTIALMETALAREA 2.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.026 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.6 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.368 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 9.65315 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 39.6892 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END cacheDataOut_B[5]
  PIN cacheDataOut_B[4] 
    ANTENNAPARTIALMETALAREA 4.42 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.354 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.2 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M3 ; 
    ANTENNAMAXAREACAR 6.04955 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 26.3559 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.900901 LAYER VL ;
  END cacheDataOut_B[4]
  PIN cacheDataOut_B[3] 
    ANTENNAPARTIALMETALAREA 2.46 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.25 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 29.2477 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 110.523 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END cacheDataOut_B[3]
  PIN cacheDataOut_B[2] 
    ANTENNAPARTIALMETALAREA 3.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.766 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 37.3559 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 138.856 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END cacheDataOut_B[2]
  PIN cacheDataOut_B[1] 
    ANTENNAPARTIALMETALAREA 2.44 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.028 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 29.0225 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 108.023 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END cacheDataOut_B[1]
  PIN cacheDataOut_B[0] 
    ANTENNAPARTIALMETALAREA 2.98 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.026 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 LAYER M2 ; 
    ANTENNAMAXAREACAR 35.1036 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 130.523 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.45045 LAYER V2 ;
  END cacheDataOut_B[0]
  PIN clk 
    ANTENNAPARTIALMETALAREA 14.52 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 53.576 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 115.84 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 383.328 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.7016 LAYER MQ ; 
    ANTENNAMAXAREACAR 68.6648 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 227.718 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.141044 LAYER VQ ;
  END clk
  PIN reset 
    ANTENNAPARTIALMETALAREA 120.32 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 398.64 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 7.116 LAYER MQ ; 
    ANTENNAMAXAREACAR 62.2748 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 223.97 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.48 LAYER VQ ;
    ANTENNAMAXCUTCAR 6.38929 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 291.2 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 964.128 LAYER MG ;
    ANTENNAGATEAREA 8.988 LAYER MG ; 
    ANTENNAMAXAREACAR 104.988 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 365.202 LAYER MG ;
    ANTENNAMAXCUTCAR 6.38929 LAYER FY ;
  END reset
  PIN readIn_NORTH 
    ANTENNAPARTIALMETALAREA 8.62 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 31.894 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.22 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.014 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M3 ; 
    ANTENNAMAXAREACAR 115.847 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 431.438 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAMAXCUTCAR 4.16667 LAYER VL ;
    ANTENNAPARTIALMETALAREA 29.76 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 98.736 LAYER MQ ;
    ANTENNAGATEAREA 0.3624 LAYER MQ ; 
    ANTENNAMAXAREACAR 197.966 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 703.888 LAYER MQ ;
    ANTENNAMAXCUTCAR 4.16667 LAYER VQ ;
  END readIn_NORTH
  PIN writeIn_NORTH 
    ANTENNAPARTIALMETALAREA 8.92 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 33.004 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 6.94 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 25.678 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 66.08 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 219.648 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 2.24 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 9.504 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3624 LAYER MG ; 
    ANTENNAMAXAREACAR 22.3755 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 94.7807 LAYER MG ;
    ANTENNAMAXCUTCAR 6.94444 LAYER FY ;
  END writeIn_NORTH
  PIN readIn_SOUTH 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.46 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.85 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 0.8 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 3.168 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 5.28 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 23.232 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3624 LAYER MG ; 
    ANTENNAMAXAREACAR 221.927 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 809.419 LAYER MG ;
    ANTENNAMAXCUTCAR 7.53968 LAYER FY ;
  END readIn_SOUTH
  PIN writeIn_SOUTH 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.56 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 53.28 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 177.408 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3624 LAYER MQ ; 
    ANTENNAMAXAREACAR 282.034 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 990.435 LAYER MQ ;
    ANTENNAMAXCUTCAR 3.6075 LAYER VQ ;
  END writeIn_SOUTH
  PIN readIn_EAST 
    ANTENNAPARTIALMETALAREA 0.12 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.444 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 7.58 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 28.046 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 33.6 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 113.52 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 4.96 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 21.12 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3624 LAYER MG ; 
    ANTENNAMAXAREACAR 144.495 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 543.863 LAYER MG ;
    ANTENNAMAXCUTCAR 6.94444 LAYER FY ;
  END readIn_EAST
  PIN writeIn_EAST 
    ANTENNAPARTIALMETALAREA 8.5 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 31.598 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 23.82 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 88.134 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 36.96 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 124.608 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3624 LAYER MQ ; 
    ANTENNAMAXAREACAR 134.658 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 465.408 LAYER MQ ;
    ANTENNAMAXCUTCAR 2.52483 LAYER VQ ;
  END writeIn_EAST
  PIN readIn_WEST 
    ANTENNAPARTIALMETALAREA 20.08 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 74.444 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 2.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.992 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3624 LAYER M3 ; 
    ANTENNAMAXAREACAR 45.9921 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 172.905 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL ;
  END readIn_WEST
  PIN writeIn_WEST 
    ANTENNAPARTIALMETALAREA 17.94 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 66.526 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.24 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.736 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3624 LAYER M3 ; 
    ANTENNAMAXAREACAR 43.1667 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 162.876 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.94246 LAYER VL ;
  END writeIn_WEST
  PIN portA_writtenTo 
  END portA_writtenTo
  PIN portB_writtenTo 
  END portB_writtenTo
  PIN readOut_NORTH 
    ANTENNAPARTIALMETALAREA 6.66 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 24.79 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.184 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 0.341908 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 1.24265 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END readOut_NORTH
  PIN writeOut_NORTH 
    ANTENNAPARTIALMETALAREA 2.88 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.656 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 12.12 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 44.992 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M3 ; 
    ANTENNAMAXAREACAR 5.32714 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 19.688 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0236267 LAYER VL ;
  END writeOut_NORTH
  PIN readOut_SOUTH 
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.26 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.962 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 2.08 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 7.392 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 35.04 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 116.16 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 16.0123 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 53.587 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END readOut_SOUTH
  PIN writeOut_SOUTH 
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.04 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.848 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 72.64 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 240.24 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 17.76 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 59.136 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 8.61716 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 29.5587 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END writeOut_SOUTH
  PIN readOut_EAST 
    ANTENNAPARTIALMETALAREA 0.2 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.74 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 4.7 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 17.39 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 40.16 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 133.584 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 13.4724 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 45.3933 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END readOut_EAST
  PIN writeOut_EAST 
    ANTENNAPARTIALMETALAREA 47.82 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 177.23 LAYER M2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER M2 ; 
    ANTENNAMAXAREACAR 14.2758 LAYER M2 ;
    ANTENNAMAXSIDEAREACAR 52.7979 LAYER M2 ;
    ANTENNAMAXCUTCAR 0.0118133 LAYER V2 ;
  END writeOut_EAST
  PIN readOut_WEST 
    ANTENNAPARTIALMETALAREA 4.04 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.096 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.22 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.814 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 77.76 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 257.664 LAYER MQ ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VQ ;
    ANTENNAPARTIALMETALAREA 4.32 LAYER MG ;
    ANTENNAPARTIALMETALSIDEAREA 14.784 LAYER MG ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MG ; 
    ANTENNAMAXAREACAR 14.4057 LAYER MG ;
    ANTENNAMAXSIDEAREACAR 48.0087 LAYER MG ;
    ANTENNAMAXCUTCAR 0.118133 LAYER FY ;
  END readOut_WEST
  PIN writeOut_WEST 
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.37 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.5 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.55 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 75.84 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 250.8 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 25.3094 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 84.8191 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END writeOut_WEST
  PIN memWrite_A 
    ANTENNAPARTIALMETALAREA 2.3 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.51 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 1.1 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.07 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 47.68 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 157.872 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 19.2492 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 65.6791 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END memWrite_A
  PIN memWrite_B 
    ANTENNAPARTIALMETALAREA 2.1 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.77 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2 ;
    ANTENNAPARTIALMETALAREA 0.78 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.886 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER VL ;
    ANTENNAPARTIALMETALAREA 46.88 LAYER MQ ;
    ANTENNAPARTIALMETALSIDEAREA 155.232 LAYER MQ ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.386 LAYER MQ ; 
    ANTENNAMAXAREACAR 14.9078 LAYER MQ ;
    ANTENNAMAXSIDEAREACAR 49.7105 LAYER MQ ;
    ANTENNAMAXCUTCAR 0.0708801 LAYER VQ ;
  END memWrite_B
END router

END LIBRARY
