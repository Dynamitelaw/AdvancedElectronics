##
## LEF for PtnCells ;
## created by Encounter v14.23-s044_1 on Tue May 14 23:25:14 2019
##

VERSION 5.5 ;

NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO cacheBank
  CLASS BLOCK ;
  SIZE 796.5000 BY 716.0000 ;
  FOREIGN cacheBank 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.28 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.584 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.7016 LAYER M3  ;
    ANTENNAMAXAREACAR 9.73625 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 36.3655 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0470146 LAYER VL  ;
    PORT
      LAYER M3 ;
        RECT 334.9000 0.0000 335.1000 0.6000 ;
    END
  END clk
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.32 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 2.14 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.178 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.078 LAYER M3  ;
    ANTENNAMAXAREACAR 159.385 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 559.415 LAYER M3  ;
    ANTENNAMAXCUTCAR 2.05128 LAYER VL  ;
    ANTENNADIFFAREA 0.32 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.72 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 3.168 LAYER MQ  ;
    ANTENNAGATEAREA 0.078 LAYER MQ  ;
    ANTENNAMAXAREACAR 168.615 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 600.031 LAYER MQ  ;
    ANTENNAMAXCUTCAR 2.05128 LAYER VQ  ;
    PORT
      LAYER M3 ;
        RECT 342.9000 0.0000 343.1000 0.6000 ;
    END
  END reset
  PIN cacheDataIn_A[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL  ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ  ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2  ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 18.4615 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 43.6923 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.72 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.368 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 40.6667 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 118.262 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 49.8974 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 158.877 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 758.9000 0.0000 759.1000 0.6000 ;
    END
  END cacheDataIn_A[31]
  PIN cacheDataIn_A[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.706 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.8202 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 129.897 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 452.21 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 139.128 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 474.979 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 148.359 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 515.595 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 733.9000 0.0000 734.1000 0.6000 ;
    END
  END cacheDataIn_A[30]
  PIN cacheDataIn_A[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL  ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ  ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2  ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 18.4615 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 43.6923 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.64 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 38.6154 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 110.672 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 47.8462 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 151.287 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 720.9000 0.0000 721.1000 0.6000 ;
    END
  END cacheDataIn_A[29]
  PIN cacheDataIn_A[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.566 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.3022 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 126.308 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 438.928 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 135.538 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 461.697 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 144.769 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 502.313 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 695.9000 0.0000 696.1000 0.6000 ;
    END
  END cacheDataIn_A[28]
  PIN cacheDataIn_A[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL  ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ  ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 3.06 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.322 LAYER M2  ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 18.4615 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 43.6923 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.76 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.516 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 68.359 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 220.723 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 77.5897 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 261.338 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 681.9000 0.0000 682.1000 0.6000 ;
    END
  END cacheDataIn_A[27]
  PIN cacheDataIn_A[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.746 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.9682 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 130.923 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 456.005 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 140.154 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 478.774 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 149.385 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 519.39 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 656.9000 0.0000 657.1000 0.6000 ;
    END
  END cacheDataIn_A[26]
  PIN cacheDataIn_A[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL  ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ  ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2  ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 18.4615 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 43.6923 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.68 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.22 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 39.641 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 114.467 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 48.8718 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 155.082 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 643.9000 0.0000 644.1000 0.6000 ;
    END
  END cacheDataIn_A[25]
  PIN cacheDataIn_A[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.626 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5242 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 127.846 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 444.621 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 137.077 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 467.39 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 146.308 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 508.005 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 618.9000 0.0000 619.1000 0.6000 ;
    END
  END cacheDataIn_A[24]
  PIN cacheDataIn_A[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.806 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.1902 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 132.462 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 461.697 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 141.692 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 484.467 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 150.923 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 525.082 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 605.9000 0.0000 606.1000 0.6000 ;
    END
  END cacheDataIn_A[23]
  PIN cacheDataIn_A[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.786 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.1162 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 131.949 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 459.8 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 141.179 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 482.569 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 150.41 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 523.185 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 579.9000 0.0000 580.1000 0.6000 ;
    END
  END cacheDataIn_A[22]
  PIN cacheDataIn_A[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL  ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ  ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2  ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 18.4615 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 43.6923 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.72 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.368 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 40.6667 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 118.262 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 49.8974 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 158.877 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 566.9000 0.0000 567.1000 0.6000 ;
    END
  END cacheDataIn_A[21]
  PIN cacheDataIn_A[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.706 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.8202 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 129.897 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 452.21 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 139.128 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 474.979 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 148.359 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 515.595 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 541.9000 0.0000 542.1000 0.6000 ;
    END
  END cacheDataIn_A[20]
  PIN cacheDataIn_A[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL  ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ  ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2  ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 18.4615 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 43.6923 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.64 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 38.6154 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 110.672 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 47.8462 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 151.287 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 528.9000 0.0000 529.1000 0.6000 ;
    END
  END cacheDataIn_A[19]
  PIN cacheDataIn_A[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL  ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ  ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.18 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.666 LAYER M2  ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 18.4615 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 43.6923 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.64 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 139.128 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 482.569 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 148.359 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 523.185 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 502.9000 0.0000 503.1000 0.6000 ;
    END
  END cacheDataIn_A[18]
  PIN cacheDataIn_A[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL  ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ  ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 3.06 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.322 LAYER M2  ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 18.4615 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 43.6923 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.76 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.516 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 68.359 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 220.723 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 77.5897 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 261.338 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 489.9000 0.0000 490.1000 0.6000 ;
    END
  END cacheDataIn_A[17]
  PIN cacheDataIn_A[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.746 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.9682 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 130.923 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 456.005 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 140.154 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 478.774 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 149.385 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 519.39 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 464.9000 0.0000 465.1000 0.6000 ;
    END
  END cacheDataIn_A[16]
  PIN cacheDataIn_A[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL  ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ  ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2  ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 18.4615 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 43.6923 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.68 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.22 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 39.641 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 114.467 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 48.8718 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 155.082 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 325.9000 0.0000 326.1000 0.6000 ;
    END
  END cacheDataIn_A[15]
  PIN cacheDataIn_A[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.61 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.465 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 127.436 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 443.103 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 136.667 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 465.872 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 145.897 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 506.487 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 300.9000 0.0000 301.1000 0.6000 ;
    END
  END cacheDataIn_A[14]
  PIN cacheDataIn_A[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.806 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.1902 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 132.462 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 461.697 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 141.692 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 484.467 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 150.923 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 525.082 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 287.9000 0.0000 288.1000 0.6000 ;
    END
  END cacheDataIn_A[13]
  PIN cacheDataIn_A[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.77 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.057 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 131.538 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 458.282 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 140.769 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 481.051 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 150 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 521.667 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 261.9000 0.0000 262.1000 0.6000 ;
    END
  END cacheDataIn_A[12]
  PIN cacheDataIn_A[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL  ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ  ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2  ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 18.4615 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 43.6923 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.72 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.368 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 40.6667 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 118.262 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 49.8974 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 158.877 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 248.9000 0.0000 249.1000 0.6000 ;
    END
  END cacheDataIn_A[11]
  PIN cacheDataIn_A[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.69 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.761 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 129.487 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 450.692 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 138.718 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 473.462 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 147.949 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 514.077 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 223.9000 0.0000 224.1000 0.6000 ;
    END
  END cacheDataIn_A[10]
  PIN cacheDataIn_A[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL  ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ  ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2  ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 18.4615 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 43.6923 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.64 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 38.6154 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 110.672 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 47.8462 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 151.287 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 210.9000 0.0000 211.1000 0.6000 ;
    END
  END cacheDataIn_A[9]
  PIN cacheDataIn_A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.566 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.3022 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 126.308 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 438.928 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 135.538 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 461.697 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 144.769 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 502.313 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 185.9000 0.0000 186.1000 0.6000 ;
    END
  END cacheDataIn_A[8]
  PIN cacheDataIn_A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 127.333 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 446.518 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 136.564 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 469.287 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 145.795 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 509.903 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 171.9000 0.0000 172.1000 0.6000 ;
    END
  END cacheDataIn_A[7]
  PIN cacheDataIn_A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.73 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.909 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 130.513 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 454.487 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 139.744 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 477.256 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 148.974 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 517.872 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 146.9000 0.0000 147.1000 0.6000 ;
    END
  END cacheDataIn_A[6]
  PIN cacheDataIn_A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL  ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ  ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2  ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 18.4615 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 43.6923 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.68 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.22 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 39.641 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 114.467 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 48.8718 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 155.082 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 133.9000 0.0000 134.1000 0.6000 ;
    END
  END cacheDataIn_A[5]
  PIN cacheDataIn_A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 127.333 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 446.518 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 136.564 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 469.287 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 145.795 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 509.903 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 107.9000 0.0000 108.1000 0.6000 ;
    END
  END cacheDataIn_A[4]
  PIN cacheDataIn_A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 127.333 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 446.518 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 136.564 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 469.287 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 145.795 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 509.903 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 94.9000 0.0000 95.1000 0.6000 ;
    END
  END cacheDataIn_A[3]
  PIN cacheDataIn_A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.77 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.057 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 131.538 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 458.282 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 140.769 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 481.051 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 150 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 521.667 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 69.9000 0.0000 70.1000 0.6000 ;
    END
  END cacheDataIn_A[2]
  PIN cacheDataIn_A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL  ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ  ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2  ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 18.4615 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 43.6923 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.72 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.368 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 40.6667 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 118.262 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 49.8974 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 158.877 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 56.9000 0.0000 57.1000 0.6000 ;
    END
  END cacheDataIn_A[1]
  PIN cacheDataIn_A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.69 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.761 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 129.487 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 450.692 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 138.718 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 473.462 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 147.949 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 514.077 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 31.9000 0.0000 32.1000 0.6000 ;
    END
  END cacheDataIn_A[0]
  PIN cacheAddressIn_A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 127.333 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 446.518 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 136.564 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 469.287 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 145.795 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 509.903 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 409.9000 0.0000 410.1000 0.6000 ;
    END
  END cacheAddressIn_A[7]
  PIN cacheAddressIn_A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL  ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ  ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2  ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 18.4615 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 43.6923 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.72 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.368 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 40.6667 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 118.262 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 49.8974 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 158.877 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 412.9000 0.0000 413.1000 0.6000 ;
    END
  END cacheAddressIn_A[6]
  PIN cacheAddressIn_A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL  ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ  ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2  ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 18.4615 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 43.6923 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.4 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.884 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 58.1026 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 182.774 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 67.3333 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 223.39 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 415.9000 0.0000 416.1000 0.6000 ;
    END
  END cacheAddressIn_A[5]
  PIN cacheAddressIn_A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 127.333 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 446.518 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 136.564 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 469.287 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 145.795 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 509.903 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 418.9000 0.0000 419.1000 0.6000 ;
    END
  END cacheAddressIn_A[4]
  PIN cacheAddressIn_A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL  ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ  ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2  ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 18.4615 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 43.6923 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 1.48 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.18 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 60.1538 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 190.364 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 69.3846 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 230.979 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 421.9000 0.0000 422.1000 0.6000 ;
    END
  END cacheAddressIn_A[3]
  PIN cacheAddressIn_A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 127.333 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 446.518 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 136.564 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 469.287 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 145.795 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 509.903 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 424.9000 0.0000 425.1000 0.6000 ;
    END
  END cacheAddressIn_A[2]
  PIN cacheAddressIn_A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL  ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ  ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2  ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 18.4615 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 43.6923 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 2.12 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.548 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 76.5641 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 251.082 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 85.7949 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 291.697 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 427.9000 0.0000 428.1000 0.6000 ;
    END
  END cacheAddressIn_A[1]
  PIN cacheAddressIn_A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL  ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ  ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 3.06 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.322 LAYER M2  ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 18.4615 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 43.6923 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 2.8 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.064 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 120.667 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 414.262 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 129.897 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 454.877 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 430.9000 0.0000 431.1000 0.6000 ;
    END
  END cacheAddressIn_A[0]
  PIN memWrite_A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 127.333 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 446.518 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 136.564 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 469.287 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 145.795 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 509.903 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 433.9000 0.0000 434.1000 0.6000 ;
    END
  END memWrite_A
  PIN cacheDataOut_A[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 756.9000 0.0000 757.1000 0.6000 ;
    END
  END cacheDataOut_A[31]
  PIN cacheDataOut_A[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.726 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.8942 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 735.9000 0.0000 736.1000 0.6000 ;
    END
  END cacheDataOut_A[30]
  PIN cacheDataOut_A[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.37 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.64 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 718.9000 0.0000 719.1000 0.6000 ;
    END
  END cacheDataOut_A[29]
  PIN cacheDataOut_A[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.4502 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 697.9000 0.0000 698.1000 0.6000 ;
    END
  END cacheDataOut_A[28]
  PIN cacheDataOut_A[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.85 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.701 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 679.9000 0.0000 680.1000 0.6000 ;
    END
  END cacheDataOut_A[27]
  PIN cacheDataOut_A[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.766 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.0422 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 658.9000 0.0000 659.1000 0.6000 ;
    END
  END cacheDataOut_A[26]
  PIN cacheDataOut_A[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 641.9000 0.0000 642.1000 0.6000 ;
    END
  END cacheDataOut_A[25]
  PIN cacheDataOut_A[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.646 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 620.9000 0.0000 621.1000 0.6000 ;
    END
  END cacheDataOut_A[24]
  PIN cacheDataOut_A[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.79 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.131 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 603.9000 0.0000 604.1000 0.6000 ;
    END
  END cacheDataOut_A[23]
  PIN cacheDataOut_A[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.806 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.1902 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 581.9000 0.0000 582.1000 0.6000 ;
    END
  END cacheDataOut_A[22]
  PIN cacheDataOut_A[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 564.9000 0.0000 565.1000 0.6000 ;
    END
  END cacheDataOut_A[21]
  PIN cacheDataOut_A[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.726 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.8942 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 543.9000 0.0000 544.1000 0.6000 ;
    END
  END cacheDataOut_A[20]
  PIN cacheDataOut_A[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.37 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.64 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 526.9000 0.0000 527.1000 0.6000 ;
    END
  END cacheDataOut_A[19]
  PIN cacheDataOut_A[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.64 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 504.9000 0.0000 505.1000 0.6000 ;
    END
  END cacheDataOut_A[18]
  PIN cacheDataOut_A[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.85 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.701 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 487.9000 0.0000 488.1000 0.6000 ;
    END
  END cacheDataOut_A[17]
  PIN cacheDataOut_A[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.766 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.0422 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 466.9000 0.0000 467.1000 0.6000 ;
    END
  END cacheDataOut_A[16]
  PIN cacheDataOut_A[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 323.9000 0.0000 324.1000 0.6000 ;
    END
  END cacheDataOut_A[15]
  PIN cacheDataOut_A[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.646 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 302.9000 0.0000 303.1000 0.6000 ;
    END
  END cacheDataOut_A[14]
  PIN cacheDataOut_A[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.774 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.0718 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 285.9000 0.0000 286.1000 0.6000 ;
    END
  END cacheDataOut_A[13]
  PIN cacheDataOut_A[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.806 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.1902 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 263.9000 0.0000 264.1000 0.6000 ;
    END
  END cacheDataOut_A[12]
  PIN cacheDataOut_A[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 246.9000 0.0000 247.1000 0.6000 ;
    END
  END cacheDataOut_A[11]
  PIN cacheDataOut_A[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.726 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.8942 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 225.9000 0.0000 226.1000 0.6000 ;
    END
  END cacheDataOut_A[10]
  PIN cacheDataOut_A[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 208.9000 0.0000 209.1000 0.6000 ;
    END
  END cacheDataOut_A[9]
  PIN cacheDataOut_A[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.4502 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 187.9000 0.0000 188.1000 0.6000 ;
    END
  END cacheDataOut_A[8]
  PIN cacheDataOut_A[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 169.9000 0.0000 170.1000 0.6000 ;
    END
  END cacheDataOut_A[7]
  PIN cacheDataOut_A[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.766 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.0422 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 148.9000 0.0000 149.1000 0.6000 ;
    END
  END cacheDataOut_A[6]
  PIN cacheDataOut_A[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 131.9000 0.0000 132.1000 0.6000 ;
    END
  END cacheDataOut_A[5]
  PIN cacheDataOut_A[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.68 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.22 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 109.9000 0.0000 110.1000 0.6000 ;
    END
  END cacheDataOut_A[4]
  PIN cacheDataOut_A[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 1.94 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.178 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.8 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.664 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 92.9000 0.0000 93.1000 0.6000 ;
    END
  END cacheDataOut_A[3]
  PIN cacheDataOut_A[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.806 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.1902 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 71.9000 0.0000 72.1000 0.6000 ;
    END
  END cacheDataOut_A[2]
  PIN cacheDataOut_A[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 54.9000 0.0000 55.1000 0.6000 ;
    END
  END cacheDataOut_A[1]
  PIN cacheDataOut_A[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.726 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.8942 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 33.9000 0.0000 34.1000 0.6000 ;
    END
  END cacheDataOut_A[0]
  PIN portA_writtenTo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 760.9000 0.0000 761.1000 0.6000 ;
    END
  END portA_writtenTo
  PIN cacheDataIn_B[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.746 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.9682 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 130.923 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 456.005 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 140.154 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 478.774 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 149.385 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 519.39 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 752.9000 0.0000 753.1000 0.6000 ;
    END
  END cacheDataIn_B[31]
  PIN cacheDataIn_B[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL  ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ  ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2  ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 18.4615 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 43.6923 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.68 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.22 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 39.641 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 114.467 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 48.8718 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 155.082 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 739.9000 0.0000 740.1000 0.6000 ;
    END
  END cacheDataIn_B[30]
  PIN cacheDataIn_B[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.626 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5242 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 127.846 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 444.621 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 137.077 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 467.39 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 146.308 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 508.005 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 714.9000 0.0000 715.1000 0.6000 ;
    END
  END cacheDataIn_B[29]
  PIN cacheDataIn_B[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.806 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.1902 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 132.462 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 461.697 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 141.692 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 484.467 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 150.923 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 525.082 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 701.9000 0.0000 702.1000 0.6000 ;
    END
  END cacheDataIn_B[28]
  PIN cacheDataIn_B[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.786 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.1162 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 131.949 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 459.8 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 141.179 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 482.569 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 150.41 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 523.185 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 675.9000 0.0000 676.1000 0.6000 ;
    END
  END cacheDataIn_B[27]
  PIN cacheDataIn_B[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL  ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ  ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2  ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 18.4615 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 43.6923 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.72 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.368 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 40.6667 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 118.262 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 49.8974 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 158.877 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 662.9000 0.0000 663.1000 0.6000 ;
    END
  END cacheDataIn_B[26]
  PIN cacheDataIn_B[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.706 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.8202 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 129.897 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 452.21 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 139.128 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 474.979 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 148.359 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 515.595 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 637.9000 0.0000 638.1000 0.6000 ;
    END
  END cacheDataIn_B[25]
  PIN cacheDataIn_B[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL  ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ  ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2  ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 18.4615 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 43.6923 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.64 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 38.6154 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 110.672 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 47.8462 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 151.287 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 624.9000 0.0000 625.1000 0.6000 ;
    END
  END cacheDataIn_B[24]
  PIN cacheDataIn_B[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.566 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.3022 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 126.308 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 438.928 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 135.538 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 461.697 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 144.769 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 502.313 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 599.9000 0.0000 600.1000 0.6000 ;
    END
  END cacheDataIn_B[23]
  PIN cacheDataIn_B[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL  ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ  ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 3.06 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.322 LAYER M2  ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 18.4615 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 43.6923 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.76 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.516 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 68.359 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 220.723 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 77.5897 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 261.338 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 585.9000 0.0000 586.1000 0.6000 ;
    END
  END cacheDataIn_B[22]
  PIN cacheDataIn_B[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.746 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.9682 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 130.923 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 456.005 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 140.154 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 478.774 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 149.385 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 519.39 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 560.9000 0.0000 561.1000 0.6000 ;
    END
  END cacheDataIn_B[21]
  PIN cacheDataIn_B[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL  ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ  ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2  ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 18.4615 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 43.6923 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.68 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.22 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 39.641 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 114.467 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 48.8718 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 155.082 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 547.9000 0.0000 548.1000 0.6000 ;
    END
  END cacheDataIn_B[20]
  PIN cacheDataIn_B[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.626 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5242 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 127.846 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 444.621 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 137.077 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 467.39 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 146.308 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 508.005 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 522.9000 0.0000 523.1000 0.6000 ;
    END
  END cacheDataIn_B[19]
  PIN cacheDataIn_B[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL  ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ  ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.98 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.626 LAYER M2  ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 18.4615 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 43.6923 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.8 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.664 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 122.718 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 421.851 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 131.949 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 462.467 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 508.9000 0.0000 509.1000 0.6000 ;
    END
  END cacheDataIn_B[18]
  PIN cacheDataIn_B[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.786 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.1162 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 131.949 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 459.8 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 141.179 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 482.569 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 150.41 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 523.185 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 483.9000 0.0000 484.1000 0.6000 ;
    END
  END cacheDataIn_B[17]
  PIN cacheDataIn_B[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL  ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ  ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2  ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 18.4615 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 43.6923 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.72 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.368 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 40.6667 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 118.262 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 49.8974 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 158.877 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 470.9000 0.0000 471.1000 0.6000 ;
    END
  END cacheDataIn_B[16]
  PIN cacheDataIn_B[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.69 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.761 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 129.487 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 450.692 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 138.718 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 473.462 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 147.949 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 514.077 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 319.9000 0.0000 320.1000 0.6000 ;
    END
  END cacheDataIn_B[15]
  PIN cacheDataIn_B[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL  ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ  ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2  ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 18.4615 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 43.6923 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.64 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 38.6154 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 110.672 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 47.8462 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 151.287 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 306.9000 0.0000 307.1000 0.6000 ;
    END
  END cacheDataIn_B[14]
  PIN cacheDataIn_B[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.566 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.3022 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 126.308 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 438.928 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 135.538 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 461.697 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 144.769 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 502.313 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 281.9000 0.0000 282.1000 0.6000 ;
    END
  END cacheDataIn_B[13]
  PIN cacheDataIn_B[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 127.333 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 446.518 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 136.564 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 469.287 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 145.795 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 509.903 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 267.9000 0.0000 268.1000 0.6000 ;
    END
  END cacheDataIn_B[12]
  PIN cacheDataIn_B[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.73 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.909 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 130.513 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 454.487 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 139.744 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 477.256 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 148.974 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 517.872 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 242.9000 0.0000 243.1000 0.6000 ;
    END
  END cacheDataIn_B[11]
  PIN cacheDataIn_B[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL  ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ  ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2  ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 18.4615 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 43.6923 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.68 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.22 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 39.641 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 114.467 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 48.8718 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 155.082 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 229.9000 0.0000 230.1000 0.6000 ;
    END
  END cacheDataIn_B[10]
  PIN cacheDataIn_B[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.61 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.465 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 127.436 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 443.103 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 136.667 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 465.872 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 145.897 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 506.487 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 204.9000 0.0000 205.1000 0.6000 ;
    END
  END cacheDataIn_B[9]
  PIN cacheDataIn_B[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.806 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.1902 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 132.462 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 461.697 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 141.692 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 484.467 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 150.923 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 525.082 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 191.9000 0.0000 192.1000 0.6000 ;
    END
  END cacheDataIn_B[8]
  PIN cacheDataIn_B[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.77 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.057 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 131.538 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 458.282 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 140.769 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 481.051 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 150 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 521.667 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 165.9000 0.0000 166.1000 0.6000 ;
    END
  END cacheDataIn_B[7]
  PIN cacheDataIn_B[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL  ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ  ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2  ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 18.4615 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 43.6923 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.72 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.368 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 40.6667 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 118.262 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 49.8974 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 158.877 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 152.9000 0.0000 153.1000 0.6000 ;
    END
  END cacheDataIn_B[6]
  PIN cacheDataIn_B[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.69 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.761 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 129.487 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 450.692 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 138.718 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 473.462 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 147.949 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 514.077 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 127.9000 0.0000 128.1000 0.6000 ;
    END
  END cacheDataIn_B[5]
  PIN cacheDataIn_B[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 127.333 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 446.518 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 136.564 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 469.287 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 145.795 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 509.903 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 113.9000 0.0000 114.1000 0.6000 ;
    END
  END cacheDataIn_B[4]
  PIN cacheDataIn_B[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 127.333 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 446.518 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 136.564 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 469.287 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 145.795 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 509.903 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 88.9000 0.0000 89.1000 0.6000 ;
    END
  END cacheDataIn_B[3]
  PIN cacheDataIn_B[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 127.333 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 446.518 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 136.564 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 469.287 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 145.795 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 509.903 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 75.9000 0.0000 76.1000 0.6000 ;
    END
  END cacheDataIn_B[2]
  PIN cacheDataIn_B[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.73 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.909 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 130.513 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 454.487 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 139.744 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 477.256 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 148.974 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 517.872 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 50.9000 0.0000 51.1000 0.6000 ;
    END
  END cacheDataIn_B[1]
  PIN cacheDataIn_B[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL  ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ  ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2  ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 18.4615 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 43.6923 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.68 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.22 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 39.641 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 114.467 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 48.8718 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 155.082 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 37.9000 0.0000 38.1000 0.6000 ;
    END
  END cacheDataIn_B[0]
  PIN cacheAddressIn_B[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL  ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ  ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2  ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 18.4615 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 43.6923 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 2.76 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.916 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 92.9744 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 311.8 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 102.205 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 352.415 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 369.9000 0.0000 370.1000 0.6000 ;
    END
  END cacheAddressIn_B[7]
  PIN cacheAddressIn_B[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 127.333 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 446.518 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 136.564 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 469.287 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 145.795 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 509.903 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 366.9000 0.0000 367.1000 0.6000 ;
    END
  END cacheAddressIn_B[6]
  PIN cacheAddressIn_B[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 127.333 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 446.518 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 136.564 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 469.287 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 145.795 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 509.903 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 363.9000 0.0000 364.1000 0.6000 ;
    END
  END cacheAddressIn_B[5]
  PIN cacheAddressIn_B[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VL  ;
    ANTENNAMAXCUTCAR 1.02564 LAYER VQ  ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2  ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 18.4615 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 43.6923 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 2 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.104 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 73.4872 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 239.697 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 82.7179 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 280.313 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 360.9000 0.0000 361.1000 0.6000 ;
    END
  END cacheAddressIn_B[4]
  PIN cacheAddressIn_B[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 127.333 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 446.518 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 136.564 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 469.287 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 145.795 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 509.903 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 357.9000 0.0000 358.1000 0.6000 ;
    END
  END cacheAddressIn_B[3]
  PIN cacheAddressIn_B[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 127.333 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 446.518 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 136.564 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 469.287 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 145.795 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 509.903 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 354.9000 0.0000 355.1000 0.6000 ;
    END
  END cacheAddressIn_B[2]
  PIN cacheAddressIn_B[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 127.333 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 446.518 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 136.564 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 469.287 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 145.795 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 509.903 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 351.9000 0.0000 352.1000 0.6000 ;
    END
  END cacheAddressIn_B[1]
  PIN cacheAddressIn_B[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 127.333 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 446.518 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 136.564 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 469.287 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 145.795 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 509.903 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 348.9000 0.0000 349.1000 0.6000 ;
    END
  END cacheAddressIn_B[0]
  PIN memWrite_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.754 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.9978 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.039 LAYER M2  ;
    ANTENNAMAXAREACAR 131.128 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 456.764 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNAGATEAREA 0.039 LAYER M3  ;
    ANTENNAMAXAREACAR 140.359 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 479.533 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    ANTENNAGATEAREA 0.039 LAYER MQ  ;
    ANTENNAMAXAREACAR 149.59 LAYER MQ  ;
    ANTENNAMAXSIDEAREACAR 520.149 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 340.9000 0.0000 341.1000 0.6000 ;
    END
  END memWrite_B
  PIN cacheDataOut_B[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.766 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.0422 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 754.9000 0.0000 755.1000 0.6000 ;
    END
  END cacheDataOut_B[31]
  PIN cacheDataOut_B[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 737.9000 0.0000 738.1000 0.6000 ;
    END
  END cacheDataOut_B[30]
  PIN cacheDataOut_B[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.646 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 716.9000 0.0000 717.1000 0.6000 ;
    END
  END cacheDataOut_B[29]
  PIN cacheDataOut_B[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.79 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.131 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 699.9000 0.0000 700.1000 0.6000 ;
    END
  END cacheDataOut_B[28]
  PIN cacheDataOut_B[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.806 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.1902 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 677.9000 0.0000 678.1000 0.6000 ;
    END
  END cacheDataOut_B[27]
  PIN cacheDataOut_B[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 660.9000 0.0000 661.1000 0.6000 ;
    END
  END cacheDataOut_B[26]
  PIN cacheDataOut_B[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.726 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.8942 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 639.9000 0.0000 640.1000 0.6000 ;
    END
  END cacheDataOut_B[25]
  PIN cacheDataOut_B[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.37 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.64 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 622.9000 0.0000 623.1000 0.6000 ;
    END
  END cacheDataOut_B[24]
  PIN cacheDataOut_B[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.4502 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 601.9000 0.0000 602.1000 0.6000 ;
    END
  END cacheDataOut_B[23]
  PIN cacheDataOut_B[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.85 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.701 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 583.9000 0.0000 584.1000 0.6000 ;
    END
  END cacheDataOut_B[22]
  PIN cacheDataOut_B[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.766 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.0422 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 562.9000 0.0000 563.1000 0.6000 ;
    END
  END cacheDataOut_B[21]
  PIN cacheDataOut_B[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 545.9000 0.0000 546.1000 0.6000 ;
    END
  END cacheDataOut_B[20]
  PIN cacheDataOut_B[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.646 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 524.9000 0.0000 525.1000 0.6000 ;
    END
  END cacheDataOut_B[19]
  PIN cacheDataOut_B[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 1.86 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.882 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.8 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.664 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 506.9000 0.0000 507.1000 0.6000 ;
    END
  END cacheDataOut_B[18]
  PIN cacheDataOut_B[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.806 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.1902 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 485.9000 0.0000 486.1000 0.6000 ;
    END
  END cacheDataOut_B[17]
  PIN cacheDataOut_B[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 468.9000 0.0000 469.1000 0.6000 ;
    END
  END cacheDataOut_B[16]
  PIN cacheDataOut_B[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.726 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.8942 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 321.9000 0.0000 322.1000 0.6000 ;
    END
  END cacheDataOut_B[15]
  PIN cacheDataOut_B[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 304.9000 0.0000 305.1000 0.6000 ;
    END
  END cacheDataOut_B[14]
  PIN cacheDataOut_B[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.4502 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 283.9000 0.0000 284.1000 0.6000 ;
    END
  END cacheDataOut_B[13]
  PIN cacheDataOut_B[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 265.9000 0.0000 266.1000 0.6000 ;
    END
  END cacheDataOut_B[12]
  PIN cacheDataOut_B[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.766 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.0422 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 244.9000 0.0000 245.1000 0.6000 ;
    END
  END cacheDataOut_B[11]
  PIN cacheDataOut_B[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 227.9000 0.0000 228.1000 0.6000 ;
    END
  END cacheDataOut_B[10]
  PIN cacheDataOut_B[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.646 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 206.9000 0.0000 207.1000 0.6000 ;
    END
  END cacheDataOut_B[9]
  PIN cacheDataOut_B[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.774 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.0718 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 189.9000 0.0000 190.1000 0.6000 ;
    END
  END cacheDataOut_B[8]
  PIN cacheDataOut_B[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.806 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.1902 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 167.9000 0.0000 168.1000 0.6000 ;
    END
  END cacheDataOut_B[7]
  PIN cacheDataOut_B[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 150.9000 0.0000 151.1000 0.6000 ;
    END
  END cacheDataOut_B[6]
  PIN cacheDataOut_B[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.726 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.8942 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 129.9000 0.0000 130.1000 0.6000 ;
    END
  END cacheDataOut_B[5]
  PIN cacheDataOut_B[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 111.9000 0.0000 112.1000 0.6000 ;
    END
  END cacheDataOut_B[4]
  PIN cacheDataOut_B[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.1 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.17 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.64 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 90.9000 0.0000 91.1000 0.6000 ;
    END
  END cacheDataOut_B[3]
  PIN cacheDataOut_B[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 73.9000 0.0000 74.1000 0.6000 ;
    END
  END cacheDataOut_B[2]
  PIN cacheDataOut_B[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.766 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.0422 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 52.9000 0.0000 53.1000 0.6000 ;
    END
  END cacheDataOut_B[1]
  PIN cacheDataOut_B[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16 LAYER M2  ;
    ANTENNAPARTIALMETALAREA 4.606 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5982 LAYER M2  ;
    ANTENNADIFFAREA 0.16 LAYER M3  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.888 LAYER M3  ;
    ANTENNADIFFAREA 0.16 LAYER MQ  ;
    ANTENNAPARTIALMETALAREA 0.36 LAYER MQ  ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER MQ  ;
    PORT
      LAYER M2 ;
        RECT 35.9000 0.0000 36.1000 0.6000 ;
    END
  END cacheDataOut_B[0]
  PIN portB_writtenTo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 762.9000 0.0000 763.1000 0.6000 ;
    END
  END portB_writtenTo
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER MQ ;
        RECT 17.8800 27.7200 21.8800 28.2800 ;
        RECT 17.8800 42.1200 21.8800 42.5700 ;
        RECT 17.8800 34.9200 21.8800 35.4800 ;
        RECT 17.8800 70.9200 21.8800 71.4800 ;
        RECT 17.8800 63.7200 21.8800 64.2800 ;
        RECT 17.8800 78.1200 21.8800 78.6800 ;
        RECT 17.8800 85.3200 21.8800 85.8800 ;
        RECT 17.8800 236.5200 21.8800 237.0800 ;
        RECT 771.2800 27.7200 775.2800 28.2800 ;
        RECT 771.2800 42.1200 775.2800 42.5700 ;
        RECT 771.2800 34.9200 775.2800 35.4800 ;
        RECT 771.2800 78.1200 775.2800 78.6800 ;
        RECT 771.2800 70.9200 775.2800 71.4800 ;
        RECT 771.2800 63.7200 775.2800 64.2800 ;
        RECT 771.2800 85.3200 775.2800 85.8800 ;
        RECT 771.2800 236.5200 775.2800 237.0800 ;
        RECT 17.8800 452.5200 21.8800 453.0800 ;
        RECT 17.8800 675.7200 21.8800 676.2800 ;
        RECT 771.2800 452.5200 775.2800 453.0800 ;
        RECT 771.2800 675.7200 775.2800 676.2800 ;
    END
# end of P/G power stripe data as pin

  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER MQ ;
        RECT 18.5000 6.0000 22.5000 15.3900 ;
        RECT 18.5000 6.0000 22.5000 9.0000 ;
        RECT 18.5000 11.3900 22.5000 15.3900 ;
        RECT 18.5000 9.7200 22.5000 10.2800 ;
        RECT 12.7600 31.3200 16.7600 31.8800 ;
        RECT 12.7600 45.7200 16.7600 46.2800 ;
        RECT 12.7600 38.5200 16.7600 39.0800 ;
        RECT 12.7600 52.9200 16.7600 53.4800 ;
        RECT 12.7600 67.3200 16.7600 67.8800 ;
        RECT 12.7600 60.1200 16.7600 60.6800 ;
        RECT 12.7600 74.5200 16.7600 75.0800 ;
        RECT 12.7600 96.1200 16.7600 96.6800 ;
        RECT 12.7600 88.9200 16.7600 89.4800 ;
        RECT 12.7600 103.3200 16.7600 103.8800 ;
        RECT 12.7600 117.7200 16.7600 118.2800 ;
        RECT 12.7600 110.5200 16.7600 111.0800 ;
        RECT 12.7600 132.1200 16.7600 132.6800 ;
        RECT 12.7600 124.9200 16.7600 125.4800 ;
        RECT 12.7600 139.3200 16.7600 139.8800 ;
        RECT 12.7600 153.7200 16.7600 154.2800 ;
        RECT 12.7600 146.5200 16.7600 147.0800 ;
        RECT 12.7600 168.1200 16.7600 168.6800 ;
        RECT 12.7600 160.9200 16.7600 161.4800 ;
        RECT 12.7600 182.5200 16.7600 183.0800 ;
        RECT 12.7600 175.3200 16.7600 175.8800 ;
        RECT 12.7600 189.7200 16.7600 190.2800 ;
        RECT 12.7600 204.1200 16.7600 204.6800 ;
        RECT 12.7600 196.9200 16.7600 197.4800 ;
        RECT 12.7600 218.5200 16.7600 219.0800 ;
        RECT 12.7600 211.3200 16.7600 211.8800 ;
        RECT 12.7600 232.9200 16.7600 233.4800 ;
        RECT 12.7600 225.7200 16.7600 226.2800 ;
        RECT 12.7600 240.1200 16.7600 240.6800 ;
        RECT 12.7600 254.5200 16.7600 255.0800 ;
        RECT 12.7600 247.3200 16.7600 247.8800 ;
        RECT 12.7600 283.3200 16.7600 283.8800 ;
        RECT 12.7600 268.9200 16.7600 269.4800 ;
        RECT 12.7600 261.7200 16.7600 262.2800 ;
        RECT 12.7600 276.1200 16.7600 276.6800 ;
        RECT 12.7600 290.5200 16.7600 291.0800 ;
        RECT 12.7600 304.9200 16.7600 305.4800 ;
        RECT 12.7600 297.7200 16.7600 298.2800 ;
        RECT 12.7600 319.3200 16.7600 319.8800 ;
        RECT 12.7600 312.1200 16.7600 312.6800 ;
        RECT 12.7600 326.5200 16.7600 327.0800 ;
        RECT 12.7600 340.9200 16.7600 341.4800 ;
        RECT 12.7600 333.7200 16.7600 334.2800 ;
        RECT 12.7600 355.3200 16.7600 355.8800 ;
        RECT 12.7600 348.1200 16.7600 348.6800 ;
        RECT 776.4000 16.9200 780.4000 17.4800 ;
        RECT 776.4000 31.3200 780.4000 31.8800 ;
        RECT 776.4000 45.7200 780.4000 46.2800 ;
        RECT 776.4000 38.5200 780.4000 39.0800 ;
        RECT 776.4000 52.9200 780.4000 53.4800 ;
        RECT 776.4000 67.3200 780.4000 67.8800 ;
        RECT 776.4000 60.1200 780.4000 60.6800 ;
        RECT 776.4000 74.5200 780.4000 75.0800 ;
        RECT 776.4000 96.1200 780.4000 96.6800 ;
        RECT 776.4000 88.9200 780.4000 89.4800 ;
        RECT 776.4000 103.3200 780.4000 103.8800 ;
        RECT 776.4000 117.7200 780.4000 118.2800 ;
        RECT 776.4000 110.5200 780.4000 111.0800 ;
        RECT 776.4000 132.1200 780.4000 132.6800 ;
        RECT 776.4000 124.9200 780.4000 125.4800 ;
        RECT 776.4000 139.3200 780.4000 139.8800 ;
        RECT 776.4000 153.7200 780.4000 154.2800 ;
        RECT 776.4000 146.5200 780.4000 147.0800 ;
        RECT 776.4000 168.1200 780.4000 168.6800 ;
        RECT 776.4000 160.9200 780.4000 161.4800 ;
        RECT 776.4000 182.5200 780.4000 183.0800 ;
        RECT 776.4000 175.3200 780.4000 175.8800 ;
        RECT 776.4000 189.7200 780.4000 190.2800 ;
        RECT 776.4000 204.1200 780.4000 204.6800 ;
        RECT 776.4000 196.9200 780.4000 197.4800 ;
        RECT 776.4000 218.5200 780.4000 219.0800 ;
        RECT 776.4000 211.3200 780.4000 211.8800 ;
        RECT 776.4000 232.9200 780.4000 233.4800 ;
        RECT 776.4000 225.7200 780.4000 226.2800 ;
        RECT 776.4000 240.1200 780.4000 240.6800 ;
        RECT 776.4000 254.5200 780.4000 255.0800 ;
        RECT 776.4000 247.3200 780.4000 247.8800 ;
        RECT 776.4000 283.3200 780.4000 283.8800 ;
        RECT 776.4000 268.9200 780.4000 269.4800 ;
        RECT 776.4000 261.7200 780.4000 262.2800 ;
        RECT 776.4000 276.1200 780.4000 276.6800 ;
        RECT 776.4000 290.5200 780.4000 291.0800 ;
        RECT 776.4000 304.9200 780.4000 305.4800 ;
        RECT 776.4000 297.7200 780.4000 298.2800 ;
        RECT 776.4000 319.3200 780.4000 319.8800 ;
        RECT 776.4000 312.1200 780.4000 312.6800 ;
        RECT 776.4000 326.5200 780.4000 327.0800 ;
        RECT 776.4000 340.9200 780.4000 341.4800 ;
        RECT 776.4000 333.7200 780.4000 334.2800 ;
        RECT 776.4000 355.3200 780.4000 355.8800 ;
        RECT 776.4000 348.1200 780.4000 348.6800 ;
        RECT 12.7600 556.9200 16.7600 557.4800 ;
        RECT 12.7600 369.7200 16.7600 370.2800 ;
        RECT 12.7600 362.5200 16.7600 363.0800 ;
        RECT 12.7600 376.9200 16.7600 377.4800 ;
        RECT 12.7600 391.3200 16.7600 391.8800 ;
        RECT 12.7600 384.1200 16.7600 384.6800 ;
        RECT 12.7600 405.7200 16.7600 406.2800 ;
        RECT 12.7600 398.5200 16.7600 399.0800 ;
        RECT 12.7600 420.1200 16.7600 420.6800 ;
        RECT 12.7600 412.9200 16.7600 413.4800 ;
        RECT 12.7600 427.3200 16.7600 427.8800 ;
        RECT 12.7600 441.7200 16.7600 442.2800 ;
        RECT 12.7600 434.5200 16.7600 435.0800 ;
        RECT 12.7600 456.1200 16.7600 456.6800 ;
        RECT 12.7600 448.9200 16.7600 449.4800 ;
        RECT 12.7600 463.3200 16.7600 463.8800 ;
        RECT 12.7600 477.7200 16.7600 478.2800 ;
        RECT 12.7600 470.5200 16.7600 471.0800 ;
        RECT 12.7600 492.1200 16.7600 492.6800 ;
        RECT 12.7600 484.9200 16.7600 485.4800 ;
        RECT 12.7600 506.5200 16.7600 507.0800 ;
        RECT 12.7600 499.3200 16.7600 499.8800 ;
        RECT 12.7600 513.7200 16.7600 514.2800 ;
        RECT 12.7600 528.1200 16.7600 528.6800 ;
        RECT 12.7600 520.9200 16.7600 521.4800 ;
        RECT 12.7600 542.5200 16.7600 543.0800 ;
        RECT 12.7600 535.3200 16.7600 535.8800 ;
        RECT 12.7600 549.7200 16.7600 550.2800 ;
        RECT 12.7600 564.1200 16.7600 564.6800 ;
        RECT 12.7600 578.5200 16.7600 579.0800 ;
        RECT 12.7600 571.3200 16.7600 571.8800 ;
        RECT 12.7600 592.9200 16.7600 593.4800 ;
        RECT 12.7600 585.7200 16.7600 586.2800 ;
        RECT 12.7600 600.1200 16.7600 600.6800 ;
        RECT 12.7600 614.5200 16.7600 615.0800 ;
        RECT 12.7600 607.3200 16.7600 607.8800 ;
        RECT 12.7600 628.9200 16.7600 629.4800 ;
        RECT 12.7600 621.7200 16.7600 622.2800 ;
        RECT 12.7600 643.3200 16.7600 643.8800 ;
        RECT 12.7600 636.1200 16.7600 636.6800 ;
        RECT 12.7600 650.5200 16.7600 651.0800 ;
        RECT 12.7600 664.9200 16.7600 665.4800 ;
        RECT 12.7600 657.7200 16.7600 658.2800 ;
        RECT 12.7600 672.1200 16.7600 672.6800 ;
        RECT 776.4000 556.9200 780.4000 557.4800 ;
        RECT 776.4000 369.7200 780.4000 370.2800 ;
        RECT 776.4000 362.5200 780.4000 363.0800 ;
        RECT 776.4000 376.9200 780.4000 377.4800 ;
        RECT 776.4000 391.3200 780.4000 391.8800 ;
        RECT 776.4000 384.1200 780.4000 384.6800 ;
        RECT 776.4000 405.7200 780.4000 406.2800 ;
        RECT 776.4000 398.5200 780.4000 399.0800 ;
        RECT 776.4000 420.1200 780.4000 420.6800 ;
        RECT 776.4000 412.9200 780.4000 413.4800 ;
        RECT 776.4000 427.3200 780.4000 427.8800 ;
        RECT 776.4000 441.7200 780.4000 442.2800 ;
        RECT 776.4000 434.5200 780.4000 435.0800 ;
        RECT 776.4000 456.1200 780.4000 456.6800 ;
        RECT 776.4000 448.9200 780.4000 449.4800 ;
        RECT 776.4000 463.3200 780.4000 463.8800 ;
        RECT 776.4000 477.7200 780.4000 478.2800 ;
        RECT 776.4000 470.5200 780.4000 471.0800 ;
        RECT 776.4000 492.1200 780.4000 492.6800 ;
        RECT 776.4000 484.9200 780.4000 485.4800 ;
        RECT 776.4000 506.5200 780.4000 507.0800 ;
        RECT 776.4000 499.3200 780.4000 499.8800 ;
        RECT 776.4000 513.7200 780.4000 514.2800 ;
        RECT 776.4000 528.1200 780.4000 528.6800 ;
        RECT 776.4000 520.9200 780.4000 521.4800 ;
        RECT 776.4000 542.5200 780.4000 543.0800 ;
        RECT 776.4000 535.3200 780.4000 535.8800 ;
        RECT 776.4000 549.7200 780.4000 550.2800 ;
        RECT 776.4000 564.1200 780.4000 564.6800 ;
        RECT 776.4000 578.5200 780.4000 579.0800 ;
        RECT 776.4000 571.3200 780.4000 571.8800 ;
        RECT 776.4000 592.9200 780.4000 593.4800 ;
        RECT 776.4000 585.7200 780.4000 586.2800 ;
        RECT 776.4000 600.1200 780.4000 600.6800 ;
        RECT 776.4000 614.5200 780.4000 615.0800 ;
        RECT 776.4000 607.3200 780.4000 607.8800 ;
        RECT 776.4000 628.9200 780.4000 629.4800 ;
        RECT 776.4000 621.7200 780.4000 622.2800 ;
        RECT 776.4000 643.3200 780.4000 643.8800 ;
        RECT 776.4000 636.1200 780.4000 636.6800 ;
        RECT 776.4000 650.5200 780.4000 651.0800 ;
        RECT 776.4000 664.9200 780.4000 665.4800 ;
        RECT 776.4000 657.7200 780.4000 658.2800 ;
        RECT 776.4000 679.3200 780.4000 679.8800 ;
        RECT 776.4000 672.1200 780.4000 672.6800 ;
    END
# end of P/G power stripe data as pin

  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 796.5000 716.0000 ;
    LAYER M2 ;
      RECT 0.0000 2.5200 796.5000 716.0000 ;
      RECT 765.0200 0.0000 796.5000 2.5200 ;
      RECT 742.0200 0.0000 750.9800 2.5200 ;
      RECT 723.0200 0.0000 731.9800 2.5200 ;
      RECT 704.0200 0.0000 712.9800 2.5200 ;
      RECT 684.0200 0.0000 693.9800 2.5200 ;
      RECT 665.0200 0.0000 673.9800 2.5200 ;
      RECT 646.0200 0.0000 654.9800 2.5200 ;
      RECT 627.0200 0.0000 635.9800 2.5200 ;
      RECT 608.0200 0.0000 616.9800 2.5200 ;
      RECT 588.0200 0.0000 597.9800 2.5200 ;
      RECT 569.0200 0.0000 577.9800 2.5200 ;
      RECT 550.0200 0.0000 558.9800 2.5200 ;
      RECT 531.0200 0.0000 539.9800 2.5200 ;
      RECT 511.0200 0.0000 520.9800 2.5200 ;
      RECT 492.0200 0.0000 500.9800 2.5200 ;
      RECT 473.0200 0.0000 481.9800 2.5200 ;
      RECT 436.0200 0.0000 462.9800 2.5200 ;
      RECT 372.0200 0.0000 407.9800 2.5200 ;
      RECT 343.0200 0.0000 346.9800 2.5200 ;
      RECT 328.0200 0.0000 338.9800 2.5200 ;
      RECT 309.0200 0.0000 317.9800 2.5200 ;
      RECT 290.0200 0.0000 298.9800 2.5200 ;
      RECT 270.0200 0.0000 279.9800 2.5200 ;
      RECT 251.0200 0.0000 259.9800 2.5200 ;
      RECT 232.0200 0.0000 240.9800 2.5200 ;
      RECT 213.0200 0.0000 221.9800 2.5200 ;
      RECT 194.0200 0.0000 202.9800 2.5200 ;
      RECT 174.0200 0.0000 183.9800 2.5200 ;
      RECT 155.0200 0.0000 163.9800 2.5200 ;
      RECT 136.0200 0.0000 144.9800 2.5200 ;
      RECT 116.0200 0.0000 125.9800 2.5200 ;
      RECT 97.0200 0.0000 105.9800 2.5200 ;
      RECT 78.0200 0.0000 86.9800 2.5200 ;
      RECT 59.0200 0.0000 67.9800 2.5200 ;
      RECT 40.0200 0.0000 48.9800 2.5200 ;
      RECT 0.0000 0.0000 29.9800 2.5200 ;
    LAYER M3 ;
      RECT 0.0000 2.5200 796.5000 716.0000 ;
      RECT 345.0200 0.0000 796.5000 2.5200 ;
      RECT 337.0200 0.0000 340.9800 2.5200 ;
      RECT 0.0000 0.0000 332.9800 2.5200 ;
    LAYER MQ ;
      RECT 0.0000 681.8000 796.5000 716.0000 ;
      RECT 0.0000 678.2000 774.4800 681.8000 ;
      RECT 782.3200 677.4000 796.5000 681.8000 ;
      RECT 777.2000 674.6000 796.5000 677.4000 ;
      RECT 0.0000 674.6000 15.9600 678.2000 ;
      RECT 23.8000 673.8000 769.3600 678.2000 ;
      RECT 782.3200 670.2000 796.5000 674.6000 ;
      RECT 18.6800 670.2000 774.4800 673.8000 ;
      RECT 0.0000 670.2000 10.8400 674.6000 ;
      RECT 0.0000 667.4000 796.5000 670.2000 ;
      RECT 782.3200 663.0000 796.5000 667.4000 ;
      RECT 18.6800 663.0000 774.4800 667.4000 ;
      RECT 0.0000 663.0000 10.8400 667.4000 ;
      RECT 0.0000 660.2000 796.5000 663.0000 ;
      RECT 782.3200 655.8000 796.5000 660.2000 ;
      RECT 18.6800 655.8000 774.4800 660.2000 ;
      RECT 0.0000 655.8000 10.8400 660.2000 ;
      RECT 0.0000 653.0000 796.5000 655.8000 ;
      RECT 782.3200 648.6000 796.5000 653.0000 ;
      RECT 18.6800 648.6000 774.4800 653.0000 ;
      RECT 0.0000 648.6000 10.8400 653.0000 ;
      RECT 0.0000 645.8000 796.5000 648.6000 ;
      RECT 782.3200 641.4000 796.5000 645.8000 ;
      RECT 18.6800 641.4000 774.4800 645.8000 ;
      RECT 0.0000 641.4000 10.8400 645.8000 ;
      RECT 0.0000 638.6000 796.5000 641.4000 ;
      RECT 782.3200 634.2000 796.5000 638.6000 ;
      RECT 18.6800 634.2000 774.4800 638.6000 ;
      RECT 0.0000 634.2000 10.8400 638.6000 ;
      RECT 0.0000 631.4000 796.5000 634.2000 ;
      RECT 782.3200 627.0000 796.5000 631.4000 ;
      RECT 18.6800 627.0000 774.4800 631.4000 ;
      RECT 0.0000 627.0000 10.8400 631.4000 ;
      RECT 0.0000 624.2000 796.5000 627.0000 ;
      RECT 782.3200 619.8000 796.5000 624.2000 ;
      RECT 18.6800 619.8000 774.4800 624.2000 ;
      RECT 0.0000 619.8000 10.8400 624.2000 ;
      RECT 0.0000 617.0000 796.5000 619.8000 ;
      RECT 782.3200 612.6000 796.5000 617.0000 ;
      RECT 18.6800 612.6000 774.4800 617.0000 ;
      RECT 0.0000 612.6000 10.8400 617.0000 ;
      RECT 0.0000 609.8000 796.5000 612.6000 ;
      RECT 782.3200 605.4000 796.5000 609.8000 ;
      RECT 18.6800 605.4000 774.4800 609.8000 ;
      RECT 0.0000 605.4000 10.8400 609.8000 ;
      RECT 0.0000 602.6000 796.5000 605.4000 ;
      RECT 782.3200 598.2000 796.5000 602.6000 ;
      RECT 18.6800 598.2000 774.4800 602.6000 ;
      RECT 0.0000 598.2000 10.8400 602.6000 ;
      RECT 0.0000 595.4000 796.5000 598.2000 ;
      RECT 782.3200 591.0000 796.5000 595.4000 ;
      RECT 18.6800 591.0000 774.4800 595.4000 ;
      RECT 0.0000 591.0000 10.8400 595.4000 ;
      RECT 0.0000 588.2000 796.5000 591.0000 ;
      RECT 782.3200 583.8000 796.5000 588.2000 ;
      RECT 18.6800 583.8000 774.4800 588.2000 ;
      RECT 0.0000 583.8000 10.8400 588.2000 ;
      RECT 0.0000 581.0000 796.5000 583.8000 ;
      RECT 782.3200 576.6000 796.5000 581.0000 ;
      RECT 18.6800 576.6000 774.4800 581.0000 ;
      RECT 0.0000 576.6000 10.8400 581.0000 ;
      RECT 0.0000 573.8000 796.5000 576.6000 ;
      RECT 782.3200 569.4000 796.5000 573.8000 ;
      RECT 18.6800 569.4000 774.4800 573.8000 ;
      RECT 0.0000 569.4000 10.8400 573.8000 ;
      RECT 0.0000 566.6000 796.5000 569.4000 ;
      RECT 782.3200 562.2000 796.5000 566.6000 ;
      RECT 18.6800 562.2000 774.4800 566.6000 ;
      RECT 0.0000 562.2000 10.8400 566.6000 ;
      RECT 0.0000 559.4000 796.5000 562.2000 ;
      RECT 782.3200 555.0000 796.5000 559.4000 ;
      RECT 18.6800 555.0000 774.4800 559.4000 ;
      RECT 0.0000 555.0000 10.8400 559.4000 ;
      RECT 0.0000 552.2000 796.5000 555.0000 ;
      RECT 782.3200 547.8000 796.5000 552.2000 ;
      RECT 18.6800 547.8000 774.4800 552.2000 ;
      RECT 0.0000 547.8000 10.8400 552.2000 ;
      RECT 0.0000 545.0000 796.5000 547.8000 ;
      RECT 782.3200 540.6000 796.5000 545.0000 ;
      RECT 18.6800 540.6000 774.4800 545.0000 ;
      RECT 0.0000 540.6000 10.8400 545.0000 ;
      RECT 0.0000 537.8000 796.5000 540.6000 ;
      RECT 782.3200 533.4000 796.5000 537.8000 ;
      RECT 18.6800 533.4000 774.4800 537.8000 ;
      RECT 0.0000 533.4000 10.8400 537.8000 ;
      RECT 0.0000 530.6000 796.5000 533.4000 ;
      RECT 782.3200 526.2000 796.5000 530.6000 ;
      RECT 18.6800 526.2000 774.4800 530.6000 ;
      RECT 0.0000 526.2000 10.8400 530.6000 ;
      RECT 0.0000 523.4000 796.5000 526.2000 ;
      RECT 782.3200 519.0000 796.5000 523.4000 ;
      RECT 18.6800 519.0000 774.4800 523.4000 ;
      RECT 0.0000 519.0000 10.8400 523.4000 ;
      RECT 0.0000 516.2000 796.5000 519.0000 ;
      RECT 782.3200 511.8000 796.5000 516.2000 ;
      RECT 18.6800 511.8000 774.4800 516.2000 ;
      RECT 0.0000 511.8000 10.8400 516.2000 ;
      RECT 0.0000 509.0000 796.5000 511.8000 ;
      RECT 782.3200 504.6000 796.5000 509.0000 ;
      RECT 18.6800 504.6000 774.4800 509.0000 ;
      RECT 0.0000 504.6000 10.8400 509.0000 ;
      RECT 0.0000 501.8000 796.5000 504.6000 ;
      RECT 782.3200 497.4000 796.5000 501.8000 ;
      RECT 18.6800 497.4000 774.4800 501.8000 ;
      RECT 0.0000 497.4000 10.8400 501.8000 ;
      RECT 0.0000 494.6000 796.5000 497.4000 ;
      RECT 782.3200 490.2000 796.5000 494.6000 ;
      RECT 18.6800 490.2000 774.4800 494.6000 ;
      RECT 0.0000 490.2000 10.8400 494.6000 ;
      RECT 0.0000 487.4000 796.5000 490.2000 ;
      RECT 782.3200 483.0000 796.5000 487.4000 ;
      RECT 18.6800 483.0000 774.4800 487.4000 ;
      RECT 0.0000 483.0000 10.8400 487.4000 ;
      RECT 0.0000 480.2000 796.5000 483.0000 ;
      RECT 782.3200 475.8000 796.5000 480.2000 ;
      RECT 18.6800 475.8000 774.4800 480.2000 ;
      RECT 0.0000 475.8000 10.8400 480.2000 ;
      RECT 0.0000 473.0000 796.5000 475.8000 ;
      RECT 782.3200 468.6000 796.5000 473.0000 ;
      RECT 18.6800 468.6000 774.4800 473.0000 ;
      RECT 0.0000 468.6000 10.8400 473.0000 ;
      RECT 0.0000 465.8000 796.5000 468.6000 ;
      RECT 782.3200 461.4000 796.5000 465.8000 ;
      RECT 18.6800 461.4000 774.4800 465.8000 ;
      RECT 0.0000 461.4000 10.8400 465.8000 ;
      RECT 0.0000 458.6000 796.5000 461.4000 ;
      RECT 18.6800 455.0000 774.4800 458.6000 ;
      RECT 782.3200 454.2000 796.5000 458.6000 ;
      RECT 0.0000 454.2000 10.8400 458.6000 ;
      RECT 777.2000 451.4000 796.5000 454.2000 ;
      RECT 0.0000 451.4000 15.9600 454.2000 ;
      RECT 23.8000 450.6000 769.3600 455.0000 ;
      RECT 782.3200 447.0000 796.5000 451.4000 ;
      RECT 18.6800 447.0000 774.4800 450.6000 ;
      RECT 0.0000 447.0000 10.8400 451.4000 ;
      RECT 0.0000 444.2000 796.5000 447.0000 ;
      RECT 782.3200 439.8000 796.5000 444.2000 ;
      RECT 18.6800 439.8000 774.4800 444.2000 ;
      RECT 0.0000 439.8000 10.8400 444.2000 ;
      RECT 0.0000 437.0000 796.5000 439.8000 ;
      RECT 782.3200 432.6000 796.5000 437.0000 ;
      RECT 18.6800 432.6000 774.4800 437.0000 ;
      RECT 0.0000 432.6000 10.8400 437.0000 ;
      RECT 0.0000 429.8000 796.5000 432.6000 ;
      RECT 782.3200 425.4000 796.5000 429.8000 ;
      RECT 18.6800 425.4000 774.4800 429.8000 ;
      RECT 0.0000 425.4000 10.8400 429.8000 ;
      RECT 0.0000 422.6000 796.5000 425.4000 ;
      RECT 782.3200 418.2000 796.5000 422.6000 ;
      RECT 18.6800 418.2000 774.4800 422.6000 ;
      RECT 0.0000 418.2000 10.8400 422.6000 ;
      RECT 0.0000 415.4000 796.5000 418.2000 ;
      RECT 782.3200 411.0000 796.5000 415.4000 ;
      RECT 18.6800 411.0000 774.4800 415.4000 ;
      RECT 0.0000 411.0000 10.8400 415.4000 ;
      RECT 0.0000 408.2000 796.5000 411.0000 ;
      RECT 782.3200 403.8000 796.5000 408.2000 ;
      RECT 18.6800 403.8000 774.4800 408.2000 ;
      RECT 0.0000 403.8000 10.8400 408.2000 ;
      RECT 0.0000 401.0000 796.5000 403.8000 ;
      RECT 782.3200 396.6000 796.5000 401.0000 ;
      RECT 18.6800 396.6000 774.4800 401.0000 ;
      RECT 0.0000 396.6000 10.8400 401.0000 ;
      RECT 0.0000 393.8000 796.5000 396.6000 ;
      RECT 782.3200 389.4000 796.5000 393.8000 ;
      RECT 18.6800 389.4000 774.4800 393.8000 ;
      RECT 0.0000 389.4000 10.8400 393.8000 ;
      RECT 0.0000 386.6000 796.5000 389.4000 ;
      RECT 782.3200 382.2000 796.5000 386.6000 ;
      RECT 18.6800 382.2000 774.4800 386.6000 ;
      RECT 0.0000 382.2000 10.8400 386.6000 ;
      RECT 0.0000 379.4000 796.5000 382.2000 ;
      RECT 782.3200 375.0000 796.5000 379.4000 ;
      RECT 18.6800 375.0000 774.4800 379.4000 ;
      RECT 0.0000 375.0000 10.8400 379.4000 ;
      RECT 0.0000 372.2000 796.5000 375.0000 ;
      RECT 782.3200 367.8000 796.5000 372.2000 ;
      RECT 18.6800 367.8000 774.4800 372.2000 ;
      RECT 0.0000 367.8000 10.8400 372.2000 ;
      RECT 0.0000 365.0000 796.5000 367.8000 ;
      RECT 782.3200 360.6000 796.5000 365.0000 ;
      RECT 18.6800 360.6000 774.4800 365.0000 ;
      RECT 0.0000 360.6000 10.8400 365.0000 ;
      RECT 0.0000 357.8000 796.5000 360.6000 ;
      RECT 782.3200 353.4000 796.5000 357.8000 ;
      RECT 18.6800 353.4000 774.4800 357.8000 ;
      RECT 0.0000 353.4000 10.8400 357.8000 ;
      RECT 0.0000 350.6000 796.5000 353.4000 ;
      RECT 782.3200 346.2000 796.5000 350.6000 ;
      RECT 18.6800 346.2000 774.4800 350.6000 ;
      RECT 0.0000 346.2000 10.8400 350.6000 ;
      RECT 0.0000 343.4000 796.5000 346.2000 ;
      RECT 782.3200 339.0000 796.5000 343.4000 ;
      RECT 18.6800 339.0000 774.4800 343.4000 ;
      RECT 0.0000 339.0000 10.8400 343.4000 ;
      RECT 0.0000 336.2000 796.5000 339.0000 ;
      RECT 782.3200 331.8000 796.5000 336.2000 ;
      RECT 18.6800 331.8000 774.4800 336.2000 ;
      RECT 0.0000 331.8000 10.8400 336.2000 ;
      RECT 0.0000 329.0000 796.5000 331.8000 ;
      RECT 782.3200 324.6000 796.5000 329.0000 ;
      RECT 18.6800 324.6000 774.4800 329.0000 ;
      RECT 0.0000 324.6000 10.8400 329.0000 ;
      RECT 0.0000 321.8000 796.5000 324.6000 ;
      RECT 782.3200 317.4000 796.5000 321.8000 ;
      RECT 18.6800 317.4000 774.4800 321.8000 ;
      RECT 0.0000 317.4000 10.8400 321.8000 ;
      RECT 0.0000 314.6000 796.5000 317.4000 ;
      RECT 782.3200 310.2000 796.5000 314.6000 ;
      RECT 18.6800 310.2000 774.4800 314.6000 ;
      RECT 0.0000 310.2000 10.8400 314.6000 ;
      RECT 0.0000 307.4000 796.5000 310.2000 ;
      RECT 782.3200 303.0000 796.5000 307.4000 ;
      RECT 18.6800 303.0000 774.4800 307.4000 ;
      RECT 0.0000 303.0000 10.8400 307.4000 ;
      RECT 0.0000 300.2000 796.5000 303.0000 ;
      RECT 782.3200 295.8000 796.5000 300.2000 ;
      RECT 18.6800 295.8000 774.4800 300.2000 ;
      RECT 0.0000 295.8000 10.8400 300.2000 ;
      RECT 0.0000 293.0000 796.5000 295.8000 ;
      RECT 782.3200 288.6000 796.5000 293.0000 ;
      RECT 18.6800 288.6000 774.4800 293.0000 ;
      RECT 0.0000 288.6000 10.8400 293.0000 ;
      RECT 0.0000 285.8000 796.5000 288.6000 ;
      RECT 782.3200 281.4000 796.5000 285.8000 ;
      RECT 18.6800 281.4000 774.4800 285.8000 ;
      RECT 0.0000 281.4000 10.8400 285.8000 ;
      RECT 0.0000 278.6000 796.5000 281.4000 ;
      RECT 782.3200 274.2000 796.5000 278.6000 ;
      RECT 18.6800 274.2000 774.4800 278.6000 ;
      RECT 0.0000 274.2000 10.8400 278.6000 ;
      RECT 0.0000 271.4000 796.5000 274.2000 ;
      RECT 782.3200 267.0000 796.5000 271.4000 ;
      RECT 18.6800 267.0000 774.4800 271.4000 ;
      RECT 0.0000 267.0000 10.8400 271.4000 ;
      RECT 0.0000 264.2000 796.5000 267.0000 ;
      RECT 782.3200 259.8000 796.5000 264.2000 ;
      RECT 18.6800 259.8000 774.4800 264.2000 ;
      RECT 0.0000 259.8000 10.8400 264.2000 ;
      RECT 0.0000 257.0000 796.5000 259.8000 ;
      RECT 782.3200 252.6000 796.5000 257.0000 ;
      RECT 18.6800 252.6000 774.4800 257.0000 ;
      RECT 0.0000 252.6000 10.8400 257.0000 ;
      RECT 0.0000 249.8000 796.5000 252.6000 ;
      RECT 782.3200 245.4000 796.5000 249.8000 ;
      RECT 18.6800 245.4000 774.4800 249.8000 ;
      RECT 0.0000 245.4000 10.8400 249.8000 ;
      RECT 0.0000 242.6000 796.5000 245.4000 ;
      RECT 18.6800 239.0000 774.4800 242.6000 ;
      RECT 782.3200 238.2000 796.5000 242.6000 ;
      RECT 0.0000 238.2000 10.8400 242.6000 ;
      RECT 777.2000 235.4000 796.5000 238.2000 ;
      RECT 0.0000 235.4000 15.9600 238.2000 ;
      RECT 23.8000 234.6000 769.3600 239.0000 ;
      RECT 782.3200 231.0000 796.5000 235.4000 ;
      RECT 18.6800 231.0000 774.4800 234.6000 ;
      RECT 0.0000 231.0000 10.8400 235.4000 ;
      RECT 0.0000 228.2000 796.5000 231.0000 ;
      RECT 782.3200 223.8000 796.5000 228.2000 ;
      RECT 18.6800 223.8000 774.4800 228.2000 ;
      RECT 0.0000 223.8000 10.8400 228.2000 ;
      RECT 0.0000 221.0000 796.5000 223.8000 ;
      RECT 782.3200 216.6000 796.5000 221.0000 ;
      RECT 18.6800 216.6000 774.4800 221.0000 ;
      RECT 0.0000 216.6000 10.8400 221.0000 ;
      RECT 0.0000 213.8000 796.5000 216.6000 ;
      RECT 782.3200 209.4000 796.5000 213.8000 ;
      RECT 18.6800 209.4000 774.4800 213.8000 ;
      RECT 0.0000 209.4000 10.8400 213.8000 ;
      RECT 0.0000 206.6000 796.5000 209.4000 ;
      RECT 782.3200 202.2000 796.5000 206.6000 ;
      RECT 18.6800 202.2000 774.4800 206.6000 ;
      RECT 0.0000 202.2000 10.8400 206.6000 ;
      RECT 0.0000 199.4000 796.5000 202.2000 ;
      RECT 782.3200 195.0000 796.5000 199.4000 ;
      RECT 18.6800 195.0000 774.4800 199.4000 ;
      RECT 0.0000 195.0000 10.8400 199.4000 ;
      RECT 0.0000 192.2000 796.5000 195.0000 ;
      RECT 782.3200 187.8000 796.5000 192.2000 ;
      RECT 18.6800 187.8000 774.4800 192.2000 ;
      RECT 0.0000 187.8000 10.8400 192.2000 ;
      RECT 0.0000 185.0000 796.5000 187.8000 ;
      RECT 782.3200 180.6000 796.5000 185.0000 ;
      RECT 18.6800 180.6000 774.4800 185.0000 ;
      RECT 0.0000 180.6000 10.8400 185.0000 ;
      RECT 0.0000 177.8000 796.5000 180.6000 ;
      RECT 782.3200 173.4000 796.5000 177.8000 ;
      RECT 18.6800 173.4000 774.4800 177.8000 ;
      RECT 0.0000 173.4000 10.8400 177.8000 ;
      RECT 0.0000 170.6000 796.5000 173.4000 ;
      RECT 782.3200 166.2000 796.5000 170.6000 ;
      RECT 18.6800 166.2000 774.4800 170.6000 ;
      RECT 0.0000 166.2000 10.8400 170.6000 ;
      RECT 0.0000 163.4000 796.5000 166.2000 ;
      RECT 782.3200 159.0000 796.5000 163.4000 ;
      RECT 18.6800 159.0000 774.4800 163.4000 ;
      RECT 0.0000 159.0000 10.8400 163.4000 ;
      RECT 0.0000 156.2000 796.5000 159.0000 ;
      RECT 782.3200 151.8000 796.5000 156.2000 ;
      RECT 18.6800 151.8000 774.4800 156.2000 ;
      RECT 0.0000 151.8000 10.8400 156.2000 ;
      RECT 0.0000 149.0000 796.5000 151.8000 ;
      RECT 782.3200 144.6000 796.5000 149.0000 ;
      RECT 18.6800 144.6000 774.4800 149.0000 ;
      RECT 0.0000 144.6000 10.8400 149.0000 ;
      RECT 0.0000 141.8000 796.5000 144.6000 ;
      RECT 782.3200 137.4000 796.5000 141.8000 ;
      RECT 18.6800 137.4000 774.4800 141.8000 ;
      RECT 0.0000 137.4000 10.8400 141.8000 ;
      RECT 0.0000 134.6000 796.5000 137.4000 ;
      RECT 782.3200 130.2000 796.5000 134.6000 ;
      RECT 18.6800 130.2000 774.4800 134.6000 ;
      RECT 0.0000 130.2000 10.8400 134.6000 ;
      RECT 0.0000 127.4000 796.5000 130.2000 ;
      RECT 782.3200 123.0000 796.5000 127.4000 ;
      RECT 18.6800 123.0000 774.4800 127.4000 ;
      RECT 0.0000 123.0000 10.8400 127.4000 ;
      RECT 0.0000 120.2000 796.5000 123.0000 ;
      RECT 782.3200 115.8000 796.5000 120.2000 ;
      RECT 18.6800 115.8000 774.4800 120.2000 ;
      RECT 0.0000 115.8000 10.8400 120.2000 ;
      RECT 0.0000 113.0000 796.5000 115.8000 ;
      RECT 782.3200 108.6000 796.5000 113.0000 ;
      RECT 18.6800 108.6000 774.4800 113.0000 ;
      RECT 0.0000 108.6000 10.8400 113.0000 ;
      RECT 0.0000 105.8000 796.5000 108.6000 ;
      RECT 782.3200 101.4000 796.5000 105.8000 ;
      RECT 18.6800 101.4000 774.4800 105.8000 ;
      RECT 0.0000 101.4000 10.8400 105.8000 ;
      RECT 0.0000 98.6000 796.5000 101.4000 ;
      RECT 782.3200 94.2000 796.5000 98.6000 ;
      RECT 18.6800 94.2000 774.4800 98.6000 ;
      RECT 0.0000 94.2000 10.8400 98.6000 ;
      RECT 0.0000 91.4000 796.5000 94.2000 ;
      RECT 18.6800 87.8000 774.4800 91.4000 ;
      RECT 782.3200 87.0000 796.5000 91.4000 ;
      RECT 0.0000 87.0000 10.8400 91.4000 ;
      RECT 777.2000 83.4000 796.5000 87.0000 ;
      RECT 23.8000 83.4000 769.3600 87.8000 ;
      RECT 0.0000 83.4000 15.9600 87.0000 ;
      RECT 0.0000 80.6000 796.5000 83.4000 ;
      RECT 777.2000 77.0000 796.5000 80.6000 ;
      RECT 0.0000 77.0000 15.9600 80.6000 ;
      RECT 23.8000 76.2000 769.3600 80.6000 ;
      RECT 18.6800 73.4000 774.4800 76.2000 ;
      RECT 782.3200 72.6000 796.5000 77.0000 ;
      RECT 0.0000 72.6000 10.8400 77.0000 ;
      RECT 777.2000 69.8000 796.5000 72.6000 ;
      RECT 0.0000 69.8000 15.9600 72.6000 ;
      RECT 23.8000 69.0000 769.3600 73.4000 ;
      RECT 18.6800 66.2000 774.4800 69.0000 ;
      RECT 782.3200 65.4000 796.5000 69.8000 ;
      RECT 0.0000 65.4000 10.8400 69.8000 ;
      RECT 777.2000 62.6000 796.5000 65.4000 ;
      RECT 0.0000 62.6000 15.9600 65.4000 ;
      RECT 23.8000 61.8000 769.3600 66.2000 ;
      RECT 782.3200 58.2000 796.5000 62.6000 ;
      RECT 18.6800 58.2000 774.4800 61.8000 ;
      RECT 0.0000 58.2000 10.8400 62.6000 ;
      RECT 0.0000 55.4000 796.5000 58.2000 ;
      RECT 782.3200 51.0000 796.5000 55.4000 ;
      RECT 18.6800 51.0000 774.4800 55.4000 ;
      RECT 0.0000 51.0000 10.8400 55.4000 ;
      RECT 0.0000 48.2000 796.5000 51.0000 ;
      RECT 18.6800 44.4900 774.4800 48.2000 ;
      RECT 782.3200 43.8000 796.5000 48.2000 ;
      RECT 0.0000 43.8000 10.8400 48.2000 ;
      RECT 777.2000 41.0000 796.5000 43.8000 ;
      RECT 0.0000 41.0000 15.9600 43.8000 ;
      RECT 23.8000 40.2000 769.3600 44.4900 ;
      RECT 18.6800 37.4000 774.4800 40.2000 ;
      RECT 782.3200 36.6000 796.5000 41.0000 ;
      RECT 0.0000 36.6000 10.8400 41.0000 ;
      RECT 777.2000 33.8000 796.5000 36.6000 ;
      RECT 0.0000 33.8000 15.9600 36.6000 ;
      RECT 23.8000 33.0000 769.3600 37.4000 ;
      RECT 18.6800 30.2000 774.4800 33.0000 ;
      RECT 782.3200 29.4000 796.5000 33.8000 ;
      RECT 0.0000 29.4000 10.8400 33.8000 ;
      RECT 777.2000 25.8000 796.5000 29.4000 ;
      RECT 23.8000 25.8000 769.3600 30.2000 ;
      RECT 0.0000 25.8000 15.9600 29.4000 ;
      RECT 0.0000 19.4000 796.5000 25.8000 ;
      RECT 0.0000 17.3100 774.4800 19.4000 ;
      RECT 782.3200 15.0000 796.5000 19.4000 ;
      RECT 24.4200 15.0000 774.4800 17.3100 ;
      RECT 24.4200 4.0800 796.5000 15.0000 ;
      RECT 0.0000 4.0800 16.5800 17.3100 ;
      RECT 0.0000 0.0000 796.5000 4.0800 ;
  END
END cacheBank

END LIBRARY
