
module cacheAccessArbiter ( clk, reset, cacheAddressIn_NORTH, 
        requesterAddressIn_NORTH, memRead_NORTH, memWrite_NORTH, dataIn_NORTH, 
        readReady_NORTH, requesterAddressOut_NORTH, cacheDataOut_NORTH, 
        cacheAddressIn_SOUTH, requesterAddressIn_SOUTH, memRead_SOUTH, 
        memWrite_SOUTH, dataIn_SOUTH, readReady_SOUTH, 
        requesterAddressOut_SOUTH, cacheDataOut_SOUTH, cacheAddressIn_EAST, 
        requesterAddressIn_EAST, memRead_EAST, memWrite_EAST, dataIn_EAST, 
        readReady_EAST, requesterAddressOut_EAST, cacheDataOut_EAST, 
        cacheAddressIn_WEST, requesterAddressIn_WEST, memRead_WEST, 
        memWrite_WEST, dataIn_WEST, readReady_WEST, requesterAddressOut_WEST, 
        cacheDataOut_WEST, cacheDataIn_A, cacheAddressIn_A, cacheDataOut_A, 
        memWrite_A, cacheDataIn_B, cacheAddressIn_B, cacheDataOut_B, 
        memWrite_B );
  input [7:0] cacheAddressIn_NORTH;
  input [5:0] requesterAddressIn_NORTH;
  input [31:0] dataIn_NORTH;
  output [5:0] requesterAddressOut_NORTH;
  output [31:0] cacheDataOut_NORTH;
  input [7:0] cacheAddressIn_SOUTH;
  input [5:0] requesterAddressIn_SOUTH;
  input [31:0] dataIn_SOUTH;
  output [5:0] requesterAddressOut_SOUTH;
  output [31:0] cacheDataOut_SOUTH;
  input [7:0] cacheAddressIn_EAST;
  input [5:0] requesterAddressIn_EAST;
  input [31:0] dataIn_EAST;
  output [5:0] requesterAddressOut_EAST;
  output [31:0] cacheDataOut_EAST;
  input [7:0] cacheAddressIn_WEST;
  input [5:0] requesterAddressIn_WEST;
  input [31:0] dataIn_WEST;
  output [5:0] requesterAddressOut_WEST;
  output [31:0] cacheDataOut_WEST;
  output [31:0] cacheDataIn_A;
  output [7:0] cacheAddressIn_A;
  input [31:0] cacheDataOut_A;
  output [31:0] cacheDataIn_B;
  output [7:0] cacheAddressIn_B;
  input [31:0] cacheDataOut_B;
  input clk, reset, memRead_NORTH, memWrite_NORTH, memRead_SOUTH,
         memWrite_SOUTH, memRead_EAST, memWrite_EAST, memRead_WEST,
         memWrite_WEST;
  output readReady_NORTH, readReady_SOUTH, readReady_EAST, readReady_WEST,
         memWrite_A, memWrite_B;
  wire   N589, \indexIncrementer_EAST[1] , N605, N606, N607, N608, N609, N610,
         N615, N616, N617, N650, N651, N6314, N6316, N6318, N6371, N6372,
         N6373, N6374, N6375, N6618, N6619, N6620, N6621, N6622, N6699, N6701,
         N8209, \dataToWriteBuffer[2][31] , \dataToWriteBuffer[2][30] ,
         \dataToWriteBuffer[2][29] , \dataToWriteBuffer[2][28] ,
         \dataToWriteBuffer[2][27] , \dataToWriteBuffer[2][26] ,
         \dataToWriteBuffer[2][25] , \dataToWriteBuffer[2][24] ,
         \dataToWriteBuffer[2][23] , \dataToWriteBuffer[2][22] ,
         \dataToWriteBuffer[2][21] , \dataToWriteBuffer[2][20] ,
         \dataToWriteBuffer[2][19] , \dataToWriteBuffer[2][18] ,
         \dataToWriteBuffer[2][17] , \dataToWriteBuffer[2][16] ,
         \dataToWriteBuffer[2][15] , \dataToWriteBuffer[2][14] ,
         \dataToWriteBuffer[2][13] , \dataToWriteBuffer[2][12] ,
         \dataToWriteBuffer[2][11] , \dataToWriteBuffer[2][10] ,
         \dataToWriteBuffer[2][9] , \dataToWriteBuffer[2][8] ,
         \dataToWriteBuffer[2][7] , \dataToWriteBuffer[2][6] ,
         \dataToWriteBuffer[2][5] , \dataToWriteBuffer[2][4] ,
         \dataToWriteBuffer[2][3] , \dataToWriteBuffer[2][2] ,
         \dataToWriteBuffer[2][1] , \dataToWriteBuffer[2][0] ,
         \dataToWriteBuffer[0][31] , \dataToWriteBuffer[0][30] ,
         \dataToWriteBuffer[0][29] , \dataToWriteBuffer[0][28] ,
         \dataToWriteBuffer[0][27] , \dataToWriteBuffer[0][26] ,
         \dataToWriteBuffer[0][25] , \dataToWriteBuffer[0][24] ,
         \dataToWriteBuffer[0][23] , \dataToWriteBuffer[0][22] ,
         \dataToWriteBuffer[0][21] , \dataToWriteBuffer[0][20] ,
         \dataToWriteBuffer[0][19] , \dataToWriteBuffer[0][18] ,
         \dataToWriteBuffer[0][17] , \dataToWriteBuffer[0][16] ,
         \dataToWriteBuffer[0][15] , \dataToWriteBuffer[0][14] ,
         \dataToWriteBuffer[0][13] , \dataToWriteBuffer[0][12] ,
         \dataToWriteBuffer[0][11] , \dataToWriteBuffer[0][10] ,
         \dataToWriteBuffer[0][9] , \dataToWriteBuffer[0][8] ,
         \dataToWriteBuffer[0][7] , \dataToWriteBuffer[0][6] ,
         \dataToWriteBuffer[0][5] , \dataToWriteBuffer[0][4] ,
         \dataToWriteBuffer[0][3] , \dataToWriteBuffer[0][2] ,
         \dataToWriteBuffer[0][1] , \dataToWriteBuffer[0][0] ,
         \addressToWriteBuffer[2][7] , \addressToWriteBuffer[2][6] ,
         \addressToWriteBuffer[2][5] , \addressToWriteBuffer[2][4] ,
         \addressToWriteBuffer[2][3] , \addressToWriteBuffer[2][2] ,
         \addressToWriteBuffer[2][1] , \addressToWriteBuffer[2][0] ,
         \addressToWriteBuffer[0][7] , \addressToWriteBuffer[0][6] ,
         \addressToWriteBuffer[0][5] , \addressToWriteBuffer[0][4] ,
         \addressToWriteBuffer[0][3] , \addressToWriteBuffer[0][2] ,
         \addressToWriteBuffer[0][1] , \addressToWriteBuffer[0][0] ,
         \requesterAddressBuffer[0][5] , \requesterAddressBuffer[0][4] ,
         \requesterAddressBuffer[0][3] , \requesterAddressBuffer[0][2] ,
         \requesterAddressBuffer[0][1] , \requesterAddressBuffer[0][0] ,
         \requesterPortBuffer[7][1] , \requesterPortBuffer[7][0] ,
         \requesterPortBuffer[6][1] , \requesterPortBuffer[6][0] ,
         \requesterPortBuffer[5][1] , \requesterPortBuffer[5][0] ,
         \requesterPortBuffer[4][1] , \requesterPortBuffer[4][0] ,
         \requesterPortBuffer[2][0] , \requesterPortBuffer[0][1] ,
         \requesterPortBuffer[0][0] , N10004, prevMemRead_B, prevMemRead_A,
         N10076, N10077, N10078, N10079, N10087, N10088, N10089, N10090,
         N10091, N10092, N10093, N10094, N10095, N10096, N10097, N10098,
         N10099, N10100, N10101, N10102, N10103, N10104, N10105, N10106,
         N10107, N10108, N10109, N10110, N10111, N10112, N10113, N10114,
         N10115, N10116, N10117, N10118, N10121, N10122, N10123, N10124,
         N10125, N10126, N10127, N10128, N10129, N10130, N10131, N10132,
         N10133, N10134, N10135, N10136, N10137, N10138, N10139, N10140,
         N10141, N10142, N10143, N10144, N10145, N10146, N10147, N10148,
         N10149, N10150, N10151, N10152, N10155, N10156, N10157, N10158,
         N10159, N10160, N10161, N10162, N10163, N10164, N10165, N10166,
         N10167, N10168, N10169, N10170, N10171, N10172, N10173, N10174,
         N10175, N10176, N10177, N10178, N10179, N10180, N10181, N10182,
         N10183, N10184, N10185, N10186, N10189, N10190, N10191, N10192,
         N10193, N10194, N10195, N10196, N10197, N10198, N10199, N10200,
         N10201, N10202, N10203, N10204, N10205, N10206, N10207, N10208,
         N10209, N10210, N10211, N10212, N10213, N10214, N10215, N10216,
         N10217, N10218, N10219, N10220, n880, n910, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1571, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1588, n1589, n1590, n1592, n1593, n1594, n1595, n1596,
         n1598, n1599, n1600, n1601, n1603, n1604, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1618, n1619, n1620,
         n1621, n1622, n1624, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1830, n1831, n1832, n1834, n1835, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1875, n1876, n1877, n1879, n1880,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1919, n1920, n1921, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1964, n1965,
         n1966, n1968, n1969, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
         n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
         n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
         n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2008,
         n2009, n2010, n2012, n2013, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2252, n2253, n2255, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, N614, \add_0_root_sub_278_I2/B[2] ,
         \add_0_root_sub_278_I2/A[0] , \r1472/carry[3] , \r1471/carry[3] ,
         \r1470/carry[3] , \r1467/carry[3] , \add_0_root_r1463/SUM[0] ,
         \add_0_root_r1463/SUM[1] , \add_0_root_r1463/SUM[2] ,
         \add_0_root_r1463/SUM[3] , \add_0_root_r1463/SUM[4] ,
         \add_0_root_r1463/B[4] , \add_0_root_r1459/SUM[0] ,
         \add_0_root_r1459/SUM[1] , \add_0_root_r1459/SUM[2] ,
         \add_0_root_r1459/SUM[3] , \add_0_root_r1459/SUM[4] ,
         \add_0_root_r1459/B[0] , \add_0_root_r1459/B[4] ,
         \add_0_root_sub_0_root_sub_231/B[2] , n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981;
  wire   [2:0] totalAccesses;
  wire   [7:0] isWrite;
  wire   [1:0] prevRequesterPort_B;
  wire   [5:0] prevRequesterAddress_B;
  wire   [5:0] prevRequesterAddress_A;
  wire   [4:1] \add_0_root_sub_278_I2/carry ;
  wire   [4:1] \add_0_root_sub_277_I2/carry ;
  wire   [4:1] \add_0_root_r1463/carry ;
  wire   [4:1] \add_0_root_r1459/carry ;
  wire   [4:1] \add_0_root_sub_0_root_sub_231/carry ;

  DFFNSRX2TS \isRead_reg[1]  ( .D(n3345), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .QN(n1175) );
  DFFNSRX2TS \isRead_reg[0]  ( .D(n3343), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .QN(n1176) );
  DFFNSRX2TS \dataToWriteBuffer_reg[2][31]  ( .D(n3546), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[2][31] ), .QN(n1072) );
  DFFNSRX2TS \dataToWriteBuffer_reg[2][30]  ( .D(n3547), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[2][30] ), .QN(n1073) );
  DFFNSRX2TS \dataToWriteBuffer_reg[2][29]  ( .D(n3548), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[2][29] ), .QN(n1074) );
  DFFNSRX2TS \dataToWriteBuffer_reg[2][28]  ( .D(n3549), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[2][28] ), .QN(n1075) );
  DFFNSRX2TS \dataToWriteBuffer_reg[2][27]  ( .D(n3550), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[2][27] ), .QN(n1076) );
  DFFNSRX2TS \dataToWriteBuffer_reg[2][26]  ( .D(n3551), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[2][26] ), .QN(n1077) );
  DFFNSRX2TS \dataToWriteBuffer_reg[2][25]  ( .D(n3552), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[2][25] ), .QN(n1078) );
  DFFNSRX2TS \dataToWriteBuffer_reg[2][24]  ( .D(n3553), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[2][24] ), .QN(n1079) );
  DFFNSRX2TS \dataToWriteBuffer_reg[2][23]  ( .D(n3554), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[2][23] ), .QN(n1080) );
  DFFNSRX2TS \dataToWriteBuffer_reg[2][22]  ( .D(n3555), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[2][22] ), .QN(n1081) );
  DFFNSRX2TS \dataToWriteBuffer_reg[2][21]  ( .D(n3556), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[2][21] ), .QN(n1082) );
  DFFNSRX2TS \dataToWriteBuffer_reg[2][20]  ( .D(n3557), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[2][20] ), .QN(n1083) );
  DFFNSRX2TS \dataToWriteBuffer_reg[2][19]  ( .D(n3558), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[2][19] ), .QN(n1084) );
  DFFNSRX2TS \dataToWriteBuffer_reg[2][18]  ( .D(n3559), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[2][18] ), .QN(n1085) );
  DFFNSRX2TS \dataToWriteBuffer_reg[2][17]  ( .D(n3560), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[2][17] ), .QN(n1086) );
  DFFNSRX2TS \dataToWriteBuffer_reg[2][16]  ( .D(n3561), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[2][16] ), .QN(n1087) );
  DFFNSRX2TS \dataToWriteBuffer_reg[2][15]  ( .D(n3562), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[2][15] ), .QN(n1088) );
  DFFNSRX2TS \dataToWriteBuffer_reg[2][14]  ( .D(n3563), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[2][14] ), .QN(n1089) );
  DFFNSRX2TS \dataToWriteBuffer_reg[2][13]  ( .D(n3564), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[2][13] ), .QN(n1090) );
  DFFNSRX2TS \dataToWriteBuffer_reg[2][12]  ( .D(n3565), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[2][12] ), .QN(n1091) );
  DFFNSRX2TS \dataToWriteBuffer_reg[2][11]  ( .D(n3566), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[2][11] ), .QN(n1092) );
  DFFNSRX2TS \dataToWriteBuffer_reg[2][10]  ( .D(n3567), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[2][10] ), .QN(n1093) );
  DFFNSRX2TS \dataToWriteBuffer_reg[2][9]  ( .D(n3568), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[2][9] ), .QN(n1094) );
  DFFNSRX2TS \dataToWriteBuffer_reg[2][8]  ( .D(n3569), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[2][8] ), .QN(n1095) );
  DFFNSRX2TS \dataToWriteBuffer_reg[2][7]  ( .D(n3570), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[2][7] ), .QN(n1096) );
  DFFNSRX2TS \dataToWriteBuffer_reg[2][6]  ( .D(n3571), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[2][6] ), .QN(n1097) );
  DFFNSRX2TS \dataToWriteBuffer_reg[2][5]  ( .D(n3572), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[2][5] ), .QN(n1098) );
  DFFNSRX2TS \dataToWriteBuffer_reg[2][4]  ( .D(n3573), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[2][4] ), .QN(n1099) );
  DFFNSRX2TS \dataToWriteBuffer_reg[2][3]  ( .D(n3574), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[2][3] ), .QN(n1100) );
  DFFNSRX2TS \dataToWriteBuffer_reg[2][2]  ( .D(n3575), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[2][2] ), .QN(n1101) );
  DFFNSRX2TS \dataToWriteBuffer_reg[2][1]  ( .D(n3576), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[2][1] ), .QN(n1102) );
  DFFNSRX2TS \dataToWriteBuffer_reg[2][0]  ( .D(n3577), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[2][0] ), .QN(n1103) );
  DFFNSRX2TS \requesterPortBuffer_reg[7][0]  ( .D(n3253), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[7][0] ) );
  DFFNSRX2TS \requesterPortBuffer_reg[1][1]  ( .D(n3266), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1261) );
  DFFNSRX2TS \dataToWriteBuffer_reg[1][31]  ( .D(n3578), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1104) );
  DFFNSRX2TS \dataToWriteBuffer_reg[1][30]  ( .D(n3579), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1105) );
  DFFNSRX2TS \dataToWriteBuffer_reg[1][29]  ( .D(n3580), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1106) );
  DFFNSRX2TS \dataToWriteBuffer_reg[1][28]  ( .D(n3581), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1107) );
  DFFNSRX2TS \dataToWriteBuffer_reg[1][27]  ( .D(n3582), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1108) );
  DFFNSRX2TS \dataToWriteBuffer_reg[1][26]  ( .D(n3583), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1109) );
  DFFNSRX2TS \dataToWriteBuffer_reg[1][25]  ( .D(n3584), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1110) );
  DFFNSRX2TS \dataToWriteBuffer_reg[1][24]  ( .D(n3585), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1111) );
  DFFNSRX2TS \dataToWriteBuffer_reg[1][23]  ( .D(n3586), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1112) );
  DFFNSRX2TS \dataToWriteBuffer_reg[1][22]  ( .D(n3587), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1113) );
  DFFNSRX2TS \dataToWriteBuffer_reg[1][21]  ( .D(n3588), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1114) );
  DFFNSRX2TS \dataToWriteBuffer_reg[1][20]  ( .D(n3589), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1115) );
  DFFNSRX2TS \dataToWriteBuffer_reg[1][19]  ( .D(n3590), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1116) );
  DFFNSRX2TS \dataToWriteBuffer_reg[1][18]  ( .D(n3591), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1117) );
  DFFNSRX2TS \dataToWriteBuffer_reg[1][17]  ( .D(n3592), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1118) );
  DFFNSRX2TS \dataToWriteBuffer_reg[1][16]  ( .D(n3593), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1119) );
  DFFNSRX2TS \dataToWriteBuffer_reg[1][15]  ( .D(n3594), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1120) );
  DFFNSRX2TS \dataToWriteBuffer_reg[1][14]  ( .D(n3595), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1121) );
  DFFNSRX2TS \dataToWriteBuffer_reg[1][13]  ( .D(n3596), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1122) );
  DFFNSRX2TS \dataToWriteBuffer_reg[1][12]  ( .D(n3597), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1123) );
  DFFNSRX2TS \dataToWriteBuffer_reg[1][11]  ( .D(n3598), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1124) );
  DFFNSRX2TS \dataToWriteBuffer_reg[1][10]  ( .D(n3599), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1125) );
  DFFNSRX2TS \dataToWriteBuffer_reg[1][9]  ( .D(n3600), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1126) );
  DFFNSRX2TS \dataToWriteBuffer_reg[1][8]  ( .D(n3601), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1127) );
  DFFNSRX2TS \dataToWriteBuffer_reg[1][7]  ( .D(n3602), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1128) );
  DFFNSRX2TS \dataToWriteBuffer_reg[1][6]  ( .D(n3603), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1129) );
  DFFNSRX2TS \dataToWriteBuffer_reg[1][5]  ( .D(n3604), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1130) );
  DFFNSRX2TS \dataToWriteBuffer_reg[1][4]  ( .D(n3605), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1131) );
  DFFNSRX2TS \dataToWriteBuffer_reg[1][3]  ( .D(n3606), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1132) );
  DFFNSRX2TS \dataToWriteBuffer_reg[1][2]  ( .D(n3607), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1133) );
  DFFNSRX2TS \dataToWriteBuffer_reg[1][1]  ( .D(n3608), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1134) );
  DFFNSRX2TS \dataToWriteBuffer_reg[1][0]  ( .D(n3609), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1135) );
  DFFNSRX2TS \addressToWriteBuffer_reg[1][7]  ( .D(n3326), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1225) );
  DFFNSRX2TS \addressToWriteBuffer_reg[1][6]  ( .D(n3327), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1226) );
  DFFNSRX2TS \addressToWriteBuffer_reg[1][5]  ( .D(n3328), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1227) );
  DFFNSRX2TS \addressToWriteBuffer_reg[1][4]  ( .D(n3329), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1228) );
  DFFNSRX2TS \addressToWriteBuffer_reg[1][3]  ( .D(n3330), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1229) );
  DFFNSRX2TS \addressToWriteBuffer_reg[1][2]  ( .D(n3331), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1230) );
  DFFNSRX2TS \addressToWriteBuffer_reg[1][1]  ( .D(n3332), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1231) );
  DFFNSRX2TS \addressToWriteBuffer_reg[1][0]  ( .D(n3333), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1232) );
  DFFNSRX2TS \requesterAddressBuffer_reg[1][5]  ( .D(n3208), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n1273) );
  DFFNSRX2TS \requesterAddressBuffer_reg[1][4]  ( .D(n3207), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n1274) );
  DFFNSRX2TS \requesterAddressBuffer_reg[1][3]  ( .D(n3206), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n1275) );
  DFFNSRX2TS \requesterAddressBuffer_reg[1][2]  ( .D(n3205), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n1276) );
  DFFNSRX2TS \requesterAddressBuffer_reg[1][1]  ( .D(n3204), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n1277) );
  DFFNSRX2TS \requesterAddressBuffer_reg[1][0]  ( .D(n3203), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n1278) );
  DFFNSRX2TS \requesterPortBuffer_reg[0][0]  ( .D(n3269), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[0][0] ) );
  DFFNSRX2TS \requesterPortBuffer_reg[0][1]  ( .D(n3268), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[0][1] ) );
  DFFNSRX2TS \isWrite_reg[3]  ( .D(n3382), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(isWrite[3]), .QN(n1171) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][31]  ( .D(n3386), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n912) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][30]  ( .D(n3387), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n913) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][29]  ( .D(n3388), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n914) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][28]  ( .D(n3389), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n915) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][27]  ( .D(n3390), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n916) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][26]  ( .D(n3391), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n917) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][25]  ( .D(n3392), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n918) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][24]  ( .D(n3393), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n919) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][23]  ( .D(n3394), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n920) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][22]  ( .D(n3395), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n921) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][21]  ( .D(n3396), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n922) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][20]  ( .D(n3397), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n923) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][19]  ( .D(n3398), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n924) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][18]  ( .D(n3399), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n925) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][17]  ( .D(n3400), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n926) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][16]  ( .D(n3401), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n927) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][15]  ( .D(n3402), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n928) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][14]  ( .D(n3403), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n929) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][13]  ( .D(n3404), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n930) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][12]  ( .D(n3405), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n931) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][11]  ( .D(n3406), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n932) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][10]  ( .D(n3407), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n933) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][9]  ( .D(n3408), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n934) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][8]  ( .D(n3409), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n935) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][7]  ( .D(n3410), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n936) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][6]  ( .D(n3411), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n937) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][5]  ( .D(n3412), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n938) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][4]  ( .D(n3413), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n939) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][3]  ( .D(n3414), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n940) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][2]  ( .D(n3415), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n941) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][1]  ( .D(n3416), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n942) );
  DFFNSRX2TS \dataToWriteBuffer_reg[7][0]  ( .D(n3417), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n943) );
  DFFNSRX2TS \requesterPortBuffer_reg[3][0]  ( .D(n3261), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1258) );
  DFFNSRX2TS \addressToWriteBuffer_reg[7][7]  ( .D(n3278), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1177) );
  DFFNSRX2TS \addressToWriteBuffer_reg[7][6]  ( .D(n3279), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1178) );
  DFFNSRX2TS \addressToWriteBuffer_reg[7][5]  ( .D(n3280), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1179) );
  DFFNSRX2TS \addressToWriteBuffer_reg[7][4]  ( .D(n3281), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1180) );
  DFFNSRX2TS \addressToWriteBuffer_reg[7][3]  ( .D(n3282), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1181) );
  DFFNSRX2TS \addressToWriteBuffer_reg[7][2]  ( .D(n3283), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1182) );
  DFFNSRX2TS \addressToWriteBuffer_reg[7][1]  ( .D(n3284), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1183) );
  DFFNSRX2TS \addressToWriteBuffer_reg[7][0]  ( .D(n3285), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1184) );
  DFFNSRX2TS \requesterPortBuffer_reg[2][1]  ( .D(n3262), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1259) );
  DFFNSRX2TS \isWrite_reg[7]  ( .D(n3378), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(isWrite[7]) );
  DFFNSRX2TS \requesterPortBuffer_reg[1][0]  ( .D(n3267), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1262) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][31]  ( .D(n3450), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n976) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][30]  ( .D(n3451), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n977) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][29]  ( .D(n3452), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n978) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][28]  ( .D(n3453), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n979) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][27]  ( .D(n3454), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n980) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][26]  ( .D(n3455), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n981) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][25]  ( .D(n3456), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n982) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][24]  ( .D(n3457), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n983) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][23]  ( .D(n3458), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n984) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][22]  ( .D(n3459), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n985) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][21]  ( .D(n3460), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n986) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][20]  ( .D(n3461), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n987) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][19]  ( .D(n3462), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n988) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][18]  ( .D(n3463), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n989) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][17]  ( .D(n3464), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n990) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][16]  ( .D(n3465), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n991) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][15]  ( .D(n3466), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n992) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][14]  ( .D(n3467), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n993) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][13]  ( .D(n3468), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n994) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][12]  ( .D(n3469), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n995) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][11]  ( .D(n3470), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n996) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][10]  ( .D(n3471), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n997) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][9]  ( .D(n3472), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n998) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][8]  ( .D(n3473), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n999) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][7]  ( .D(n3474), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1000) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][6]  ( .D(n3475), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1001) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][5]  ( .D(n3476), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1002) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][4]  ( .D(n3477), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1003) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][3]  ( .D(n3478), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1004) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][2]  ( .D(n3479), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1005) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][1]  ( .D(n3480), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1006) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][0]  ( .D(n3481), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1007) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][31]  ( .D(n3418), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n944) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][31]  ( .D(n3482), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1008) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][30]  ( .D(n3419), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n945) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][30]  ( .D(n3483), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1009) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][29]  ( .D(n3420), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n946) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][29]  ( .D(n3484), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1010) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][28]  ( .D(n3421), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n947) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][28]  ( .D(n3485), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1011) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][27]  ( .D(n3422), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n948) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][27]  ( .D(n3486), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1012) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][26]  ( .D(n3423), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n949) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][26]  ( .D(n3487), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1013) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][25]  ( .D(n3424), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n950) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][25]  ( .D(n3488), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1014) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][24]  ( .D(n3425), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n951) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][24]  ( .D(n3489), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1015) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][23]  ( .D(n3426), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n952) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][23]  ( .D(n3490), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1016) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][22]  ( .D(n3427), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n953) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][22]  ( .D(n3491), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1017) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][21]  ( .D(n3428), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n954) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][21]  ( .D(n3492), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1018) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][20]  ( .D(n3429), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n955) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][20]  ( .D(n3493), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1019) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][19]  ( .D(n3430), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n956) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][19]  ( .D(n3494), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1020) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][18]  ( .D(n3431), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n957) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][18]  ( .D(n3495), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1021) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][17]  ( .D(n3432), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n958) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][17]  ( .D(n3496), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1022) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][16]  ( .D(n3433), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n959) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][16]  ( .D(n3497), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1023) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][15]  ( .D(n3434), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n960) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][15]  ( .D(n3498), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1024) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][14]  ( .D(n3435), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n961) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][14]  ( .D(n3499), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1025) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][13]  ( .D(n3436), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n962) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][13]  ( .D(n3500), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1026) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][12]  ( .D(n3437), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n963) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][12]  ( .D(n3501), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1027) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][11]  ( .D(n3438), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n964) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][11]  ( .D(n3502), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1028) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][10]  ( .D(n3439), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n965) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][10]  ( .D(n3503), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1029) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][9]  ( .D(n3440), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n966) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][9]  ( .D(n3504), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1030) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][8]  ( .D(n3441), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n967) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][8]  ( .D(n3505), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1031) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][7]  ( .D(n3442), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n968) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][7]  ( .D(n3506), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1032) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][6]  ( .D(n3443), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n969) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][6]  ( .D(n3507), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1033) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][5]  ( .D(n3444), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n970) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][5]  ( .D(n3508), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1034) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][4]  ( .D(n3445), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n971) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][4]  ( .D(n3509), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1035) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][3]  ( .D(n3446), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n972) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][3]  ( .D(n3510), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1036) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][2]  ( .D(n3447), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n973) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][2]  ( .D(n3511), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1037) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][1]  ( .D(n3448), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n974) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][1]  ( .D(n3512), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1038) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][0]  ( .D(n3449), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n975) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][0]  ( .D(n3513), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1039) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][31]  ( .D(n3514), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1040) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][30]  ( .D(n3515), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1041) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][29]  ( .D(n3516), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1042) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][28]  ( .D(n3517), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1043) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][27]  ( .D(n3518), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1044) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][26]  ( .D(n3519), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1045) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][25]  ( .D(n3520), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1046) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][24]  ( .D(n3521), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1047) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][23]  ( .D(n3522), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1048) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][22]  ( .D(n3523), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1049) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][21]  ( .D(n3524), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1050) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][20]  ( .D(n3525), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1051) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][19]  ( .D(n3526), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1052) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][18]  ( .D(n3527), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1053) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][17]  ( .D(n3528), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1054) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][16]  ( .D(n3529), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1055) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][15]  ( .D(n3530), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1056) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][14]  ( .D(n3531), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1057) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][13]  ( .D(n3532), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1058) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][12]  ( .D(n3533), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1059) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][11]  ( .D(n3534), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1060) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][10]  ( .D(n3535), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1061) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][9]  ( .D(n3536), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1062) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][8]  ( .D(n3537), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1063) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][7]  ( .D(n3538), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1064) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][6]  ( .D(n3539), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1065) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][5]  ( .D(n3540), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1066) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][4]  ( .D(n3541), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1067) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][3]  ( .D(n3542), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1068) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][2]  ( .D(n3543), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1069) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][1]  ( .D(n3544), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1070) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][0]  ( .D(n3545), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1071) );
  DFFNSRX2TS \addressToWriteBuffer_reg[5][7]  ( .D(n3294), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1193) );
  DFFNSRX2TS \addressToWriteBuffer_reg[5][6]  ( .D(n3295), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1194) );
  DFFNSRX2TS \addressToWriteBuffer_reg[5][5]  ( .D(n3296), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1195) );
  DFFNSRX2TS \addressToWriteBuffer_reg[5][4]  ( .D(n3297), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1196) );
  DFFNSRX2TS \addressToWriteBuffer_reg[5][3]  ( .D(n3298), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1197) );
  DFFNSRX2TS \addressToWriteBuffer_reg[5][2]  ( .D(n3299), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1198) );
  DFFNSRX2TS \addressToWriteBuffer_reg[5][1]  ( .D(n3300), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1199) );
  DFFNSRX2TS \addressToWriteBuffer_reg[5][0]  ( .D(n3301), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1200) );
  DFFNSRX2TS \addressToWriteBuffer_reg[3][7]  ( .D(n3310), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1209) );
  DFFNSRX2TS \addressToWriteBuffer_reg[3][6]  ( .D(n3311), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1210) );
  DFFNSRX2TS \addressToWriteBuffer_reg[3][5]  ( .D(n3312), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1211) );
  DFFNSRX2TS \addressToWriteBuffer_reg[3][4]  ( .D(n3313), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1212) );
  DFFNSRX2TS \addressToWriteBuffer_reg[3][3]  ( .D(n3314), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1213) );
  DFFNSRX2TS \addressToWriteBuffer_reg[3][2]  ( .D(n3315), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1214) );
  DFFNSRX2TS \addressToWriteBuffer_reg[3][1]  ( .D(n3316), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1215) );
  DFFNSRX2TS \addressToWriteBuffer_reg[3][0]  ( .D(n3317), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1216) );
  DFFNSRX2TS \addressToWriteBuffer_reg[6][7]  ( .D(n3286), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1185) );
  DFFNSRX2TS \addressToWriteBuffer_reg[4][7]  ( .D(n3302), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1201) );
  DFFNSRX2TS \addressToWriteBuffer_reg[6][6]  ( .D(n3287), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1186) );
  DFFNSRX2TS \addressToWriteBuffer_reg[4][6]  ( .D(n3303), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1202) );
  DFFNSRX2TS \addressToWriteBuffer_reg[6][5]  ( .D(n3288), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1187) );
  DFFNSRX2TS \addressToWriteBuffer_reg[4][5]  ( .D(n3304), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1203) );
  DFFNSRX2TS \addressToWriteBuffer_reg[6][4]  ( .D(n3289), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1188) );
  DFFNSRX2TS \addressToWriteBuffer_reg[4][4]  ( .D(n3305), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1204) );
  DFFNSRX2TS \addressToWriteBuffer_reg[6][3]  ( .D(n3290), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1189) );
  DFFNSRX2TS \addressToWriteBuffer_reg[4][3]  ( .D(n3306), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1205) );
  DFFNSRX2TS \addressToWriteBuffer_reg[6][2]  ( .D(n3291), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1190) );
  DFFNSRX2TS \addressToWriteBuffer_reg[4][2]  ( .D(n3307), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1206) );
  DFFNSRX2TS \addressToWriteBuffer_reg[6][1]  ( .D(n3292), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1191) );
  DFFNSRX2TS \addressToWriteBuffer_reg[4][1]  ( .D(n3308), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1207) );
  DFFNSRX2TS \addressToWriteBuffer_reg[6][0]  ( .D(n3293), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1192) );
  DFFNSRX2TS \addressToWriteBuffer_reg[4][0]  ( .D(n3309), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n1208) );
  DFFNSRX2TS \requesterPortBuffer_reg[3][1]  ( .D(n3260), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1257) );
  DFFNSRX2TS \dataToWriteBuffer_reg[0][20]  ( .D(n3621), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[0][20] ), .QN(n1147) );
  DFFNSRX2TS \dataToWriteBuffer_reg[0][19]  ( .D(n3622), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[0][19] ), .QN(n1148) );
  DFFNSRX2TS \dataToWriteBuffer_reg[0][18]  ( .D(n3623), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[0][18] ), .QN(n1149) );
  DFFNSRX2TS \dataToWriteBuffer_reg[0][17]  ( .D(n3624), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[0][17] ), .QN(n1150) );
  DFFNSRX2TS \dataToWriteBuffer_reg[0][16]  ( .D(n3625), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[0][16] ), .QN(n1151) );
  DFFNSRX2TS \dataToWriteBuffer_reg[0][15]  ( .D(n3626), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[0][15] ), .QN(n1152) );
  DFFNSRX2TS \dataToWriteBuffer_reg[0][14]  ( .D(n3627), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[0][14] ), .QN(n1153) );
  DFFNSRX2TS \dataToWriteBuffer_reg[0][13]  ( .D(n3628), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[0][13] ), .QN(n1154) );
  DFFNSRX2TS \dataToWriteBuffer_reg[0][12]  ( .D(n3629), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[0][12] ), .QN(n1155) );
  DFFNSRX2TS \dataToWriteBuffer_reg[0][11]  ( .D(n3630), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[0][11] ), .QN(n1156) );
  DFFNSRX2TS \dataToWriteBuffer_reg[0][10]  ( .D(n3631), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[0][10] ), .QN(n1157) );
  DFFNSRX2TS \dataToWriteBuffer_reg[0][9]  ( .D(n3632), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[0][9] ), .QN(n1158) );
  DFFNSRX2TS \dataToWriteBuffer_reg[0][8]  ( .D(n3633), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[0][8] ), .QN(n1159) );
  DFFNSRX2TS \dataToWriteBuffer_reg[0][7]  ( .D(n3634), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[0][7] ), .QN(n1160) );
  DFFNSRX2TS \dataToWriteBuffer_reg[0][6]  ( .D(n3635), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[0][6] ), .QN(n1161) );
  DFFNSRX2TS \dataToWriteBuffer_reg[0][5]  ( .D(n3636), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[0][5] ), .QN(n1162) );
  DFFNSRX2TS \dataToWriteBuffer_reg[0][4]  ( .D(n3637), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[0][4] ), .QN(n1163) );
  DFFNSRX2TS \dataToWriteBuffer_reg[0][3]  ( .D(n3638), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[0][3] ), .QN(n1164) );
  DFFNSRX2TS \dataToWriteBuffer_reg[0][2]  ( .D(n3639), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[0][2] ), .QN(n1165) );
  DFFNSRX2TS \dataToWriteBuffer_reg[0][1]  ( .D(n3640), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[0][1] ), .QN(n1166) );
  DFFNSRX2TS \dataToWriteBuffer_reg[0][0]  ( .D(n3641), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[0][0] ), .QN(n1167) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[0][5]  ( .D(n3165), .CK(clk), 
        .Q(requesterAddressOut_NORTH[5]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[0][4]  ( .D(n3164), .CK(clk), 
        .Q(requesterAddressOut_NORTH[4]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[0][3]  ( .D(n3163), .CK(clk), 
        .Q(requesterAddressOut_NORTH[3]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[0][2]  ( .D(n3162), .CK(clk), 
        .Q(requesterAddressOut_NORTH[2]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[0][1]  ( .D(n3161), .CK(clk), 
        .Q(requesterAddressOut_NORTH[1]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[0][0]  ( .D(n3160), .CK(clk), 
        .Q(requesterAddressOut_NORTH[0]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[3][5]  ( .D(n3183), .CK(clk), 
        .Q(requesterAddressOut_WEST[5]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[3][4]  ( .D(n3182), .CK(clk), 
        .Q(requesterAddressOut_WEST[4]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[3][3]  ( .D(n3181), .CK(clk), 
        .Q(requesterAddressOut_WEST[3]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[3][2]  ( .D(n3180), .CK(clk), 
        .Q(requesterAddressOut_WEST[2]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[3][1]  ( .D(n3179), .CK(clk), 
        .Q(requesterAddressOut_WEST[1]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[3][0]  ( .D(n3178), .CK(clk), 
        .Q(requesterAddressOut_WEST[0]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[2][5]  ( .D(n3177), .CK(clk), 
        .Q(requesterAddressOut_EAST[5]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[2][4]  ( .D(n3176), .CK(clk), 
        .Q(requesterAddressOut_EAST[4]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[2][3]  ( .D(n3175), .CK(clk), 
        .Q(requesterAddressOut_EAST[3]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[2][2]  ( .D(n3174), .CK(clk), 
        .Q(requesterAddressOut_EAST[2]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[2][1]  ( .D(n3173), .CK(clk), 
        .Q(requesterAddressOut_EAST[1]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[2][0]  ( .D(n3172), .CK(clk), 
        .Q(requesterAddressOut_EAST[0]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[1][5]  ( .D(n3171), .CK(clk), 
        .Q(requesterAddressOut_SOUTH[5]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[1][4]  ( .D(n3170), .CK(clk), 
        .Q(requesterAddressOut_SOUTH[4]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[1][3]  ( .D(n3169), .CK(clk), 
        .Q(requesterAddressOut_SOUTH[3]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[1][2]  ( .D(n3168), .CK(clk), 
        .Q(requesterAddressOut_SOUTH[2]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[1][1]  ( .D(n3167), .CK(clk), 
        .Q(requesterAddressOut_SOUTH[1]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[1][0]  ( .D(n3166), .CK(clk), 
        .Q(requesterAddressOut_SOUTH[0]) );
  DFFNSRX2TS prevMemRead_B_reg ( .D(n3344), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(prevMemRead_B) );
  DFFNSRX2TS prevMemRead_A_reg ( .D(n3342), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(prevMemRead_A) );
  DFFNSRX2TS \prevRequesterPort_A_reg[0]  ( .D(n3250), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3645), .QN(n3677) );
  DFFNSRX2TS \prevRequesterPort_A_reg[1]  ( .D(n3251), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3646), .QN(n3678) );
  DFFNSRX2TS \cacheAddressIn_A_reg[7]  ( .D(n3277), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_A[7]) );
  DFFNSRX2TS \cacheAddressIn_A_reg[6]  ( .D(n3276), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_A[6]) );
  DFFNSRX2TS \cacheAddressIn_A_reg[5]  ( .D(n3275), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_A[5]) );
  DFFNSRX2TS \cacheAddressIn_A_reg[4]  ( .D(n3274), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_A[4]) );
  DFFNSRX2TS \cacheAddressIn_A_reg[3]  ( .D(n3273), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_A[3]) );
  DFFNSRX2TS \cacheAddressIn_A_reg[2]  ( .D(n3272), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_A[2]) );
  DFFNSRX2TS \cacheAddressIn_A_reg[1]  ( .D(n3271), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_A[1]) );
  DFFNSRX2TS \cacheAddressIn_A_reg[0]  ( .D(n3270), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_A[0]) );
  DFFNSRX2TS \cacheDataIn_A_reg[31]  ( .D(n3249), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[31]) );
  DFFNSRX2TS \cacheDataIn_A_reg[30]  ( .D(n3248), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[30]) );
  DFFNSRX2TS \cacheDataIn_A_reg[29]  ( .D(n3247), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[29]) );
  DFFNSRX2TS \cacheDataIn_A_reg[28]  ( .D(n3246), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[28]) );
  DFFNSRX2TS \cacheDataIn_A_reg[27]  ( .D(n3245), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[27]) );
  DFFNSRX2TS \cacheDataIn_A_reg[26]  ( .D(n3244), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[26]) );
  DFFNSRX2TS \cacheDataIn_A_reg[25]  ( .D(n3243), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[25]) );
  DFFNSRX2TS \cacheDataIn_A_reg[24]  ( .D(n3242), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[24]) );
  DFFNSRX2TS \cacheDataIn_A_reg[23]  ( .D(n3241), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[23]) );
  DFFNSRX2TS \cacheDataIn_A_reg[22]  ( .D(n3240), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[22]) );
  DFFNSRX2TS \cacheDataIn_A_reg[21]  ( .D(n3239), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[21]) );
  DFFNSRX2TS \cacheDataIn_A_reg[20]  ( .D(n3238), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[20]) );
  DFFNSRX2TS \cacheDataIn_A_reg[19]  ( .D(n3237), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[19]) );
  DFFNSRX2TS \cacheDataIn_A_reg[18]  ( .D(n3236), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[18]) );
  DFFNSRX2TS \cacheDataIn_A_reg[17]  ( .D(n3235), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[17]) );
  DFFNSRX2TS \cacheDataIn_A_reg[16]  ( .D(n3234), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[16]) );
  DFFNSRX2TS \cacheDataIn_A_reg[15]  ( .D(n3233), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[15]) );
  DFFNSRX2TS \cacheDataIn_A_reg[14]  ( .D(n3232), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[14]) );
  DFFNSRX2TS \cacheDataIn_A_reg[13]  ( .D(n3231), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[13]) );
  DFFNSRX2TS \cacheDataIn_A_reg[12]  ( .D(n3230), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[12]) );
  DFFNSRX2TS \cacheDataIn_A_reg[11]  ( .D(n3229), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[11]) );
  DFFNSRX2TS \cacheDataIn_A_reg[10]  ( .D(n3228), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[10]) );
  DFFNSRX2TS \cacheDataIn_A_reg[9]  ( .D(n3227), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[9]) );
  DFFNSRX2TS \cacheDataIn_A_reg[8]  ( .D(n3226), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[8]) );
  DFFNSRX2TS \cacheDataIn_A_reg[7]  ( .D(n3225), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[7]) );
  DFFNSRX2TS \cacheDataIn_A_reg[6]  ( .D(n3224), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[6]) );
  DFFNSRX2TS \cacheDataIn_A_reg[5]  ( .D(n3223), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[5]) );
  DFFNSRX2TS \cacheDataIn_A_reg[4]  ( .D(n3222), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[4]) );
  DFFNSRX2TS \cacheDataIn_A_reg[3]  ( .D(n3221), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[3]) );
  DFFNSRX2TS \cacheDataIn_A_reg[2]  ( .D(n3220), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[2]) );
  DFFNSRX2TS \cacheDataIn_A_reg[1]  ( .D(n3219), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[1]) );
  DFFNSRX2TS \cacheDataIn_A_reg[0]  ( .D(n3218), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[0]) );
  DFFNSRX2TS memWrite_A_reg ( .D(n3184), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        memWrite_A) );
  DFFNSRX2TS memWrite_B_reg ( .D(n3217), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        memWrite_B) );
  DFFNSRX2TS \cacheDataIn_B_reg[31]  ( .D(n3377), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[31]) );
  DFFNSRX2TS \cacheDataIn_B_reg[30]  ( .D(n3376), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[30]) );
  DFFNSRX2TS \cacheDataIn_B_reg[29]  ( .D(n3375), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[29]) );
  DFFNSRX2TS \cacheDataIn_B_reg[28]  ( .D(n3374), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[28]) );
  DFFNSRX2TS \cacheDataIn_B_reg[27]  ( .D(n3373), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[27]) );
  DFFNSRX2TS \cacheDataIn_B_reg[26]  ( .D(n3372), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[26]) );
  DFFNSRX2TS \cacheDataIn_B_reg[25]  ( .D(n3371), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[25]) );
  DFFNSRX2TS \cacheDataIn_B_reg[24]  ( .D(n3370), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[24]) );
  DFFNSRX2TS \cacheDataIn_B_reg[23]  ( .D(n3369), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[23]) );
  DFFNSRX2TS \cacheDataIn_B_reg[22]  ( .D(n3368), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[22]) );
  DFFNSRX2TS \cacheDataIn_B_reg[21]  ( .D(n3367), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[21]) );
  DFFNSRX2TS \cacheDataIn_B_reg[20]  ( .D(n3366), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[20]) );
  DFFNSRX2TS \cacheDataIn_B_reg[19]  ( .D(n3365), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[19]) );
  DFFNSRX2TS \cacheDataIn_B_reg[18]  ( .D(n3364), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[18]) );
  DFFNSRX2TS \cacheDataIn_B_reg[17]  ( .D(n3363), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[17]) );
  DFFNSRX2TS \cacheDataIn_B_reg[16]  ( .D(n3362), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[16]) );
  DFFNSRX2TS \cacheDataIn_B_reg[15]  ( .D(n3361), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[15]) );
  DFFNSRX2TS \cacheDataIn_B_reg[14]  ( .D(n3360), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[14]) );
  DFFNSRX2TS \cacheDataIn_B_reg[13]  ( .D(n3359), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[13]) );
  DFFNSRX2TS \cacheDataIn_B_reg[12]  ( .D(n3358), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[12]) );
  DFFNSRX2TS \cacheDataIn_B_reg[11]  ( .D(n3357), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[11]) );
  DFFNSRX2TS \cacheDataIn_B_reg[10]  ( .D(n3356), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[10]) );
  DFFNSRX2TS \cacheDataIn_B_reg[9]  ( .D(n3355), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[9]) );
  DFFNSRX2TS \cacheDataIn_B_reg[8]  ( .D(n3354), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[8]) );
  DFFNSRX2TS \cacheDataIn_B_reg[7]  ( .D(n3353), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[7]) );
  DFFNSRX2TS \cacheDataIn_B_reg[6]  ( .D(n3352), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[6]) );
  DFFNSRX2TS \cacheDataIn_B_reg[5]  ( .D(n3351), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[5]) );
  DFFNSRX2TS \cacheDataIn_B_reg[4]  ( .D(n3350), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[4]) );
  DFFNSRX2TS \cacheDataIn_B_reg[3]  ( .D(n3349), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[3]) );
  DFFNSRX2TS \cacheDataIn_B_reg[2]  ( .D(n3348), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[2]) );
  DFFNSRX2TS \cacheDataIn_B_reg[1]  ( .D(n3347), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[1]) );
  DFFNSRX2TS \cacheDataIn_B_reg[0]  ( .D(n3346), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[0]) );
  DFFNSRX2TS \cacheAddressIn_B_reg[7]  ( .D(n3216), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_B[7]) );
  DFFNSRX2TS \cacheAddressIn_B_reg[6]  ( .D(n3215), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_B[6]) );
  DFFNSRX2TS \cacheAddressIn_B_reg[5]  ( .D(n3214), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_B[5]) );
  DFFNSRX2TS \cacheAddressIn_B_reg[4]  ( .D(n3213), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_B[4]) );
  DFFNSRX2TS \cacheAddressIn_B_reg[3]  ( .D(n3212), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_B[3]) );
  DFFNSRX2TS \cacheAddressIn_B_reg[2]  ( .D(n3211), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_B[2]) );
  DFFNSRX2TS \cacheAddressIn_B_reg[1]  ( .D(n3210), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_B[1]) );
  DFFNSRX2TS \cacheAddressIn_B_reg[0]  ( .D(n3209), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_B[0]) );
  TLATXLTS \dataOut_Concatenated_reg[3][31]  ( .G(clk), .D(N10220), .Q(
        cacheDataOut_WEST[31]) );
  TLATXLTS \dataOut_Concatenated_reg[3][30]  ( .G(clk), .D(N10219), .Q(
        cacheDataOut_WEST[30]) );
  TLATXLTS \dataOut_Concatenated_reg[3][29]  ( .G(clk), .D(N10218), .Q(
        cacheDataOut_WEST[29]) );
  TLATXLTS \dataOut_Concatenated_reg[3][28]  ( .G(clk), .D(N10217), .Q(
        cacheDataOut_WEST[28]) );
  TLATXLTS \dataOut_Concatenated_reg[3][27]  ( .G(clk), .D(N10216), .Q(
        cacheDataOut_WEST[27]) );
  TLATXLTS \dataOut_Concatenated_reg[3][26]  ( .G(clk), .D(N10215), .Q(
        cacheDataOut_WEST[26]) );
  TLATXLTS \dataOut_Concatenated_reg[3][25]  ( .G(clk), .D(N10214), .Q(
        cacheDataOut_WEST[25]) );
  TLATXLTS \dataOut_Concatenated_reg[3][24]  ( .G(clk), .D(N10213), .Q(
        cacheDataOut_WEST[24]) );
  TLATXLTS \dataOut_Concatenated_reg[3][23]  ( .G(clk), .D(N10212), .Q(
        cacheDataOut_WEST[23]) );
  TLATXLTS \dataOut_Concatenated_reg[3][22]  ( .G(clk), .D(N10211), .Q(
        cacheDataOut_WEST[22]) );
  TLATXLTS \dataOut_Concatenated_reg[3][21]  ( .G(clk), .D(N10210), .Q(
        cacheDataOut_WEST[21]) );
  TLATXLTS \dataOut_Concatenated_reg[3][20]  ( .G(clk), .D(N10209), .Q(
        cacheDataOut_WEST[20]) );
  TLATXLTS \dataOut_Concatenated_reg[3][19]  ( .G(clk), .D(N10208), .Q(
        cacheDataOut_WEST[19]) );
  TLATXLTS \dataOut_Concatenated_reg[3][18]  ( .G(clk), .D(N10207), .Q(
        cacheDataOut_WEST[18]) );
  TLATXLTS \dataOut_Concatenated_reg[3][17]  ( .G(clk), .D(N10206), .Q(
        cacheDataOut_WEST[17]) );
  TLATXLTS \dataOut_Concatenated_reg[3][16]  ( .G(clk), .D(N10205), .Q(
        cacheDataOut_WEST[16]) );
  TLATXLTS \dataOut_Concatenated_reg[3][15]  ( .G(clk), .D(N10204), .Q(
        cacheDataOut_WEST[15]) );
  TLATXLTS \dataOut_Concatenated_reg[3][14]  ( .G(clk), .D(N10203), .Q(
        cacheDataOut_WEST[14]) );
  TLATXLTS \dataOut_Concatenated_reg[3][13]  ( .G(clk), .D(N10202), .Q(
        cacheDataOut_WEST[13]) );
  TLATXLTS \dataOut_Concatenated_reg[3][12]  ( .G(clk), .D(N10201), .Q(
        cacheDataOut_WEST[12]) );
  TLATXLTS \dataOut_Concatenated_reg[3][11]  ( .G(clk), .D(N10200), .Q(
        cacheDataOut_WEST[11]) );
  TLATXLTS \dataOut_Concatenated_reg[3][10]  ( .G(clk), .D(N10199), .Q(
        cacheDataOut_WEST[10]) );
  TLATXLTS \dataOut_Concatenated_reg[3][9]  ( .G(clk), .D(N10198), .Q(
        cacheDataOut_WEST[9]) );
  TLATXLTS \dataOut_Concatenated_reg[3][8]  ( .G(clk), .D(N10197), .Q(
        cacheDataOut_WEST[8]) );
  TLATXLTS \dataOut_Concatenated_reg[3][7]  ( .G(clk), .D(N10196), .Q(
        cacheDataOut_WEST[7]) );
  TLATXLTS \dataOut_Concatenated_reg[3][6]  ( .G(clk), .D(N10195), .Q(
        cacheDataOut_WEST[6]) );
  TLATXLTS \dataOut_Concatenated_reg[3][5]  ( .G(clk), .D(N10194), .Q(
        cacheDataOut_WEST[5]) );
  TLATXLTS \dataOut_Concatenated_reg[3][4]  ( .G(clk), .D(N10193), .Q(
        cacheDataOut_WEST[4]) );
  TLATXLTS \dataOut_Concatenated_reg[3][3]  ( .G(clk), .D(N10192), .Q(
        cacheDataOut_WEST[3]) );
  TLATXLTS \dataOut_Concatenated_reg[3][2]  ( .G(clk), .D(N10191), .Q(
        cacheDataOut_WEST[2]) );
  TLATXLTS \dataOut_Concatenated_reg[3][1]  ( .G(clk), .D(N10190), .Q(
        cacheDataOut_WEST[1]) );
  TLATXLTS \dataOut_Concatenated_reg[3][0]  ( .G(clk), .D(N10189), .Q(
        cacheDataOut_WEST[0]) );
  TLATXLTS \dataOut_Concatenated_reg[2][31]  ( .G(clk), .D(N10186), .Q(
        cacheDataOut_EAST[31]) );
  TLATXLTS \dataOut_Concatenated_reg[2][30]  ( .G(clk), .D(N10185), .Q(
        cacheDataOut_EAST[30]) );
  TLATXLTS \dataOut_Concatenated_reg[2][29]  ( .G(clk), .D(N10184), .Q(
        cacheDataOut_EAST[29]) );
  TLATXLTS \dataOut_Concatenated_reg[2][28]  ( .G(clk), .D(N10183), .Q(
        cacheDataOut_EAST[28]) );
  TLATXLTS \dataOut_Concatenated_reg[2][27]  ( .G(clk), .D(N10182), .Q(
        cacheDataOut_EAST[27]) );
  TLATXLTS \dataOut_Concatenated_reg[2][26]  ( .G(clk), .D(N10181), .Q(
        cacheDataOut_EAST[26]) );
  TLATXLTS \dataOut_Concatenated_reg[2][25]  ( .G(clk), .D(N10180), .Q(
        cacheDataOut_EAST[25]) );
  TLATXLTS \dataOut_Concatenated_reg[2][24]  ( .G(clk), .D(N10179), .Q(
        cacheDataOut_EAST[24]) );
  TLATXLTS \dataOut_Concatenated_reg[2][23]  ( .G(clk), .D(N10178), .Q(
        cacheDataOut_EAST[23]) );
  TLATXLTS \dataOut_Concatenated_reg[2][22]  ( .G(clk), .D(N10177), .Q(
        cacheDataOut_EAST[22]) );
  TLATXLTS \dataOut_Concatenated_reg[2][21]  ( .G(clk), .D(N10176), .Q(
        cacheDataOut_EAST[21]) );
  TLATXLTS \dataOut_Concatenated_reg[2][20]  ( .G(clk), .D(N10175), .Q(
        cacheDataOut_EAST[20]) );
  TLATXLTS \dataOut_Concatenated_reg[2][19]  ( .G(clk), .D(N10174), .Q(
        cacheDataOut_EAST[19]) );
  TLATXLTS \dataOut_Concatenated_reg[2][18]  ( .G(clk), .D(N10173), .Q(
        cacheDataOut_EAST[18]) );
  TLATXLTS \dataOut_Concatenated_reg[2][17]  ( .G(clk), .D(N10172), .Q(
        cacheDataOut_EAST[17]) );
  TLATXLTS \dataOut_Concatenated_reg[2][16]  ( .G(clk), .D(N10171), .Q(
        cacheDataOut_EAST[16]) );
  TLATXLTS \dataOut_Concatenated_reg[2][15]  ( .G(clk), .D(N10170), .Q(
        cacheDataOut_EAST[15]) );
  TLATXLTS \dataOut_Concatenated_reg[2][14]  ( .G(clk), .D(N10169), .Q(
        cacheDataOut_EAST[14]) );
  TLATXLTS \dataOut_Concatenated_reg[2][13]  ( .G(clk), .D(N10168), .Q(
        cacheDataOut_EAST[13]) );
  TLATXLTS \dataOut_Concatenated_reg[2][12]  ( .G(clk), .D(N10167), .Q(
        cacheDataOut_EAST[12]) );
  TLATXLTS \dataOut_Concatenated_reg[2][11]  ( .G(clk), .D(N10166), .Q(
        cacheDataOut_EAST[11]) );
  TLATXLTS \dataOut_Concatenated_reg[2][10]  ( .G(clk), .D(N10165), .Q(
        cacheDataOut_EAST[10]) );
  TLATXLTS \dataOut_Concatenated_reg[2][9]  ( .G(clk), .D(N10164), .Q(
        cacheDataOut_EAST[9]) );
  TLATXLTS \dataOut_Concatenated_reg[2][8]  ( .G(clk), .D(N10163), .Q(
        cacheDataOut_EAST[8]) );
  TLATXLTS \dataOut_Concatenated_reg[2][7]  ( .G(clk), .D(N10162), .Q(
        cacheDataOut_EAST[7]) );
  TLATXLTS \dataOut_Concatenated_reg[2][6]  ( .G(clk), .D(N10161), .Q(
        cacheDataOut_EAST[6]) );
  TLATXLTS \dataOut_Concatenated_reg[2][5]  ( .G(clk), .D(N10160), .Q(
        cacheDataOut_EAST[5]) );
  TLATXLTS \dataOut_Concatenated_reg[2][4]  ( .G(clk), .D(N10159), .Q(
        cacheDataOut_EAST[4]) );
  TLATXLTS \dataOut_Concatenated_reg[2][3]  ( .G(clk), .D(N10158), .Q(
        cacheDataOut_EAST[3]) );
  TLATXLTS \dataOut_Concatenated_reg[2][2]  ( .G(clk), .D(N10157), .Q(
        cacheDataOut_EAST[2]) );
  TLATXLTS \dataOut_Concatenated_reg[2][1]  ( .G(clk), .D(N10156), .Q(
        cacheDataOut_EAST[1]) );
  TLATXLTS \dataOut_Concatenated_reg[2][0]  ( .G(clk), .D(N10155), .Q(
        cacheDataOut_EAST[0]) );
  TLATXLTS \dataOut_Concatenated_reg[1][31]  ( .G(clk), .D(N10152), .Q(
        cacheDataOut_SOUTH[31]) );
  TLATXLTS \dataOut_Concatenated_reg[1][30]  ( .G(clk), .D(N10151), .Q(
        cacheDataOut_SOUTH[30]) );
  TLATXLTS \dataOut_Concatenated_reg[1][29]  ( .G(clk), .D(N10150), .Q(
        cacheDataOut_SOUTH[29]) );
  TLATXLTS \dataOut_Concatenated_reg[1][28]  ( .G(clk), .D(N10149), .Q(
        cacheDataOut_SOUTH[28]) );
  TLATXLTS \dataOut_Concatenated_reg[1][27]  ( .G(clk), .D(N10148), .Q(
        cacheDataOut_SOUTH[27]) );
  TLATXLTS \dataOut_Concatenated_reg[1][26]  ( .G(clk), .D(N10147), .Q(
        cacheDataOut_SOUTH[26]) );
  TLATXLTS \dataOut_Concatenated_reg[1][25]  ( .G(clk), .D(N10146), .Q(
        cacheDataOut_SOUTH[25]) );
  TLATXLTS \dataOut_Concatenated_reg[1][24]  ( .G(clk), .D(N10145), .Q(
        cacheDataOut_SOUTH[24]) );
  TLATXLTS \dataOut_Concatenated_reg[1][23]  ( .G(clk), .D(N10144), .Q(
        cacheDataOut_SOUTH[23]) );
  TLATXLTS \dataOut_Concatenated_reg[1][22]  ( .G(clk), .D(N10143), .Q(
        cacheDataOut_SOUTH[22]) );
  TLATXLTS \dataOut_Concatenated_reg[1][21]  ( .G(clk), .D(N10142), .Q(
        cacheDataOut_SOUTH[21]) );
  TLATXLTS \dataOut_Concatenated_reg[1][20]  ( .G(clk), .D(N10141), .Q(
        cacheDataOut_SOUTH[20]) );
  TLATXLTS \dataOut_Concatenated_reg[1][19]  ( .G(clk), .D(N10140), .Q(
        cacheDataOut_SOUTH[19]) );
  TLATXLTS \dataOut_Concatenated_reg[1][18]  ( .G(clk), .D(N10139), .Q(
        cacheDataOut_SOUTH[18]) );
  TLATXLTS \dataOut_Concatenated_reg[1][17]  ( .G(clk), .D(N10138), .Q(
        cacheDataOut_SOUTH[17]) );
  TLATXLTS \dataOut_Concatenated_reg[1][16]  ( .G(clk), .D(N10137), .Q(
        cacheDataOut_SOUTH[16]) );
  TLATXLTS \dataOut_Concatenated_reg[1][15]  ( .G(clk), .D(N10136), .Q(
        cacheDataOut_SOUTH[15]) );
  TLATXLTS \dataOut_Concatenated_reg[1][14]  ( .G(clk), .D(N10135), .Q(
        cacheDataOut_SOUTH[14]) );
  TLATXLTS \dataOut_Concatenated_reg[1][13]  ( .G(clk), .D(N10134), .Q(
        cacheDataOut_SOUTH[13]) );
  TLATXLTS \dataOut_Concatenated_reg[1][12]  ( .G(clk), .D(N10133), .Q(
        cacheDataOut_SOUTH[12]) );
  TLATXLTS \dataOut_Concatenated_reg[1][11]  ( .G(clk), .D(N10132), .Q(
        cacheDataOut_SOUTH[11]) );
  TLATXLTS \dataOut_Concatenated_reg[1][10]  ( .G(clk), .D(N10131), .Q(
        cacheDataOut_SOUTH[10]) );
  TLATXLTS \dataOut_Concatenated_reg[1][9]  ( .G(clk), .D(N10130), .Q(
        cacheDataOut_SOUTH[9]) );
  TLATXLTS \dataOut_Concatenated_reg[1][8]  ( .G(clk), .D(N10129), .Q(
        cacheDataOut_SOUTH[8]) );
  TLATXLTS \dataOut_Concatenated_reg[1][7]  ( .G(clk), .D(N10128), .Q(
        cacheDataOut_SOUTH[7]) );
  TLATXLTS \dataOut_Concatenated_reg[1][6]  ( .G(clk), .D(N10127), .Q(
        cacheDataOut_SOUTH[6]) );
  TLATXLTS \dataOut_Concatenated_reg[1][5]  ( .G(clk), .D(N10126), .Q(
        cacheDataOut_SOUTH[5]) );
  TLATXLTS \dataOut_Concatenated_reg[1][4]  ( .G(clk), .D(N10125), .Q(
        cacheDataOut_SOUTH[4]) );
  TLATXLTS \dataOut_Concatenated_reg[1][3]  ( .G(clk), .D(N10124), .Q(
        cacheDataOut_SOUTH[3]) );
  TLATXLTS \dataOut_Concatenated_reg[1][2]  ( .G(clk), .D(N10123), .Q(
        cacheDataOut_SOUTH[2]) );
  TLATXLTS \dataOut_Concatenated_reg[1][1]  ( .G(clk), .D(N10122), .Q(
        cacheDataOut_SOUTH[1]) );
  TLATXLTS \dataOut_Concatenated_reg[1][0]  ( .G(clk), .D(N10121), .Q(
        cacheDataOut_SOUTH[0]) );
  TLATXLTS \dataOut_Concatenated_reg[0][31]  ( .G(clk), .D(N10118), .Q(
        cacheDataOut_NORTH[31]) );
  TLATXLTS \dataOut_Concatenated_reg[0][30]  ( .G(clk), .D(N10117), .Q(
        cacheDataOut_NORTH[30]) );
  TLATXLTS \dataOut_Concatenated_reg[0][29]  ( .G(clk), .D(N10116), .Q(
        cacheDataOut_NORTH[29]) );
  TLATXLTS \dataOut_Concatenated_reg[0][28]  ( .G(clk), .D(N10115), .Q(
        cacheDataOut_NORTH[28]) );
  TLATXLTS \dataOut_Concatenated_reg[0][27]  ( .G(clk), .D(N10114), .Q(
        cacheDataOut_NORTH[27]) );
  TLATXLTS \dataOut_Concatenated_reg[0][26]  ( .G(clk), .D(N10113), .Q(
        cacheDataOut_NORTH[26]) );
  TLATXLTS \dataOut_Concatenated_reg[0][25]  ( .G(clk), .D(N10112), .Q(
        cacheDataOut_NORTH[25]) );
  TLATXLTS \dataOut_Concatenated_reg[0][24]  ( .G(clk), .D(N10111), .Q(
        cacheDataOut_NORTH[24]) );
  TLATXLTS \dataOut_Concatenated_reg[0][23]  ( .G(clk), .D(N10110), .Q(
        cacheDataOut_NORTH[23]) );
  TLATXLTS \dataOut_Concatenated_reg[0][22]  ( .G(clk), .D(N10109), .Q(
        cacheDataOut_NORTH[22]) );
  TLATXLTS \dataOut_Concatenated_reg[0][21]  ( .G(clk), .D(N10108), .Q(
        cacheDataOut_NORTH[21]) );
  TLATXLTS \dataOut_Concatenated_reg[0][20]  ( .G(clk), .D(N10107), .Q(
        cacheDataOut_NORTH[20]) );
  TLATXLTS \dataOut_Concatenated_reg[0][19]  ( .G(clk), .D(N10106), .Q(
        cacheDataOut_NORTH[19]) );
  TLATXLTS \dataOut_Concatenated_reg[0][18]  ( .G(clk), .D(N10105), .Q(
        cacheDataOut_NORTH[18]) );
  TLATXLTS \dataOut_Concatenated_reg[0][17]  ( .G(clk), .D(N10104), .Q(
        cacheDataOut_NORTH[17]) );
  TLATXLTS \dataOut_Concatenated_reg[0][16]  ( .G(clk), .D(N10103), .Q(
        cacheDataOut_NORTH[16]) );
  TLATXLTS \dataOut_Concatenated_reg[0][15]  ( .G(clk), .D(N10102), .Q(
        cacheDataOut_NORTH[15]) );
  TLATXLTS \dataOut_Concatenated_reg[0][14]  ( .G(clk), .D(N10101), .Q(
        cacheDataOut_NORTH[14]) );
  TLATXLTS \dataOut_Concatenated_reg[0][13]  ( .G(clk), .D(N10100), .Q(
        cacheDataOut_NORTH[13]) );
  TLATXLTS \dataOut_Concatenated_reg[0][12]  ( .G(clk), .D(N10099), .Q(
        cacheDataOut_NORTH[12]) );
  TLATXLTS \dataOut_Concatenated_reg[0][11]  ( .G(clk), .D(N10098), .Q(
        cacheDataOut_NORTH[11]) );
  TLATXLTS \dataOut_Concatenated_reg[0][10]  ( .G(clk), .D(N10097), .Q(
        cacheDataOut_NORTH[10]) );
  TLATXLTS \dataOut_Concatenated_reg[0][9]  ( .G(clk), .D(N10096), .Q(
        cacheDataOut_NORTH[9]) );
  TLATXLTS \dataOut_Concatenated_reg[0][8]  ( .G(clk), .D(N10095), .Q(
        cacheDataOut_NORTH[8]) );
  TLATXLTS \dataOut_Concatenated_reg[0][7]  ( .G(clk), .D(N10094), .Q(
        cacheDataOut_NORTH[7]) );
  TLATXLTS \dataOut_Concatenated_reg[0][6]  ( .G(clk), .D(N10093), .Q(
        cacheDataOut_NORTH[6]) );
  TLATXLTS \dataOut_Concatenated_reg[0][5]  ( .G(clk), .D(N10092), .Q(
        cacheDataOut_NORTH[5]) );
  TLATXLTS \dataOut_Concatenated_reg[0][4]  ( .G(clk), .D(N10091), .Q(
        cacheDataOut_NORTH[4]) );
  TLATXLTS \dataOut_Concatenated_reg[0][3]  ( .G(clk), .D(N10090), .Q(
        cacheDataOut_NORTH[3]) );
  TLATXLTS \dataOut_Concatenated_reg[0][2]  ( .G(clk), .D(N10089), .Q(
        cacheDataOut_NORTH[2]) );
  TLATXLTS \dataOut_Concatenated_reg[0][1]  ( .G(clk), .D(N10088), .Q(
        cacheDataOut_NORTH[1]) );
  TLATXLTS \dataOut_Concatenated_reg[0][0]  ( .G(clk), .D(N10087), .Q(
        cacheDataOut_NORTH[0]) );
  DFFQX1TS \readReady_Concatenated_reg[3]  ( .D(N10079), .CK(clk), .Q(
        readReady_WEST) );
  DFFQX1TS \readReady_Concatenated_reg[2]  ( .D(N10078), .CK(clk), .Q(
        readReady_EAST) );
  DFFQX1TS \readReady_Concatenated_reg[1]  ( .D(N10077), .CK(clk), .Q(
        readReady_SOUTH) );
  DFFQX1TS \readReady_Concatenated_reg[0]  ( .D(N10076), .CK(clk), .Q(
        readReady_NORTH) );
  DFFNSRXLTS \prevRequesterPort_B_reg[1]  ( .D(n3264), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterPort_B[1]), .QN(n1241) );
  DFFNSRXLTS \prevRequesterPort_B_reg[0]  ( .D(n3265), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterPort_B[0]), .QN(n1243) );
  DFFNSRXLTS \prevRequesterAddress_B_reg[5]  ( .D(n3197), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_B[5]), .QN(n1244) );
  DFFNSRXLTS \prevRequesterAddress_B_reg[4]  ( .D(n3198), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_B[4]), .QN(n1245) );
  DFFNSRXLTS \prevRequesterAddress_B_reg[3]  ( .D(n3199), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_B[3]), .QN(n1246) );
  DFFNSRXLTS \prevRequesterAddress_B_reg[2]  ( .D(n3200), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_B[2]), .QN(n1247) );
  DFFNSRXLTS \prevRequesterAddress_B_reg[1]  ( .D(n3201), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_B[1]), .QN(n1248) );
  DFFNSRXLTS \prevRequesterAddress_B_reg[0]  ( .D(n3202), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_B[0]), .QN(n1249) );
  DFFNSRXLTS \prevRequesterAddress_A_reg[5]  ( .D(n3185), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_A[5]), .QN(n1267) );
  DFFNSRXLTS \prevRequesterAddress_A_reg[4]  ( .D(n3186), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_A[4]), .QN(n1268) );
  DFFNSRXLTS \prevRequesterAddress_A_reg[3]  ( .D(n3187), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_A[3]), .QN(n1269) );
  DFFNSRXLTS \prevRequesterAddress_A_reg[2]  ( .D(n3188), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_A[2]), .QN(n1270) );
  DFFNSRXLTS \prevRequesterAddress_A_reg[1]  ( .D(n3189), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_A[1]), .QN(n1271) );
  DFFNSRXLTS \prevRequesterAddress_A_reg[0]  ( .D(n3190), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_A[0]), .QN(n1272) );
  DFFNSRXLTS \requesterPortBuffer_reg[4][1]  ( .D(n3258), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[4][1] ), .QN(n1255) );
  DFFNSRXLTS \requesterPortBuffer_reg[4][0]  ( .D(n3259), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[4][0] ), .QN(n1256) );
  DFFNSRXLTS \requesterPortBuffer_reg[2][0]  ( .D(n3263), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[2][0] ), .QN(n1260) );
  DFFNSRXLTS \requesterPortBuffer_reg[5][1]  ( .D(n3256), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[5][1] ), .QN(n1253) );
  DFFNSRXLTS \requesterPortBuffer_reg[5][0]  ( .D(n3257), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[5][0] ), .QN(n1254) );
  DFFNSRXLTS \requesterPortBuffer_reg[6][1]  ( .D(n3254), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[6][1] ), .QN(n1251) );
  DFFNSRXLTS \requesterPortBuffer_reg[6][0]  ( .D(n3255), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[6][0] ), .QN(n1252) );
  DFFNSRXLTS \requesterPortBuffer_reg[7][1]  ( .D(n3252), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[7][1] ), .QN(n1250) );
  DFFNSRXLTS \isWrite_reg[6]  ( .D(n3379), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(isWrite[6]), .QN(n1168) );
  DFFNSRXLTS \addressToWriteBuffer_reg[2][7]  ( .D(n3318), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[2][7] ), .QN(n1217) );
  DFFNSRXLTS \addressToWriteBuffer_reg[2][6]  ( .D(n3319), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[2][6] ), .QN(n1218) );
  DFFNSRXLTS \addressToWriteBuffer_reg[2][5]  ( .D(n3320), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[2][5] ), .QN(n1219) );
  DFFNSRXLTS \addressToWriteBuffer_reg[2][4]  ( .D(n3321), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[2][4] ), .QN(n1220) );
  DFFNSRXLTS \addressToWriteBuffer_reg[2][3]  ( .D(n3322), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[2][3] ), .QN(n1221) );
  DFFNSRXLTS \addressToWriteBuffer_reg[2][2]  ( .D(n3323), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[2][2] ), .QN(n1222) );
  DFFNSRXLTS \addressToWriteBuffer_reg[2][1]  ( .D(n3324), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[2][1] ), .QN(n1223) );
  DFFNSRXLTS \addressToWriteBuffer_reg[2][0]  ( .D(n3325), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[2][0] ), .QN(n1224) );
  DFFNSRXLTS \isWrite_reg[1]  ( .D(n3384), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(isWrite[1]), .QN(n1173) );
  DFFNSRXLTS \isWrite_reg[2]  ( .D(n3383), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(isWrite[2]), .QN(n1172) );
  DFFNSRXLTS \isWrite_reg[4]  ( .D(n3381), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(isWrite[4]), .QN(n1170) );
  DFFNSRXLTS \requesterAddressBuffer_reg[0][5]  ( .D(n3196), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressBuffer[0][5] ), .QN(n1279) );
  DFFNSRXLTS \requesterAddressBuffer_reg[0][4]  ( .D(n3195), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressBuffer[0][4] ), .QN(n1280) );
  DFFNSRXLTS \requesterAddressBuffer_reg[0][2]  ( .D(n3193), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressBuffer[0][2] ), .QN(n1282) );
  DFFNSRXLTS \requesterAddressBuffer_reg[0][3]  ( .D(n3194), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressBuffer[0][3] ), .QN(n1281) );
  DFFNSRXLTS \requesterAddressBuffer_reg[0][1]  ( .D(n3192), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressBuffer[0][1] ), .QN(n1283) );
  DFFNSRXLTS \requesterAddressBuffer_reg[0][0]  ( .D(n3191), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressBuffer[0][0] ), .QN(n1284) );
  DFFNSRXLTS \addressToWriteBuffer_reg[0][7]  ( .D(n3334), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[0][7] ), .QN(n1233) );
  DFFNSRXLTS \addressToWriteBuffer_reg[0][6]  ( .D(n3335), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[0][6] ), .QN(n1234) );
  DFFNSRXLTS \addressToWriteBuffer_reg[0][5]  ( .D(n3336), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[0][5] ), .QN(n1235) );
  DFFNSRXLTS \addressToWriteBuffer_reg[0][4]  ( .D(n3337), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[0][4] ), .QN(n1236) );
  DFFNSRXLTS \addressToWriteBuffer_reg[0][3]  ( .D(n3338), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[0][3] ), .QN(n1237) );
  DFFNSRXLTS \addressToWriteBuffer_reg[0][2]  ( .D(n3339), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[0][2] ), .QN(n1238) );
  DFFNSRXLTS \addressToWriteBuffer_reg[0][1]  ( .D(n3340), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[0][1] ), .QN(n1239) );
  DFFNSRXLTS \addressToWriteBuffer_reg[0][0]  ( .D(n3341), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(\addressToWriteBuffer[0][0] ), .QN(n1240) );
  DFFNSRXLTS \isWrite_reg[5]  ( .D(n3380), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(isWrite[5]), .QN(n1169) );
  DFFNSRXLTS \isWrite_reg[0]  ( .D(n3385), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(isWrite[0]), .QN(n1174) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][31]  ( .D(n3610), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[0][31] ), .QN(n1136) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][30]  ( .D(n3611), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[0][30] ), .QN(n1137) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][29]  ( .D(n3612), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[0][29] ), .QN(n1138) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][28]  ( .D(n3613), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[0][28] ), .QN(n1139) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][27]  ( .D(n3614), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[0][27] ), .QN(n1140) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][26]  ( .D(n3615), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[0][26] ), .QN(n1141) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][25]  ( .D(n3616), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[0][25] ), .QN(n1142) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][24]  ( .D(n3617), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[0][24] ), .QN(n1143) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][23]  ( .D(n3618), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[0][23] ), .QN(n1144) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][22]  ( .D(n3619), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[0][22] ), .QN(n1145) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][21]  ( .D(n3620), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\dataToWriteBuffer[0][21] ), .QN(n1146) );
  DFFNSRX2TS \nextEmptyBuffer_reg[1]  ( .D(n3643), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(N650), .QN(n910) );
  DFFNSRX2TS \nextEmptyBuffer_reg[0]  ( .D(n3644), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3680), .QN(n4621) );
  DFFNSRX2TS \nextEmptyBuffer_reg[2]  ( .D(n3642), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(N651), .QN(n880) );
  AND3X2TS U3082 ( .A(n2425), .B(n5759), .C(\add_0_root_r1459/SUM[2] ), .Y(
        n2701) );
  NOR2BX2TS U3083 ( .AN(n3112), .B(\add_0_root_r1459/SUM[0] ), .Y(n2425) );
  AOI221X1TS U3084 ( .A0(n5211), .A1(n4172), .B0(n4848), .B1(n4308), .C0(n2958), .Y(n2957) );
  AOI221X1TS U3085 ( .A0(n5211), .A1(n4168), .B0(n4848), .B1(n4303), .C0(n2962), .Y(n2961) );
  OAI22XLTS U3086 ( .A0(n2840), .A1(n1090), .B0(n2917), .B1(n4860), .Y(n3564)
         );
  BUFX4TS U3087 ( .A(n2840), .Y(n4877) );
  OAI22XLTS U3088 ( .A0(n4874), .A1(n1086), .B0(n2901), .B1(n4861), .Y(n3560)
         );
  AOI221X1TS U3089 ( .A0(n5204), .A1(n4228), .B0(n4850), .B1(n4378), .C0(n2902), .Y(n2901) );
  OAI22XLTS U3090 ( .A0(n4868), .A1(n1102), .B0(n2965), .B1(n4858), .Y(n3576)
         );
  AOI221X1TS U3091 ( .A0(n2009), .A1(n4164), .B0(n4848), .B1(n4298), .C0(n2966), .Y(n2965) );
  OAI22XLTS U3092 ( .A0(n4873), .A1(n1075), .B0(n2857), .B1(n4864), .Y(n3549)
         );
  AOI221X1TS U3093 ( .A0(n5207), .A1(n4272), .B0(n4853), .B1(n4433), .C0(n2858), .Y(n2857) );
  OAI22XLTS U3094 ( .A0(n4869), .A1(n1099), .B0(n2953), .B1(n4867), .Y(n3573)
         );
  AOI221X1TS U3095 ( .A0(n5214), .A1(n4176), .B0(n4849), .B1(n4313), .C0(n2954), .Y(n2953) );
  OAI22XLTS U3096 ( .A0(n4868), .A1(n1103), .B0(n2969), .B1(n4858), .Y(n3577)
         );
  AOI221X1TS U3097 ( .A0(n5213), .A1(n4160), .B0(n4848), .B1(n4293), .C0(n2970), .Y(n2969) );
  NAND2X1TS U3098 ( .A(n4609), .B(n5224), .Y(n2002) );
  OAI31X1TS U3099 ( .A0(n5776), .A1(n5705), .A2(n2424), .B0(n5263), .Y(n1958)
         );
  AND2X2TS U3100 ( .A(n4593), .B(n4603), .Y(\add_0_root_r1463/carry [1]) );
  NOR2X1TS U3101 ( .A(\add_0_root_r1459/SUM[3] ), .B(\add_0_root_r1459/SUM[4] ), .Y(n3112) );
  XOR2X1TS U3102 ( .A(n4604), .B(n4605), .Y(\add_0_root_r1459/SUM[4] ) );
  AND3X2TS U3103 ( .A(n2426), .B(n5772), .C(n3697), .Y(n3659) );
  CMPR32X2TS U3104 ( .A(n5696), .B(\add_0_root_r1459/B[4] ), .C(
        \add_0_root_r1459/carry [2]), .CO(\add_0_root_r1459/carry [3]), .S(
        \add_0_root_r1459/SUM[2] ) );
  NOR2X1TS U3105 ( .A(n4618), .B(\add_0_root_sub_278_I2/A[0] ), .Y(n1573) );
  AOI21X1TS U3106 ( .A0(\add_0_root_sub_278_I2/A[0] ), .A1(n4618), .B0(n1573), 
        .Y(n3149) );
  NOR4XLTS U3107 ( .A(n5696), .B(n4878), .C(n2834), .D(n2002), .Y(n2836) );
  AND3X2TS U3108 ( .A(n2425), .B(n3699), .C(\add_0_root_r1459/SUM[1] ), .Y(
        n2423) );
  AND3X2TS U3109 ( .A(n2425), .B(n5758), .C(n3703), .Y(n2975) );
  NOR4XLTS U3110 ( .A(n4940), .B(n2698), .C(n5295), .D(n1958), .Y(n2700) );
  NOR4XLTS U3111 ( .A(n3806), .B(n5003), .C(n2560), .D(n1913), .Y(n2562) );
  NOR2X1TS U3112 ( .A(n3692), .B(n3688), .Y(n1748) );
  INVX2TS U3113 ( .A(n1823), .Y(\add_0_root_sub_278_I2/A[0] ) );
  OAI32XLTS U3114 ( .A0(n2217), .A1(n1752), .A2(n2218), .B0(n3791), .B1(n3689), 
        .Y(n2216) );
  OAI22XLTS U3115 ( .A0(n2270), .A1(n1641), .B0(n3810), .B1(n3689), .Y(n2269)
         );
  NAND2X2TS U3116 ( .A(\add_0_root_r1459/carry [3]), .B(n5807), .Y(n4605) );
  INVX1TS U3117 ( .A(n3689), .Y(n3690) );
  INVX1TS U3118 ( .A(n3687), .Y(n3688) );
  CLKINVX1TS U3119 ( .A(n1823), .Y(n4607) );
  NOR2X2TS U3120 ( .A(n3684), .B(n3682), .Y(n1823) );
  OAI211X1TS U3121 ( .A0(n5587), .A1(n2562), .B0(n1755), .C0(n2223), .Y(n2428)
         );
  NOR2X2TS U3122 ( .A(n3690), .B(n3686), .Y(n2255) );
  INVXLTS U3123 ( .A(n4603), .Y(n3151) );
  OR3XLTS U3124 ( .A(n4600), .B(n3695), .C(n4603), .Y(n3661) );
  AND4XLTS U3125 ( .A(n3763), .B(n2425), .C(n5758), .D(n5759), .Y(n3671) );
  OAI211XLTS U3126 ( .A0(n5599), .A1(n2836), .B0(n1775), .C0(n2249), .Y(n2702)
         );
  INVX1TS U3127 ( .A(N589), .Y(\add_0_root_r1463/B[4] ) );
  OAI31X1TS U3128 ( .A0(n5713), .A1(n2424), .A2(n5776), .B0(n5357), .Y(n1869)
         );
  OAI31X1TS U3129 ( .A0(n5713), .A1(n4578), .A2(n2424), .B0(n5185), .Y(n2046)
         );
  CMPR32X2TS U3130 ( .A(n5711), .B(\add_0_root_r1463/B[4] ), .C(
        \add_0_root_r1463/carry [1]), .CO(\add_0_root_r1463/carry [2]), .S(
        \add_0_root_r1463/SUM[1] ) );
  XNOR2X1TS U3131 ( .A(n3156), .B(n4607), .Y(n4603) );
  CMPR32X2TS U3132 ( .A(n5711), .B(\add_0_root_r1459/B[4] ), .C(
        \add_0_root_r1459/carry [1]), .CO(\add_0_root_r1459/carry [2]), .S(
        \add_0_root_r1459/SUM[1] ) );
  NAND2X1TS U3133 ( .A(n4992), .B(n5722), .Y(n2568) );
  NAND2X1TS U3134 ( .A(n5116), .B(n5722), .Y(n2289) );
  CMPR32X2TS U3135 ( .A(n5696), .B(\add_0_root_r1463/B[4] ), .C(
        \add_0_root_r1463/carry [2]), .CO(\add_0_root_r1463/carry [3]), .S(
        \add_0_root_r1463/SUM[2] ) );
  NAND2X1TS U3136 ( .A(n4868), .B(n5723), .Y(n2842) );
  CLKBUFX2TS U3137 ( .A(n5280), .Y(n5279) );
  CLKBUFX2TS U3138 ( .A(n5374), .Y(n5373) );
  NOR4X1TS U3139 ( .A(n1740), .B(n5064), .C(n2419), .D(n1869), .Y(n2422) );
  NOR4X1TS U3140 ( .A(n1783), .B(n4816), .C(n2972), .D(n2046), .Y(n2974) );
  NAND2X1TS U3141 ( .A(n5766), .B(n4544), .Y(n2274) );
  NAND2X1TS U3142 ( .A(n2701), .B(n4590), .Y(n1924) );
  NAND2X1TS U3143 ( .A(n4620), .B(n5718), .Y(n1620) );
  CLKBUFX2TS U3144 ( .A(n1618), .Y(n4620) );
  OAI21X1TS U3145 ( .A0(n4567), .A1(n2275), .B0(n2274), .Y(n2126) );
  NOR3XLTS U3146 ( .A(\indexIncrementer_EAST[1] ), .B(\add_0_root_r1459/B[0] ), 
        .C(n3745), .Y(n1585) );
  INVX2TS U3147 ( .A(n3683), .Y(n3684) );
  OAI211X1TS U3148 ( .A0(n5586), .A1(n2974), .B0(n1786), .C0(n2265), .Y(n2840)
         );
  OAI211X1TS U3149 ( .A0(n5593), .A1(n2700), .B0(n1765), .C0(n2236), .Y(n2566)
         );
  OAI211X1TS U3150 ( .A0(n5588), .A1(n2422), .B0(n1743), .C0(n2211), .Y(n2287)
         );
  OAI21X1TS U3151 ( .A0(n5763), .A1(n5570), .B0(n2205), .Y(n3647) );
  OAI21X1TS U3152 ( .A0(n5762), .A1(n5570), .B0(n2205), .Y(n3648) );
  OAI21X1TS U3153 ( .A0(n5768), .A1(n5569), .B0(n2205), .Y(n3649) );
  AND2X2TS U3154 ( .A(n3666), .B(n2426), .Y(n3650) );
  AO21X1TS U3155 ( .A0(n5907), .A1(n5763), .B0(n5292), .Y(n3651) );
  AO21X1TS U3156 ( .A0(n5907), .A1(n5762), .B0(n1783), .Y(n3652) );
  AND3X2TS U3157 ( .A(n4597), .B(n5775), .C(n1914), .Y(n3653) );
  NAND2X1TS U3158 ( .A(n2563), .B(n4591), .Y(n1879) );
  AND3X2TS U3159 ( .A(n4599), .B(n5785), .C(n2228), .Y(n3654) );
  INVX1TS U3160 ( .A(n3691), .Y(n3692) );
  OR2X2TS U3161 ( .A(n5591), .B(n5728), .Y(n3655) );
  OA21XLTS U3162 ( .A0(n2280), .A1(n5566), .B0(n3749), .Y(n3656) );
  OAI21X1TS U3163 ( .A0(n5765), .A1(n5569), .B0(n3749), .Y(n3657) );
  OAI21X1TS U3164 ( .A0(n5770), .A1(n5569), .B0(n3749), .Y(n3658) );
  OA21XLTS U3165 ( .A0(n5766), .A1(n5566), .B0(n3749), .Y(n3660) );
  OR3X1TS U3166 ( .A(n4600), .B(n3695), .C(n3151), .Y(n3662) );
  AO21X1TS U3167 ( .A0(n3754), .A1(n5765), .B0(n1740), .Y(n3663) );
  AO21X1TS U3168 ( .A0(n3754), .A1(n5768), .B0(n5697), .Y(n3664) );
  AO21X1TS U3169 ( .A0(n3754), .A1(n5770), .B0(n3806), .Y(n3665) );
  AND2X2TS U3170 ( .A(\add_0_root_r1463/SUM[1] ), .B(n3701), .Y(n3666) );
  AND3X2TS U3171 ( .A(N6620), .B(n4599), .C(n1914), .Y(n3667) );
  AND3X2TS U3172 ( .A(n1870), .B(n3718), .C(N6619), .Y(n3668) );
  AND3X2TS U3173 ( .A(N6618), .B(n4597), .C(n2003), .Y(n3669) );
  AND3X2TS U3174 ( .A(n3719), .B(n5796), .C(n2003), .Y(n3670) );
  NAND2X1TS U3175 ( .A(n1584), .B(n1585), .Y(n3672) );
  NAND2X1TS U3176 ( .A(n1584), .B(n3721), .Y(n3673) );
  OR2X2TS U3177 ( .A(n1733), .B(n5592), .Y(n3674) );
  OR2X2TS U3178 ( .A(n1616), .B(n3728), .Y(n3675) );
  OR3X1TS U3179 ( .A(n1585), .B(n5527), .C(n3745), .Y(n3676) );
  NAND2X1TS U3180 ( .A(n2423), .B(n4592), .Y(n1834) );
  INVX2TS U3181 ( .A(n2255), .Y(n3744) );
  AND2X2TS U3182 ( .A(n3684), .B(n4617), .Y(n3679) );
  INVX1TS U3183 ( .A(n3685), .Y(n3686) );
  INVX1TS U3184 ( .A(n3681), .Y(n3682) );
  INVXLTS U3185 ( .A(memRead_NORTH), .Y(n3681) );
  INVXLTS U3186 ( .A(memWrite_NORTH), .Y(n3683) );
  INVXLTS U3187 ( .A(memRead_EAST), .Y(n3685) );
  INVXLTS U3188 ( .A(memRead_SOUTH), .Y(n3687) );
  INVXLTS U3189 ( .A(memWrite_EAST), .Y(n3689) );
  INVXLTS U3190 ( .A(memWrite_SOUTH), .Y(n3691) );
  INVXLTS U3191 ( .A(n3678), .Y(n3693) );
  INVXLTS U3192 ( .A(n3677), .Y(n3694) );
  INVXLTS U3193 ( .A(n4548), .Y(n3695) );
  INVXLTS U3194 ( .A(\add_0_root_r1463/SUM[1] ), .Y(n3696) );
  INVXLTS U3195 ( .A(n3696), .Y(n3697) );
  INVXLTS U3196 ( .A(\add_0_root_r1459/SUM[2] ), .Y(n3698) );
  INVXLTS U3197 ( .A(n3698), .Y(n3699) );
  INVXLTS U3198 ( .A(\add_0_root_r1463/SUM[2] ), .Y(n3700) );
  INVXLTS U3199 ( .A(n3700), .Y(n3701) );
  INVXLTS U3200 ( .A(\add_0_root_r1459/SUM[1] ), .Y(n3702) );
  INVXLTS U3201 ( .A(n3702), .Y(n3703) );
  INVXLTS U3202 ( .A(n1585), .Y(n3704) );
  INVXLTS U3203 ( .A(n1955), .Y(n3705) );
  INVXLTS U3204 ( .A(n3705), .Y(n3706) );
  INVX1TS U3205 ( .A(n1910), .Y(n3707) );
  CLKINVX1TS U3206 ( .A(n3707), .Y(n3708) );
  INVXLTS U3207 ( .A(n3659), .Y(n3709) );
  INVXLTS U3208 ( .A(n3659), .Y(n3710) );
  INVX1TS U3209 ( .A(n1999), .Y(n3711) );
  INVXLTS U3210 ( .A(n3711), .Y(n3712) );
  INVXLTS U3211 ( .A(n3650), .Y(n3713) );
  INVXLTS U3212 ( .A(n3650), .Y(n3714) );
  INVXLTS U3213 ( .A(n3679), .Y(n3715) );
  INVXLTS U3214 ( .A(n3679), .Y(n3716) );
  INVXLTS U3215 ( .A(n4598), .Y(n3717) );
  INVXLTS U3216 ( .A(n3717), .Y(n3718) );
  INVXLTS U3217 ( .A(n3717), .Y(n3719) );
  INVXLTS U3218 ( .A(n3704), .Y(n3720) );
  INVXLTS U3219 ( .A(n3720), .Y(n3721) );
  INVXLTS U3220 ( .A(n4619), .Y(n3722) );
  INVXLTS U3221 ( .A(n3722), .Y(n3723) );
  INVXLTS U3222 ( .A(n3722), .Y(n3724) );
  INVXLTS U3223 ( .A(n3671), .Y(n3725) );
  INVXLTS U3224 ( .A(n3671), .Y(n3726) );
  INVXLTS U3225 ( .A(n3662), .Y(n3727) );
  INVXLTS U3226 ( .A(n3662), .Y(n3728) );
  INVXLTS U3227 ( .A(n3661), .Y(n3729) );
  INVXLTS U3228 ( .A(n3661), .Y(n3730) );
  INVXLTS U3229 ( .A(n1865), .Y(n3731) );
  INVXLTS U3230 ( .A(n3731), .Y(n3732) );
  INVXLTS U3231 ( .A(n3673), .Y(n3733) );
  INVXLTS U3232 ( .A(n3673), .Y(n3734) );
  INVXLTS U3233 ( .A(n3675), .Y(n3735) );
  INVXLTS U3234 ( .A(n3675), .Y(n3736) );
  INVXLTS U3235 ( .A(n3672), .Y(n3737) );
  INVXLTS U3236 ( .A(n3672), .Y(n3738) );
  INVXLTS U3237 ( .A(n1641), .Y(n3739) );
  INVXLTS U3238 ( .A(n1641), .Y(n3740) );
  INVXLTS U3239 ( .A(n3684), .Y(n3741) );
  INVXLTS U3240 ( .A(n1554), .Y(n3742) );
  INVXLTS U3241 ( .A(n3742), .Y(n3743) );
  INVXLTS U3242 ( .A(n3744), .Y(n3745) );
  INVXLTS U3243 ( .A(n1621), .Y(n3746) );
  INVXLTS U3244 ( .A(n3746), .Y(n3747) );
  INVXLTS U3245 ( .A(n2205), .Y(n3748) );
  INVXLTS U3246 ( .A(n3748), .Y(n3749) );
  INVXLTS U3247 ( .A(n1604), .Y(n3750) );
  INVXLTS U3248 ( .A(n3750), .Y(n3751) );
  INVXLTS U3249 ( .A(n3692), .Y(n3752) );
  INVXLTS U3250 ( .A(n3692), .Y(n3753) );
  INVXLTS U3251 ( .A(n4539), .Y(n3754) );
  INVXLTS U3252 ( .A(n3660), .Y(n3755) );
  INVXLTS U3253 ( .A(n3660), .Y(n3756) );
  INVXLTS U3254 ( .A(n3651), .Y(n3757) );
  INVXLTS U3255 ( .A(n3651), .Y(n3758) );
  INVXLTS U3256 ( .A(n3652), .Y(n3759) );
  INVXLTS U3257 ( .A(n3652), .Y(n3760) );
  INVXLTS U3258 ( .A(n3663), .Y(n3761) );
  INVXLTS U3259 ( .A(n3663), .Y(n3762) );
  INVXLTS U3260 ( .A(n3676), .Y(n3763) );
  INVXLTS U3261 ( .A(n3676), .Y(n3764) );
  INVXLTS U3262 ( .A(n3664), .Y(n3765) );
  INVXLTS U3263 ( .A(n3664), .Y(n3766) );
  INVXLTS U3264 ( .A(n3665), .Y(n3767) );
  INVXLTS U3265 ( .A(n3665), .Y(n3768) );
  INVXLTS U3266 ( .A(n3674), .Y(n3769) );
  INVXLTS U3267 ( .A(n3674), .Y(n3770) );
  INVXLTS U3268 ( .A(n3807), .Y(n3771) );
  INVXLTS U3269 ( .A(n3808), .Y(n3772) );
  INVXLTS U3270 ( .A(n3823), .Y(n3773) );
  INVXLTS U3271 ( .A(n3824), .Y(n3774) );
  INVXLTS U3272 ( .A(n3829), .Y(n3775) );
  INVXLTS U3273 ( .A(n3830), .Y(n3776) );
  INVXLTS U3274 ( .A(n3648), .Y(n3777) );
  INVXLTS U3275 ( .A(n3648), .Y(n3778) );
  INVXLTS U3276 ( .A(n3648), .Y(n3779) );
  INVXLTS U3277 ( .A(n3647), .Y(n3780) );
  INVXLTS U3278 ( .A(n3647), .Y(n3781) );
  INVXLTS U3279 ( .A(n3647), .Y(n3782) );
  INVXLTS U3280 ( .A(n3657), .Y(n3783) );
  INVXLTS U3281 ( .A(n3657), .Y(n3784) );
  INVXLTS U3282 ( .A(n3657), .Y(n3785) );
  INVXLTS U3283 ( .A(n3649), .Y(n3786) );
  INVXLTS U3284 ( .A(n3649), .Y(n3787) );
  INVXLTS U3285 ( .A(n3649), .Y(n3788) );
  INVXLTS U3286 ( .A(n3658), .Y(n3789) );
  INVXLTS U3287 ( .A(n3658), .Y(n3790) );
  INVXLTS U3288 ( .A(n3658), .Y(n3791) );
  INVXLTS U3289 ( .A(n3667), .Y(n3792) );
  INVXLTS U3290 ( .A(n3667), .Y(n3793) );
  INVXLTS U3291 ( .A(n3667), .Y(n3794) );
  INVXLTS U3292 ( .A(n3668), .Y(n3795) );
  INVXLTS U3293 ( .A(n3668), .Y(n3796) );
  INVXLTS U3294 ( .A(n3668), .Y(n3797) );
  INVXLTS U3295 ( .A(n3670), .Y(n3798) );
  INVXLTS U3296 ( .A(n3670), .Y(n3799) );
  INVXLTS U3297 ( .A(n3670), .Y(n3800) );
  INVXLTS U3298 ( .A(n3669), .Y(n3801) );
  INVXLTS U3299 ( .A(n3669), .Y(n3802) );
  INVXLTS U3300 ( .A(n3669), .Y(n3803) );
  INVXLTS U3301 ( .A(n1752), .Y(n3804) );
  INVXLTS U3302 ( .A(n3804), .Y(n3805) );
  INVXLTS U3303 ( .A(n3804), .Y(n3806) );
  INVXLTS U3304 ( .A(n3690), .Y(n3807) );
  INVXLTS U3305 ( .A(n3690), .Y(n3808) );
  INVXLTS U3306 ( .A(n3660), .Y(n3809) );
  INVXLTS U3307 ( .A(n3809), .Y(n3810) );
  INVXLTS U3308 ( .A(n3809), .Y(n3811) );
  INVXLTS U3309 ( .A(n3792), .Y(n3812) );
  INVXLTS U3310 ( .A(n3794), .Y(n3813) );
  INVXLTS U3311 ( .A(n3796), .Y(n3814) );
  INVXLTS U3312 ( .A(n3797), .Y(n3815) );
  INVXLTS U3313 ( .A(n3799), .Y(n3816) );
  INVXLTS U3314 ( .A(n3800), .Y(n3817) );
  INVXLTS U3315 ( .A(n3802), .Y(n3818) );
  INVXLTS U3316 ( .A(n3803), .Y(n3819) );
  INVXLTS U3317 ( .A(n3827), .Y(n3820) );
  INVXLTS U3318 ( .A(n3825), .Y(n3821) );
  INVXLTS U3319 ( .A(n3653), .Y(n3822) );
  INVXLTS U3320 ( .A(n3653), .Y(n3823) );
  INVXLTS U3321 ( .A(n3653), .Y(n3824) );
  INVXLTS U3322 ( .A(n3654), .Y(n3825) );
  INVXLTS U3323 ( .A(n3654), .Y(n3826) );
  INVXLTS U3324 ( .A(n3654), .Y(n3827) );
  INVXLTS U3325 ( .A(n1926), .Y(n3828) );
  INVXLTS U3326 ( .A(n3828), .Y(n3829) );
  INVXLTS U3327 ( .A(n3828), .Y(n3830) );
  INVXLTS U3328 ( .A(n4043), .Y(n3831) );
  INVXLTS U3329 ( .A(n3831), .Y(n3832) );
  INVXLTS U3330 ( .A(n3831), .Y(n3833) );
  INVXLTS U3331 ( .A(n3831), .Y(n3834) );
  INVXLTS U3332 ( .A(n4045), .Y(n3835) );
  INVXLTS U3333 ( .A(n3835), .Y(n3836) );
  INVXLTS U3334 ( .A(n3835), .Y(n3837) );
  INVXLTS U3335 ( .A(n3835), .Y(n3838) );
  INVXLTS U3336 ( .A(n4047), .Y(n3839) );
  INVXLTS U3337 ( .A(n3839), .Y(n3840) );
  INVXLTS U3338 ( .A(n3839), .Y(n3841) );
  INVXLTS U3339 ( .A(n3839), .Y(n3842) );
  INVXLTS U3340 ( .A(n4049), .Y(n3843) );
  INVXLTS U3341 ( .A(n3843), .Y(n3844) );
  INVXLTS U3342 ( .A(n3843), .Y(n3845) );
  INVXLTS U3343 ( .A(n3843), .Y(n3846) );
  INVXLTS U3344 ( .A(n4051), .Y(n3847) );
  INVXLTS U3345 ( .A(n3847), .Y(n3848) );
  INVXLTS U3346 ( .A(n3847), .Y(n3849) );
  INVXLTS U3347 ( .A(n3847), .Y(n3850) );
  INVXLTS U3348 ( .A(n4053), .Y(n3851) );
  INVXLTS U3349 ( .A(n3851), .Y(n3852) );
  INVXLTS U3350 ( .A(n3851), .Y(n3853) );
  INVXLTS U3351 ( .A(n3851), .Y(n3854) );
  INVXLTS U3352 ( .A(n4055), .Y(n3855) );
  INVXLTS U3353 ( .A(n3855), .Y(n3856) );
  INVXLTS U3354 ( .A(n3855), .Y(n3857) );
  INVXLTS U3355 ( .A(n3855), .Y(n3858) );
  INVXLTS U3356 ( .A(n4057), .Y(n3859) );
  INVXLTS U3357 ( .A(n3859), .Y(n3860) );
  INVXLTS U3358 ( .A(n3859), .Y(n3861) );
  INVXLTS U3359 ( .A(n3859), .Y(n3862) );
  INVXLTS U3360 ( .A(n3656), .Y(n3863) );
  INVXLTS U3361 ( .A(n3656), .Y(n3864) );
  INVXLTS U3362 ( .A(n3656), .Y(n3865) );
  INVXLTS U3363 ( .A(n3656), .Y(n3866) );
  INVXLTS U3364 ( .A(n5786), .Y(n3867) );
  INVXLTS U3365 ( .A(n3867), .Y(n3868) );
  INVXLTS U3366 ( .A(n3867), .Y(n3869) );
  INVXLTS U3367 ( .A(n3867), .Y(n3870) );
  INVXLTS U3368 ( .A(n3867), .Y(n3871) );
  INVXLTS U3369 ( .A(n4621), .Y(n3872) );
  INVXLTS U3370 ( .A(n3872), .Y(n3873) );
  INVXLTS U3371 ( .A(n3872), .Y(n3874) );
  INVXLTS U3372 ( .A(reset), .Y(n3875) );
  INVXLTS U3373 ( .A(n3875), .Y(n3876) );
  INVXLTS U3374 ( .A(requesterAddressIn_NORTH[0]), .Y(n3877) );
  INVXLTS U3375 ( .A(n3877), .Y(n3878) );
  INVXLTS U3376 ( .A(requesterAddressIn_NORTH[1]), .Y(n3879) );
  INVXLTS U3377 ( .A(n3879), .Y(n3880) );
  INVXLTS U3378 ( .A(requesterAddressIn_NORTH[2]), .Y(n3881) );
  INVXLTS U3379 ( .A(n3881), .Y(n3882) );
  INVXLTS U3380 ( .A(requesterAddressIn_NORTH[3]), .Y(n3883) );
  INVXLTS U3381 ( .A(n3883), .Y(n3884) );
  INVXLTS U3382 ( .A(requesterAddressIn_NORTH[4]), .Y(n3885) );
  INVXLTS U3383 ( .A(n3885), .Y(n3886) );
  INVXLTS U3384 ( .A(requesterAddressIn_NORTH[5]), .Y(n3887) );
  INVXLTS U3385 ( .A(n3887), .Y(n3888) );
  INVXLTS U3386 ( .A(dataIn_NORTH[0]), .Y(n3889) );
  INVXLTS U3387 ( .A(n3889), .Y(n3890) );
  INVXLTS U3388 ( .A(dataIn_NORTH[1]), .Y(n3891) );
  INVXLTS U3389 ( .A(n3891), .Y(n3892) );
  INVXLTS U3390 ( .A(dataIn_NORTH[2]), .Y(n3893) );
  INVXLTS U3391 ( .A(n3893), .Y(n3894) );
  INVXLTS U3392 ( .A(dataIn_NORTH[3]), .Y(n3895) );
  INVXLTS U3393 ( .A(n3895), .Y(n3896) );
  INVXLTS U3394 ( .A(dataIn_NORTH[4]), .Y(n3897) );
  INVXLTS U3395 ( .A(n3897), .Y(n3898) );
  INVXLTS U3396 ( .A(dataIn_NORTH[5]), .Y(n3899) );
  INVXLTS U3397 ( .A(n3899), .Y(n3900) );
  INVXLTS U3398 ( .A(dataIn_NORTH[6]), .Y(n3901) );
  INVXLTS U3399 ( .A(n3901), .Y(n3902) );
  INVXLTS U3400 ( .A(dataIn_NORTH[7]), .Y(n3903) );
  INVXLTS U3401 ( .A(n3903), .Y(n3904) );
  INVXLTS U3402 ( .A(dataIn_NORTH[8]), .Y(n3905) );
  INVXLTS U3403 ( .A(n3905), .Y(n3906) );
  INVXLTS U3404 ( .A(dataIn_NORTH[9]), .Y(n3907) );
  INVXLTS U3405 ( .A(n3907), .Y(n3908) );
  INVXLTS U3406 ( .A(dataIn_NORTH[10]), .Y(n3909) );
  INVXLTS U3407 ( .A(n3909), .Y(n3910) );
  INVXLTS U3408 ( .A(dataIn_NORTH[11]), .Y(n3911) );
  INVXLTS U3409 ( .A(n3911), .Y(n3912) );
  INVXLTS U3410 ( .A(dataIn_NORTH[12]), .Y(n3913) );
  INVXLTS U3411 ( .A(n3913), .Y(n3914) );
  INVXLTS U3412 ( .A(dataIn_NORTH[13]), .Y(n3915) );
  INVXLTS U3413 ( .A(n3915), .Y(n3916) );
  INVXLTS U3414 ( .A(dataIn_NORTH[14]), .Y(n3917) );
  INVXLTS U3415 ( .A(n3917), .Y(n3918) );
  INVXLTS U3416 ( .A(dataIn_NORTH[15]), .Y(n3919) );
  INVXLTS U3417 ( .A(n3919), .Y(n3920) );
  INVXLTS U3418 ( .A(dataIn_NORTH[16]), .Y(n3921) );
  INVXLTS U3419 ( .A(n3921), .Y(n3922) );
  INVXLTS U3420 ( .A(dataIn_NORTH[17]), .Y(n3923) );
  INVXLTS U3421 ( .A(n3923), .Y(n3924) );
  INVXLTS U3422 ( .A(dataIn_NORTH[18]), .Y(n3925) );
  INVXLTS U3423 ( .A(n3925), .Y(n3926) );
  INVXLTS U3424 ( .A(dataIn_NORTH[19]), .Y(n3927) );
  INVXLTS U3425 ( .A(n3927), .Y(n3928) );
  INVXLTS U3426 ( .A(dataIn_NORTH[20]), .Y(n3929) );
  INVXLTS U3427 ( .A(n3929), .Y(n3930) );
  INVXLTS U3428 ( .A(dataIn_NORTH[21]), .Y(n3931) );
  INVXLTS U3429 ( .A(n3931), .Y(n3932) );
  INVXLTS U3430 ( .A(dataIn_NORTH[22]), .Y(n3933) );
  INVXLTS U3431 ( .A(n3933), .Y(n3934) );
  INVXLTS U3432 ( .A(dataIn_NORTH[23]), .Y(n3935) );
  INVXLTS U3433 ( .A(n3935), .Y(n3936) );
  INVXLTS U3434 ( .A(dataIn_NORTH[24]), .Y(n3937) );
  INVXLTS U3435 ( .A(n3937), .Y(n3938) );
  INVXLTS U3436 ( .A(dataIn_NORTH[25]), .Y(n3939) );
  INVXLTS U3437 ( .A(n3939), .Y(n3940) );
  INVXLTS U3438 ( .A(dataIn_NORTH[26]), .Y(n3941) );
  INVXLTS U3439 ( .A(n3941), .Y(n3942) );
  INVXLTS U3440 ( .A(dataIn_NORTH[27]), .Y(n3943) );
  INVXLTS U3441 ( .A(n3943), .Y(n3944) );
  INVXLTS U3442 ( .A(dataIn_NORTH[28]), .Y(n3945) );
  INVXLTS U3443 ( .A(n3945), .Y(n3946) );
  INVXLTS U3444 ( .A(dataIn_NORTH[29]), .Y(n3947) );
  INVXLTS U3445 ( .A(n3947), .Y(n3948) );
  INVXLTS U3446 ( .A(dataIn_NORTH[30]), .Y(n3949) );
  INVXLTS U3447 ( .A(n3949), .Y(n3950) );
  INVXLTS U3448 ( .A(dataIn_NORTH[31]), .Y(n3951) );
  INVXLTS U3449 ( .A(n3951), .Y(n3952) );
  INVXLTS U3450 ( .A(requesterAddressIn_SOUTH[0]), .Y(n3953) );
  INVXLTS U3451 ( .A(n3953), .Y(n3954) );
  INVXLTS U3452 ( .A(requesterAddressIn_SOUTH[1]), .Y(n3955) );
  INVXLTS U3453 ( .A(n3955), .Y(n3956) );
  INVXLTS U3454 ( .A(requesterAddressIn_SOUTH[2]), .Y(n3957) );
  INVXLTS U3455 ( .A(n3957), .Y(n3958) );
  INVXLTS U3456 ( .A(requesterAddressIn_SOUTH[3]), .Y(n3959) );
  INVXLTS U3457 ( .A(n3959), .Y(n3960) );
  INVXLTS U3458 ( .A(requesterAddressIn_SOUTH[4]), .Y(n3961) );
  INVXLTS U3459 ( .A(n3961), .Y(n3962) );
  INVXLTS U3460 ( .A(requesterAddressIn_SOUTH[5]), .Y(n3963) );
  INVXLTS U3461 ( .A(n3963), .Y(n3964) );
  INVXLTS U3462 ( .A(memRead_WEST), .Y(n3965) );
  INVXLTS U3463 ( .A(n3965), .Y(n3966) );
  INVXLTS U3464 ( .A(dataIn_SOUTH[0]), .Y(n3967) );
  INVXLTS U3465 ( .A(n3967), .Y(n3968) );
  INVXLTS U3466 ( .A(dataIn_SOUTH[1]), .Y(n3969) );
  INVXLTS U3467 ( .A(n3969), .Y(n3970) );
  INVXLTS U3468 ( .A(dataIn_SOUTH[2]), .Y(n3971) );
  INVXLTS U3469 ( .A(n3971), .Y(n3972) );
  INVXLTS U3470 ( .A(dataIn_SOUTH[3]), .Y(n3973) );
  INVXLTS U3471 ( .A(n3973), .Y(n3974) );
  INVXLTS U3472 ( .A(dataIn_SOUTH[4]), .Y(n3975) );
  INVXLTS U3473 ( .A(n3975), .Y(n3976) );
  INVXLTS U3474 ( .A(dataIn_SOUTH[5]), .Y(n3977) );
  INVXLTS U3475 ( .A(n3977), .Y(n3978) );
  INVXLTS U3476 ( .A(dataIn_SOUTH[6]), .Y(n3979) );
  INVXLTS U3477 ( .A(n3979), .Y(n3980) );
  INVXLTS U3478 ( .A(dataIn_SOUTH[7]), .Y(n3981) );
  INVXLTS U3479 ( .A(n3981), .Y(n3982) );
  INVXLTS U3480 ( .A(dataIn_SOUTH[8]), .Y(n3983) );
  INVXLTS U3481 ( .A(n3983), .Y(n3984) );
  INVXLTS U3482 ( .A(dataIn_SOUTH[9]), .Y(n3985) );
  INVXLTS U3483 ( .A(n3985), .Y(n3986) );
  INVXLTS U3484 ( .A(dataIn_SOUTH[10]), .Y(n3987) );
  INVXLTS U3485 ( .A(n3987), .Y(n3988) );
  INVXLTS U3486 ( .A(dataIn_SOUTH[11]), .Y(n3989) );
  INVXLTS U3487 ( .A(n3989), .Y(n3990) );
  INVXLTS U3488 ( .A(dataIn_SOUTH[12]), .Y(n3991) );
  INVXLTS U3489 ( .A(n3991), .Y(n3992) );
  INVXLTS U3490 ( .A(dataIn_SOUTH[13]), .Y(n3993) );
  INVXLTS U3491 ( .A(n3993), .Y(n3994) );
  INVXLTS U3492 ( .A(dataIn_SOUTH[14]), .Y(n3995) );
  INVXLTS U3493 ( .A(n3995), .Y(n3996) );
  INVXLTS U3494 ( .A(dataIn_SOUTH[15]), .Y(n3997) );
  INVXLTS U3495 ( .A(n3997), .Y(n3998) );
  INVXLTS U3496 ( .A(dataIn_SOUTH[16]), .Y(n3999) );
  INVXLTS U3497 ( .A(n3999), .Y(n4000) );
  INVXLTS U3498 ( .A(dataIn_SOUTH[17]), .Y(n4001) );
  INVXLTS U3499 ( .A(n4001), .Y(n4002) );
  INVXLTS U3500 ( .A(dataIn_SOUTH[18]), .Y(n4003) );
  INVXLTS U3501 ( .A(n4003), .Y(n4004) );
  INVXLTS U3502 ( .A(dataIn_SOUTH[19]), .Y(n4005) );
  INVXLTS U3503 ( .A(n4005), .Y(n4006) );
  INVXLTS U3504 ( .A(dataIn_SOUTH[20]), .Y(n4007) );
  INVXLTS U3505 ( .A(n4007), .Y(n4008) );
  INVXLTS U3506 ( .A(dataIn_SOUTH[21]), .Y(n4009) );
  INVXLTS U3507 ( .A(n4009), .Y(n4010) );
  INVXLTS U3508 ( .A(dataIn_SOUTH[22]), .Y(n4011) );
  INVXLTS U3509 ( .A(n4011), .Y(n4012) );
  INVXLTS U3510 ( .A(dataIn_SOUTH[23]), .Y(n4013) );
  INVXLTS U3511 ( .A(n4013), .Y(n4014) );
  INVXLTS U3512 ( .A(dataIn_SOUTH[24]), .Y(n4015) );
  INVXLTS U3513 ( .A(n4015), .Y(n4016) );
  INVXLTS U3514 ( .A(dataIn_SOUTH[25]), .Y(n4017) );
  INVXLTS U3515 ( .A(n4017), .Y(n4018) );
  INVXLTS U3516 ( .A(dataIn_SOUTH[26]), .Y(n4019) );
  INVXLTS U3517 ( .A(n4019), .Y(n4020) );
  INVXLTS U3518 ( .A(dataIn_SOUTH[27]), .Y(n4021) );
  INVXLTS U3519 ( .A(n4021), .Y(n4022) );
  INVXLTS U3520 ( .A(dataIn_SOUTH[28]), .Y(n4023) );
  INVXLTS U3521 ( .A(n4023), .Y(n4024) );
  INVXLTS U3522 ( .A(dataIn_SOUTH[29]), .Y(n4025) );
  INVXLTS U3523 ( .A(n4025), .Y(n4026) );
  INVXLTS U3524 ( .A(dataIn_SOUTH[30]), .Y(n4027) );
  INVXLTS U3525 ( .A(n4027), .Y(n4028) );
  INVXLTS U3526 ( .A(dataIn_SOUTH[31]), .Y(n4029) );
  INVXLTS U3527 ( .A(n4029), .Y(n4030) );
  INVXLTS U3528 ( .A(requesterAddressIn_WEST[0]), .Y(n4031) );
  INVXLTS U3529 ( .A(n4031), .Y(n4032) );
  INVXLTS U3530 ( .A(requesterAddressIn_WEST[1]), .Y(n4033) );
  INVXLTS U3531 ( .A(n4033), .Y(n4034) );
  INVXLTS U3532 ( .A(requesterAddressIn_WEST[2]), .Y(n4035) );
  INVXLTS U3533 ( .A(n4035), .Y(n4036) );
  INVXLTS U3534 ( .A(requesterAddressIn_WEST[3]), .Y(n4037) );
  INVXLTS U3535 ( .A(n4037), .Y(n4038) );
  INVXLTS U3536 ( .A(requesterAddressIn_WEST[4]), .Y(n4039) );
  INVXLTS U3537 ( .A(n4039), .Y(n4040) );
  INVXLTS U3538 ( .A(requesterAddressIn_WEST[5]), .Y(n4041) );
  INVXLTS U3539 ( .A(n4041), .Y(n4042) );
  INVXLTS U3540 ( .A(cacheAddressIn_EAST[0]), .Y(n4043) );
  INVXLTS U3541 ( .A(n4043), .Y(n4044) );
  INVXLTS U3542 ( .A(cacheAddressIn_EAST[1]), .Y(n4045) );
  INVXLTS U3543 ( .A(n4045), .Y(n4046) );
  INVXLTS U3544 ( .A(cacheAddressIn_EAST[2]), .Y(n4047) );
  INVXLTS U3545 ( .A(n4047), .Y(n4048) );
  INVXLTS U3546 ( .A(cacheAddressIn_EAST[3]), .Y(n4049) );
  INVXLTS U3547 ( .A(n4049), .Y(n4050) );
  INVXLTS U3548 ( .A(cacheAddressIn_EAST[4]), .Y(n4051) );
  INVXLTS U3549 ( .A(n4051), .Y(n4052) );
  INVXLTS U3550 ( .A(cacheAddressIn_EAST[5]), .Y(n4053) );
  INVXLTS U3551 ( .A(n4053), .Y(n4054) );
  INVXLTS U3552 ( .A(cacheAddressIn_EAST[6]), .Y(n4055) );
  INVXLTS U3553 ( .A(n4055), .Y(n4056) );
  INVXLTS U3554 ( .A(cacheAddressIn_EAST[7]), .Y(n4057) );
  INVXLTS U3555 ( .A(n4057), .Y(n4058) );
  INVXLTS U3556 ( .A(requesterAddressIn_EAST[0]), .Y(n4059) );
  INVXLTS U3557 ( .A(n4059), .Y(n4060) );
  INVXLTS U3558 ( .A(n4059), .Y(n4061) );
  INVXLTS U3559 ( .A(requesterAddressIn_EAST[1]), .Y(n4062) );
  INVXLTS U3560 ( .A(n4062), .Y(n4063) );
  INVXLTS U3561 ( .A(n4062), .Y(n4064) );
  INVXLTS U3562 ( .A(requesterAddressIn_EAST[2]), .Y(n4065) );
  INVXLTS U3563 ( .A(n4065), .Y(n4066) );
  INVXLTS U3564 ( .A(n4065), .Y(n4067) );
  INVXLTS U3565 ( .A(requesterAddressIn_EAST[3]), .Y(n4068) );
  INVXLTS U3566 ( .A(n4068), .Y(n4069) );
  INVXLTS U3567 ( .A(n4068), .Y(n4070) );
  INVXLTS U3568 ( .A(requesterAddressIn_EAST[4]), .Y(n4071) );
  INVXLTS U3569 ( .A(n4071), .Y(n4072) );
  INVXLTS U3570 ( .A(n4071), .Y(n4073) );
  INVXLTS U3571 ( .A(requesterAddressIn_EAST[5]), .Y(n4074) );
  INVXLTS U3572 ( .A(n4074), .Y(n4075) );
  INVXLTS U3573 ( .A(n4074), .Y(n4076) );
  INVXLTS U3574 ( .A(cacheAddressIn_NORTH[0]), .Y(n4077) );
  INVXLTS U3575 ( .A(n4077), .Y(n4078) );
  INVXLTS U3576 ( .A(n4077), .Y(n4079) );
  INVXLTS U3577 ( .A(cacheAddressIn_NORTH[1]), .Y(n4080) );
  INVXLTS U3578 ( .A(n4080), .Y(n4081) );
  INVXLTS U3579 ( .A(n4080), .Y(n4082) );
  INVXLTS U3580 ( .A(cacheAddressIn_NORTH[2]), .Y(n4083) );
  INVXLTS U3581 ( .A(n4083), .Y(n4084) );
  INVXLTS U3582 ( .A(n4083), .Y(n4085) );
  INVXLTS U3583 ( .A(cacheAddressIn_NORTH[3]), .Y(n4086) );
  INVXLTS U3584 ( .A(n4086), .Y(n4087) );
  INVXLTS U3585 ( .A(n4086), .Y(n4088) );
  INVXLTS U3586 ( .A(cacheAddressIn_NORTH[4]), .Y(n4089) );
  INVXLTS U3587 ( .A(n4089), .Y(n4090) );
  INVXLTS U3588 ( .A(n4089), .Y(n4091) );
  INVXLTS U3589 ( .A(cacheAddressIn_NORTH[5]), .Y(n4092) );
  INVXLTS U3590 ( .A(n4092), .Y(n4093) );
  INVXLTS U3591 ( .A(n4092), .Y(n4094) );
  INVXLTS U3592 ( .A(cacheAddressIn_NORTH[6]), .Y(n4095) );
  INVXLTS U3593 ( .A(n4095), .Y(n4096) );
  INVXLTS U3594 ( .A(n4095), .Y(n4097) );
  INVXLTS U3595 ( .A(cacheAddressIn_NORTH[7]), .Y(n4098) );
  INVXLTS U3596 ( .A(n4098), .Y(n4099) );
  INVXLTS U3597 ( .A(n4098), .Y(n4100) );
  INVXLTS U3598 ( .A(cacheAddressIn_SOUTH[0]), .Y(n4101) );
  INVXLTS U3599 ( .A(n4101), .Y(n4102) );
  INVXLTS U3600 ( .A(n4101), .Y(n4103) );
  INVXLTS U3601 ( .A(cacheAddressIn_SOUTH[1]), .Y(n4104) );
  INVXLTS U3602 ( .A(n4104), .Y(n4105) );
  INVXLTS U3603 ( .A(n4104), .Y(n4106) );
  INVXLTS U3604 ( .A(cacheAddressIn_SOUTH[2]), .Y(n4107) );
  INVXLTS U3605 ( .A(n4107), .Y(n4108) );
  INVXLTS U3606 ( .A(n4107), .Y(n4109) );
  INVXLTS U3607 ( .A(cacheAddressIn_SOUTH[3]), .Y(n4110) );
  INVXLTS U3608 ( .A(n4110), .Y(n4111) );
  INVXLTS U3609 ( .A(n4110), .Y(n4112) );
  INVXLTS U3610 ( .A(cacheAddressIn_SOUTH[4]), .Y(n4113) );
  INVXLTS U3611 ( .A(n4113), .Y(n4114) );
  INVXLTS U3612 ( .A(n4113), .Y(n4115) );
  INVXLTS U3613 ( .A(cacheAddressIn_SOUTH[5]), .Y(n4116) );
  INVXLTS U3614 ( .A(n4116), .Y(n4117) );
  INVXLTS U3615 ( .A(n4116), .Y(n4118) );
  INVXLTS U3616 ( .A(cacheAddressIn_SOUTH[6]), .Y(n4119) );
  INVXLTS U3617 ( .A(n4119), .Y(n4120) );
  INVXLTS U3618 ( .A(n4119), .Y(n4121) );
  INVXLTS U3619 ( .A(cacheAddressIn_SOUTH[7]), .Y(n4122) );
  INVXLTS U3620 ( .A(n4122), .Y(n4123) );
  INVXLTS U3621 ( .A(n4122), .Y(n4124) );
  INVXLTS U3622 ( .A(cacheAddressIn_WEST[0]), .Y(n4125) );
  INVXLTS U3623 ( .A(n4125), .Y(n4126) );
  INVXLTS U3624 ( .A(n4125), .Y(n4127) );
  INVXLTS U3625 ( .A(n4125), .Y(n4128) );
  INVXLTS U3626 ( .A(cacheAddressIn_WEST[1]), .Y(n4129) );
  INVXLTS U3627 ( .A(n4129), .Y(n4130) );
  INVXLTS U3628 ( .A(n4129), .Y(n4131) );
  INVXLTS U3629 ( .A(n4129), .Y(n4132) );
  INVXLTS U3630 ( .A(cacheAddressIn_WEST[2]), .Y(n4133) );
  INVXLTS U3631 ( .A(n4133), .Y(n4134) );
  INVXLTS U3632 ( .A(n4133), .Y(n4135) );
  INVXLTS U3633 ( .A(n4133), .Y(n4136) );
  INVXLTS U3634 ( .A(cacheAddressIn_WEST[3]), .Y(n4137) );
  INVXLTS U3635 ( .A(n4137), .Y(n4138) );
  INVXLTS U3636 ( .A(n4137), .Y(n4139) );
  INVXLTS U3637 ( .A(n4137), .Y(n4140) );
  INVXLTS U3638 ( .A(cacheAddressIn_WEST[4]), .Y(n4141) );
  INVXLTS U3639 ( .A(n4141), .Y(n4142) );
  INVXLTS U3640 ( .A(n4141), .Y(n4143) );
  INVXLTS U3641 ( .A(n4141), .Y(n4144) );
  INVXLTS U3642 ( .A(cacheAddressIn_WEST[5]), .Y(n4145) );
  INVXLTS U3643 ( .A(n4145), .Y(n4146) );
  INVXLTS U3644 ( .A(n4145), .Y(n4147) );
  INVXLTS U3645 ( .A(n4145), .Y(n4148) );
  INVXLTS U3646 ( .A(cacheAddressIn_WEST[6]), .Y(n4149) );
  INVXLTS U3647 ( .A(n4149), .Y(n4150) );
  INVXLTS U3648 ( .A(n4149), .Y(n4151) );
  INVXLTS U3649 ( .A(n4149), .Y(n4152) );
  INVXLTS U3650 ( .A(cacheAddressIn_WEST[7]), .Y(n4153) );
  INVXLTS U3651 ( .A(n4153), .Y(n4154) );
  INVXLTS U3652 ( .A(n4153), .Y(n4155) );
  INVXLTS U3653 ( .A(n4153), .Y(n4156) );
  INVXLTS U3654 ( .A(dataIn_WEST[0]), .Y(n4157) );
  INVXLTS U3655 ( .A(n4157), .Y(n4158) );
  INVXLTS U3656 ( .A(n4157), .Y(n4159) );
  INVXLTS U3657 ( .A(n4157), .Y(n4160) );
  INVXLTS U3658 ( .A(dataIn_WEST[1]), .Y(n4161) );
  INVXLTS U3659 ( .A(n4161), .Y(n4162) );
  INVXLTS U3660 ( .A(n4161), .Y(n4163) );
  INVXLTS U3661 ( .A(n4161), .Y(n4164) );
  INVXLTS U3662 ( .A(dataIn_WEST[2]), .Y(n4165) );
  INVXLTS U3663 ( .A(n4165), .Y(n4166) );
  INVXLTS U3664 ( .A(n4165), .Y(n4167) );
  INVXLTS U3665 ( .A(n4165), .Y(n4168) );
  INVXLTS U3666 ( .A(dataIn_WEST[3]), .Y(n4169) );
  INVXLTS U3667 ( .A(n4169), .Y(n4170) );
  INVXLTS U3668 ( .A(n4169), .Y(n4171) );
  INVXLTS U3669 ( .A(n4169), .Y(n4172) );
  INVXLTS U3670 ( .A(dataIn_WEST[4]), .Y(n4173) );
  INVXLTS U3671 ( .A(n4173), .Y(n4174) );
  INVXLTS U3672 ( .A(n4173), .Y(n4175) );
  INVXLTS U3673 ( .A(n4173), .Y(n4176) );
  INVXLTS U3674 ( .A(dataIn_WEST[5]), .Y(n4177) );
  INVXLTS U3675 ( .A(n4177), .Y(n4178) );
  INVXLTS U3676 ( .A(n4177), .Y(n4179) );
  INVXLTS U3677 ( .A(n4177), .Y(n4180) );
  INVXLTS U3678 ( .A(dataIn_WEST[6]), .Y(n4181) );
  INVXLTS U3679 ( .A(n4181), .Y(n4182) );
  INVXLTS U3680 ( .A(n4181), .Y(n4183) );
  INVXLTS U3681 ( .A(n4181), .Y(n4184) );
  INVXLTS U3682 ( .A(dataIn_WEST[7]), .Y(n4185) );
  INVXLTS U3683 ( .A(n4185), .Y(n4186) );
  INVXLTS U3684 ( .A(n4185), .Y(n4187) );
  INVXLTS U3685 ( .A(n4185), .Y(n4188) );
  INVXLTS U3686 ( .A(dataIn_WEST[8]), .Y(n4189) );
  INVXLTS U3687 ( .A(n4189), .Y(n4190) );
  INVXLTS U3688 ( .A(n4189), .Y(n4191) );
  INVXLTS U3689 ( .A(n4189), .Y(n4192) );
  INVXLTS U3690 ( .A(dataIn_WEST[9]), .Y(n4193) );
  INVXLTS U3691 ( .A(n4193), .Y(n4194) );
  INVXLTS U3692 ( .A(n4193), .Y(n4195) );
  INVXLTS U3693 ( .A(n4193), .Y(n4196) );
  INVXLTS U3694 ( .A(dataIn_WEST[10]), .Y(n4197) );
  INVXLTS U3695 ( .A(n4197), .Y(n4198) );
  INVXLTS U3696 ( .A(n4197), .Y(n4199) );
  INVXLTS U3697 ( .A(n4197), .Y(n4200) );
  INVXLTS U3698 ( .A(dataIn_WEST[11]), .Y(n4201) );
  INVXLTS U3699 ( .A(n4201), .Y(n4202) );
  INVXLTS U3700 ( .A(n4201), .Y(n4203) );
  INVXLTS U3701 ( .A(n4201), .Y(n4204) );
  INVXLTS U3702 ( .A(dataIn_WEST[12]), .Y(n4205) );
  INVXLTS U3703 ( .A(n4205), .Y(n4206) );
  INVXLTS U3704 ( .A(n4205), .Y(n4207) );
  INVXLTS U3705 ( .A(n4205), .Y(n4208) );
  INVXLTS U3706 ( .A(dataIn_WEST[13]), .Y(n4209) );
  INVXLTS U3707 ( .A(n4209), .Y(n4210) );
  INVXLTS U3708 ( .A(n4209), .Y(n4211) );
  INVXLTS U3709 ( .A(n4209), .Y(n4212) );
  INVXLTS U3710 ( .A(dataIn_WEST[14]), .Y(n4213) );
  INVXLTS U3711 ( .A(n4213), .Y(n4214) );
  INVXLTS U3712 ( .A(n4213), .Y(n4215) );
  INVXLTS U3713 ( .A(n4213), .Y(n4216) );
  INVXLTS U3714 ( .A(dataIn_WEST[15]), .Y(n4217) );
  INVXLTS U3715 ( .A(n4217), .Y(n4218) );
  INVXLTS U3716 ( .A(n4217), .Y(n4219) );
  INVXLTS U3717 ( .A(n4217), .Y(n4220) );
  INVXLTS U3718 ( .A(dataIn_WEST[16]), .Y(n4221) );
  INVXLTS U3719 ( .A(n4221), .Y(n4222) );
  INVXLTS U3720 ( .A(n4221), .Y(n4223) );
  INVXLTS U3721 ( .A(n4221), .Y(n4224) );
  INVXLTS U3722 ( .A(dataIn_WEST[17]), .Y(n4225) );
  INVXLTS U3723 ( .A(n4225), .Y(n4226) );
  INVXLTS U3724 ( .A(n4225), .Y(n4227) );
  INVXLTS U3725 ( .A(n4225), .Y(n4228) );
  INVXLTS U3726 ( .A(dataIn_WEST[18]), .Y(n4229) );
  INVXLTS U3727 ( .A(n4229), .Y(n4230) );
  INVXLTS U3728 ( .A(n4229), .Y(n4231) );
  INVXLTS U3729 ( .A(n4229), .Y(n4232) );
  INVXLTS U3730 ( .A(dataIn_WEST[19]), .Y(n4233) );
  INVXLTS U3731 ( .A(n4233), .Y(n4234) );
  INVXLTS U3732 ( .A(n4233), .Y(n4235) );
  INVXLTS U3733 ( .A(n4233), .Y(n4236) );
  INVXLTS U3734 ( .A(dataIn_WEST[20]), .Y(n4237) );
  INVXLTS U3735 ( .A(n4237), .Y(n4238) );
  INVXLTS U3736 ( .A(n4237), .Y(n4239) );
  INVXLTS U3737 ( .A(n4237), .Y(n4240) );
  INVXLTS U3738 ( .A(dataIn_WEST[21]), .Y(n4241) );
  INVXLTS U3739 ( .A(n4241), .Y(n4242) );
  INVXLTS U3740 ( .A(n4241), .Y(n4243) );
  INVXLTS U3741 ( .A(n4241), .Y(n4244) );
  INVXLTS U3742 ( .A(dataIn_WEST[22]), .Y(n4245) );
  INVXLTS U3743 ( .A(n4245), .Y(n4246) );
  INVXLTS U3744 ( .A(n4245), .Y(n4247) );
  INVXLTS U3745 ( .A(n4245), .Y(n4248) );
  INVXLTS U3746 ( .A(dataIn_WEST[23]), .Y(n4249) );
  INVXLTS U3747 ( .A(n4249), .Y(n4250) );
  INVXLTS U3748 ( .A(n4249), .Y(n4251) );
  INVXLTS U3749 ( .A(n4249), .Y(n4252) );
  INVXLTS U3750 ( .A(dataIn_WEST[24]), .Y(n4253) );
  INVXLTS U3751 ( .A(n4253), .Y(n4254) );
  INVXLTS U3752 ( .A(n4253), .Y(n4255) );
  INVXLTS U3753 ( .A(n4253), .Y(n4256) );
  INVXLTS U3754 ( .A(dataIn_WEST[25]), .Y(n4257) );
  INVXLTS U3755 ( .A(n4257), .Y(n4258) );
  INVXLTS U3756 ( .A(n4257), .Y(n4259) );
  INVXLTS U3757 ( .A(n4257), .Y(n4260) );
  INVXLTS U3758 ( .A(dataIn_WEST[26]), .Y(n4261) );
  INVXLTS U3759 ( .A(n4261), .Y(n4262) );
  INVXLTS U3760 ( .A(n4261), .Y(n4263) );
  INVXLTS U3761 ( .A(n4261), .Y(n4264) );
  INVXLTS U3762 ( .A(dataIn_WEST[27]), .Y(n4265) );
  INVXLTS U3763 ( .A(n4265), .Y(n4266) );
  INVXLTS U3764 ( .A(n4265), .Y(n4267) );
  INVXLTS U3765 ( .A(n4265), .Y(n4268) );
  INVXLTS U3766 ( .A(dataIn_WEST[28]), .Y(n4269) );
  INVXLTS U3767 ( .A(n4269), .Y(n4270) );
  INVXLTS U3768 ( .A(n4269), .Y(n4271) );
  INVXLTS U3769 ( .A(n4269), .Y(n4272) );
  INVXLTS U3770 ( .A(dataIn_WEST[29]), .Y(n4273) );
  INVXLTS U3771 ( .A(n4273), .Y(n4274) );
  INVXLTS U3772 ( .A(n4273), .Y(n4275) );
  INVXLTS U3773 ( .A(n4273), .Y(n4276) );
  INVXLTS U3774 ( .A(dataIn_WEST[30]), .Y(n4277) );
  INVXLTS U3775 ( .A(n4277), .Y(n4278) );
  INVXLTS U3776 ( .A(n4277), .Y(n4279) );
  INVXLTS U3777 ( .A(n4277), .Y(n4280) );
  INVXLTS U3778 ( .A(dataIn_WEST[31]), .Y(n4281) );
  INVXLTS U3779 ( .A(n4281), .Y(n4282) );
  INVXLTS U3780 ( .A(n4281), .Y(n4283) );
  INVXLTS U3781 ( .A(n4281), .Y(n4284) );
  INVXLTS U3782 ( .A(memWrite_WEST), .Y(n4285) );
  INVXLTS U3783 ( .A(n4285), .Y(n4286) );
  INVXLTS U3784 ( .A(n4285), .Y(n4287) );
  INVXLTS U3785 ( .A(n4285), .Y(n4288) );
  INVXLTS U3786 ( .A(dataIn_EAST[0]), .Y(n4289) );
  INVXLTS U3787 ( .A(n4289), .Y(n4290) );
  INVXLTS U3788 ( .A(n4289), .Y(n4291) );
  INVXLTS U3789 ( .A(n4289), .Y(n4292) );
  INVXLTS U3790 ( .A(n4289), .Y(n4293) );
  INVXLTS U3791 ( .A(dataIn_EAST[1]), .Y(n4294) );
  INVXLTS U3792 ( .A(n4294), .Y(n4295) );
  INVXLTS U3793 ( .A(n4294), .Y(n4296) );
  INVXLTS U3794 ( .A(n4294), .Y(n4297) );
  INVXLTS U3795 ( .A(n4294), .Y(n4298) );
  INVXLTS U3796 ( .A(dataIn_EAST[2]), .Y(n4299) );
  INVXLTS U3797 ( .A(n4299), .Y(n4300) );
  INVXLTS U3798 ( .A(n4299), .Y(n4301) );
  INVXLTS U3799 ( .A(n4299), .Y(n4302) );
  INVXLTS U3800 ( .A(n4299), .Y(n4303) );
  INVXLTS U3801 ( .A(dataIn_EAST[3]), .Y(n4304) );
  INVXLTS U3802 ( .A(n4304), .Y(n4305) );
  INVXLTS U3803 ( .A(n4304), .Y(n4306) );
  INVXLTS U3804 ( .A(n4304), .Y(n4307) );
  INVXLTS U3805 ( .A(n4304), .Y(n4308) );
  INVXLTS U3806 ( .A(dataIn_EAST[4]), .Y(n4309) );
  INVXLTS U3807 ( .A(n4309), .Y(n4310) );
  INVXLTS U3808 ( .A(n4309), .Y(n4311) );
  INVXLTS U3809 ( .A(n4309), .Y(n4312) );
  INVXLTS U3810 ( .A(n4309), .Y(n4313) );
  INVXLTS U3811 ( .A(dataIn_EAST[5]), .Y(n4314) );
  INVXLTS U3812 ( .A(n4314), .Y(n4315) );
  INVXLTS U3813 ( .A(n4314), .Y(n4316) );
  INVXLTS U3814 ( .A(n4314), .Y(n4317) );
  INVXLTS U3815 ( .A(n4314), .Y(n4318) );
  INVXLTS U3816 ( .A(dataIn_EAST[6]), .Y(n4319) );
  INVXLTS U3817 ( .A(n4319), .Y(n4320) );
  INVXLTS U3818 ( .A(n4319), .Y(n4321) );
  INVXLTS U3819 ( .A(n4319), .Y(n4322) );
  INVXLTS U3820 ( .A(n4319), .Y(n4323) );
  INVXLTS U3821 ( .A(dataIn_EAST[7]), .Y(n4324) );
  INVXLTS U3822 ( .A(n4324), .Y(n4325) );
  INVXLTS U3823 ( .A(n4324), .Y(n4326) );
  INVXLTS U3824 ( .A(n4324), .Y(n4327) );
  INVXLTS U3825 ( .A(n4324), .Y(n4328) );
  INVXLTS U3826 ( .A(dataIn_EAST[8]), .Y(n4329) );
  INVXLTS U3827 ( .A(n4329), .Y(n4330) );
  INVXLTS U3828 ( .A(n4329), .Y(n4331) );
  INVXLTS U3829 ( .A(n4329), .Y(n4332) );
  INVXLTS U3830 ( .A(n4329), .Y(n4333) );
  INVXLTS U3831 ( .A(dataIn_EAST[9]), .Y(n4334) );
  INVXLTS U3832 ( .A(n4334), .Y(n4335) );
  INVXLTS U3833 ( .A(n4334), .Y(n4336) );
  INVXLTS U3834 ( .A(n4334), .Y(n4337) );
  INVXLTS U3835 ( .A(n4334), .Y(n4338) );
  INVXLTS U3836 ( .A(dataIn_EAST[10]), .Y(n4339) );
  INVXLTS U3837 ( .A(n4339), .Y(n4340) );
  INVXLTS U3838 ( .A(n4339), .Y(n4341) );
  INVXLTS U3839 ( .A(n4339), .Y(n4342) );
  INVXLTS U3840 ( .A(n4339), .Y(n4343) );
  INVXLTS U3841 ( .A(dataIn_EAST[11]), .Y(n4344) );
  INVXLTS U3842 ( .A(n4344), .Y(n4345) );
  INVXLTS U3843 ( .A(n4344), .Y(n4346) );
  INVXLTS U3844 ( .A(n4344), .Y(n4347) );
  INVXLTS U3845 ( .A(n4344), .Y(n4348) );
  INVXLTS U3846 ( .A(dataIn_EAST[12]), .Y(n4349) );
  INVXLTS U3847 ( .A(n4349), .Y(n4350) );
  INVXLTS U3848 ( .A(n4349), .Y(n4351) );
  INVXLTS U3849 ( .A(n4349), .Y(n4352) );
  INVXLTS U3850 ( .A(n4349), .Y(n4353) );
  INVXLTS U3851 ( .A(dataIn_EAST[13]), .Y(n4354) );
  INVXLTS U3852 ( .A(n4354), .Y(n4355) );
  INVXLTS U3853 ( .A(n4354), .Y(n4356) );
  INVXLTS U3854 ( .A(n4354), .Y(n4357) );
  INVXLTS U3855 ( .A(n4354), .Y(n4358) );
  INVXLTS U3856 ( .A(dataIn_EAST[14]), .Y(n4359) );
  INVXLTS U3857 ( .A(n4359), .Y(n4360) );
  INVXLTS U3858 ( .A(n4359), .Y(n4361) );
  INVXLTS U3859 ( .A(n4359), .Y(n4362) );
  INVXLTS U3860 ( .A(n4359), .Y(n4363) );
  INVXLTS U3861 ( .A(dataIn_EAST[15]), .Y(n4364) );
  INVXLTS U3862 ( .A(n4364), .Y(n4365) );
  INVXLTS U3863 ( .A(n4364), .Y(n4366) );
  INVXLTS U3864 ( .A(n4364), .Y(n4367) );
  INVXLTS U3865 ( .A(n4364), .Y(n4368) );
  INVXLTS U3866 ( .A(dataIn_EAST[16]), .Y(n4369) );
  INVXLTS U3867 ( .A(n4369), .Y(n4370) );
  INVXLTS U3868 ( .A(n4369), .Y(n4371) );
  INVXLTS U3869 ( .A(n4369), .Y(n4372) );
  INVXLTS U3870 ( .A(n4369), .Y(n4373) );
  INVXLTS U3871 ( .A(dataIn_EAST[17]), .Y(n4374) );
  INVXLTS U3872 ( .A(n4374), .Y(n4375) );
  INVXLTS U3873 ( .A(n4374), .Y(n4376) );
  INVXLTS U3874 ( .A(n4374), .Y(n4377) );
  INVXLTS U3875 ( .A(n4374), .Y(n4378) );
  INVXLTS U3876 ( .A(dataIn_EAST[18]), .Y(n4379) );
  INVXLTS U3877 ( .A(n4379), .Y(n4380) );
  INVXLTS U3878 ( .A(n4379), .Y(n4381) );
  INVXLTS U3879 ( .A(n4379), .Y(n4382) );
  INVXLTS U3880 ( .A(n4379), .Y(n4383) );
  INVXLTS U3881 ( .A(dataIn_EAST[19]), .Y(n4384) );
  INVXLTS U3882 ( .A(n4384), .Y(n4385) );
  INVXLTS U3883 ( .A(n4384), .Y(n4386) );
  INVXLTS U3884 ( .A(n4384), .Y(n4387) );
  INVXLTS U3885 ( .A(n4384), .Y(n4388) );
  INVXLTS U3886 ( .A(dataIn_EAST[20]), .Y(n4389) );
  INVXLTS U3887 ( .A(n4389), .Y(n4390) );
  INVXLTS U3888 ( .A(n4389), .Y(n4391) );
  INVXLTS U3889 ( .A(n4389), .Y(n4392) );
  INVXLTS U3890 ( .A(n4389), .Y(n4393) );
  INVXLTS U3891 ( .A(dataIn_EAST[21]), .Y(n4394) );
  INVXLTS U3892 ( .A(n4394), .Y(n4395) );
  INVXLTS U3893 ( .A(n4394), .Y(n4396) );
  INVXLTS U3894 ( .A(n4394), .Y(n4397) );
  INVXLTS U3895 ( .A(n4394), .Y(n4398) );
  INVXLTS U3896 ( .A(dataIn_EAST[22]), .Y(n4399) );
  INVXLTS U3897 ( .A(n4399), .Y(n4400) );
  INVXLTS U3898 ( .A(n4399), .Y(n4401) );
  INVXLTS U3899 ( .A(n4399), .Y(n4402) );
  INVXLTS U3900 ( .A(n4399), .Y(n4403) );
  INVXLTS U3901 ( .A(dataIn_EAST[23]), .Y(n4404) );
  INVXLTS U3902 ( .A(n4404), .Y(n4405) );
  INVXLTS U3903 ( .A(n4404), .Y(n4406) );
  INVXLTS U3904 ( .A(n4404), .Y(n4407) );
  INVXLTS U3905 ( .A(n4404), .Y(n4408) );
  INVXLTS U3906 ( .A(dataIn_EAST[24]), .Y(n4409) );
  INVXLTS U3907 ( .A(n4409), .Y(n4410) );
  INVXLTS U3908 ( .A(n4409), .Y(n4411) );
  INVXLTS U3909 ( .A(n4409), .Y(n4412) );
  INVXLTS U3910 ( .A(n4409), .Y(n4413) );
  INVXLTS U3911 ( .A(dataIn_EAST[25]), .Y(n4414) );
  INVXLTS U3912 ( .A(n4414), .Y(n4415) );
  INVXLTS U3913 ( .A(n4414), .Y(n4416) );
  INVXLTS U3914 ( .A(n4414), .Y(n4417) );
  INVXLTS U3915 ( .A(n4414), .Y(n4418) );
  INVXLTS U3916 ( .A(dataIn_EAST[26]), .Y(n4419) );
  INVXLTS U3917 ( .A(n4419), .Y(n4420) );
  INVXLTS U3918 ( .A(n4419), .Y(n4421) );
  INVXLTS U3919 ( .A(n4419), .Y(n4422) );
  INVXLTS U3920 ( .A(n4419), .Y(n4423) );
  INVXLTS U3921 ( .A(dataIn_EAST[27]), .Y(n4424) );
  INVXLTS U3922 ( .A(n4424), .Y(n4425) );
  INVXLTS U3923 ( .A(n4424), .Y(n4426) );
  INVXLTS U3924 ( .A(n4424), .Y(n4427) );
  INVXLTS U3925 ( .A(n4424), .Y(n4428) );
  INVXLTS U3926 ( .A(dataIn_EAST[28]), .Y(n4429) );
  INVXLTS U3927 ( .A(n4429), .Y(n4430) );
  INVXLTS U3928 ( .A(n4429), .Y(n4431) );
  INVXLTS U3929 ( .A(n4429), .Y(n4432) );
  INVXLTS U3930 ( .A(n4429), .Y(n4433) );
  INVXLTS U3931 ( .A(dataIn_EAST[29]), .Y(n4434) );
  INVXLTS U3932 ( .A(n4434), .Y(n4435) );
  INVXLTS U3933 ( .A(n4434), .Y(n4436) );
  INVXLTS U3934 ( .A(n4434), .Y(n4437) );
  INVXLTS U3935 ( .A(n4434), .Y(n4438) );
  INVXLTS U3936 ( .A(dataIn_EAST[30]), .Y(n4439) );
  INVXLTS U3937 ( .A(n4439), .Y(n4440) );
  INVXLTS U3938 ( .A(n4439), .Y(n4441) );
  INVXLTS U3939 ( .A(n4439), .Y(n4442) );
  INVXLTS U3940 ( .A(n4439), .Y(n4443) );
  INVXLTS U3941 ( .A(dataIn_EAST[31]), .Y(n4444) );
  INVXLTS U3942 ( .A(n4444), .Y(n4445) );
  INVXLTS U3943 ( .A(n4444), .Y(n4446) );
  INVXLTS U3944 ( .A(n4444), .Y(n4447) );
  INVXLTS U3945 ( .A(n4444), .Y(n4448) );
  CLKBUFX2TS U4010 ( .A(n1871), .Y(n4513) );
  CLKBUFX2TS U4011 ( .A(n1871), .Y(n4514) );
  OAI211XLTS U4012 ( .A0(n3732), .A1(n3708), .B0(n1911), .C0(n1912), .Y(n1871)
         );
  CLKBUFX2TS U4013 ( .A(n1826), .Y(n4515) );
  CLKBUFX2TS U4014 ( .A(n1826), .Y(n4516) );
  CLKBUFX2TS U4015 ( .A(n2004), .Y(n4517) );
  CLKBUFX2TS U4016 ( .A(n2004), .Y(n4518) );
  INVX2TS U4017 ( .A(n5760), .Y(n4519) );
  AND3XLTS U4018 ( .A(n2426), .B(n5772), .C(n5773), .Y(n2280) );
  CLKBUFX2TS U4019 ( .A(prevRequesterPort_B[0]), .Y(n4520) );
  CLKBUFX2TS U4020 ( .A(n2047), .Y(n4521) );
  CLKBUFX2TS U4021 ( .A(n2047), .Y(n4522) );
  OAI211XLTS U4022 ( .A0(n3732), .A1(n2085), .B0(n5410), .C0(n2086), .Y(n2047)
         );
  CLKBUFX2TS U4023 ( .A(prevRequesterPort_B[1]), .Y(n4523) );
  CLKBUFX2TS U4024 ( .A(n1590), .Y(n4524) );
  CLKBUFX2TS U4025 ( .A(totalAccesses[1]), .Y(n4525) );
  AND2X2TS U4026 ( .A(n1960), .B(n5720), .Y(n1962) );
  INVX2TS U4027 ( .A(n1962), .Y(n4526) );
  INVX2TS U4028 ( .A(n1962), .Y(n4527) );
  CLKBUFX2TS U4029 ( .A(n1915), .Y(n4528) );
  CLKBUFX2TS U4030 ( .A(n1915), .Y(n4529) );
  OAI211XLTS U4031 ( .A0(n1865), .A1(n3706), .B0(n5291), .C0(n1956), .Y(n1915)
         );
  CLKBUFX2TS U4032 ( .A(n1545), .Y(n4530) );
  INVX2TS U4033 ( .A(n5806), .Y(n4531) );
  INVX2TS U4034 ( .A(n4561), .Y(n4532) );
  CLKBUFX2TS U4035 ( .A(n1588), .Y(n4533) );
  INVX2TS U4036 ( .A(n5973), .Y(n4534) );
  NOR2X1TS U4037 ( .A(n3873), .B(n4691), .Y(n1740) );
  CLKBUFX2TS U4038 ( .A(n1960), .Y(n4535) );
  CLKBUFX2TS U4039 ( .A(n1960), .Y(n4536) );
  OAI22XLTS U4040 ( .A0(n4536), .A1(n1209), .B0(n1961), .B1(n4527), .Y(n3310)
         );
  OAI22XLTS U4041 ( .A0(n4535), .A1(n1210), .B0(n1971), .B1(n4527), .Y(n3311)
         );
  OAI22XLTS U4042 ( .A0(n4535), .A1(n1211), .B0(n1975), .B1(n4527), .Y(n3312)
         );
  OAI22XLTS U4043 ( .A0(n4536), .A1(n1212), .B0(n1979), .B1(n4527), .Y(n3313)
         );
  OAI22XLTS U4044 ( .A0(n4535), .A1(n1213), .B0(n1983), .B1(n4526), .Y(n3314)
         );
  OAI22XLTS U4045 ( .A0(n4536), .A1(n1214), .B0(n1987), .B1(n4526), .Y(n3315)
         );
  OAI22XLTS U4046 ( .A0(n4536), .A1(n1215), .B0(n1991), .B1(n4526), .Y(n3316)
         );
  OAI22XLTS U4047 ( .A0(n4535), .A1(n1216), .B0(n1995), .B1(n4526), .Y(n3317)
         );
  CLKBUFX2TS U4048 ( .A(n1528), .Y(n4537) );
  CLKBUFX2TS U4049 ( .A(N10004), .Y(n4538) );
  CLKBUFX2TS U4050 ( .A(n2130), .Y(n4539) );
  CLKBUFX2TS U4051 ( .A(n5797), .Y(n4540) );
  AND2X2TS U4052 ( .A(n2047), .B(n5720), .Y(n2049) );
  INVX2TS U4053 ( .A(n2049), .Y(n4541) );
  INVX2TS U4054 ( .A(n2049), .Y(n4542) );
  INVX2TS U4055 ( .A(n5972), .Y(n4543) );
  AOI21X1TS U4056 ( .A0(n5690), .A1(N6314), .B0(n5409), .Y(n1783) );
  INVX2TS U4057 ( .A(n4610), .Y(n4544) );
  INVX2TS U4058 ( .A(n4610), .Y(n4545) );
  AOI21XLTS U4059 ( .A0(n4545), .A1(n5768), .B0(n5740), .Y(n2249) );
  INVX1TS U4060 ( .A(n1823), .Y(n4546) );
  CLKBUFX2TS U4061 ( .A(n1748), .Y(n4547) );
  CLKBUFX2TS U4062 ( .A(\add_0_root_r1463/B[4] ), .Y(n4548) );
  OAI22X1TS U4063 ( .A0(n4617), .A1(n3745), .B0(n4608), .B1(n3156), .Y(N589)
         );
  CLKBUFX2TS U4064 ( .A(n1620), .Y(n4549) );
  CLKBUFX2TS U4065 ( .A(n5799), .Y(n4550) );
  INVX2TS U4066 ( .A(n5975), .Y(n4551) );
  AND2X2TS U4067 ( .A(n4514), .B(n5719), .Y(n1873) );
  INVX2TS U4068 ( .A(n1873), .Y(n4552) );
  INVX2TS U4069 ( .A(n1873), .Y(n4553) );
  AND2X2TS U4070 ( .A(n4585), .B(n5721), .Y(n2093) );
  INVX2TS U4071 ( .A(n2093), .Y(n4554) );
  INVX2TS U4072 ( .A(n2093), .Y(n4555) );
  AND2X2TS U4073 ( .A(n1915), .B(n5720), .Y(n1917) );
  INVX2TS U4074 ( .A(n1917), .Y(n4556) );
  INVX2TS U4075 ( .A(n1917), .Y(n4557) );
  AND2X2TS U4076 ( .A(n4582), .B(n5561), .Y(n1599) );
  INVX2TS U4077 ( .A(n1599), .Y(n4558) );
  INVX2TS U4078 ( .A(n1599), .Y(n4559) );
  INVX2TS U4079 ( .A(n5804), .Y(n4560) );
  CLKBUFX2TS U4080 ( .A(n1573), .Y(n5801) );
  INVX2TS U4081 ( .A(n5801), .Y(n4561) );
  INVX2TS U4082 ( .A(n5801), .Y(n4562) );
  INVX2TS U4083 ( .A(n5801), .Y(n4563) );
  CLKBUFX2TS U4084 ( .A(n3874), .Y(N6314) );
  INVX2TS U4085 ( .A(N6314), .Y(n4564) );
  INVX2TS U4086 ( .A(N6314), .Y(n4565) );
  NOR2BX1TS U4087 ( .AN(\r1472/carry[3] ), .B(n3680), .Y(n2117) );
  NOR2BX1TS U4088 ( .AN(\r1471/carry[3] ), .B(n3680), .Y(n2120) );
  NOR2BX1TS U4089 ( .AN(\r1470/carry[3] ), .B(n4564), .Y(n2121) );
  AND2X2TS U4090 ( .A(n5560), .B(n3724), .Y(n2089) );
  INVX2TS U4091 ( .A(n2089), .Y(n4566) );
  INVX2TS U4092 ( .A(n2089), .Y(n4567) );
  INVX2TS U4093 ( .A(n2089), .Y(n4568) );
  INVX2TS U4094 ( .A(n2089), .Y(n4569) );
  CLKBUFX2TS U4095 ( .A(n1555), .Y(n4570) );
  CLKBUFX2TS U4096 ( .A(n1536), .Y(n4571) );
  AND2X2TS U4097 ( .A(n1826), .B(n5719), .Y(n1828) );
  INVX2TS U4098 ( .A(n1828), .Y(n4572) );
  INVX2TS U4099 ( .A(n1828), .Y(n4573) );
  AND2X2TS U4100 ( .A(n2004), .B(n5720), .Y(n2006) );
  INVX2TS U4101 ( .A(n2006), .Y(n4574) );
  INVX2TS U4102 ( .A(n2006), .Y(n4575) );
  NOR2X1TS U4103 ( .A(n1586), .B(n5802), .Y(n1567) );
  INVX2TS U4104 ( .A(n1567), .Y(n4576) );
  INVX2TS U4105 ( .A(n1567), .Y(n4577) );
  INVX2TS U4106 ( .A(n5776), .Y(n4578) );
  OR2X2TS U4107 ( .A(n3693), .B(n3645), .Y(n1530) );
  INVX2TS U4108 ( .A(n1530), .Y(n4579) );
  INVX2TS U4109 ( .A(n1530), .Y(n4580) );
  INVX2TS U4110 ( .A(n1530), .Y(n4581) );
  OR2X2TS U4111 ( .A(n1794), .B(n5733), .Y(n1600) );
  INVX2TS U4112 ( .A(n1600), .Y(n4582) );
  INVX2TS U4113 ( .A(n1600), .Y(n4583) );
  INVX2TS U4114 ( .A(n1600), .Y(n4584) );
  AND3X2TS U4115 ( .A(n2281), .B(n3726), .C(N10004), .Y(n2091) );
  INVX2TS U4116 ( .A(n2091), .Y(n4585) );
  INVX2TS U4117 ( .A(n2091), .Y(n4586) );
  INVX2TS U4118 ( .A(n2091), .Y(n4587) );
  CLKBUFX2TS U4119 ( .A(n1618), .Y(n4588) );
  CLKBUFX2TS U4120 ( .A(n1618), .Y(n4589) );
  CLKBUFX2TS U4121 ( .A(n2255), .Y(n5874) );
  INVX2TS U4122 ( .A(n5874), .Y(n4590) );
  INVX2TS U4123 ( .A(n5874), .Y(n4591) );
  INVX2TS U4124 ( .A(n5874), .Y(n4592) );
  INVX2TS U4125 ( .A(n3873), .Y(n4593) );
  INVX2TS U4126 ( .A(n3874), .Y(n4594) );
  INVX2TS U4127 ( .A(N6314), .Y(n4595) );
  INVX2TS U4128 ( .A(n3873), .Y(n4596) );
  CLKBUFX2TS U4129 ( .A(n4547), .Y(n5840) );
  INVX2TS U4130 ( .A(n5840), .Y(n4597) );
  INVX2TS U4131 ( .A(n5840), .Y(n4598) );
  INVX2TS U4132 ( .A(n5840), .Y(n4599) );
  INVX2TS U4133 ( .A(n2421), .Y(n4619) );
  INVX2TS U4134 ( .A(n4619), .Y(n4600) );
  INVX2TS U4135 ( .A(n4619), .Y(n4601) );
  INVX2TS U4136 ( .A(n4619), .Y(n4602) );
  NAND2X1TS U4137 ( .A(n2702), .B(n5723), .Y(n2704) );
  CLKBUFX2TS U4138 ( .A(n2702), .Y(n4938) );
  NOR2X1TS U4139 ( .A(n3713), .B(n3722), .Y(n2419) );
  CLKBUFX2TS U4140 ( .A(n1748), .Y(n4618) );
  INVX2TS U4141 ( .A(n5807), .Y(n4604) );
  NAND2X1TS U4142 ( .A(n2975), .B(n4590), .Y(n2012) );
  CLKINVX1TS U4143 ( .A(n3713), .Y(n5765) );
  CLKBUFX2TS U4144 ( .A(n2428), .Y(n5054) );
  NAND2X1TS U4145 ( .A(n2837), .B(n3744), .Y(n1968) );
  NOR2X1TS U4146 ( .A(n3709), .B(n4602), .Y(n2972) );
  NOR2X1TS U4147 ( .A(n1955), .B(n4602), .Y(n2698) );
  CLKBUFX2TS U4148 ( .A(n4532), .Y(n4606) );
  INVX2TS U4149 ( .A(n4607), .Y(n4608) );
  NOR2BX1TS U4150 ( .AN(n3113), .B(\add_0_root_r1463/SUM[0] ), .Y(n2426) );
  OR3X1TS U4151 ( .A(n2564), .B(n4578), .C(n5713), .Y(n4609) );
  NOR3X1TS U4152 ( .A(n3730), .B(n3727), .C(n2421), .Y(n2286) );
  INVXLTS U4153 ( .A(cacheDataOut_A[0]), .Y(n5939) );
  INVXLTS U4154 ( .A(cacheDataOut_A[1]), .Y(n5938) );
  INVXLTS U4155 ( .A(cacheDataOut_A[2]), .Y(n5937) );
  INVXLTS U4156 ( .A(cacheDataOut_A[3]), .Y(n5936) );
  INVXLTS U4157 ( .A(cacheDataOut_A[4]), .Y(n5935) );
  INVXLTS U4158 ( .A(cacheDataOut_A[5]), .Y(n5934) );
  INVXLTS U4159 ( .A(cacheDataOut_A[6]), .Y(n5933) );
  INVXLTS U4160 ( .A(cacheDataOut_A[7]), .Y(n5932) );
  INVXLTS U4161 ( .A(cacheDataOut_A[8]), .Y(n5931) );
  INVXLTS U4162 ( .A(cacheDataOut_A[9]), .Y(n5930) );
  INVXLTS U4163 ( .A(cacheDataOut_A[10]), .Y(n5929) );
  INVXLTS U4164 ( .A(cacheDataOut_A[11]), .Y(n5928) );
  INVXLTS U4165 ( .A(cacheDataOut_A[12]), .Y(n5927) );
  INVXLTS U4166 ( .A(cacheDataOut_A[13]), .Y(n5926) );
  INVXLTS U4167 ( .A(cacheDataOut_A[14]), .Y(n5925) );
  INVXLTS U4168 ( .A(cacheDataOut_A[15]), .Y(n5924) );
  INVXLTS U4169 ( .A(cacheDataOut_A[16]), .Y(n5923) );
  INVXLTS U4170 ( .A(cacheDataOut_A[17]), .Y(n5922) );
  INVXLTS U4171 ( .A(cacheDataOut_A[18]), .Y(n5921) );
  INVXLTS U4172 ( .A(cacheDataOut_A[19]), .Y(n5920) );
  INVXLTS U4173 ( .A(cacheDataOut_A[20]), .Y(n5919) );
  INVXLTS U4174 ( .A(cacheDataOut_A[21]), .Y(n5918) );
  INVXLTS U4175 ( .A(cacheDataOut_A[22]), .Y(n5917) );
  INVXLTS U4176 ( .A(cacheDataOut_A[23]), .Y(n5916) );
  INVXLTS U4177 ( .A(cacheDataOut_A[24]), .Y(n5915) );
  INVXLTS U4178 ( .A(cacheDataOut_A[25]), .Y(n5914) );
  INVXLTS U4179 ( .A(cacheDataOut_A[26]), .Y(n5913) );
  INVXLTS U4180 ( .A(cacheDataOut_A[27]), .Y(n5912) );
  INVXLTS U4181 ( .A(cacheDataOut_A[28]), .Y(n5911) );
  INVXLTS U4182 ( .A(cacheDataOut_A[29]), .Y(n5910) );
  INVXLTS U4183 ( .A(cacheDataOut_A[30]), .Y(n5909) );
  INVXLTS U4184 ( .A(cacheDataOut_A[31]), .Y(n5908) );
  INVXLTS U4185 ( .A(n3952), .Y(n5808) );
  INVXLTS U4186 ( .A(n3890), .Y(n5839) );
  INVXLTS U4187 ( .A(n3892), .Y(n5838) );
  INVXLTS U4188 ( .A(n3894), .Y(n5837) );
  INVXLTS U4189 ( .A(n3896), .Y(n5836) );
  INVXLTS U4190 ( .A(n3898), .Y(n5835) );
  INVXLTS U4191 ( .A(n3900), .Y(n5834) );
  INVXLTS U4192 ( .A(n3902), .Y(n5833) );
  INVXLTS U4193 ( .A(n3904), .Y(n5832) );
  INVXLTS U4194 ( .A(n3906), .Y(n5831) );
  INVXLTS U4195 ( .A(n3908), .Y(n5830) );
  INVXLTS U4196 ( .A(n3910), .Y(n5829) );
  INVXLTS U4197 ( .A(n3912), .Y(n5828) );
  INVXLTS U4198 ( .A(n3914), .Y(n5827) );
  INVXLTS U4199 ( .A(n3916), .Y(n5826) );
  INVXLTS U4200 ( .A(n3918), .Y(n5825) );
  INVXLTS U4201 ( .A(n3920), .Y(n5824) );
  INVXLTS U4202 ( .A(n3922), .Y(n5823) );
  INVXLTS U4203 ( .A(n3924), .Y(n5822) );
  INVXLTS U4204 ( .A(n3926), .Y(n5821) );
  INVXLTS U4205 ( .A(n3928), .Y(n5820) );
  INVXLTS U4206 ( .A(n3930), .Y(n5819) );
  INVXLTS U4207 ( .A(n3932), .Y(n5818) );
  INVXLTS U4208 ( .A(n3934), .Y(n5817) );
  INVXLTS U4209 ( .A(n3936), .Y(n5816) );
  INVXLTS U4210 ( .A(n3938), .Y(n5815) );
  INVXLTS U4211 ( .A(n3940), .Y(n5814) );
  INVXLTS U4212 ( .A(n3942), .Y(n5813) );
  INVXLTS U4213 ( .A(n3944), .Y(n5812) );
  INVXLTS U4214 ( .A(n3946), .Y(n5811) );
  INVXLTS U4215 ( .A(n3948), .Y(n5810) );
  INVXLTS U4216 ( .A(n3950), .Y(n5809) );
  INVXLTS U4217 ( .A(n4030), .Y(n5841) );
  INVXLTS U4218 ( .A(n3968), .Y(n5872) );
  INVXLTS U4219 ( .A(n3970), .Y(n5871) );
  INVXLTS U4220 ( .A(n3972), .Y(n5870) );
  INVXLTS U4221 ( .A(n3974), .Y(n5869) );
  INVXLTS U4222 ( .A(n3976), .Y(n5868) );
  INVXLTS U4223 ( .A(n3978), .Y(n5867) );
  INVXLTS U4224 ( .A(n3980), .Y(n5866) );
  INVXLTS U4225 ( .A(n3982), .Y(n5865) );
  INVXLTS U4226 ( .A(n3984), .Y(n5864) );
  INVXLTS U4227 ( .A(n3986), .Y(n5863) );
  INVXLTS U4228 ( .A(n3988), .Y(n5862) );
  INVXLTS U4229 ( .A(n3990), .Y(n5861) );
  INVXLTS U4230 ( .A(n3992), .Y(n5860) );
  INVXLTS U4231 ( .A(n3994), .Y(n5859) );
  INVXLTS U4232 ( .A(n3996), .Y(n5858) );
  INVXLTS U4233 ( .A(n3998), .Y(n5857) );
  INVXLTS U4234 ( .A(n4000), .Y(n5856) );
  INVXLTS U4235 ( .A(n4002), .Y(n5855) );
  INVXLTS U4236 ( .A(n4004), .Y(n5854) );
  INVXLTS U4237 ( .A(n4006), .Y(n5853) );
  INVXLTS U4238 ( .A(n4008), .Y(n5852) );
  INVXLTS U4239 ( .A(n4010), .Y(n5851) );
  INVXLTS U4240 ( .A(n4012), .Y(n5850) );
  INVXLTS U4241 ( .A(n4014), .Y(n5849) );
  INVXLTS U4242 ( .A(n4016), .Y(n5848) );
  INVXLTS U4243 ( .A(n4018), .Y(n5847) );
  INVXLTS U4244 ( .A(n4020), .Y(n5846) );
  INVXLTS U4245 ( .A(n4022), .Y(n5845) );
  INVXLTS U4246 ( .A(n4024), .Y(n5844) );
  INVXLTS U4247 ( .A(n4026), .Y(n5843) );
  INVXLTS U4248 ( .A(n4028), .Y(n5842) );
  CLKBUFX2TS U4249 ( .A(n4783), .Y(n4773) );
  CLKBUFX2TS U4250 ( .A(n5428), .Y(n5425) );
  CLKBUFX2TS U4251 ( .A(n5428), .Y(n5426) );
  CLKBUFX2TS U4252 ( .A(n5597), .Y(n5590) );
  CLKBUFX2TS U4253 ( .A(n5598), .Y(n5587) );
  CLKBUFX2TS U4254 ( .A(n5597), .Y(n5589) );
  CLKBUFX2TS U4255 ( .A(n5414), .Y(n5411) );
  CLKBUFX2TS U4256 ( .A(n5599), .Y(n5586) );
  CLKBUFX2TS U4257 ( .A(n5598), .Y(n5588) );
  OAI32XLTS U4258 ( .A0(n2233), .A1(n4568), .A2(n5295), .B0(n5803), .B1(n3706), 
        .Y(n1764) );
  OAI211XLTS U4259 ( .A0(n3732), .A1(n3710), .B0(n2044), .C0(n2045), .Y(n2004)
         );
  OAI21XLTS U4260 ( .A0(n3670), .A1(n2046), .B0(n5569), .Y(n2044) );
  OAI211XLTS U4261 ( .A0(n1865), .A1(n3714), .B0(n1867), .C0(n1868), .Y(n1826)
         );
  OAI21XLTS U4262 ( .A0(n3668), .A1(n1869), .B0(n5568), .Y(n1867) );
  OAI211XLTS U4263 ( .A0(n1865), .A1(n3712), .B0(n2000), .C0(n2001), .Y(n1960)
         );
  OAI21XLTS U4264 ( .A0(n5974), .A1(n2272), .B0(n2274), .Y(n1797) );
  OAI21XLTS U4265 ( .A0(n5804), .A1(n2085), .B0(n5598), .Y(n2981) );
  NAND4XLTS U4266 ( .A(n3109), .B(n2274), .C(n2132), .D(n5718), .Y(n2976) );
  INVX1TS U4267 ( .A(n3149), .Y(\add_0_root_r1459/B[0] ) );
  INVXLTS U4268 ( .A(n1999), .Y(n5768) );
  AND2XLTS U4269 ( .A(n3108), .B(n2271), .Y(n2051) );
  NAND4X1TS U4270 ( .A(N6372), .B(n2427), .C(n3719), .D(n5774), .Y(n2848) );
  NAND4X1TS U4271 ( .A(n4598), .B(n5774), .C(n2838), .D(n2839), .Y(n2710) );
  AND2XLTS U4272 ( .A(n1821), .B(n4532), .Y(n1666) );
  CLKBUFX2TS U4273 ( .A(n5296), .Y(n5295) );
  CLKBUFX2TS U4274 ( .A(n5296), .Y(n5293) );
  CLKBUFX2TS U4275 ( .A(n5296), .Y(n5294) );
  OAI211XLTS U4276 ( .A0(n5593), .A1(n2264), .B0(n2265), .C0(n2266), .Y(n2263)
         );
  OAI211XLTS U4277 ( .A0(n5590), .A1(n2210), .B0(n2211), .C0(n2212), .Y(n2209)
         );
  NAND2XLTS U4278 ( .A(n2701), .B(n3764), .Y(n1765) );
  NAND2XLTS U4279 ( .A(n2563), .B(n3763), .Y(n1755) );
  AOI21XLTS U4280 ( .A0(n2286), .A1(n5762), .B0(n5567), .Y(n2843) );
  AOI21XLTS U4281 ( .A0(n4560), .A1(n5763), .B0(n5567), .Y(n2569) );
  AOI21XLTS U4282 ( .A0(n4560), .A1(n5765), .B0(n5567), .Y(n2290) );
  AOI21X1TS U4283 ( .A0(n4560), .A1(n5768), .B0(n5567), .Y(n2705) );
  AOI21X1TS U4284 ( .A0(n4560), .A1(n5770), .B0(n5568), .Y(n2431) );
  CLKINVX2TS U4285 ( .A(n5186), .Y(n5185) );
  CLKINVX2TS U4286 ( .A(n5374), .Y(n5357) );
  CLKINVX2TS U4287 ( .A(n5280), .Y(n5263) );
  AND2XLTS U4288 ( .A(\add_0_root_r1463/SUM[0] ), .B(n3113), .Y(n2285) );
  CLKAND2X2TS U4289 ( .A(\add_0_root_r1459/SUM[0] ), .B(n3112), .Y(n2283) );
  NAND2X1TS U4290 ( .A(n3110), .B(n4591), .Y(n2054) );
  OAI32XLTS U4291 ( .A0(n2246), .A1(n5699), .A2(n4569), .B0(n5803), .B1(n3712), 
        .Y(n1774) );
  NOR4XLTS U4292 ( .A(n5559), .B(n3728), .C(n5527), .D(
        \indexIncrementer_EAST[1] ), .Y(n1794) );
  NAND4XLTS U4293 ( .A(n3703), .B(\add_0_root_r1459/SUM[2] ), .C(n2283), .D(
        n3763), .Y(n1736) );
  CLKBUFX2TS U4294 ( .A(n5629), .Y(n5625) );
  NOR2X1TS U4295 ( .A(n3724), .B(n5592), .Y(n2130) );
  CLKBUFX2TS U4296 ( .A(n4614), .Y(n5292) );
  AND3XLTS U4297 ( .A(n2236), .B(n5291), .C(n2237), .Y(n2235) );
  NOR2X1TS U4298 ( .A(n4618), .B(n1823), .Y(\indexIncrementer_EAST[1] ) );
  OAI21XLTS U4299 ( .A0(n5563), .A1(n2132), .B0(n2276), .Y(n1618) );
  OAI32XLTS U4300 ( .A0(n2208), .A1(n1740), .A2(n4569), .B0(n5803), .B1(n3714), 
        .Y(n1742) );
  OAI32XLTS U4301 ( .A0(n2262), .A1(n1783), .A2(n4568), .B0(n5803), .B1(n3709), 
        .Y(n1785) );
  AOI211XLTS U4302 ( .A0(n1788), .A1(n5584), .B0(n4602), .C0(n3709), .Y(n2009)
         );
  AOI211XLTS U4303 ( .A0(n1745), .A1(n5583), .B0(n4601), .C0(n3714), .Y(n1831)
         );
  AOI211XLTS U4304 ( .A0(n1777), .A1(n5585), .B0(n2421), .C0(n3712), .Y(n1965)
         );
  AOI211XLTS U4305 ( .A0(n1767), .A1(n5583), .B0(n4602), .C0(n3706), .Y(n1920)
         );
  AOI211XLTS U4306 ( .A0(n5974), .A1(n5584), .B0(n2421), .C0(n2085), .Y(n2050)
         );
  NOR2XLTS U4307 ( .A(n1910), .B(n3722), .Y(n2560) );
  OAI32XLTS U4308 ( .A0(n2220), .A1(n3805), .A2(n4567), .B0(n4610), .B1(n3708), 
        .Y(n1754) );
  OAI21XLTS U4309 ( .A0(n4600), .A1(n3151), .B0(n3695), .Y(n3152) );
  XOR2XLTS U4310 ( .A(n4603), .B(n4596), .Y(\add_0_root_r1463/SUM[0] ) );
  OR2XLTS U4311 ( .A(n3149), .B(n3745), .Y(n4613) );
  NOR3BXLTS U4312 ( .AN(n3695), .B(n4601), .C(n3151), .Y(totalAccesses[2]) );
  INVXLTS U4313 ( .A(cacheDataOut_B[0]), .Y(n5971) );
  INVXLTS U4314 ( .A(cacheDataOut_B[1]), .Y(n5970) );
  INVXLTS U4315 ( .A(cacheDataOut_B[2]), .Y(n5969) );
  INVXLTS U4316 ( .A(cacheDataOut_B[3]), .Y(n5968) );
  INVXLTS U4317 ( .A(cacheDataOut_B[4]), .Y(n5967) );
  INVXLTS U4318 ( .A(cacheDataOut_B[5]), .Y(n5966) );
  INVXLTS U4319 ( .A(cacheDataOut_B[6]), .Y(n5965) );
  INVXLTS U4320 ( .A(cacheDataOut_B[7]), .Y(n5964) );
  INVXLTS U4321 ( .A(cacheDataOut_B[8]), .Y(n5963) );
  INVXLTS U4322 ( .A(cacheDataOut_B[9]), .Y(n5962) );
  INVXLTS U4323 ( .A(cacheDataOut_B[10]), .Y(n5961) );
  INVXLTS U4324 ( .A(cacheDataOut_B[11]), .Y(n5960) );
  INVXLTS U4325 ( .A(cacheDataOut_B[12]), .Y(n5959) );
  INVXLTS U4326 ( .A(cacheDataOut_B[13]), .Y(n5958) );
  INVXLTS U4327 ( .A(cacheDataOut_B[14]), .Y(n5957) );
  INVXLTS U4328 ( .A(cacheDataOut_B[15]), .Y(n5956) );
  INVXLTS U4329 ( .A(cacheDataOut_B[16]), .Y(n5955) );
  INVXLTS U4330 ( .A(cacheDataOut_B[17]), .Y(n5954) );
  INVXLTS U4331 ( .A(cacheDataOut_B[18]), .Y(n5953) );
  INVXLTS U4332 ( .A(cacheDataOut_B[19]), .Y(n5952) );
  INVXLTS U4333 ( .A(cacheDataOut_B[20]), .Y(n5951) );
  INVXLTS U4334 ( .A(cacheDataOut_B[21]), .Y(n5950) );
  INVXLTS U4335 ( .A(cacheDataOut_B[22]), .Y(n5949) );
  INVXLTS U4336 ( .A(cacheDataOut_B[23]), .Y(n5948) );
  INVXLTS U4337 ( .A(cacheDataOut_B[24]), .Y(n5947) );
  INVXLTS U4338 ( .A(cacheDataOut_B[25]), .Y(n5946) );
  INVXLTS U4339 ( .A(cacheDataOut_B[26]), .Y(n5945) );
  INVXLTS U4340 ( .A(cacheDataOut_B[27]), .Y(n5944) );
  INVXLTS U4341 ( .A(cacheDataOut_B[28]), .Y(n5943) );
  INVXLTS U4342 ( .A(cacheDataOut_B[29]), .Y(n5942) );
  INVXLTS U4343 ( .A(cacheDataOut_B[30]), .Y(n5941) );
  INVXLTS U4344 ( .A(cacheDataOut_B[31]), .Y(n5940) );
  AOI211XLTS U4345 ( .A0(n5598), .A1(n5754), .B0(n2126), .C0(n2131), .Y(n2124)
         );
  OAI32XLTS U4346 ( .A0(n5755), .A1(n5730), .A2(n2268), .B0(n4589), .B1(n1173), 
        .Y(n3384) );
  INVXLTS U4347 ( .A(n4588), .Y(n5755) );
  OAI22XLTS U4348 ( .A0(n4678), .A1(n1240), .B0(n3783), .B1(n3832), .Y(n1863)
         );
  OAI22XLTS U4349 ( .A0(n4678), .A1(n1239), .B0(n3784), .B1(n3836), .Y(n1859)
         );
  OAI22XLTS U4350 ( .A0(n4678), .A1(n1238), .B0(n3785), .B1(n3840), .Y(n1855)
         );
  OAI22XLTS U4351 ( .A0(n4678), .A1(n1237), .B0(n3783), .B1(n3844), .Y(n1851)
         );
  OAI22XLTS U4352 ( .A0(n4677), .A1(n1236), .B0(n3784), .B1(n3848), .Y(n1847)
         );
  OAI22XLTS U4353 ( .A0(n3853), .A1(n5356), .B0(n5373), .B1(n1844), .Y(n1842)
         );
  OAI22XLTS U4354 ( .A0(n4677), .A1(n1235), .B0(n3785), .B1(n3852), .Y(n1843)
         );
  OAI22XLTS U4355 ( .A0(n3857), .A1(n5356), .B0(n5373), .B1(n1840), .Y(n1838)
         );
  OAI22XLTS U4356 ( .A0(n4677), .A1(n1234), .B0(n3783), .B1(n3856), .Y(n1839)
         );
  OAI22XLTS U4357 ( .A0(n4679), .A1(n1233), .B0(n3784), .B1(n3860), .Y(n1832)
         );
  OAI22XLTS U4358 ( .A0(n4053), .A1(n5184), .B0(n5186), .B1(n2022), .Y(n2020)
         );
  OAI22XLTS U4359 ( .A0(n3853), .A1(n5262), .B0(n5279), .B1(n1934), .Y(n1932)
         );
  OAI22XLTS U4360 ( .A0(n4055), .A1(n5184), .B0(n5186), .B1(n2018), .Y(n2016)
         );
  OAI22XLTS U4361 ( .A0(n3857), .A1(n5262), .B0(n5279), .B1(n1930), .Y(n1928)
         );
  OAI22XLTS U4362 ( .A0(n3854), .A1(n5317), .B0(n5319), .B1(n1889), .Y(n1887)
         );
  OAI22XLTS U4363 ( .A0(n3858), .A1(n5317), .B0(n5326), .B1(n1885), .Y(n1883)
         );
  OAI22XLTS U4364 ( .A0(n1277), .A1(n4588), .B0(n1626), .B1(n1620), .Y(n3204)
         );
  OAI22XLTS U4365 ( .A0(n1276), .A1(n4589), .B0(n1629), .B1(n1620), .Y(n3205)
         );
  OAI22XLTS U4366 ( .A0(n1275), .A1(n4620), .B0(n1632), .B1(n4549), .Y(n3206)
         );
  OAI22XLTS U4367 ( .A0(n1274), .A1(n4588), .B0(n1635), .B1(n4549), .Y(n3207)
         );
  OAI22XLTS U4368 ( .A0(n1273), .A1(n4589), .B0(n1638), .B1(n4549), .Y(n3208)
         );
  OAI22XLTS U4369 ( .A0(n1262), .A1(n4620), .B0(n5738), .B1(n1800), .Y(n3267)
         );
  OAI22XLTS U4370 ( .A0(n1261), .A1(n4588), .B0(n5738), .B1(n1795), .Y(n3266)
         );
  OAI22XLTS U4371 ( .A0(n4938), .A1(n1071), .B0(n2831), .B1(n4920), .Y(n3545)
         );
  OAI22XLTS U4372 ( .A0(n4935), .A1(n1070), .B0(n2827), .B1(n4920), .Y(n3544)
         );
  OAI22XLTS U4373 ( .A0(n4939), .A1(n1069), .B0(n2823), .B1(n4920), .Y(n3543)
         );
  OAI22XLTS U4374 ( .A0(n4930), .A1(n1068), .B0(n2819), .B1(n4920), .Y(n3542)
         );
  OAI22XLTS U4375 ( .A0(n4930), .A1(n1067), .B0(n2815), .B1(n4921), .Y(n3541)
         );
  OAI22XLTS U4376 ( .A0(n4930), .A1(n1066), .B0(n2811), .B1(n4921), .Y(n3540)
         );
  OAI22XLTS U4377 ( .A0(n4930), .A1(n1065), .B0(n2807), .B1(n4921), .Y(n3539)
         );
  OAI22XLTS U4378 ( .A0(n4937), .A1(n1064), .B0(n2803), .B1(n4921), .Y(n3538)
         );
  OAI22XLTS U4379 ( .A0(n4934), .A1(n1063), .B0(n2799), .B1(n4922), .Y(n3537)
         );
  OAI22XLTS U4380 ( .A0(n4937), .A1(n1062), .B0(n2795), .B1(n4922), .Y(n3536)
         );
  OAI22XLTS U4381 ( .A0(n4939), .A1(n1061), .B0(n2791), .B1(n4922), .Y(n3535)
         );
  OAI22XLTS U4382 ( .A0(n4936), .A1(n1060), .B0(n2787), .B1(n4922), .Y(n3534)
         );
  OAI22XLTS U4383 ( .A0(n4936), .A1(n1059), .B0(n2783), .B1(n4923), .Y(n3533)
         );
  OAI22XLTS U4384 ( .A0(n4937), .A1(n1058), .B0(n2779), .B1(n4923), .Y(n3532)
         );
  OAI22XLTS U4385 ( .A0(n4935), .A1(n1057), .B0(n2775), .B1(n4923), .Y(n3531)
         );
  OAI22XLTS U4386 ( .A0(n4936), .A1(n1056), .B0(n2771), .B1(n4923), .Y(n3530)
         );
  OAI22XLTS U4387 ( .A0(n4936), .A1(n1055), .B0(n2767), .B1(n4927), .Y(n3529)
         );
  OAI22XLTS U4388 ( .A0(n4938), .A1(n1054), .B0(n2763), .B1(n4929), .Y(n3528)
         );
  OAI22XLTS U4389 ( .A0(n4934), .A1(n1053), .B0(n2759), .B1(n4929), .Y(n3527)
         );
  OAI22XLTS U4390 ( .A0(n4931), .A1(n1052), .B0(n2755), .B1(n4928), .Y(n3526)
         );
  OAI22XLTS U4391 ( .A0(n4931), .A1(n1051), .B0(n2751), .B1(n4924), .Y(n3525)
         );
  OAI22XLTS U4392 ( .A0(n4931), .A1(n1050), .B0(n2747), .B1(n4924), .Y(n3524)
         );
  OAI22XLTS U4393 ( .A0(n4931), .A1(n1049), .B0(n2743), .B1(n4924), .Y(n3523)
         );
  OAI22XLTS U4394 ( .A0(n4932), .A1(n1048), .B0(n2739), .B1(n4924), .Y(n3522)
         );
  OAI22XLTS U4395 ( .A0(n4932), .A1(n1047), .B0(n2735), .B1(n4925), .Y(n3521)
         );
  OAI22XLTS U4396 ( .A0(n4932), .A1(n1046), .B0(n2731), .B1(n4925), .Y(n3520)
         );
  OAI22XLTS U4397 ( .A0(n4932), .A1(n1045), .B0(n2727), .B1(n4925), .Y(n3519)
         );
  OAI22XLTS U4398 ( .A0(n4933), .A1(n1044), .B0(n2723), .B1(n4925), .Y(n3518)
         );
  OAI22XLTS U4399 ( .A0(n4933), .A1(n1043), .B0(n2719), .B1(n4926), .Y(n3517)
         );
  OAI22XLTS U4400 ( .A0(n4933), .A1(n1042), .B0(n2715), .B1(n4926), .Y(n3516)
         );
  OAI22XLTS U4401 ( .A0(n4933), .A1(n1041), .B0(n2711), .B1(n4926), .Y(n3515)
         );
  OAI22XLTS U4402 ( .A0(n4934), .A1(n1040), .B0(n2703), .B1(n4926), .Y(n3514)
         );
  OAI22XLTS U4403 ( .A0(n2967), .A1(n4846), .B0(n4668), .B1(n1038), .Y(n2966)
         );
  OAI22XLTS U4404 ( .A0(n2963), .A1(n4845), .B0(n4670), .B1(n1037), .Y(n2962)
         );
  OAI22XLTS U4405 ( .A0(n2959), .A1(n4845), .B0(n4669), .B1(n1036), .Y(n2958)
         );
  OAI22XLTS U4406 ( .A0(n2951), .A1(n4838), .B0(n4668), .B1(n1034), .Y(n2950)
         );
  OAI22XLTS U4407 ( .A0(n2947), .A1(n4838), .B0(n4669), .B1(n1033), .Y(n2946)
         );
  OAI22XLTS U4408 ( .A0(n2943), .A1(n4838), .B0(n4669), .B1(n1032), .Y(n2942)
         );
  OAI22XLTS U4409 ( .A0(n2935), .A1(n4839), .B0(n4665), .B1(n1030), .Y(n2934)
         );
  OAI22XLTS U4410 ( .A0(n2931), .A1(n4839), .B0(n4668), .B1(n1029), .Y(n2930)
         );
  OAI22XLTS U4411 ( .A0(n2927), .A1(n4839), .B0(n4667), .B1(n1028), .Y(n2926)
         );
  OAI22XLTS U4412 ( .A0(n2919), .A1(n4840), .B0(n4667), .B1(n1026), .Y(n2918)
         );
  OAI22XLTS U4413 ( .A0(n2915), .A1(n4840), .B0(n4667), .B1(n1025), .Y(n2914)
         );
  OAI22XLTS U4414 ( .A0(n2911), .A1(n4840), .B0(n4666), .B1(n1024), .Y(n2910)
         );
  OAI22XLTS U4415 ( .A0(n2903), .A1(n4841), .B0(n4666), .B1(n1022), .Y(n2902)
         );
  OAI22XLTS U4416 ( .A0(n2899), .A1(n4841), .B0(n4666), .B1(n1021), .Y(n2898)
         );
  OAI22XLTS U4417 ( .A0(n2895), .A1(n4841), .B0(n4665), .B1(n1020), .Y(n2894)
         );
  OAI22XLTS U4418 ( .A0(n2887), .A1(n4842), .B0(n4665), .B1(n1018), .Y(n2886)
         );
  OAI22XLTS U4419 ( .A0(n2883), .A1(n4842), .B0(n4675), .B1(n1017), .Y(n2882)
         );
  OAI22XLTS U4420 ( .A0(n2879), .A1(n4842), .B0(n4671), .B1(n1016), .Y(n2878)
         );
  OAI22XLTS U4421 ( .A0(n2871), .A1(n4843), .B0(n4671), .B1(n1014), .Y(n2870)
         );
  OAI22XLTS U4422 ( .A0(n2867), .A1(n4843), .B0(n4675), .B1(n1013), .Y(n2866)
         );
  OAI22XLTS U4423 ( .A0(n2863), .A1(n4843), .B0(n4673), .B1(n1012), .Y(n2862)
         );
  OAI22XLTS U4424 ( .A0(n2855), .A1(n4844), .B0(n4676), .B1(n1010), .Y(n2854)
         );
  OAI22XLTS U4425 ( .A0(n2851), .A1(n4844), .B0(n4664), .B1(n1009), .Y(n2850)
         );
  OAI22XLTS U4426 ( .A0(n2845), .A1(n4844), .B0(n4664), .B1(n1008), .Y(n2844)
         );
  OAI22XLTS U4427 ( .A0(n2414), .A1(n5086), .B0(n1166), .B1(n4685), .Y(n2413)
         );
  OAI22XLTS U4428 ( .A0(n2410), .A1(n5086), .B0(n1165), .B1(n4690), .Y(n2409)
         );
  OAI22XLTS U4429 ( .A0(n2406), .A1(n5086), .B0(n1164), .B1(n4686), .Y(n2405)
         );
  OAI22XLTS U4430 ( .A0(n2398), .A1(n5087), .B0(n1162), .B1(n4685), .Y(n2397)
         );
  OAI22XLTS U4431 ( .A0(n2394), .A1(n5087), .B0(n1161), .B1(n4687), .Y(n2393)
         );
  OAI22XLTS U4432 ( .A0(n2390), .A1(n5087), .B0(n1160), .B1(n4689), .Y(n2389)
         );
  OAI22XLTS U4433 ( .A0(n2382), .A1(n5094), .B0(n1158), .B1(n4682), .Y(n2381)
         );
  OAI22XLTS U4434 ( .A0(n2378), .A1(n5094), .B0(n1157), .B1(n4685), .Y(n2377)
         );
  OAI22XLTS U4435 ( .A0(n2374), .A1(n5092), .B0(n1156), .B1(n4684), .Y(n2373)
         );
  OAI22XLTS U4436 ( .A0(n2366), .A1(n5094), .B0(n1154), .B1(n4684), .Y(n2365)
         );
  OAI22XLTS U4437 ( .A0(n2362), .A1(n5094), .B0(n1153), .B1(n4684), .Y(n2361)
         );
  OAI22XLTS U4438 ( .A0(n2358), .A1(n5095), .B0(n1152), .B1(n4683), .Y(n2357)
         );
  OAI22XLTS U4439 ( .A0(n2350), .A1(n5088), .B0(n1150), .B1(n4683), .Y(n2349)
         );
  OAI22XLTS U4440 ( .A0(n2346), .A1(n5088), .B0(n1149), .B1(n4683), .Y(n2345)
         );
  OAI22XLTS U4441 ( .A0(n2342), .A1(n5088), .B0(n1148), .B1(n4682), .Y(n2341)
         );
  OAI22XLTS U4442 ( .A0(n2334), .A1(n5089), .B0(n1146), .B1(n4682), .Y(n2333)
         );
  OAI22XLTS U4443 ( .A0(n2330), .A1(n5089), .B0(n1145), .B1(n4681), .Y(n2329)
         );
  OAI22XLTS U4444 ( .A0(n2326), .A1(n5089), .B0(n1144), .B1(n4681), .Y(n2325)
         );
  OAI22XLTS U4445 ( .A0(n2318), .A1(n5090), .B0(n1142), .B1(n4681), .Y(n2317)
         );
  OAI22XLTS U4446 ( .A0(n2314), .A1(n5090), .B0(n1141), .B1(n4680), .Y(n2313)
         );
  OAI22XLTS U4447 ( .A0(n2310), .A1(n5090), .B0(n1140), .B1(n4680), .Y(n2309)
         );
  OAI22XLTS U4448 ( .A0(n2302), .A1(n5091), .B0(n1138), .B1(n4680), .Y(n2301)
         );
  OAI22XLTS U4449 ( .A0(n2298), .A1(n5091), .B0(n1137), .B1(n4679), .Y(n2297)
         );
  OAI22XLTS U4450 ( .A0(n2292), .A1(n5091), .B0(n1136), .B1(n4679), .Y(n2291)
         );
  OAI22XLTS U4451 ( .A0(n2693), .A1(n4962), .B0(n5289), .B1(n974), .Y(n2692)
         );
  OAI22XLTS U4452 ( .A0(n2689), .A1(n4962), .B0(n5291), .B1(n973), .Y(n2688)
         );
  OAI22XLTS U4453 ( .A0(n2685), .A1(n4962), .B0(n5290), .B1(n972), .Y(n2684)
         );
  OAI22XLTS U4454 ( .A0(n2677), .A1(n4963), .B0(n5289), .B1(n970), .Y(n2676)
         );
  OAI22XLTS U4455 ( .A0(n2673), .A1(n4963), .B0(n5290), .B1(n969), .Y(n2672)
         );
  OAI22XLTS U4456 ( .A0(n2669), .A1(n4963), .B0(n5290), .B1(n968), .Y(n2668)
         );
  OAI22XLTS U4457 ( .A0(n2661), .A1(n4964), .B0(n5286), .B1(n966), .Y(n2660)
         );
  OAI22XLTS U4458 ( .A0(n2657), .A1(n4964), .B0(n5289), .B1(n965), .Y(n2656)
         );
  OAI22XLTS U4459 ( .A0(n2653), .A1(n4964), .B0(n5288), .B1(n964), .Y(n2652)
         );
  OAI22XLTS U4460 ( .A0(n2645), .A1(n4965), .B0(n5288), .B1(n962), .Y(n2644)
         );
  OAI22XLTS U4461 ( .A0(n2641), .A1(n4965), .B0(n5288), .B1(n961), .Y(n2640)
         );
  OAI22XLTS U4462 ( .A0(n2637), .A1(n4965), .B0(n5287), .B1(n960), .Y(n2636)
         );
  OAI22XLTS U4463 ( .A0(n2629), .A1(n4971), .B0(n5287), .B1(n958), .Y(n2628)
         );
  OAI22XLTS U4464 ( .A0(n2625), .A1(n4970), .B0(n5287), .B1(n957), .Y(n2624)
         );
  OAI22XLTS U4465 ( .A0(n2621), .A1(n4970), .B0(n5286), .B1(n956), .Y(n2620)
         );
  OAI22XLTS U4466 ( .A0(n2613), .A1(n4966), .B0(n5286), .B1(n954), .Y(n2612)
         );
  OAI22XLTS U4467 ( .A0(n2609), .A1(n4966), .B0(n5285), .B1(n953), .Y(n2608)
         );
  OAI22XLTS U4468 ( .A0(n2605), .A1(n4966), .B0(n5285), .B1(n952), .Y(n2604)
         );
  OAI22XLTS U4469 ( .A0(n2597), .A1(n4967), .B0(n5285), .B1(n950), .Y(n2596)
         );
  OAI22XLTS U4470 ( .A0(n2593), .A1(n4967), .B0(n5284), .B1(n949), .Y(n2592)
         );
  OAI22XLTS U4471 ( .A0(n2589), .A1(n4967), .B0(n5284), .B1(n948), .Y(n2588)
         );
  OAI22XLTS U4472 ( .A0(n2581), .A1(n4968), .B0(n5284), .B1(n946), .Y(n2580)
         );
  OAI22XLTS U4473 ( .A0(n2577), .A1(n4968), .B0(n5283), .B1(n945), .Y(n2576)
         );
  OAI22XLTS U4474 ( .A0(n2571), .A1(n4968), .B0(n5283), .B1(n944), .Y(n2570)
         );
  OAI22XLTS U4475 ( .A0(n5054), .A1(n1007), .B0(n2557), .B1(n5044), .Y(n3481)
         );
  OAI22XLTS U4476 ( .A0(n5054), .A1(n1006), .B0(n2553), .B1(n5044), .Y(n3480)
         );
  OAI22XLTS U4477 ( .A0(n5054), .A1(n1005), .B0(n2549), .B1(n5044), .Y(n3479)
         );
  OAI22XLTS U4478 ( .A0(n5055), .A1(n1004), .B0(n2545), .B1(n5044), .Y(n3478)
         );
  OAI22XLTS U4479 ( .A0(n5055), .A1(n1003), .B0(n2541), .B1(n5053), .Y(n3477)
         );
  OAI22XLTS U4480 ( .A0(n5055), .A1(n1002), .B0(n2537), .B1(n5051), .Y(n3476)
         );
  OAI22XLTS U4481 ( .A0(n5055), .A1(n1001), .B0(n2533), .B1(n5053), .Y(n3475)
         );
  OAI22XLTS U4482 ( .A0(n5062), .A1(n1000), .B0(n2529), .B1(n5051), .Y(n3474)
         );
  OAI22XLTS U4483 ( .A0(n5062), .A1(n999), .B0(n2525), .B1(n5045), .Y(n3473)
         );
  OAI22XLTS U4484 ( .A0(n5060), .A1(n998), .B0(n2521), .B1(n5045), .Y(n3472)
         );
  OAI22XLTS U4485 ( .A0(n2428), .A1(n997), .B0(n2517), .B1(n5045), .Y(n3471)
         );
  OAI22XLTS U4486 ( .A0(n5056), .A1(n996), .B0(n2513), .B1(n5045), .Y(n3470)
         );
  OAI22XLTS U4487 ( .A0(n5056), .A1(n995), .B0(n2509), .B1(n5046), .Y(n3469)
         );
  OAI22XLTS U4488 ( .A0(n5056), .A1(n994), .B0(n2505), .B1(n5046), .Y(n3468)
         );
  OAI22XLTS U4489 ( .A0(n5056), .A1(n993), .B0(n2501), .B1(n5046), .Y(n3467)
         );
  OAI22XLTS U4490 ( .A0(n5057), .A1(n992), .B0(n2497), .B1(n5046), .Y(n3466)
         );
  OAI22XLTS U4491 ( .A0(n5057), .A1(n991), .B0(n2493), .B1(n5047), .Y(n3465)
         );
  OAI22XLTS U4492 ( .A0(n5057), .A1(n990), .B0(n2489), .B1(n5047), .Y(n3464)
         );
  OAI22XLTS U4493 ( .A0(n5057), .A1(n989), .B0(n2485), .B1(n5047), .Y(n3463)
         );
  OAI22XLTS U4494 ( .A0(n5063), .A1(n988), .B0(n2481), .B1(n5047), .Y(n3462)
         );
  OAI22XLTS U4495 ( .A0(n5061), .A1(n987), .B0(n2477), .B1(n5048), .Y(n3461)
         );
  OAI22XLTS U4496 ( .A0(n5061), .A1(n986), .B0(n2473), .B1(n5048), .Y(n3460)
         );
  OAI22XLTS U4497 ( .A0(n5062), .A1(n985), .B0(n2469), .B1(n5048), .Y(n3459)
         );
  OAI22XLTS U4498 ( .A0(n5058), .A1(n984), .B0(n2465), .B1(n5048), .Y(n3458)
         );
  OAI22XLTS U4499 ( .A0(n5058), .A1(n983), .B0(n2461), .B1(n5049), .Y(n3457)
         );
  OAI22XLTS U4500 ( .A0(n5058), .A1(n982), .B0(n2457), .B1(n5049), .Y(n3456)
         );
  OAI22XLTS U4501 ( .A0(n5058), .A1(n981), .B0(n2453), .B1(n5049), .Y(n3455)
         );
  OAI22XLTS U4502 ( .A0(n5059), .A1(n980), .B0(n2449), .B1(n5049), .Y(n3454)
         );
  OAI22XLTS U4503 ( .A0(n5059), .A1(n979), .B0(n2445), .B1(n5050), .Y(n3453)
         );
  OAI22XLTS U4504 ( .A0(n5059), .A1(n978), .B0(n2441), .B1(n5050), .Y(n3452)
         );
  OAI22XLTS U4505 ( .A0(n5059), .A1(n977), .B0(n2437), .B1(n5050), .Y(n3451)
         );
  OAI22XLTS U4506 ( .A0(n5060), .A1(n976), .B0(n2429), .B1(n5050), .Y(n3450)
         );
  OAI22XLTS U4507 ( .A0(n1135), .A1(n2976), .B0(n3104), .B1(n4796), .Y(n3609)
         );
  OAI22XLTS U4508 ( .A0(n1134), .A1(n4814), .B0(n3100), .B1(n4796), .Y(n3608)
         );
  OAI22XLTS U4509 ( .A0(n1133), .A1(n4811), .B0(n3096), .B1(n4796), .Y(n3607)
         );
  OAI22XLTS U4510 ( .A0(n1132), .A1(n4806), .B0(n3092), .B1(n4796), .Y(n3606)
         );
  OAI22XLTS U4511 ( .A0(n1131), .A1(n4806), .B0(n3088), .B1(n4797), .Y(n3605)
         );
  OAI22XLTS U4512 ( .A0(n1130), .A1(n4806), .B0(n3084), .B1(n4797), .Y(n3604)
         );
  OAI22XLTS U4513 ( .A0(n1129), .A1(n4806), .B0(n3080), .B1(n4797), .Y(n3603)
         );
  OAI22XLTS U4514 ( .A0(n1128), .A1(n4813), .B0(n3076), .B1(n4797), .Y(n3602)
         );
  OAI22XLTS U4515 ( .A0(n1127), .A1(n4813), .B0(n3072), .B1(n4798), .Y(n3601)
         );
  OAI22XLTS U4516 ( .A0(n1126), .A1(n4815), .B0(n3068), .B1(n4798), .Y(n3600)
         );
  OAI22XLTS U4517 ( .A0(n1125), .A1(n4813), .B0(n3064), .B1(n4798), .Y(n3599)
         );
  OAI22XLTS U4518 ( .A0(n1124), .A1(n4812), .B0(n3060), .B1(n4798), .Y(n3598)
         );
  OAI22XLTS U4519 ( .A0(n1123), .A1(n4812), .B0(n3056), .B1(n4799), .Y(n3597)
         );
  OAI22XLTS U4520 ( .A0(n1122), .A1(n4814), .B0(n3052), .B1(n4799), .Y(n3596)
         );
  OAI22XLTS U4521 ( .A0(n1121), .A1(n4811), .B0(n3048), .B1(n4799), .Y(n3595)
         );
  OAI22XLTS U4522 ( .A0(n1120), .A1(n4810), .B0(n3044), .B1(n4799), .Y(n3594)
         );
  OAI22XLTS U4523 ( .A0(n1119), .A1(n4812), .B0(n3040), .B1(n4803), .Y(n3593)
         );
  OAI22XLTS U4524 ( .A0(n1118), .A1(n4810), .B0(n3036), .B1(n4805), .Y(n3592)
         );
  OAI22XLTS U4525 ( .A0(n1117), .A1(n4812), .B0(n3032), .B1(n4805), .Y(n3591)
         );
  OAI22XLTS U4526 ( .A0(n1116), .A1(n4807), .B0(n3028), .B1(n4804), .Y(n3590)
         );
  OAI22XLTS U4527 ( .A0(n1115), .A1(n4807), .B0(n3024), .B1(n4800), .Y(n3589)
         );
  OAI22XLTS U4528 ( .A0(n1114), .A1(n4807), .B0(n3020), .B1(n4800), .Y(n3588)
         );
  OAI22XLTS U4529 ( .A0(n1113), .A1(n4807), .B0(n3016), .B1(n4800), .Y(n3587)
         );
  OAI22XLTS U4530 ( .A0(n1112), .A1(n4808), .B0(n3012), .B1(n4800), .Y(n3586)
         );
  OAI22XLTS U4531 ( .A0(n1111), .A1(n4808), .B0(n3008), .B1(n4801), .Y(n3585)
         );
  OAI22XLTS U4532 ( .A0(n1110), .A1(n4808), .B0(n3004), .B1(n4801), .Y(n3584)
         );
  OAI22XLTS U4533 ( .A0(n1109), .A1(n4808), .B0(n3000), .B1(n4801), .Y(n3583)
         );
  OAI22XLTS U4534 ( .A0(n1108), .A1(n4809), .B0(n2996), .B1(n4801), .Y(n3582)
         );
  OAI22XLTS U4535 ( .A0(n1107), .A1(n4809), .B0(n2992), .B1(n4802), .Y(n3581)
         );
  OAI22XLTS U4536 ( .A0(n1106), .A1(n4809), .B0(n2988), .B1(n4802), .Y(n3580)
         );
  OAI22XLTS U4537 ( .A0(n1105), .A1(n4809), .B0(n2984), .B1(n4802), .Y(n3579)
         );
  OAI22XLTS U4538 ( .A0(n1104), .A1(n4810), .B0(n2977), .B1(n4802), .Y(n3578)
         );
  NOR3X1TS U4539 ( .A(prevRequesterPort_B[0]), .B(prevRequesterPort_B[1]), .C(
        n4579), .Y(n1529) );
  INVXLTS U4540 ( .A(\indexIncrementer_EAST[1] ), .Y(n5807) );
  AOI211X1TS U4541 ( .A0(prevRequesterPort_B[0]), .A1(prevRequesterPort_B[1]), 
        .B0(n5629), .C0(n5735), .Y(n1554) );
  AO22XLTS U4542 ( .A0(n2112), .A1(n3688), .B0(n3682), .B1(n5783), .Y(n4616)
         );
  NOR2X1TS U4543 ( .A(n5682), .B(n910), .Y(n1752) );
  NAND3BXLTS U4544 ( .AN(N6701), .B(n4607), .C(n4596), .Y(n2564) );
  CLKINVX2TS U4545 ( .A(n5225), .Y(n5224) );
  OAI21XLTS U4546 ( .A0(n3669), .A1(n2002), .B0(n5568), .Y(n2000) );
  CLKBUFX2TS U4547 ( .A(n4634), .Y(n4622) );
  CLKBUFX2TS U4548 ( .A(n4634), .Y(n4623) );
  CLKBUFX2TS U4549 ( .A(n4633), .Y(n4625) );
  CLKBUFX2TS U4550 ( .A(n4633), .Y(n4624) );
  CLKBUFX2TS U4551 ( .A(n4630), .Y(n4629) );
  CLKBUFX2TS U4552 ( .A(n4630), .Y(n4628) );
  CLKBUFX2TS U4553 ( .A(n4632), .Y(n4627) );
  CLKBUFX2TS U4554 ( .A(n4632), .Y(n4626) );
  INVX2TS U4555 ( .A(n5452), .Y(n5449) );
  INVX2TS U4556 ( .A(n5453), .Y(n5448) );
  INVX2TS U4557 ( .A(n5454), .Y(n5447) );
  INVX2TS U4558 ( .A(n5455), .Y(n5446) );
  INVX2TS U4559 ( .A(n5456), .Y(n5445) );
  INVX2TS U4560 ( .A(n5457), .Y(n5444) );
  INVX2TS U4561 ( .A(n5458), .Y(n5443) );
  INVX2TS U4562 ( .A(n5459), .Y(n5442) );
  INVX2TS U4563 ( .A(n5460), .Y(n5441) );
  INVX2TS U4564 ( .A(n5023), .Y(n5003) );
  CLKBUFX2TS U4565 ( .A(n4635), .Y(n4633) );
  CLKBUFX2TS U4566 ( .A(n4635), .Y(n4634) );
  CLKBUFX2TS U4567 ( .A(n4636), .Y(n4630) );
  CLKBUFX2TS U4568 ( .A(n4636), .Y(n4631) );
  CLKBUFX2TS U4569 ( .A(n4635), .Y(n4632) );
  CLKBUFX2TS U4570 ( .A(n4989), .Y(n4982) );
  CLKBUFX2TS U4571 ( .A(n4991), .Y(n4983) );
  CLKBUFX2TS U4572 ( .A(n4991), .Y(n4984) );
  CLKBUFX2TS U4573 ( .A(n4990), .Y(n4985) );
  CLKBUFX2TS U4574 ( .A(n4990), .Y(n4986) );
  CLKBUFX2TS U4575 ( .A(n4989), .Y(n4987) );
  CLKBUFX2TS U4576 ( .A(n4989), .Y(n4988) );
  CLKBUFX2TS U4577 ( .A(n4929), .Y(n4920) );
  CLKBUFX2TS U4578 ( .A(n4929), .Y(n4921) );
  CLKBUFX2TS U4579 ( .A(n4928), .Y(n4922) );
  CLKBUFX2TS U4580 ( .A(n4928), .Y(n4923) );
  CLKBUFX2TS U4581 ( .A(n4927), .Y(n4924) );
  CLKBUFX2TS U4582 ( .A(n4927), .Y(n4925) );
  CLKBUFX2TS U4583 ( .A(n4927), .Y(n4926) );
  CLKBUFX2TS U4584 ( .A(n4805), .Y(n4796) );
  CLKBUFX2TS U4585 ( .A(n4805), .Y(n4797) );
  CLKBUFX2TS U4586 ( .A(n4804), .Y(n4798) );
  CLKBUFX2TS U4587 ( .A(n4804), .Y(n4799) );
  CLKBUFX2TS U4588 ( .A(n4803), .Y(n4800) );
  CLKBUFX2TS U4589 ( .A(n4803), .Y(n4801) );
  CLKBUFX2TS U4590 ( .A(n4803), .Y(n4802) );
  INVX2TS U4591 ( .A(n4773), .Y(n4767) );
  INVX2TS U4592 ( .A(n4773), .Y(n4768) );
  INVX2TS U4593 ( .A(n4773), .Y(n4769) );
  INVX2TS U4594 ( .A(n4774), .Y(n4765) );
  INVX2TS U4595 ( .A(n4774), .Y(n4766) );
  CLKBUFX2TS U4596 ( .A(n5393), .Y(n5391) );
  CLKBUFX2TS U4597 ( .A(n5393), .Y(n5392) );
  CLKBUFX2TS U4598 ( .A(n5397), .Y(n5387) );
  CLKBUFX2TS U4599 ( .A(n5394), .Y(n5388) );
  CLKBUFX2TS U4600 ( .A(n5394), .Y(n5389) );
  CLKBUFX2TS U4601 ( .A(n5394), .Y(n5390) );
  CLKBUFX2TS U4602 ( .A(n4754), .Y(n4745) );
  CLKBUFX2TS U4603 ( .A(n4754), .Y(n4746) );
  CLKBUFX2TS U4604 ( .A(n4753), .Y(n4747) );
  CLKBUFX2TS U4605 ( .A(n4753), .Y(n4748) );
  CLKBUFX2TS U4606 ( .A(n4752), .Y(n4749) );
  CLKBUFX2TS U4607 ( .A(n4752), .Y(n4750) );
  CLKBUFX2TS U4608 ( .A(n4754), .Y(n4751) );
  INVX2TS U4609 ( .A(n5017), .Y(n5004) );
  INVX2TS U4610 ( .A(n5017), .Y(n5005) );
  INVX2TS U4611 ( .A(n5023), .Y(n5006) );
  INVX2TS U4612 ( .A(n5016), .Y(n5007) );
  INVX2TS U4613 ( .A(n5015), .Y(n5008) );
  INVX2TS U4614 ( .A(n5014), .Y(n5009) );
  INVX2TS U4615 ( .A(n5013), .Y(n5010) );
  CLKBUFX2TS U4616 ( .A(n4648), .Y(n4637) );
  CLKBUFX2TS U4617 ( .A(n4645), .Y(n4643) );
  CLKBUFX2TS U4618 ( .A(n4646), .Y(n4642) );
  CLKBUFX2TS U4619 ( .A(n4646), .Y(n4641) );
  CLKBUFX2TS U4620 ( .A(n4647), .Y(n4640) );
  CLKBUFX2TS U4621 ( .A(n4645), .Y(n4638) );
  CLKBUFX2TS U4622 ( .A(n4647), .Y(n4639) );
  CLKBUFX2TS U4623 ( .A(n4645), .Y(n4644) );
  CLKBUFX2TS U4624 ( .A(n4659), .Y(n4651) );
  CLKBUFX2TS U4625 ( .A(n4659), .Y(n4652) );
  CLKBUFX2TS U4626 ( .A(n4658), .Y(n4653) );
  CLKBUFX2TS U4627 ( .A(n4658), .Y(n4654) );
  CLKBUFX2TS U4628 ( .A(n4657), .Y(n4655) );
  CLKBUFX2TS U4629 ( .A(n4658), .Y(n4656) );
  CLKBUFX2TS U4630 ( .A(n5499), .Y(n5498) );
  CLKBUFX2TS U4631 ( .A(n5499), .Y(n5497) );
  CLKBUFX2TS U4632 ( .A(n5499), .Y(n5496) );
  CLKBUFX2TS U4633 ( .A(n1663), .Y(n5495) );
  CLKBUFX2TS U4634 ( .A(n5500), .Y(n5494) );
  CLKBUFX2TS U4635 ( .A(n5500), .Y(n5493) );
  CLKBUFX2TS U4636 ( .A(n5501), .Y(n5492) );
  CLKBUFX2TS U4637 ( .A(n5501), .Y(n5491) );
  CLKBUFX2TS U4638 ( .A(n5465), .Y(n5452) );
  CLKBUFX2TS U4639 ( .A(n5465), .Y(n5453) );
  CLKBUFX2TS U4640 ( .A(n5465), .Y(n5454) );
  CLKBUFX2TS U4641 ( .A(n5465), .Y(n5455) );
  CLKBUFX2TS U4642 ( .A(n5464), .Y(n5456) );
  CLKBUFX2TS U4643 ( .A(n5464), .Y(n5457) );
  CLKBUFX2TS U4644 ( .A(n5464), .Y(n5458) );
  CLKBUFX2TS U4645 ( .A(n5464), .Y(n5459) );
  CLKBUFX2TS U4646 ( .A(n5466), .Y(n5460) );
  INVX2TS U4647 ( .A(n5451), .Y(n5450) );
  CLKBUFX2TS U4648 ( .A(n5466), .Y(n5462) );
  CLKBUFX2TS U4649 ( .A(n3655), .Y(n5461) );
  CLKBUFX2TS U4650 ( .A(n5466), .Y(n5463) );
  CLKBUFX2TS U4651 ( .A(n2983), .Y(n4774) );
  INVX2TS U4652 ( .A(n2574), .Y(n4940) );
  INVX2TS U4653 ( .A(n4837), .Y(n4816) );
  INVX2TS U4654 ( .A(n5078), .Y(n5064) );
  INVX2TS U4655 ( .A(n4897), .Y(n4878) );
  CLKBUFX2TS U4656 ( .A(n2568), .Y(n4991) );
  CLKBUFX2TS U4657 ( .A(n2568), .Y(n4990) );
  CLKBUFX2TS U4658 ( .A(n2568), .Y(n4989) );
  CLKBUFX2TS U4659 ( .A(n2704), .Y(n4929) );
  CLKBUFX2TS U4660 ( .A(n2704), .Y(n4928) );
  CLKBUFX2TS U4661 ( .A(n2704), .Y(n4927) );
  CLKBUFX2TS U4662 ( .A(n2978), .Y(n4805) );
  CLKBUFX2TS U4663 ( .A(n2978), .Y(n4804) );
  CLKBUFX2TS U4664 ( .A(n2978), .Y(n4803) );
  CLKBUFX2TS U4665 ( .A(n5397), .Y(n5396) );
  CLKBUFX2TS U4666 ( .A(n5397), .Y(n5395) );
  CLKBUFX2TS U4667 ( .A(n5398), .Y(n5393) );
  CLKBUFX2TS U4668 ( .A(n5398), .Y(n5394) );
  CLKBUFX2TS U4669 ( .A(n5760), .Y(n4636) );
  CLKBUFX2TS U4670 ( .A(n5760), .Y(n4635) );
  CLKBUFX2TS U4671 ( .A(n4813), .Y(n4806) );
  CLKBUFX2TS U4672 ( .A(n4811), .Y(n4807) );
  CLKBUFX2TS U4673 ( .A(n4811), .Y(n4808) );
  CLKBUFX2TS U4674 ( .A(n4810), .Y(n4809) );
  CLKBUFX2TS U4675 ( .A(n4867), .Y(n4858) );
  CLKBUFX2TS U4676 ( .A(n5115), .Y(n5106) );
  CLKBUFX2TS U4677 ( .A(n4867), .Y(n4859) );
  CLKBUFX2TS U4678 ( .A(n5115), .Y(n5107) );
  CLKBUFX2TS U4679 ( .A(n4866), .Y(n4860) );
  CLKBUFX2TS U4680 ( .A(n5114), .Y(n5108) );
  CLKBUFX2TS U4681 ( .A(n4866), .Y(n4861) );
  CLKBUFX2TS U4682 ( .A(n5114), .Y(n5109) );
  CLKBUFX2TS U4683 ( .A(n4866), .Y(n4862) );
  CLKBUFX2TS U4684 ( .A(n5114), .Y(n5110) );
  CLKBUFX2TS U4685 ( .A(n4865), .Y(n4863) );
  CLKBUFX2TS U4686 ( .A(n5113), .Y(n5111) );
  CLKBUFX2TS U4687 ( .A(n4865), .Y(n4864) );
  CLKBUFX2TS U4688 ( .A(n5113), .Y(n5112) );
  CLKBUFX2TS U4689 ( .A(n5053), .Y(n5044) );
  CLKBUFX2TS U4690 ( .A(n5053), .Y(n5045) );
  CLKBUFX2TS U4691 ( .A(n5052), .Y(n5046) );
  CLKBUFX2TS U4692 ( .A(n5052), .Y(n5047) );
  CLKBUFX2TS U4693 ( .A(n5052), .Y(n5048) );
  CLKBUFX2TS U4694 ( .A(n5051), .Y(n5049) );
  CLKBUFX2TS U4695 ( .A(n5051), .Y(n5050) );
  INVX2TS U4696 ( .A(n4773), .Y(n4770) );
  INVX2TS U4697 ( .A(n4784), .Y(n4771) );
  INVX2TS U4698 ( .A(n4780), .Y(n4772) );
  INVX2TS U4699 ( .A(n5428), .Y(n5415) );
  CLKBUFX2TS U4700 ( .A(n5022), .Y(n5013) );
  CLKBUFX2TS U4701 ( .A(n5022), .Y(n5014) );
  CLKBUFX2TS U4702 ( .A(n5022), .Y(n5015) );
  CLKBUFX2TS U4703 ( .A(n5022), .Y(n5016) );
  CLKBUFX2TS U4704 ( .A(n2436), .Y(n5017) );
  CLKBUFX2TS U4705 ( .A(n5021), .Y(n5018) );
  CLKBUFX2TS U4706 ( .A(n5021), .Y(n5019) );
  CLKBUFX2TS U4707 ( .A(n5021), .Y(n5020) );
  CLKBUFX2TS U4708 ( .A(n3116), .Y(n4754) );
  CLKBUFX2TS U4709 ( .A(n3116), .Y(n4753) );
  CLKBUFX2TS U4710 ( .A(n3116), .Y(n4752) );
  CLKBUFX2TS U4711 ( .A(n4649), .Y(n4645) );
  CLKBUFX2TS U4712 ( .A(n4649), .Y(n4646) );
  CLKBUFX2TS U4713 ( .A(n4649), .Y(n4647) );
  CLKBUFX2TS U4714 ( .A(n4764), .Y(n4755) );
  CLKBUFX2TS U4715 ( .A(n4761), .Y(n4756) );
  CLKBUFX2TS U4716 ( .A(n4761), .Y(n4757) );
  CLKBUFX2TS U4717 ( .A(n4761), .Y(n4758) );
  CLKBUFX2TS U4718 ( .A(n4760), .Y(n4759) );
  CLKBUFX2TS U4719 ( .A(n4783), .Y(n4775) );
  CLKBUFX2TS U4720 ( .A(n4783), .Y(n4776) );
  CLKBUFX2TS U4721 ( .A(n4782), .Y(n4777) );
  CLKBUFX2TS U4722 ( .A(n4782), .Y(n4778) );
  CLKBUFX2TS U4723 ( .A(n4781), .Y(n4779) );
  INVX2TS U4724 ( .A(n4830), .Y(n4817) );
  INVX2TS U4725 ( .A(n4954), .Y(n4941) );
  INVX2TS U4726 ( .A(n5076), .Y(n5065) );
  INVX2TS U4727 ( .A(n4829), .Y(n4818) );
  INVX2TS U4728 ( .A(n4961), .Y(n4942) );
  INVX2TS U4729 ( .A(n5085), .Y(n5066) );
  INVX2TS U4730 ( .A(n4829), .Y(n4819) );
  INVX2TS U4731 ( .A(n4961), .Y(n4943) );
  INVX2TS U4732 ( .A(n5077), .Y(n5067) );
  INVX2TS U4733 ( .A(n4828), .Y(n4820) );
  INVX2TS U4734 ( .A(n4953), .Y(n4944) );
  INVX2TS U4735 ( .A(n5076), .Y(n5068) );
  INVX2TS U4736 ( .A(n4827), .Y(n4821) );
  INVX2TS U4737 ( .A(n4952), .Y(n4945) );
  INVX2TS U4738 ( .A(n5075), .Y(n5069) );
  INVX2TS U4739 ( .A(n4826), .Y(n4822) );
  INVX2TS U4740 ( .A(n4951), .Y(n4946) );
  INVX2TS U4741 ( .A(n5074), .Y(n5070) );
  INVX2TS U4742 ( .A(n4825), .Y(n4823) );
  INVX2TS U4743 ( .A(n4950), .Y(n4947) );
  INVX2TS U4744 ( .A(n5073), .Y(n5071) );
  INVX2TS U4745 ( .A(n4899), .Y(n4879) );
  INVX2TS U4746 ( .A(n4899), .Y(n4880) );
  INVX2TS U4747 ( .A(n4891), .Y(n4881) );
  INVX2TS U4748 ( .A(n4891), .Y(n4882) );
  INVX2TS U4749 ( .A(n4890), .Y(n4883) );
  INVX2TS U4750 ( .A(n4889), .Y(n4884) );
  INVX2TS U4751 ( .A(n4888), .Y(n4885) );
  INVX2TS U4752 ( .A(n5189), .Y(n5182) );
  INVX2TS U4753 ( .A(n5269), .Y(n5260) );
  INVX2TS U4754 ( .A(n5365), .Y(n5354) );
  INVX2TS U4755 ( .A(n5229), .Y(n5221) );
  INVX2TS U4756 ( .A(n5322), .Y(n5315) );
  INVX2TS U4757 ( .A(n5190), .Y(n5181) );
  INVX2TS U4758 ( .A(n5265), .Y(n5259) );
  INVX2TS U4759 ( .A(n5359), .Y(n5353) );
  INVX2TS U4760 ( .A(n5191), .Y(n5180) );
  INVX2TS U4761 ( .A(n5266), .Y(n5258) );
  INVX2TS U4762 ( .A(n5360), .Y(n5352) );
  INVX2TS U4763 ( .A(n5192), .Y(n5179) );
  INVX2TS U4764 ( .A(n5267), .Y(n5257) );
  INVX2TS U4765 ( .A(n5361), .Y(n5351) );
  INVX2TS U4766 ( .A(n5268), .Y(n5256) );
  INVX2TS U4767 ( .A(n5199), .Y(n5178) );
  INVX2TS U4768 ( .A(n5269), .Y(n5255) );
  INVX2TS U4769 ( .A(n5363), .Y(n5350) );
  INVX2TS U4770 ( .A(n5192), .Y(n5177) );
  INVX2TS U4771 ( .A(n5270), .Y(n5254) );
  INVX2TS U4772 ( .A(n5364), .Y(n5349) );
  INVX2TS U4773 ( .A(n5194), .Y(n5176) );
  INVX2TS U4774 ( .A(n5365), .Y(n5348) );
  INVX2TS U4775 ( .A(n5226), .Y(n5220) );
  INVX2TS U4776 ( .A(n5227), .Y(n5219) );
  INVX2TS U4777 ( .A(n5228), .Y(n5218) );
  INVX2TS U4778 ( .A(n5230), .Y(n5217) );
  INVX2TS U4779 ( .A(n5231), .Y(n5216) );
  INVX2TS U4780 ( .A(n5232), .Y(n5215) );
  INVX2TS U4781 ( .A(n5320), .Y(n5314) );
  INVX2TS U4782 ( .A(n5321), .Y(n5313) );
  INVX2TS U4783 ( .A(n5322), .Y(n5312) );
  INVX2TS U4784 ( .A(n5323), .Y(n5311) );
  INVX2TS U4785 ( .A(n5324), .Y(n5310) );
  INVX2TS U4786 ( .A(n5325), .Y(n5309) );
  INVX2TS U4787 ( .A(n5187), .Y(n5184) );
  INVX2TS U4788 ( .A(n5270), .Y(n5262) );
  INVX2TS U4789 ( .A(n5360), .Y(n5356) );
  INVX2TS U4790 ( .A(n5188), .Y(n5183) );
  INVX2TS U4791 ( .A(n5264), .Y(n5261) );
  INVX2TS U4792 ( .A(n5358), .Y(n5355) );
  INVX2TS U4793 ( .A(n5228), .Y(n5223) );
  INVX2TS U4794 ( .A(n5231), .Y(n5222) );
  INVX2TS U4795 ( .A(n5319), .Y(n5317) );
  INVX2TS U4796 ( .A(n5323), .Y(n5316) );
  CLKBUFX2TS U4797 ( .A(n4781), .Y(n4780) );
  CLKBUFX2TS U4798 ( .A(n5771), .Y(n4648) );
  CLKBUFX2TS U4799 ( .A(n1666), .Y(n5479) );
  CLKBUFX2TS U4800 ( .A(n5489), .Y(n5480) );
  CLKBUFX2TS U4801 ( .A(n5489), .Y(n5481) );
  CLKBUFX2TS U4802 ( .A(n5488), .Y(n5482) );
  CLKBUFX2TS U4803 ( .A(n5488), .Y(n5483) );
  CLKBUFX2TS U4804 ( .A(n5490), .Y(n5484) );
  CLKBUFX2TS U4805 ( .A(n5487), .Y(n5485) );
  CLKBUFX2TS U4806 ( .A(n5487), .Y(n5486) );
  CLKBUFX2TS U4807 ( .A(n5157), .Y(n5155) );
  CLKBUFX2TS U4808 ( .A(n5157), .Y(n5156) );
  CLKBUFX2TS U4809 ( .A(n5161), .Y(n5152) );
  CLKBUFX2TS U4810 ( .A(n5158), .Y(n5153) );
  CLKBUFX2TS U4811 ( .A(n5158), .Y(n5154) );
  INVX2TS U4812 ( .A(n5425), .Y(n5416) );
  INVX2TS U4813 ( .A(n5427), .Y(n5417) );
  INVX2TS U4814 ( .A(n5425), .Y(n5419) );
  INVX2TS U4815 ( .A(n5425), .Y(n5418) );
  INVX2TS U4816 ( .A(n5426), .Y(n5422) );
  INVX2TS U4817 ( .A(n5426), .Y(n5421) );
  INVX2TS U4818 ( .A(n5426), .Y(n5420) );
  INVX2TS U4819 ( .A(n5427), .Y(n5424) );
  INVX2TS U4820 ( .A(n5427), .Y(n5423) );
  NOR2X1TS U4821 ( .A(n4550), .B(n4650), .Y(n2197) );
  CLKBUFX2TS U4822 ( .A(n4661), .Y(n4659) );
  CLKBUFX2TS U4823 ( .A(n4661), .Y(n4658) );
  CLKBUFX2TS U4824 ( .A(n4662), .Y(n4657) );
  CLKBUFX2TS U4825 ( .A(n1663), .Y(n5500) );
  CLKBUFX2TS U4826 ( .A(n1663), .Y(n5501) );
  CLKBUFX2TS U4827 ( .A(n5502), .Y(n5499) );
  CLKBUFX2TS U4828 ( .A(n4660), .Y(n4650) );
  CLKBUFX2TS U4829 ( .A(n4661), .Y(n4660) );
  CLKBUFX2TS U4830 ( .A(n5472), .Y(n5471) );
  CLKBUFX2TS U4831 ( .A(n5472), .Y(n5470) );
  CLKBUFX2TS U4832 ( .A(n5473), .Y(n5469) );
  CLKBUFX2TS U4833 ( .A(n5473), .Y(n5468) );
  CLKBUFX2TS U4834 ( .A(n5474), .Y(n5467) );
  CLKBUFX2TS U4835 ( .A(n5520), .Y(n5519) );
  CLKBUFX2TS U4836 ( .A(n5520), .Y(n5518) );
  CLKBUFX2TS U4837 ( .A(n5521), .Y(n5517) );
  CLKBUFX2TS U4838 ( .A(n5521), .Y(n5516) );
  CLKBUFX2TS U4839 ( .A(n5522), .Y(n5515) );
  CLKBUFX2TS U4840 ( .A(n5466), .Y(n5451) );
  CLKBUFX2TS U4841 ( .A(n3655), .Y(n5466) );
  CLKBUFX2TS U4842 ( .A(n3655), .Y(n5465) );
  CLKBUFX2TS U4843 ( .A(n3655), .Y(n5464) );
  INVX2TS U4844 ( .A(n2271), .Y(n5974) );
  NAND2X1TS U4845 ( .A(n2976), .B(n5721), .Y(n2978) );
  CLKBUFX2TS U4846 ( .A(n5202), .Y(n5186) );
  CLKBUFX2TS U4847 ( .A(n5241), .Y(n5225) );
  CLKBUFX2TS U4848 ( .A(n2295), .Y(n5078) );
  CLKBUFX2TS U4849 ( .A(n2842), .Y(n4867) );
  CLKBUFX2TS U4850 ( .A(n2289), .Y(n5115) );
  CLKBUFX2TS U4851 ( .A(n2842), .Y(n4866) );
  CLKBUFX2TS U4852 ( .A(n2289), .Y(n5114) );
  CLKBUFX2TS U4853 ( .A(n2842), .Y(n4865) );
  CLKBUFX2TS U4854 ( .A(n2289), .Y(n5113) );
  CLKBUFX2TS U4855 ( .A(n2430), .Y(n5053) );
  CLKBUFX2TS U4856 ( .A(n2430), .Y(n5052) );
  CLKBUFX2TS U4857 ( .A(n2430), .Y(n5051) );
  CLKBUFX2TS U4858 ( .A(n4814), .Y(n4813) );
  CLKBUFX2TS U4859 ( .A(n4814), .Y(n4812) );
  CLKBUFX2TS U4860 ( .A(n4815), .Y(n4811) );
  CLKBUFX2TS U4861 ( .A(n4815), .Y(n4810) );
  CLKBUFX2TS U4862 ( .A(n1825), .Y(n5397) );
  CLKBUFX2TS U4863 ( .A(n5000), .Y(n4993) );
  CLKBUFX2TS U4864 ( .A(n5000), .Y(n4994) );
  CLKBUFX2TS U4865 ( .A(n4999), .Y(n4995) );
  CLKBUFX2TS U4866 ( .A(n4998), .Y(n4996) );
  CLKBUFX2TS U4867 ( .A(n4999), .Y(n4997) );
  CLKBUFX2TS U4868 ( .A(n4937), .Y(n4930) );
  CLKBUFX2TS U4869 ( .A(n4935), .Y(n4931) );
  CLKBUFX2TS U4870 ( .A(n4935), .Y(n4932) );
  CLKBUFX2TS U4871 ( .A(n4934), .Y(n4933) );
  CLKBUFX2TS U4872 ( .A(n1825), .Y(n5398) );
  INVX2TS U4873 ( .A(n1598), .Y(n5760) );
  CLKBUFX2TS U4874 ( .A(n4744), .Y(n4735) );
  CLKBUFX2TS U4875 ( .A(n4744), .Y(n4736) );
  CLKBUFX2TS U4876 ( .A(n4743), .Y(n4737) );
  CLKBUFX2TS U4877 ( .A(n4743), .Y(n4738) );
  CLKBUFX2TS U4878 ( .A(n4742), .Y(n4739) );
  CLKBUFX2TS U4879 ( .A(n3117), .Y(n4740) );
  CLKBUFX2TS U4880 ( .A(n4742), .Y(n4741) );
  NAND2X1TS U4881 ( .A(n4763), .B(n5723), .Y(n3116) );
  CLKBUFX2TS U4882 ( .A(n5190), .Y(n5189) );
  CLKBUFX2TS U4883 ( .A(n5193), .Y(n5187) );
  CLKBUFX2TS U4884 ( .A(n5193), .Y(n5188) );
  CLKBUFX2TS U4885 ( .A(n5279), .Y(n5264) );
  CLKBUFX2TS U4886 ( .A(n5373), .Y(n5358) );
  CLKBUFX2TS U4887 ( .A(n5335), .Y(n5319) );
  CLKBUFX2TS U4888 ( .A(n5201), .Y(n5190) );
  CLKBUFX2TS U4889 ( .A(n5278), .Y(n5265) );
  CLKBUFX2TS U4890 ( .A(n5372), .Y(n5359) );
  CLKBUFX2TS U4891 ( .A(n5201), .Y(n5191) );
  CLKBUFX2TS U4892 ( .A(n5278), .Y(n5266) );
  CLKBUFX2TS U4893 ( .A(n5372), .Y(n5360) );
  CLKBUFX2TS U4894 ( .A(n5201), .Y(n5192) );
  CLKBUFX2TS U4895 ( .A(n5278), .Y(n5267) );
  CLKBUFX2TS U4896 ( .A(n5372), .Y(n5361) );
  CLKBUFX2TS U4897 ( .A(n5201), .Y(n5193) );
  CLKBUFX2TS U4898 ( .A(n5278), .Y(n5268) );
  CLKBUFX2TS U4899 ( .A(n5372), .Y(n5362) );
  CLKBUFX2TS U4900 ( .A(n5267), .Y(n5269) );
  CLKBUFX2TS U4901 ( .A(n5362), .Y(n5363) );
  CLKBUFX2TS U4902 ( .A(n5266), .Y(n5270) );
  CLKBUFX2TS U4903 ( .A(n5361), .Y(n5364) );
  CLKBUFX2TS U4904 ( .A(n5187), .Y(n5194) );
  CLKBUFX2TS U4905 ( .A(n5268), .Y(n5271) );
  CLKBUFX2TS U4906 ( .A(n5362), .Y(n5365) );
  CLKBUFX2TS U4907 ( .A(n5240), .Y(n5226) );
  CLKBUFX2TS U4908 ( .A(n5240), .Y(n5227) );
  CLKBUFX2TS U4909 ( .A(n5240), .Y(n5228) );
  CLKBUFX2TS U4910 ( .A(n5240), .Y(n5229) );
  CLKBUFX2TS U4911 ( .A(n5239), .Y(n5230) );
  CLKBUFX2TS U4912 ( .A(n5239), .Y(n5231) );
  CLKBUFX2TS U4913 ( .A(n5239), .Y(n5232) );
  CLKBUFX2TS U4914 ( .A(n5334), .Y(n5320) );
  CLKBUFX2TS U4915 ( .A(n5334), .Y(n5321) );
  CLKBUFX2TS U4916 ( .A(n5334), .Y(n5322) );
  CLKBUFX2TS U4917 ( .A(n5334), .Y(n5323) );
  CLKBUFX2TS U4918 ( .A(n5333), .Y(n5324) );
  CLKBUFX2TS U4919 ( .A(n5333), .Y(n5325) );
  CLKBUFX2TS U4920 ( .A(n5333), .Y(n5326) );
  CLKBUFX2TS U4921 ( .A(n4960), .Y(n4950) );
  CLKBUFX2TS U4922 ( .A(n5084), .Y(n5073) );
  CLKBUFX2TS U4923 ( .A(n4960), .Y(n4951) );
  CLKBUFX2TS U4924 ( .A(n5084), .Y(n5074) );
  CLKBUFX2TS U4925 ( .A(n4960), .Y(n4952) );
  CLKBUFX2TS U4926 ( .A(n5084), .Y(n5075) );
  CLKBUFX2TS U4927 ( .A(n4960), .Y(n4953) );
  CLKBUFX2TS U4928 ( .A(n5084), .Y(n5076) );
  CLKBUFX2TS U4929 ( .A(n5085), .Y(n5077) );
  CLKBUFX2TS U4930 ( .A(n4951), .Y(n4954) );
  CLKBUFX2TS U4931 ( .A(n4836), .Y(n4825) );
  CLKBUFX2TS U4932 ( .A(n4836), .Y(n4826) );
  CLKBUFX2TS U4933 ( .A(n4836), .Y(n4827) );
  CLKBUFX2TS U4934 ( .A(n4836), .Y(n4828) );
  CLKBUFX2TS U4935 ( .A(n4837), .Y(n4829) );
  CLKBUFX2TS U4936 ( .A(n2848), .Y(n4830) );
  CLKBUFX2TS U4937 ( .A(n5023), .Y(n5012) );
  CLKBUFX2TS U4938 ( .A(n5002), .Y(n5023) );
  CLKBUFX2TS U4939 ( .A(n4898), .Y(n4888) );
  CLKBUFX2TS U4940 ( .A(n4898), .Y(n4889) );
  CLKBUFX2TS U4941 ( .A(n4898), .Y(n4890) );
  CLKBUFX2TS U4942 ( .A(n4898), .Y(n4891) );
  CLKBUFX2TS U4943 ( .A(n5200), .Y(n5198) );
  CLKBUFX2TS U4944 ( .A(n5277), .Y(n5275) );
  CLKBUFX2TS U4945 ( .A(n5371), .Y(n5369) );
  CLKBUFX2TS U4946 ( .A(n5202), .Y(n5195) );
  CLKBUFX2TS U4947 ( .A(n5265), .Y(n5272) );
  CLKBUFX2TS U4948 ( .A(n5359), .Y(n5366) );
  CLKBUFX2TS U4949 ( .A(n5200), .Y(n5196) );
  CLKBUFX2TS U4950 ( .A(n5277), .Y(n5273) );
  CLKBUFX2TS U4951 ( .A(n5371), .Y(n5367) );
  CLKBUFX2TS U4952 ( .A(n5200), .Y(n5197) );
  CLKBUFX2TS U4953 ( .A(n5277), .Y(n5274) );
  CLKBUFX2TS U4954 ( .A(n5371), .Y(n5368) );
  CLKBUFX2TS U4955 ( .A(n5238), .Y(n5236) );
  CLKBUFX2TS U4956 ( .A(n5239), .Y(n5233) );
  CLKBUFX2TS U4957 ( .A(n5238), .Y(n5234) );
  CLKBUFX2TS U4958 ( .A(n5238), .Y(n5235) );
  CLKBUFX2TS U4959 ( .A(n5332), .Y(n5330) );
  CLKBUFX2TS U4960 ( .A(n5333), .Y(n5327) );
  CLKBUFX2TS U4961 ( .A(n5332), .Y(n5328) );
  CLKBUFX2TS U4962 ( .A(n5332), .Y(n5329) );
  CLKBUFX2TS U4963 ( .A(n4959), .Y(n4955) );
  CLKBUFX2TS U4964 ( .A(n5083), .Y(n5079) );
  CLKBUFX2TS U4965 ( .A(n4959), .Y(n4956) );
  CLKBUFX2TS U4966 ( .A(n5083), .Y(n5080) );
  CLKBUFX2TS U4967 ( .A(n4959), .Y(n4957) );
  CLKBUFX2TS U4968 ( .A(n5083), .Y(n5081) );
  CLKBUFX2TS U4969 ( .A(n4835), .Y(n4831) );
  CLKBUFX2TS U4970 ( .A(n4835), .Y(n4832) );
  CLKBUFX2TS U4971 ( .A(n4835), .Y(n4833) );
  CLKBUFX2TS U4972 ( .A(n4896), .Y(n4892) );
  CLKBUFX2TS U4973 ( .A(n4896), .Y(n4893) );
  CLKBUFX2TS U4974 ( .A(n4896), .Y(n4894) );
  CLKBUFX2TS U4975 ( .A(n5428), .Y(n5427) );
  CLKBUFX2TS U4976 ( .A(n5200), .Y(n5199) );
  CLKBUFX2TS U4977 ( .A(n5277), .Y(n5276) );
  CLKBUFX2TS U4978 ( .A(n5371), .Y(n5370) );
  CLKBUFX2TS U4979 ( .A(n5238), .Y(n5237) );
  CLKBUFX2TS U4980 ( .A(n5332), .Y(n5331) );
  CLKBUFX2TS U4981 ( .A(n4785), .Y(n4784) );
  CLKBUFX2TS U4982 ( .A(n4785), .Y(n4783) );
  CLKBUFX2TS U4983 ( .A(n4785), .Y(n4782) );
  CLKBUFX2TS U4984 ( .A(n4785), .Y(n4781) );
  CLKBUFX2TS U4985 ( .A(n5490), .Y(n5489) );
  CLKBUFX2TS U4986 ( .A(n1666), .Y(n5488) );
  CLKBUFX2TS U4987 ( .A(n5162), .Y(n5161) );
  CLKBUFX2TS U4988 ( .A(n5162), .Y(n5160) );
  CLKBUFX2TS U4989 ( .A(n5162), .Y(n5159) );
  CLKBUFX2TS U4990 ( .A(n5490), .Y(n5487) );
  CLKBUFX2TS U4991 ( .A(n5163), .Y(n5157) );
  CLKBUFX2TS U4992 ( .A(n5163), .Y(n5158) );
  CLKBUFX2TS U4993 ( .A(n4764), .Y(n4761) );
  CLKBUFX2TS U4994 ( .A(n4764), .Y(n4760) );
  CLKBUFX2TS U4995 ( .A(n4835), .Y(n4834) );
  CLKBUFX2TS U4996 ( .A(n4959), .Y(n4958) );
  CLKBUFX2TS U4997 ( .A(n5083), .Y(n5082) );
  CLKBUFX2TS U4998 ( .A(n4896), .Y(n4895) );
  CLKBUFX2TS U4999 ( .A(n5771), .Y(n4649) );
  CLKBUFX2TS U5000 ( .A(n4763), .Y(n4762) );
  CLKBUFX2TS U5001 ( .A(n4795), .Y(n4786) );
  CLKBUFX2TS U5002 ( .A(n4795), .Y(n4787) );
  CLKBUFX2TS U5003 ( .A(n4794), .Y(n4788) );
  CLKBUFX2TS U5004 ( .A(n4794), .Y(n4789) );
  CLKBUFX2TS U5005 ( .A(n4795), .Y(n4790) );
  CLKBUFX2TS U5006 ( .A(n4793), .Y(n4791) );
  CLKBUFX2TS U5007 ( .A(n4793), .Y(n4792) );
  INVX2TS U5008 ( .A(n5137), .Y(n5135) );
  INVX2TS U5009 ( .A(n5140), .Y(n5134) );
  INVX2TS U5010 ( .A(n5142), .Y(n5126) );
  INVX2TS U5011 ( .A(n5141), .Y(n5127) );
  INVX2TS U5012 ( .A(n5140), .Y(n5128) );
  INVX2TS U5013 ( .A(n5139), .Y(n5129) );
  INVX2TS U5014 ( .A(n5138), .Y(n5130) );
  INVX2TS U5015 ( .A(n5137), .Y(n5131) );
  INVX2TS U5016 ( .A(n5136), .Y(n5132) );
  INVX2TS U5017 ( .A(n5139), .Y(n5133) );
  CLKBUFX2TS U5018 ( .A(n5002), .Y(n5022) );
  CLKBUFX2TS U5019 ( .A(n5002), .Y(n5021) );
  INVX2TS U5020 ( .A(n4613), .Y(n5527) );
  CLKBUFX2TS U5021 ( .A(n5477), .Y(n5474) );
  CLKBUFX2TS U5022 ( .A(n5477), .Y(n5475) );
  CLKBUFX2TS U5023 ( .A(n5477), .Y(n5476) );
  CLKBUFX2TS U5024 ( .A(n5525), .Y(n5522) );
  CLKBUFX2TS U5025 ( .A(n5525), .Y(n5523) );
  CLKBUFX2TS U5026 ( .A(n5525), .Y(n5524) );
  CLKBUFX2TS U5027 ( .A(n5478), .Y(n5472) );
  CLKBUFX2TS U5028 ( .A(n5478), .Y(n5473) );
  CLKBUFX2TS U5029 ( .A(n5526), .Y(n5520) );
  CLKBUFX2TS U5030 ( .A(n5526), .Y(n5521) );
  CLKBUFX2TS U5031 ( .A(n5798), .Y(n4662) );
  CLKBUFX2TS U5032 ( .A(n5798), .Y(n4661) );
  CLKBUFX2TS U5033 ( .A(n5511), .Y(n5510) );
  CLKBUFX2TS U5034 ( .A(n5511), .Y(n5509) );
  CLKBUFX2TS U5035 ( .A(n5511), .Y(n5508) );
  CLKBUFX2TS U5036 ( .A(n1645), .Y(n5507) );
  CLKBUFX2TS U5037 ( .A(n5512), .Y(n5506) );
  CLKBUFX2TS U5038 ( .A(n5512), .Y(n5505) );
  CLKBUFX2TS U5039 ( .A(n5513), .Y(n5504) );
  CLKBUFX2TS U5040 ( .A(n5513), .Y(n5503) );
  CLKBUFX2TS U5041 ( .A(n5438), .Y(n5430) );
  CLKBUFX2TS U5042 ( .A(n5438), .Y(n5429) );
  CLKBUFX2TS U5043 ( .A(n1663), .Y(n5502) );
  CLKBUFX2TS U5044 ( .A(n5436), .Y(n5435) );
  CLKBUFX2TS U5045 ( .A(n5436), .Y(n5434) );
  CLKBUFX2TS U5046 ( .A(n5437), .Y(n5433) );
  CLKBUFX2TS U5047 ( .A(n5437), .Y(n5432) );
  CLKBUFX2TS U5048 ( .A(n5439), .Y(n5431) );
  CLKBUFX2TS U5049 ( .A(n5610), .Y(n5602) );
  CLKBUFX2TS U5050 ( .A(n5610), .Y(n5603) );
  CLKBUFX2TS U5051 ( .A(n5609), .Y(n5604) );
  CLKBUFX2TS U5052 ( .A(n5609), .Y(n5605) );
  CLKBUFX2TS U5053 ( .A(n5608), .Y(n5606) );
  CLKBUFX2TS U5054 ( .A(n5608), .Y(n5607) );
  INVX2TS U5055 ( .A(N10004), .Y(n5799) );
  INVX2TS U5056 ( .A(n5546), .Y(n5533) );
  INVX2TS U5057 ( .A(n5545), .Y(n5534) );
  INVX2TS U5058 ( .A(n5544), .Y(n5535) );
  INVX2TS U5059 ( .A(n5543), .Y(n5536) );
  INVX2TS U5060 ( .A(n5547), .Y(n5528) );
  INVX2TS U5061 ( .A(n5552), .Y(n5529) );
  INVX2TS U5062 ( .A(n5558), .Y(n5530) );
  INVX2TS U5063 ( .A(n5548), .Y(n5531) );
  INVX2TS U5064 ( .A(n5547), .Y(n5532) );
  INVX2TS U5065 ( .A(n5542), .Y(n5537) );
  INVX2TS U5066 ( .A(n5541), .Y(n5538) );
  INVX2TS U5067 ( .A(n5413), .Y(n5409) );
  NOR2X1TS U5068 ( .A(n5413), .B(n5591), .Y(n2271) );
  INVX2TS U5069 ( .A(n5595), .Y(n5565) );
  INVX2TS U5070 ( .A(n5601), .Y(n5566) );
  INVX2TS U5071 ( .A(n5595), .Y(n5567) );
  INVX2TS U5072 ( .A(n5586), .Y(n5568) );
  INVX2TS U5073 ( .A(n5586), .Y(n5569) );
  INVX2TS U5074 ( .A(n5586), .Y(n5570) );
  INVX2TS U5075 ( .A(n5590), .Y(n5583) );
  INVX2TS U5076 ( .A(n5590), .Y(n5584) );
  INVX2TS U5077 ( .A(n5599), .Y(n5585) );
  INVX2TS U5078 ( .A(n5596), .Y(n5562) );
  INVX2TS U5079 ( .A(n5411), .Y(n5404) );
  INVX2TS U5080 ( .A(n5411), .Y(n5403) );
  INVX2TS U5081 ( .A(n5411), .Y(n5402) );
  INVX2TS U5082 ( .A(n5413), .Y(n5408) );
  INVX2TS U5083 ( .A(n5413), .Y(n5407) );
  INVX2TS U5084 ( .A(n5412), .Y(n5406) );
  INVX2TS U5085 ( .A(n5412), .Y(n5405) );
  INVX2TS U5086 ( .A(n5600), .Y(n5563) );
  INVX2TS U5087 ( .A(n5596), .Y(n5564) );
  INVX2TS U5088 ( .A(n5587), .Y(n5573) );
  INVX2TS U5089 ( .A(n5601), .Y(n5571) );
  INVX2TS U5090 ( .A(n5597), .Y(n5572) );
  INVX2TS U5091 ( .A(n5589), .Y(n5581) );
  INVX2TS U5092 ( .A(n5589), .Y(n5580) );
  INVX2TS U5093 ( .A(n5589), .Y(n5579) );
  INVX2TS U5094 ( .A(n5588), .Y(n5578) );
  INVX2TS U5095 ( .A(n5588), .Y(n5577) );
  INVX2TS U5096 ( .A(n5588), .Y(n5576) );
  INVX2TS U5097 ( .A(n5587), .Y(n5575) );
  INVX2TS U5098 ( .A(n5587), .Y(n5574) );
  INVX2TS U5099 ( .A(n5590), .Y(n5582) );
  INVX2TS U5100 ( .A(N6373), .Y(n5774) );
  NAND2X1TS U5101 ( .A(n2280), .B(n2090), .Y(n1598) );
  AOI21X1TS U5102 ( .A0(n4545), .A1(n5763), .B0(n5739), .Y(n2236) );
  NAND2X1TS U5103 ( .A(n5054), .B(n5722), .Y(n2430) );
  NAND2X1TS U5104 ( .A(n2199), .B(n5415), .Y(n1825) );
  AOI21X1TS U5105 ( .A0(n2090), .A1(n5762), .B0(n5740), .Y(n2265) );
  AOI21X1TS U5106 ( .A0(n4544), .A1(n5765), .B0(n5739), .Y(n2211) );
  AOI21X1TS U5107 ( .A0(n2090), .A1(n5770), .B0(n5739), .Y(n2223) );
  INVX2TS U5108 ( .A(n2085), .Y(n5766) );
  INVX2TS U5109 ( .A(n3706), .Y(n5763) );
  INVX2TS U5110 ( .A(n3708), .Y(n5770) );
  CLKBUFX2TS U5111 ( .A(n3117), .Y(n4744) );
  CLKBUFX2TS U5112 ( .A(n3117), .Y(n4743) );
  CLKBUFX2TS U5113 ( .A(n3117), .Y(n4742) );
  CLKBUFX2TS U5114 ( .A(n2566), .Y(n5000) );
  CLKBUFX2TS U5115 ( .A(n2566), .Y(n4999) );
  CLKBUFX2TS U5116 ( .A(n4938), .Y(n4937) );
  CLKBUFX2TS U5117 ( .A(n4938), .Y(n4936) );
  CLKBUFX2TS U5118 ( .A(n4999), .Y(n4998) );
  CLKBUFX2TS U5119 ( .A(n4939), .Y(n4935) );
  CLKBUFX2TS U5120 ( .A(n4939), .Y(n4934) );
  CLKBUFX2TS U5121 ( .A(n5001), .Y(n4992) );
  CLKBUFX2TS U5122 ( .A(n2566), .Y(n5001) );
  CLKBUFX2TS U5123 ( .A(n2976), .Y(n4814) );
  INVX2TS U5124 ( .A(n1737), .Y(n5428) );
  CLKBUFX2TS U5125 ( .A(n4876), .Y(n4869) );
  CLKBUFX2TS U5126 ( .A(n5124), .Y(n5117) );
  CLKBUFX2TS U5127 ( .A(n4876), .Y(n4870) );
  CLKBUFX2TS U5128 ( .A(n5124), .Y(n5118) );
  CLKBUFX2TS U5129 ( .A(n5123), .Y(n5119) );
  CLKBUFX2TS U5130 ( .A(n4874), .Y(n4871) );
  CLKBUFX2TS U5131 ( .A(n4874), .Y(n4872) );
  CLKBUFX2TS U5132 ( .A(n5122), .Y(n5120) );
  CLKBUFX2TS U5133 ( .A(n4875), .Y(n4873) );
  CLKBUFX2TS U5134 ( .A(n5123), .Y(n5121) );
  CLKBUFX2TS U5135 ( .A(n5062), .Y(n5055) );
  CLKBUFX2TS U5136 ( .A(n5061), .Y(n5056) );
  CLKBUFX2TS U5137 ( .A(n5061), .Y(n5057) );
  CLKBUFX2TS U5138 ( .A(n5060), .Y(n5058) );
  CLKBUFX2TS U5139 ( .A(n5060), .Y(n5059) );
  CLKBUFX2TS U5140 ( .A(n4971), .Y(n4962) );
  CLKBUFX2TS U5141 ( .A(n5095), .Y(n5086) );
  CLKBUFX2TS U5142 ( .A(n4846), .Y(n4838) );
  CLKBUFX2TS U5143 ( .A(n4971), .Y(n4963) );
  CLKBUFX2TS U5144 ( .A(n5095), .Y(n5087) );
  CLKBUFX2TS U5145 ( .A(n4847), .Y(n4839) );
  CLKBUFX2TS U5146 ( .A(n4970), .Y(n4964) );
  CLKBUFX2TS U5147 ( .A(n4847), .Y(n4840) );
  CLKBUFX2TS U5148 ( .A(n4970), .Y(n4965) );
  CLKBUFX2TS U5149 ( .A(n4846), .Y(n4841) );
  CLKBUFX2TS U5150 ( .A(n5093), .Y(n5088) );
  CLKBUFX2TS U5151 ( .A(n4846), .Y(n4842) );
  CLKBUFX2TS U5152 ( .A(n4971), .Y(n4966) );
  CLKBUFX2TS U5153 ( .A(n5093), .Y(n5089) );
  CLKBUFX2TS U5154 ( .A(n4845), .Y(n4843) );
  CLKBUFX2TS U5155 ( .A(n4969), .Y(n4967) );
  CLKBUFX2TS U5156 ( .A(n5092), .Y(n5090) );
  CLKBUFX2TS U5157 ( .A(n4845), .Y(n4844) );
  CLKBUFX2TS U5158 ( .A(n4969), .Y(n4968) );
  CLKBUFX2TS U5159 ( .A(n5092), .Y(n5091) );
  CLKBUFX2TS U5160 ( .A(n2976), .Y(n4815) );
  CLKBUFX2TS U5161 ( .A(n2710), .Y(n4897) );
  CLKBUFX2TS U5162 ( .A(n5306), .Y(n5297) );
  CLKBUFX2TS U5163 ( .A(n5213), .Y(n5203) );
  CLKBUFX2TS U5164 ( .A(n5382), .Y(n5375) );
  CLKBUFX2TS U5165 ( .A(n5212), .Y(n5204) );
  CLKBUFX2TS U5166 ( .A(n5384), .Y(n5376) );
  CLKBUFX2TS U5167 ( .A(n5212), .Y(n5205) );
  CLKBUFX2TS U5168 ( .A(n5384), .Y(n5377) );
  CLKBUFX2TS U5169 ( .A(n5211), .Y(n5206) );
  CLKBUFX2TS U5170 ( .A(n5303), .Y(n5298) );
  CLKBUFX2TS U5171 ( .A(n5383), .Y(n5378) );
  CLKBUFX2TS U5172 ( .A(n5211), .Y(n5207) );
  CLKBUFX2TS U5173 ( .A(n5303), .Y(n5299) );
  CLKBUFX2TS U5174 ( .A(n5383), .Y(n5379) );
  CLKBUFX2TS U5175 ( .A(n5210), .Y(n5208) );
  CLKBUFX2TS U5176 ( .A(n5302), .Y(n5300) );
  CLKBUFX2TS U5177 ( .A(n5382), .Y(n5380) );
  CLKBUFX2TS U5178 ( .A(n5210), .Y(n5209) );
  CLKBUFX2TS U5179 ( .A(n5302), .Y(n5301) );
  CLKBUFX2TS U5180 ( .A(n5382), .Y(n5381) );
  CLKBUFX2TS U5181 ( .A(n1876), .Y(n5343) );
  CLKBUFX2TS U5182 ( .A(n4857), .Y(n4848) );
  CLKBUFX2TS U5183 ( .A(n4981), .Y(n4972) );
  CLKBUFX2TS U5184 ( .A(n5105), .Y(n5096) );
  CLKBUFX2TS U5185 ( .A(n4857), .Y(n4849) );
  CLKBUFX2TS U5186 ( .A(n4981), .Y(n4973) );
  CLKBUFX2TS U5187 ( .A(n5105), .Y(n5097) );
  CLKBUFX2TS U5188 ( .A(n4980), .Y(n4974) );
  CLKBUFX2TS U5189 ( .A(n4980), .Y(n4975) );
  CLKBUFX2TS U5190 ( .A(n4855), .Y(n4850) );
  CLKBUFX2TS U5191 ( .A(n4979), .Y(n4976) );
  CLKBUFX2TS U5192 ( .A(n5103), .Y(n5098) );
  CLKBUFX2TS U5193 ( .A(n4855), .Y(n4851) );
  CLKBUFX2TS U5194 ( .A(n5103), .Y(n5099) );
  CLKBUFX2TS U5195 ( .A(n4854), .Y(n4852) );
  CLKBUFX2TS U5196 ( .A(n4981), .Y(n4977) );
  CLKBUFX2TS U5197 ( .A(n5102), .Y(n5100) );
  CLKBUFX2TS U5198 ( .A(n4854), .Y(n4853) );
  CLKBUFX2TS U5199 ( .A(n4980), .Y(n4978) );
  CLKBUFX2TS U5200 ( .A(n5102), .Y(n5101) );
  INVX2TS U5201 ( .A(N6620), .Y(n5775) );
  NAND2BX1TS U5202 ( .AN(n2126), .B(n5409), .Y(n1621) );
  NAND2X1TS U5203 ( .A(n1588), .B(n5719), .Y(n1590) );
  CLKBUFX2TS U5204 ( .A(n5149), .Y(n5142) );
  CLKBUFX2TS U5205 ( .A(n5149), .Y(n5141) );
  CLKBUFX2TS U5206 ( .A(n5149), .Y(n5140) );
  CLKBUFX2TS U5207 ( .A(n5150), .Y(n5139) );
  CLKBUFX2TS U5208 ( .A(n5150), .Y(n5138) );
  CLKBUFX2TS U5209 ( .A(n5150), .Y(n5137) );
  CLKBUFX2TS U5210 ( .A(n5150), .Y(n5136) );
  CLKBUFX2TS U5211 ( .A(n4961), .Y(n4949) );
  CLKBUFX2TS U5212 ( .A(n2574), .Y(n4961) );
  CLKBUFX2TS U5213 ( .A(n2295), .Y(n5085) );
  CLKBUFX2TS U5214 ( .A(n4899), .Y(n4887) );
  CLKBUFX2TS U5215 ( .A(n2710), .Y(n4899) );
  CLKBUFX2TS U5216 ( .A(n2848), .Y(n4837) );
  CLKBUFX2TS U5217 ( .A(n5148), .Y(n5147) );
  CLKBUFX2TS U5218 ( .A(n5148), .Y(n5146) );
  CLKBUFX2TS U5219 ( .A(n5148), .Y(n5145) );
  CLKBUFX2TS U5220 ( .A(n5148), .Y(n5144) );
  CLKBUFX2TS U5221 ( .A(n5149), .Y(n5143) );
  CLKBUFX2TS U5222 ( .A(n2436), .Y(n5002) );
  CLKBUFX2TS U5223 ( .A(n2981), .Y(n4795) );
  CLKBUFX2TS U5224 ( .A(n2981), .Y(n4794) );
  CLKBUFX2TS U5225 ( .A(n2981), .Y(n4793) );
  CLKBUFX2TS U5226 ( .A(n3114), .Y(n4763) );
  CLKBUFX2TS U5227 ( .A(n2983), .Y(n4785) );
  CLKBUFX2TS U5228 ( .A(n2051), .Y(n5162) );
  CLKBUFX2TS U5229 ( .A(n4909), .Y(n4900) );
  CLKBUFX2TS U5230 ( .A(n4909), .Y(n4901) );
  CLKBUFX2TS U5231 ( .A(n4909), .Y(n4902) );
  CLKBUFX2TS U5232 ( .A(n4908), .Y(n4903) );
  CLKBUFX2TS U5233 ( .A(n4908), .Y(n4904) );
  CLKBUFX2TS U5234 ( .A(n4907), .Y(n4905) );
  CLKBUFX2TS U5235 ( .A(n4907), .Y(n4906) );
  CLKBUFX2TS U5236 ( .A(n2434), .Y(n5024) );
  CLKBUFX2TS U5237 ( .A(n5033), .Y(n5025) );
  CLKBUFX2TS U5238 ( .A(n5033), .Y(n5026) );
  CLKBUFX2TS U5239 ( .A(n5033), .Y(n5027) );
  CLKBUFX2TS U5240 ( .A(n5032), .Y(n5028) );
  CLKBUFX2TS U5241 ( .A(n5032), .Y(n5029) );
  CLKBUFX2TS U5242 ( .A(n5031), .Y(n5030) );
  CLKBUFX2TS U5243 ( .A(n3114), .Y(n4764) );
  CLKBUFX2TS U5244 ( .A(n1666), .Y(n5490) );
  CLKBUFX2TS U5245 ( .A(n2051), .Y(n5163) );
  CLKBUFX2TS U5246 ( .A(n2574), .Y(n4960) );
  CLKBUFX2TS U5247 ( .A(n2295), .Y(n5084) );
  CLKBUFX2TS U5248 ( .A(n2574), .Y(n4959) );
  CLKBUFX2TS U5249 ( .A(n2295), .Y(n5083) );
  CLKBUFX2TS U5250 ( .A(n2848), .Y(n4836) );
  CLKBUFX2TS U5251 ( .A(n2848), .Y(n4835) );
  CLKBUFX2TS U5252 ( .A(n2710), .Y(n4898) );
  CLKBUFX2TS U5253 ( .A(n2710), .Y(n4896) );
  CLKBUFX2TS U5254 ( .A(n5202), .Y(n5201) );
  CLKBUFX2TS U5255 ( .A(n5280), .Y(n5278) );
  CLKBUFX2TS U5256 ( .A(n5374), .Y(n5372) );
  CLKBUFX2TS U5257 ( .A(n5188), .Y(n5200) );
  CLKBUFX2TS U5258 ( .A(n5264), .Y(n5277) );
  CLKBUFX2TS U5259 ( .A(n5358), .Y(n5371) );
  CLKBUFX2TS U5260 ( .A(n5241), .Y(n5240) );
  CLKBUFX2TS U5261 ( .A(n5226), .Y(n5239) );
  CLKBUFX2TS U5262 ( .A(n5227), .Y(n5238) );
  CLKBUFX2TS U5263 ( .A(n5335), .Y(n5334) );
  CLKBUFX2TS U5264 ( .A(n5320), .Y(n5333) );
  CLKBUFX2TS U5265 ( .A(n5321), .Y(n5332) );
  INVX2TS U5266 ( .A(n2200), .Y(n5771) );
  CLKBUFX2TS U5267 ( .A(n5171), .Y(n5169) );
  CLKBUFX2TS U5268 ( .A(n5171), .Y(n5170) );
  CLKBUFX2TS U5269 ( .A(n5174), .Y(n5164) );
  CLKBUFX2TS U5270 ( .A(n5173), .Y(n5165) );
  CLKBUFX2TS U5271 ( .A(n5173), .Y(n5166) );
  CLKBUFX2TS U5272 ( .A(n5172), .Y(n5167) );
  CLKBUFX2TS U5273 ( .A(n5172), .Y(n5168) );
  CLKBUFX2TS U5274 ( .A(n5251), .Y(n5242) );
  CLKBUFX2TS U5275 ( .A(n5251), .Y(n5243) );
  CLKBUFX2TS U5276 ( .A(n5250), .Y(n5244) );
  CLKBUFX2TS U5277 ( .A(n5250), .Y(n5245) );
  CLKBUFX2TS U5278 ( .A(n5249), .Y(n5246) );
  CLKBUFX2TS U5279 ( .A(n5249), .Y(n5247) );
  CLKBUFX2TS U5280 ( .A(n5253), .Y(n5248) );
  CLKBUFX2TS U5281 ( .A(n5346), .Y(n5336) );
  CLKBUFX2TS U5282 ( .A(n5346), .Y(n5337) );
  CLKBUFX2TS U5283 ( .A(n1876), .Y(n5338) );
  CLKBUFX2TS U5284 ( .A(n5345), .Y(n5339) );
  CLKBUFX2TS U5285 ( .A(n5345), .Y(n5340) );
  CLKBUFX2TS U5286 ( .A(n5344), .Y(n5341) );
  CLKBUFX2TS U5287 ( .A(n5344), .Y(n5342) );
  CLKBUFX2TS U5288 ( .A(n4919), .Y(n4910) );
  CLKBUFX2TS U5289 ( .A(n4919), .Y(n4911) );
  CLKBUFX2TS U5290 ( .A(n4918), .Y(n4912) );
  CLKBUFX2TS U5291 ( .A(n4918), .Y(n4913) );
  CLKBUFX2TS U5292 ( .A(n4917), .Y(n4914) );
  CLKBUFX2TS U5293 ( .A(n4917), .Y(n4915) );
  CLKBUFX2TS U5294 ( .A(n4917), .Y(n4916) );
  CLKBUFX2TS U5295 ( .A(n5043), .Y(n5034) );
  CLKBUFX2TS U5296 ( .A(n5043), .Y(n5035) );
  CLKBUFX2TS U5297 ( .A(n5042), .Y(n5036) );
  CLKBUFX2TS U5298 ( .A(n5042), .Y(n5037) );
  CLKBUFX2TS U5299 ( .A(n5041), .Y(n5038) );
  CLKBUFX2TS U5300 ( .A(n5043), .Y(n5039) );
  CLKBUFX2TS U5301 ( .A(n5042), .Y(n5040) );
  NAND2X1TS U5302 ( .A(n4582), .B(n5592), .Y(n1616) );
  NAND2X1TS U5303 ( .A(n5797), .B(n5592), .Y(n1586) );
  NAND2X1TS U5304 ( .A(n1821), .B(n4562), .Y(n1663) );
  CLKBUFX2TS U5305 ( .A(n5613), .Y(n5612) );
  CLKBUFX2TS U5306 ( .A(n5613), .Y(n5611) );
  CLKBUFX2TS U5307 ( .A(n5614), .Y(n5610) );
  CLKBUFX2TS U5308 ( .A(n5614), .Y(n5609) );
  CLKBUFX2TS U5309 ( .A(n5614), .Y(n5608) );
  CLKBUFX2TS U5310 ( .A(n5439), .Y(n5438) );
  CLKBUFX2TS U5311 ( .A(n1645), .Y(n5512) );
  CLKBUFX2TS U5312 ( .A(n1645), .Y(n5513) );
  CLKBUFX2TS U5313 ( .A(n5440), .Y(n5436) );
  CLKBUFX2TS U5314 ( .A(n5440), .Y(n5437) );
  CLKBUFX2TS U5315 ( .A(n5514), .Y(n5511) );
  CLKBUFX2TS U5316 ( .A(n1643), .Y(n5525) );
  CLKBUFX2TS U5317 ( .A(n1667), .Y(n5477) );
  CLKBUFX2TS U5318 ( .A(n4710), .Y(n4706) );
  CLKBUFX2TS U5319 ( .A(n4710), .Y(n4707) );
  CLKBUFX2TS U5320 ( .A(n4709), .Y(n4708) );
  CLKBUFX2TS U5321 ( .A(n1643), .Y(n5526) );
  CLKBUFX2TS U5322 ( .A(n1667), .Y(n5478) );
  INVX2TS U5323 ( .A(n1661), .Y(n5798) );
  INVX2TS U5324 ( .A(n4545), .Y(n5803) );
  NOR2X1TS U5325 ( .A(n5559), .B(n3876), .Y(N10004) );
  CLKBUFX2TS U5326 ( .A(n5555), .Y(n5541) );
  CLKBUFX2TS U5327 ( .A(n5555), .Y(n5542) );
  CLKBUFX2TS U5328 ( .A(n5554), .Y(n5546) );
  CLKBUFX2TS U5329 ( .A(n5554), .Y(n5545) );
  CLKBUFX2TS U5330 ( .A(n5555), .Y(n5544) );
  CLKBUFX2TS U5331 ( .A(n5555), .Y(n5543) );
  CLKBUFX2TS U5332 ( .A(n5554), .Y(n5547) );
  CLKBUFX2TS U5333 ( .A(n5554), .Y(n5548) );
  INVX2TS U5334 ( .A(n5745), .Y(n5721) );
  INVX2TS U5335 ( .A(n5733), .Y(n5719) );
  CLKBUFX2TS U5336 ( .A(n4719), .Y(n4718) );
  CLKBUFX2TS U5337 ( .A(n4720), .Y(n4717) );
  CLKBUFX2TS U5338 ( .A(n4720), .Y(n4716) );
  CLKBUFX2TS U5339 ( .A(n4721), .Y(n4715) );
  OAI21X1TS U5340 ( .A0(n5793), .A1(n5593), .B0(n3754), .Y(n2127) );
  INVX2TS U5341 ( .A(n5743), .Y(n5718) );
  INVX2TS U5342 ( .A(n5732), .Y(n5722) );
  INVX2TS U5343 ( .A(n5729), .Y(n5720) );
  INVX2TS U5344 ( .A(n5731), .Y(n5723) );
  INVX2TS U5345 ( .A(n5730), .Y(n5724) );
  INVX2TS U5346 ( .A(n5733), .Y(n5727) );
  INVX2TS U5347 ( .A(n5728), .Y(n5726) );
  NAND2X1TS U5348 ( .A(n5559), .B(n4663), .Y(n1788) );
  NAND2X1TS U5349 ( .A(n5560), .B(n4677), .Y(n1745) );
  INVX2TS U5350 ( .A(n1565), .Y(n5559) );
  INVX2TS U5351 ( .A(n5601), .Y(n5560) );
  INVX2TS U5352 ( .A(n1565), .Y(n5561) );
  NAND2X1TS U5353 ( .A(n5281), .B(n5561), .Y(n1767) );
  NAND2X1TS U5354 ( .A(n5559), .B(n4691), .Y(n1757) );
  CLKBUFX2TS U5355 ( .A(n5596), .Y(n5591) );
  CLKBUFX2TS U5356 ( .A(n5596), .Y(n5592) );
  CLKBUFX2TS U5357 ( .A(n4698), .Y(n4697) );
  CLKBUFX2TS U5358 ( .A(n4671), .Y(n4670) );
  CLKBUFX2TS U5359 ( .A(n5414), .Y(n5412) );
  CLKBUFX2TS U5360 ( .A(n4688), .Y(n4678) );
  CLKBUFX2TS U5361 ( .A(n4675), .Y(n4664) );
  CLKBUFX2TS U5362 ( .A(n4671), .Y(n4669) );
  CLKBUFX2TS U5363 ( .A(n4672), .Y(n4668) );
  CLKBUFX2TS U5364 ( .A(n4672), .Y(n4667) );
  CLKBUFX2TS U5365 ( .A(n4673), .Y(n4666) );
  CLKBUFX2TS U5366 ( .A(n4673), .Y(n4665) );
  CLKBUFX2TS U5367 ( .A(n4698), .Y(n4696) );
  CLKBUFX2TS U5368 ( .A(n4699), .Y(n4695) );
  CLKBUFX2TS U5369 ( .A(n4699), .Y(n4694) );
  CLKBUFX2TS U5370 ( .A(n4700), .Y(n4693) );
  CLKBUFX2TS U5371 ( .A(n4700), .Y(n4692) );
  CLKBUFX2TS U5372 ( .A(n4688), .Y(n4679) );
  CLKBUFX2TS U5373 ( .A(n4686), .Y(n4685) );
  CLKBUFX2TS U5374 ( .A(n4686), .Y(n4684) );
  CLKBUFX2TS U5375 ( .A(n4687), .Y(n4683) );
  CLKBUFX2TS U5376 ( .A(n4687), .Y(n4682) );
  CLKBUFX2TS U5377 ( .A(n4687), .Y(n4681) );
  CLKBUFX2TS U5378 ( .A(n4686), .Y(n4680) );
  INVX2TS U5379 ( .A(n5412), .Y(n5400) );
  INVX2TS U5380 ( .A(n5414), .Y(n5399) );
  INVX2TS U5381 ( .A(n5414), .Y(n5401) );
  INVX2TS U5382 ( .A(n5293), .Y(n5285) );
  INVX2TS U5383 ( .A(n5293), .Y(n5284) );
  INVX2TS U5384 ( .A(n5294), .Y(n5288) );
  INVX2TS U5385 ( .A(n5294), .Y(n5287) );
  INVX2TS U5386 ( .A(n5294), .Y(n5286) );
  INVX2TS U5387 ( .A(n5295), .Y(n5290) );
  INVX2TS U5388 ( .A(n5295), .Y(n5289) );
  INVX2TS U5389 ( .A(n5293), .Y(n5291) );
  INVX2TS U5390 ( .A(n5729), .Y(n5725) );
  NAND4X1TS U5391 ( .A(N6373), .B(n2427), .C(n3718), .D(n5777), .Y(n2574) );
  NAND4X1TS U5392 ( .A(N6373), .B(N6372), .C(n2427), .D(n3719), .Y(n2295) );
  NAND3XLTS U5393 ( .A(N6373), .B(n4598), .C(n2565), .Y(n2436) );
  AOI211X1TS U5394 ( .A0(n1957), .A1(n5584), .B0(n5731), .C0(n5750), .Y(n1956)
         );
  INVX2TS U5395 ( .A(n1765), .Y(n5750) );
  NAND2BX1TS U5396 ( .AN(n1958), .B(n3829), .Y(n1957) );
  NOR2BX1TS U5397 ( .AN(n2282), .B(n5799), .Y(n2199) );
  CLKINVX1TS U5398 ( .A(N6372), .Y(n5777) );
  NOR2X1TS U5399 ( .A(n5777), .B(n5795), .Y(n2839) );
  NAND3X1TS U5400 ( .A(n2426), .B(n5773), .C(\add_0_root_r1463/SUM[2] ), .Y(
        n1955) );
  NAND3X1TS U5401 ( .A(n2285), .B(n5773), .C(n3701), .Y(n1910) );
  NAND3X1TS U5402 ( .A(n4597), .B(n5774), .C(n2565), .Y(n2983) );
  NAND3X1TS U5403 ( .A(n5772), .B(n5773), .C(n2285), .Y(n2085) );
  NAND2X1TS U5404 ( .A(n2199), .B(n1736), .Y(n1737) );
  OAI31X1TS U5405 ( .A0(n3111), .A1(n5411), .A2(n2088), .B0(n5585), .Y(n3109)
         );
  NAND2X1TS U5406 ( .A(n4774), .B(n3108), .Y(n3111) );
  NOR2X1TS U5407 ( .A(\add_0_root_r1463/SUM[3] ), .B(\add_0_root_r1463/SUM[4] ), .Y(n3113) );
  AND3X2TS U5408 ( .A(n2283), .B(n5759), .C(n3699), .Y(n2563) );
  AND3X2TS U5409 ( .A(n2283), .B(n5758), .C(n5759), .Y(n3110) );
  AND3X2TS U5410 ( .A(n1786), .B(n5724), .C(n4670), .Y(n2045) );
  AND3X2TS U5411 ( .A(n1743), .B(n5724), .C(n4690), .Y(n1868) );
  AND3X2TS U5412 ( .A(n1775), .B(n5723), .C(n5690), .Y(n2001) );
  AND3X2TS U5413 ( .A(n1755), .B(n5724), .C(n4697), .Y(n1912) );
  OAI21X1TS U5414 ( .A0(n3812), .A1(n1913), .B0(n5568), .Y(n1911) );
  AND2X2TS U5415 ( .A(n2281), .B(n5599), .Y(n3117) );
  INVX2TS U5416 ( .A(\add_0_root_r1459/SUM[2] ), .Y(n5758) );
  INVX2TS U5417 ( .A(n3710), .Y(n5762) );
  CLKBUFX2TS U5418 ( .A(n2843), .Y(n4857) );
  CLKBUFX2TS U5419 ( .A(n2569), .Y(n4981) );
  CLKBUFX2TS U5420 ( .A(n2290), .Y(n5105) );
  CLKBUFX2TS U5421 ( .A(n2843), .Y(n4856) );
  CLKBUFX2TS U5422 ( .A(n2569), .Y(n4980) );
  CLKBUFX2TS U5423 ( .A(n2290), .Y(n5104) );
  CLKBUFX2TS U5424 ( .A(n2843), .Y(n4855) );
  CLKBUFX2TS U5425 ( .A(n2569), .Y(n4979) );
  CLKBUFX2TS U5426 ( .A(n2290), .Y(n5103) );
  CLKBUFX2TS U5427 ( .A(n2843), .Y(n4854) );
  CLKBUFX2TS U5428 ( .A(n2290), .Y(n5102) );
  CLKBUFX2TS U5429 ( .A(n2572), .Y(n4971) );
  CLKBUFX2TS U5430 ( .A(n2293), .Y(n5095) );
  CLKBUFX2TS U5431 ( .A(n2846), .Y(n4847) );
  CLKBUFX2TS U5432 ( .A(n2572), .Y(n4970) );
  CLKBUFX2TS U5433 ( .A(n2293), .Y(n5094) );
  CLKBUFX2TS U5434 ( .A(n2846), .Y(n4846) );
  CLKBUFX2TS U5435 ( .A(n2293), .Y(n5093) );
  CLKBUFX2TS U5436 ( .A(n2846), .Y(n4845) );
  CLKBUFX2TS U5437 ( .A(n2572), .Y(n4969) );
  CLKBUFX2TS U5438 ( .A(n2293), .Y(n5092) );
  CLKBUFX2TS U5439 ( .A(n5307), .Y(n5306) );
  CLKBUFX2TS U5440 ( .A(n5307), .Y(n5305) );
  CLKBUFX2TS U5441 ( .A(n5213), .Y(n5212) );
  CLKBUFX2TS U5442 ( .A(n5307), .Y(n5304) );
  CLKBUFX2TS U5443 ( .A(n5385), .Y(n5384) );
  CLKBUFX2TS U5444 ( .A(n2840), .Y(n4876) );
  CLKBUFX2TS U5445 ( .A(n2287), .Y(n5124) );
  CLKBUFX2TS U5446 ( .A(n2840), .Y(n4875) );
  CLKBUFX2TS U5447 ( .A(n2287), .Y(n5123) );
  CLKBUFX2TS U5448 ( .A(n5063), .Y(n5062) );
  CLKBUFX2TS U5449 ( .A(n5063), .Y(n5061) );
  CLKBUFX2TS U5450 ( .A(n5214), .Y(n5210) );
  CLKBUFX2TS U5451 ( .A(n5308), .Y(n5302) );
  CLKBUFX2TS U5452 ( .A(n5386), .Y(n5382) );
  CLKBUFX2TS U5453 ( .A(n5214), .Y(n5211) );
  CLKBUFX2TS U5454 ( .A(n5308), .Y(n5303) );
  CLKBUFX2TS U5455 ( .A(n5386), .Y(n5383) );
  CLKBUFX2TS U5456 ( .A(n4875), .Y(n4874) );
  CLKBUFX2TS U5457 ( .A(n5123), .Y(n5122) );
  CLKBUFX2TS U5458 ( .A(n5063), .Y(n5060) );
  CLKBUFX2TS U5459 ( .A(n4877), .Y(n4868) );
  CLKBUFX2TS U5460 ( .A(n5125), .Y(n5116) );
  CLKBUFX2TS U5461 ( .A(n2287), .Y(n5125) );
  INVX2TS U5462 ( .A(n2012), .Y(n5202) );
  INVX2TS U5463 ( .A(n1924), .Y(n5280) );
  INVX2TS U5464 ( .A(n1834), .Y(n5374) );
  INVX2TS U5465 ( .A(n1968), .Y(n5241) );
  INVX2TS U5466 ( .A(n1879), .Y(n5335) );
  CLKBUFX2TS U5467 ( .A(n2702), .Y(n4939) );
  INVX2TS U5468 ( .A(n5412), .Y(n5410) );
  AOI211X1TS U5469 ( .A0(n2087), .A1(n5584), .B0(n5728), .C0(n5754), .Y(n2086)
         );
  NAND2BX1TS U5470 ( .AN(n2088), .B(n3823), .Y(n2087) );
  CLKBUFX2TS U5471 ( .A(n2054), .Y(n5151) );
  NOR3BX1TS U5472 ( .AN(n1959), .B(N6619), .C(n5796), .Y(n1914) );
  NAND3X1TS U5473 ( .A(n3725), .B(n1598), .C(N10004), .Y(n1588) );
  NOR2X1TS U5474 ( .A(N6375), .B(N6374), .Y(n2838) );
  AND2X2TS U5475 ( .A(n2838), .B(n5795), .Y(n2427) );
  NOR2X1TS U5476 ( .A(n2282), .B(n4550), .Y(n2200) );
  OAI21X1TS U5477 ( .A0(n4567), .A1(n2114), .B0(n1598), .Y(n2106) );
  NOR2X1TS U5478 ( .A(N6622), .B(N6621), .Y(n1959) );
  NAND4X1TS U5479 ( .A(n5591), .B(n3725), .C(n4519), .D(n5718), .Y(n3114) );
  INVX2TS U5480 ( .A(\add_0_root_r1463/SUM[2] ), .Y(n5772) );
  AND3XLTS U5481 ( .A(n1959), .B(n5796), .C(N6620), .Y(n1870) );
  NAND2X1TS U5482 ( .A(n5591), .B(n5804), .Y(n2205) );
  OR2X2TS U5483 ( .A(n5804), .B(n5560), .Y(n4610) );
  INVX2TS U5484 ( .A(n4610), .Y(n2090) );
  NAND3BXLTS U5485 ( .AN(N6619), .B(n1870), .C(n3719), .Y(n1926) );
  AND2X2TS U5486 ( .A(n1822), .B(n3704), .Y(n1821) );
  CLKBUFX2TS U5487 ( .A(n2705), .Y(n4919) );
  CLKBUFX2TS U5488 ( .A(n2705), .Y(n4918) );
  CLKBUFX2TS U5489 ( .A(n2705), .Y(n4917) );
  CLKBUFX2TS U5490 ( .A(n2431), .Y(n5043) );
  CLKBUFX2TS U5491 ( .A(n2431), .Y(n5042) );
  CLKBUFX2TS U5492 ( .A(n2431), .Y(n5041) );
  CLKBUFX2TS U5493 ( .A(n2708), .Y(n4909) );
  CLKBUFX2TS U5494 ( .A(n2708), .Y(n4908) );
  CLKBUFX2TS U5495 ( .A(n2708), .Y(n4907) );
  CLKBUFX2TS U5496 ( .A(n2434), .Y(n5033) );
  CLKBUFX2TS U5497 ( .A(n2434), .Y(n5032) );
  CLKBUFX2TS U5498 ( .A(n2434), .Y(n5031) );
  CLKBUFX2TS U5499 ( .A(n5174), .Y(n5173) );
  CLKBUFX2TS U5500 ( .A(n5252), .Y(n5251) );
  CLKBUFX2TS U5501 ( .A(n5252), .Y(n5250) );
  CLKBUFX2TS U5502 ( .A(n5252), .Y(n5249) );
  CLKBUFX2TS U5503 ( .A(n5347), .Y(n5346) );
  CLKBUFX2TS U5504 ( .A(n5347), .Y(n5345) );
  CLKBUFX2TS U5505 ( .A(n5175), .Y(n5171) );
  CLKBUFX2TS U5506 ( .A(n5175), .Y(n5172) );
  CLKBUFX2TS U5507 ( .A(n1876), .Y(n5344) );
  CLKBUFX2TS U5508 ( .A(n1563), .Y(n5613) );
  CLKBUFX2TS U5509 ( .A(n2054), .Y(n5148) );
  CLKBUFX2TS U5510 ( .A(n2054), .Y(n5149) );
  CLKBUFX2TS U5511 ( .A(n2054), .Y(n5150) );
  INVX2TS U5512 ( .A(n2132), .Y(n5754) );
  NOR2X1TS U5513 ( .A(n5805), .B(n1616), .Y(n1604) );
  NOR2BX1TS U5514 ( .AN(n4566), .B(n4544), .Y(n1865) );
  AND3XLTS U5515 ( .A(n1959), .B(n5775), .C(N6619), .Y(n2003) );
  NOR2X1TS U5516 ( .A(n5799), .B(n5802), .Y(n1667) );
  NAND2X1TS U5517 ( .A(n1794), .B(n5721), .Y(n1661) );
  NAND2X1TS U5518 ( .A(n2197), .B(n5805), .Y(n1643) );
  CLKBUFX2TS U5519 ( .A(n4713), .Y(n4711) );
  CLKBUFX2TS U5520 ( .A(n4714), .Y(n4710) );
  CLKBUFX2TS U5521 ( .A(n4714), .Y(n4709) );
  CLKBUFX2TS U5522 ( .A(n1669), .Y(n5439) );
  CLKBUFX2TS U5523 ( .A(n1563), .Y(n5614) );
  INVX2TS U5524 ( .A(n1733), .Y(n5797) );
  CLKBUFX2TS U5525 ( .A(n5665), .Y(n5656) );
  CLKBUFX2TS U5526 ( .A(n4712), .Y(n4705) );
  CLKBUFX2TS U5527 ( .A(n4713), .Y(n4712) );
  CLKBUFX2TS U5528 ( .A(n5662), .Y(n5657) );
  CLKBUFX2TS U5529 ( .A(n5662), .Y(n5658) );
  CLKBUFX2TS U5530 ( .A(n1548), .Y(n5630) );
  CLKBUFX2TS U5531 ( .A(n5640), .Y(n5631) );
  CLKBUFX2TS U5532 ( .A(n5640), .Y(n5632) );
  CLKBUFX2TS U5533 ( .A(n5639), .Y(n5633) );
  CLKBUFX2TS U5534 ( .A(n5639), .Y(n5634) );
  CLKBUFX2TS U5535 ( .A(n5638), .Y(n5635) );
  CLKBUFX2TS U5536 ( .A(n5638), .Y(n5636) );
  CLKBUFX2TS U5537 ( .A(n5661), .Y(n5659) );
  CLKBUFX2TS U5538 ( .A(n1669), .Y(n5440) );
  CLKBUFX2TS U5539 ( .A(n1645), .Y(n5514) );
  AND2X2TS U5540 ( .A(n3725), .B(n4538), .Y(n1802) );
  INVX2TS U5541 ( .A(n1744), .Y(n5790) );
  INVX2TS U5542 ( .A(n1766), .Y(n5789) );
  INVX2TS U5543 ( .A(n1799), .Y(n5786) );
  CLKBUFX2TS U5544 ( .A(n5744), .Y(n5728) );
  CLKBUFX2TS U5545 ( .A(n5744), .Y(n5733) );
  CLKBUFX2TS U5546 ( .A(n5556), .Y(n5540) );
  CLKBUFX2TS U5547 ( .A(n5557), .Y(n5556) );
  CLKBUFX2TS U5548 ( .A(n5741), .Y(n5739) );
  INVX2TS U5549 ( .A(n1756), .Y(n5787) );
  CLKBUFX2TS U5550 ( .A(n5553), .Y(n5549) );
  CLKBUFX2TS U5551 ( .A(n5553), .Y(n5550) );
  CLKBUFX2TS U5552 ( .A(n5553), .Y(n5551) );
  CLKBUFX2TS U5553 ( .A(n5741), .Y(n5740) );
  CLKBUFX2TS U5554 ( .A(n5553), .Y(n5552) );
  INVX2TS U5555 ( .A(n1787), .Y(n5788) );
  CLKBUFX2TS U5556 ( .A(n4723), .Y(n4721) );
  CLKBUFX2TS U5557 ( .A(n4723), .Y(n4722) );
  CLKBUFX2TS U5558 ( .A(n4724), .Y(n4719) );
  CLKBUFX2TS U5559 ( .A(n4724), .Y(n4720) );
  CLKBUFX2TS U5560 ( .A(n3157), .Y(n4726) );
  CLKBUFX2TS U5561 ( .A(n3157), .Y(n4727) );
  CLKBUFX2TS U5562 ( .A(n4732), .Y(n4728) );
  CLKBUFX2TS U5563 ( .A(n4732), .Y(n4729) );
  CLKBUFX2TS U5564 ( .A(n4731), .Y(n4730) );
  INVX2TS U5565 ( .A(n5625), .Y(n5622) );
  INVX2TS U5566 ( .A(n5625), .Y(n5621) );
  INVX2TS U5567 ( .A(n5625), .Y(n5620) );
  INVX2TS U5568 ( .A(n5628), .Y(n5619) );
  INVX2TS U5569 ( .A(n5629), .Y(n5618) );
  INVX2TS U5570 ( .A(n5626), .Y(n5623) );
  INVX2TS U5571 ( .A(n5627), .Y(n5624) );
  INVX2TS U5572 ( .A(n5678), .Y(n5677) );
  INVX2TS U5573 ( .A(n5652), .Y(n5651) );
  CLKBUFX2TS U5574 ( .A(n5661), .Y(n5660) );
  CLKBUFX2TS U5575 ( .A(n5641), .Y(n5637) );
  CLKBUFX2TS U5576 ( .A(n5556), .Y(n5554) );
  CLKBUFX2TS U5577 ( .A(n5557), .Y(n5555) );
  CLKBUFX2TS U5578 ( .A(n5744), .Y(n5729) );
  CLKBUFX2TS U5579 ( .A(n5743), .Y(n5730) );
  CLKBUFX2TS U5580 ( .A(n5743), .Y(n5731) );
  CLKBUFX2TS U5581 ( .A(n5743), .Y(n5732) );
  NAND2X1TS U5582 ( .A(n2271), .B(n2272), .Y(n1641) );
  INVX2TS U5583 ( .A(n2130), .Y(n5907) );
  AOI21X1TS U5584 ( .A0(n5565), .A1(n2220), .B0(n2130), .Y(n2217) );
  AOI21X1TS U5585 ( .A0(n5565), .A1(n2208), .B0(n4539), .Y(n2203) );
  AOI21X1TS U5586 ( .A0(n5566), .A1(n2262), .B0(n4539), .Y(n2259) );
  AOI21X1TS U5587 ( .A0(n5566), .A1(n2233), .B0(n2130), .Y(n2232) );
  OAI2BB1X1TS U5588 ( .A0N(n2114), .A1N(n5570), .B0(n5907), .Y(n2107) );
  INVX2TS U5589 ( .A(n2112), .Y(n5783) );
  INVX2TS U5590 ( .A(\add_0_root_sub_0_root_sub_231/B[2] ), .Y(n5792) );
  INVX2TS U5591 ( .A(N6699), .Y(n5785) );
  CLKBUFX2TS U5592 ( .A(n5742), .Y(n5734) );
  CLKBUFX2TS U5593 ( .A(n5742), .Y(n5737) );
  CLKBUFX2TS U5594 ( .A(n5742), .Y(n5736) );
  CLKBUFX2TS U5595 ( .A(n5742), .Y(n5735) );
  CLKBUFX2TS U5596 ( .A(n5741), .Y(n5738) );
  INVX2TS U5597 ( .A(n1760), .Y(n5779) );
  INVX2TS U5598 ( .A(n1749), .Y(n5782) );
  INVX2TS U5599 ( .A(n1791), .Y(n5780) );
  INVX2TS U5600 ( .A(N8209), .Y(n5794) );
  CLKBUFX2TS U5601 ( .A(n4611), .Y(n5413) );
  INVX2TS U5602 ( .A(n2275), .Y(n5793) );
  CLKBUFX2TS U5603 ( .A(n4674), .Y(n4663) );
  CLKBUFX2TS U5604 ( .A(n4675), .Y(n4674) );
  CLKBUFX2TS U5605 ( .A(n4689), .Y(n4677) );
  CLKBUFX2TS U5606 ( .A(n4690), .Y(n4689) );
  CLKBUFX2TS U5607 ( .A(n4702), .Y(n4691) );
  CLKBUFX2TS U5608 ( .A(n4703), .Y(n4702) );
  INVX2TS U5609 ( .A(\add_0_root_sub_278_I2/B[2] ), .Y(n5776) );
  NAND2X1TS U5610 ( .A(n5560), .B(n5682), .Y(n1777) );
  CLKBUFX2TS U5611 ( .A(n5600), .Y(n5596) );
  CLKBUFX2TS U5612 ( .A(n5600), .Y(n5597) );
  CLKBUFX2TS U5613 ( .A(n5597), .Y(n5599) );
  CLKBUFX2TS U5614 ( .A(n5600), .Y(n5598) );
  CLKBUFX2TS U5615 ( .A(n4676), .Y(n4671) );
  CLKBUFX2TS U5616 ( .A(n4704), .Y(n4698) );
  INVX2TS U5617 ( .A(n5292), .Y(n5281) );
  CLKBUFX2TS U5618 ( .A(n5595), .Y(n5593) );
  CLKBUFX2TS U5619 ( .A(n4676), .Y(n4672) );
  CLKBUFX2TS U5620 ( .A(n4688), .Y(n4686) );
  CLKBUFX2TS U5621 ( .A(n4676), .Y(n4673) );
  CLKBUFX2TS U5622 ( .A(n5973), .Y(n4687) );
  CLKBUFX2TS U5623 ( .A(n4690), .Y(n4688) );
  CLKBUFX2TS U5624 ( .A(n4704), .Y(n4699) );
  CLKBUFX2TS U5625 ( .A(n4704), .Y(n4700) );
  CLKBUFX2TS U5626 ( .A(n4703), .Y(n4701) );
  CLKBUFX2TS U5627 ( .A(n4611), .Y(n5414) );
  INVX2TS U5628 ( .A(n5292), .Y(n5282) );
  INVX2TS U5629 ( .A(n5292), .Y(n5283) );
  CLKBUFX2TS U5630 ( .A(n5595), .Y(n5594) );
  NAND3X1TS U5631 ( .A(n2285), .B(n5772), .C(\add_0_root_r1463/SUM[1] ), .Y(
        n1999) );
  OAI31X1TS U5632 ( .A0(n2564), .A1(n5705), .A2(n5776), .B0(n5318), .Y(n1913)
         );
  INVX2TS U5633 ( .A(n5335), .Y(n5318) );
  NAND4X1TS U5634 ( .A(n3697), .B(\add_0_root_r1463/SUM[2] ), .C(n2285), .D(
        n2286), .Y(n2282) );
  AND3X2TS U5635 ( .A(n2838), .B(n5777), .C(N6371), .Y(n2565) );
  AND3X2TS U5636 ( .A(n2283), .B(n5758), .C(\add_0_root_r1459/SUM[1] ), .Y(
        n2837) );
  OR2X2TS U5637 ( .A(n2972), .B(n1788), .Y(n2846) );
  OR2X2TS U5638 ( .A(n2698), .B(n1767), .Y(n2572) );
  OR2X2TS U5639 ( .A(n2419), .B(n1745), .Y(n2293) );
  NAND2X1TS U5640 ( .A(n2280), .B(n2286), .Y(n2281) );
  INVX2TS U5641 ( .A(\indexIncrementer_EAST[1] ), .Y(\add_0_root_r1459/B[4] )
         );
  NAND2X1TS U5642 ( .A(n5766), .B(n3723), .Y(n3108) );
  CLKBUFX2TS U5643 ( .A(n2009), .Y(n5213) );
  CLKBUFX2TS U5644 ( .A(n1920), .Y(n5307) );
  CLKBUFX2TS U5645 ( .A(n1831), .Y(n5385) );
  OAI31XLTS U5646 ( .A0(n2564), .A1(n5705), .A2(n4578), .B0(n5151), .Y(n2088)
         );
  CLKBUFX2TS U5647 ( .A(n2428), .Y(n5063) );
  CLKBUFX2TS U5648 ( .A(n2009), .Y(n5214) );
  CLKBUFX2TS U5649 ( .A(n1920), .Y(n5308) );
  CLKBUFX2TS U5650 ( .A(n1831), .Y(n5386) );
  CLKBUFX2TS U5651 ( .A(n1965), .Y(n5253) );
  XNOR2X1TS U5652 ( .A(n3151), .B(n3723), .Y(totalAccesses[0]) );
  OAI21X1TS U5653 ( .A0(n5564), .A1(n1786), .B0(n5761), .Y(n1781) );
  INVX2TS U5654 ( .A(n2263), .Y(n5761) );
  OA21XLTS U5655 ( .A0(n2262), .A1(n4567), .B0(n4670), .Y(n2266) );
  OAI21X1TS U5656 ( .A0(n5563), .A1(n1743), .B0(n5764), .Y(n1738) );
  INVX2TS U5657 ( .A(n2209), .Y(n5764) );
  OA21XLTS U5658 ( .A0(n2208), .A1(n4569), .B0(n5973), .Y(n2212) );
  NAND2X1TS U5659 ( .A(n3110), .B(n3764), .Y(n2132) );
  NOR3X1TS U5660 ( .A(n1563), .B(n3729), .C(n5799), .Y(n1822) );
  NAND2X1TS U5661 ( .A(n2975), .B(n3764), .Y(n1786) );
  NAND2X1TS U5662 ( .A(n2423), .B(n3763), .Y(n1743) );
  NAND2X1TS U5663 ( .A(n2837), .B(n3764), .Y(n1775) );
  AOI211X1TS U5664 ( .A0(n4538), .A1(n2101), .B0(n5729), .C0(n5747), .Y(n3150)
         );
  INVX2TS U5665 ( .A(N610), .Y(n5747) );
  INVX2TS U5666 ( .A(n2286), .Y(n5804) );
  INVX2TS U5667 ( .A(n3727), .Y(n5805) );
  INVX2TS U5668 ( .A(n3697), .Y(n5773) );
  NOR2X1TS U5669 ( .A(n1735), .B(n3876), .Y(n1563) );
  OR2X2TS U5670 ( .A(n2834), .B(n1777), .Y(n2708) );
  OR2X2TS U5671 ( .A(n2560), .B(n1757), .Y(n2434) );
  INVX2TS U5672 ( .A(n3703), .Y(n5759) );
  CLKBUFX2TS U5673 ( .A(n2050), .Y(n5174) );
  CLKBUFX2TS U5674 ( .A(n1965), .Y(n5252) );
  CLKBUFX2TS U5675 ( .A(n1876), .Y(n5347) );
  CMPR32X2TS U5676 ( .A(totalAccesses[2]), .B(
        \add_0_root_sub_0_root_sub_231/B[2] ), .C(
        \add_0_root_sub_0_root_sub_231/carry [2]), .CO(
        \add_0_root_sub_0_root_sub_231/carry [3]), .S(N607) );
  CLKBUFX2TS U5677 ( .A(n2050), .Y(n5175) );
  AND2X2TS U5678 ( .A(N616), .B(n3150), .Y(n3643) );
  XNOR2X1TS U5679 ( .A(n5979), .B(n5981), .Y(N616) );
  XNOR2X1TS U5680 ( .A(n4525), .B(n5704), .Y(n5981) );
  AND2X2TS U5681 ( .A(N617), .B(n3150), .Y(n3642) );
  XOR2X1TS U5682 ( .A(n5977), .B(n5978), .Y(N617) );
  XNOR2X1TS U5683 ( .A(N614), .B(totalAccesses[2]), .Y(n5977) );
  AOI21X1TS U5684 ( .A0(n4525), .A1(n5979), .B0(n5980), .Y(n5978) );
  INVX2TS U5685 ( .A(N6618), .Y(n5796) );
  INVX2TS U5686 ( .A(N6371), .Y(n5795) );
  NAND2X1TS U5687 ( .A(n1735), .B(n5719), .Y(n1733) );
  INVX2TS U5688 ( .A(n3730), .Y(n5802) );
  NOR2X1TS U5689 ( .A(n1586), .B(n3729), .Y(n1584) );
  INVX2TS U5690 ( .A(n5681), .Y(n5668) );
  INVX2TS U5691 ( .A(n5655), .Y(n5642) );
  AND2X2TS U5692 ( .A(n2197), .B(n3728), .Y(n1645) );
  AND2X2TS U5693 ( .A(n1822), .B(n1585), .Y(n1669) );
  CLKBUFX2TS U5694 ( .A(n5666), .Y(n5665) );
  CLKBUFX2TS U5695 ( .A(n5666), .Y(n5664) );
  CLKBUFX2TS U5696 ( .A(n5666), .Y(n5663) );
  CLKBUFX2TS U5697 ( .A(n5641), .Y(n5640) );
  CLKBUFX2TS U5698 ( .A(n1548), .Y(n5639) );
  CLKBUFX2TS U5699 ( .A(n5667), .Y(n5661) );
  CLKBUFX2TS U5700 ( .A(n5667), .Y(n5662) );
  CLKBUFX2TS U5701 ( .A(n5641), .Y(n5638) );
  CLKBUFX2TS U5702 ( .A(n5975), .Y(n4713) );
  CLKBUFX2TS U5703 ( .A(n5975), .Y(n4714) );
  NAND4X1TS U5704 ( .A(\add_0_root_sub_0_root_sub_231/B[2] ), .B(n2120), .C(
        n4590), .D(n5709), .Y(n1766) );
  NAND4XLTS U5705 ( .A(N6316), .B(n5703), .C(n2120), .D(n4591), .Y(n1744) );
  NAND3XLTS U5706 ( .A(n2227), .B(n4592), .C(
        \add_0_root_sub_0_root_sub_231/B[2] ), .Y(n1756) );
  NAND3X1TS U5707 ( .A(n4592), .B(n5792), .C(n2227), .Y(n1799) );
  NAND3X1TS U5708 ( .A(\r1471/carry[3] ), .B(n4546), .C(N6316), .Y(n2214) );
  NAND4X1TS U5709 ( .A(n5702), .B(n2120), .C(n4592), .D(n5792), .Y(n1787) );
  NOR3X1TS U5710 ( .A(totalAccesses[1]), .B(totalAccesses[2]), .C(n4531), .Y(
        n2101) );
  INVX2TS U5711 ( .A(n2119), .Y(n5778) );
  OA21XLTS U5712 ( .A0(totalAccesses[1]), .A1(n5979), .B0(n5704), .Y(n5980) );
  CLKBUFX2TS U5713 ( .A(n5680), .Y(n5678) );
  CLKBUFX2TS U5714 ( .A(n5654), .Y(n5652) );
  INVX2TS U5715 ( .A(n5680), .Y(n5675) );
  INVX2TS U5716 ( .A(n5679), .Y(n5674) );
  INVX2TS U5717 ( .A(n5679), .Y(n5673) );
  INVX2TS U5718 ( .A(n5680), .Y(n5672) );
  INVX2TS U5719 ( .A(n5678), .Y(n5671) );
  INVX2TS U5720 ( .A(n5679), .Y(n5670) );
  INVX2TS U5721 ( .A(n5678), .Y(n5669) );
  INVX2TS U5722 ( .A(n5653), .Y(n5649) );
  INVX2TS U5723 ( .A(n5653), .Y(n5648) );
  INVX2TS U5724 ( .A(n5653), .Y(n5647) );
  INVX2TS U5725 ( .A(n5653), .Y(n5646) );
  INVX2TS U5726 ( .A(n5654), .Y(n5645) );
  INVX2TS U5727 ( .A(n5652), .Y(n5644) );
  INVX2TS U5728 ( .A(n5654), .Y(n5643) );
  CLKBUFX2TS U5729 ( .A(n5628), .Y(n5626) );
  INVX2TS U5730 ( .A(n1776), .Y(n5791) );
  CLKBUFX2TS U5731 ( .A(n4734), .Y(n4732) );
  CLKBUFX2TS U5732 ( .A(n4734), .Y(n4731) );
  CLKBUFX2TS U5733 ( .A(n4613), .Y(n5557) );
  CLKBUFX2TS U5734 ( .A(n5976), .Y(n4723) );
  INVX2TS U5735 ( .A(n4615), .Y(n5615) );
  CLKBUFX2TS U5736 ( .A(n4733), .Y(n4725) );
  CLKBUFX2TS U5737 ( .A(n4734), .Y(n4733) );
  CLKBUFX2TS U5738 ( .A(n5976), .Y(n4724) );
  INVX2TS U5739 ( .A(n5625), .Y(n5617) );
  INVX2TS U5740 ( .A(n5628), .Y(n5616) );
  INVX2TS U5741 ( .A(n5679), .Y(n5676) );
  CLKBUFX2TS U5742 ( .A(n5680), .Y(n5679) );
  INVX2TS U5743 ( .A(n5654), .Y(n5650) );
  CLKBUFX2TS U5744 ( .A(n5628), .Y(n5627) );
  CLKBUFX2TS U5745 ( .A(n5558), .Y(n5553) );
  CLKBUFX2TS U5746 ( .A(n4613), .Y(n5558) );
  CLKBUFX2TS U5747 ( .A(n5745), .Y(n5741) );
  NOR2X1TS U5748 ( .A(n2113), .B(n4617), .Y(n2112) );
  NAND2X1TS U5749 ( .A(n5793), .B(n3723), .Y(n2272) );
  AOI21X1TS U5750 ( .A0(n5565), .A1(n2246), .B0(n4539), .Y(n2243) );
  CLKBUFX2TS U5751 ( .A(n5744), .Y(n5743) );
  NAND2X1TS U5752 ( .A(N6699), .B(n2228), .Y(n1760) );
  NAND3XLTS U5753 ( .A(n2121), .B(n5711), .C(N6699), .Y(n1770) );
  NAND3XLTS U5754 ( .A(n910), .B(n2121), .C(N6699), .Y(n1749) );
  NAND3X1TS U5755 ( .A(n2121), .B(n5785), .C(n910), .Y(n1791) );
  AND3X2TS U5756 ( .A(n2120), .B(n5707), .C(n5792), .Y(n2111) );
  INVX2TS U5757 ( .A(n1780), .Y(n5784) );
  INVX2TS U5758 ( .A(n5709), .Y(n5704) );
  CLKBUFX2TS U5759 ( .A(n5745), .Y(n5742) );
  INVX2TS U5760 ( .A(n5707), .Y(n5706) );
  NAND2X1TS U5761 ( .A(N8209), .B(n2225), .Y(n2220) );
  NAND3XLTS U5762 ( .A(n2117), .B(n5711), .C(N8209), .Y(n2233) );
  NAND3XLTS U5763 ( .A(n5706), .B(n2117), .C(N8209), .Y(n2208) );
  OR2X2TS U5764 ( .A(n5710), .B(n5696), .Y(n4611) );
  NAND3X1TS U5765 ( .A(n2117), .B(n5794), .C(n910), .Y(n2262) );
  NAND3X1TS U5766 ( .A(N650), .B(n5785), .C(n2121), .Y(n2113) );
  NAND2X1TS U5767 ( .A(n2225), .B(n5794), .Y(n2275) );
  NAND3X1TS U5768 ( .A(n5707), .B(n5794), .C(n2117), .Y(n2114) );
  CLKBUFX2TS U5769 ( .A(n5694), .Y(n5682) );
  CLKBUFX2TS U5770 ( .A(n5972), .Y(n4675) );
  CLKBUFX2TS U5771 ( .A(n5973), .Y(n4690) );
  CLKBUFX2TS U5772 ( .A(n3804), .Y(n4703) );
  INVX2TS U5773 ( .A(\r1470/carry[3] ), .Y(N6701) );
  INVX2TS U5774 ( .A(n5708), .Y(n5705) );
  INVX2TS U5775 ( .A(n5710), .Y(n5702) );
  INVX2TS U5776 ( .A(N650), .Y(n5703) );
  NOR2X1TS U5777 ( .A(n5701), .B(n5714), .Y(n4612) );
  CLKBUFX2TS U5778 ( .A(n4614), .Y(n5296) );
  CLKBUFX2TS U5779 ( .A(n5972), .Y(n4676) );
  CLKBUFX2TS U5780 ( .A(n3804), .Y(n4704) );
  CLKBUFX2TS U5781 ( .A(n1565), .Y(n5600) );
  CLKBUFX2TS U5782 ( .A(n5695), .Y(n5690) );
  INVX2TS U5783 ( .A(\r1467/carry[3] ), .Y(N6318) );
  CLKBUFX2TS U5784 ( .A(n5601), .Y(n5595) );
  CLKBUFX2TS U5785 ( .A(n1565), .Y(n5601) );
  XOR2X1TS U5786 ( .A(n5704), .B(n5697), .Y(N614) );
  CLKBUFX2TS U5787 ( .A(n5694), .Y(n5683) );
  CLKBUFX2TS U5788 ( .A(n5691), .Y(n5689) );
  CLKBUFX2TS U5789 ( .A(n5691), .Y(n5688) );
  CLKBUFX2TS U5790 ( .A(n5692), .Y(n5687) );
  CLKBUFX2TS U5791 ( .A(n5692), .Y(n5686) );
  CLKBUFX2TS U5792 ( .A(n5693), .Y(n5685) );
  CLKBUFX2TS U5793 ( .A(n5693), .Y(n5684) );
  XNOR2X1TS U5794 ( .A(n1748), .B(n2255), .Y(n3156) );
  OAI22X1TS U5795 ( .A0(n4718), .A1(n5939), .B0(n4705), .B1(n5971), .Y(N10087)
         );
  OAI22X1TS U5796 ( .A0(n4718), .A1(n5938), .B0(n4705), .B1(n5970), .Y(N10088)
         );
  OAI22X1TS U5797 ( .A0(n4718), .A1(n5937), .B0(n4705), .B1(n5969), .Y(N10089)
         );
  OAI22X1TS U5798 ( .A0(n4718), .A1(n5936), .B0(n4711), .B1(n5968), .Y(N10090)
         );
  OAI22X1TS U5799 ( .A0(n4717), .A1(n5935), .B0(n4713), .B1(n5967), .Y(N10091)
         );
  OAI22X1TS U5800 ( .A0(n4717), .A1(n5934), .B0(n4713), .B1(n5966), .Y(N10092)
         );
  OAI22X1TS U5801 ( .A0(n4717), .A1(n5933), .B0(n4714), .B1(n5965), .Y(N10093)
         );
  OAI22X1TS U5802 ( .A0(n4717), .A1(n5932), .B0(n4711), .B1(n5964), .Y(N10094)
         );
  OAI22X1TS U5803 ( .A0(n4716), .A1(n5931), .B0(n4709), .B1(n5963), .Y(N10095)
         );
  OAI22X1TS U5804 ( .A0(n4716), .A1(n5930), .B0(n4714), .B1(n5962), .Y(N10096)
         );
  OAI22X1TS U5805 ( .A0(n4716), .A1(n5929), .B0(n5975), .B1(n5961), .Y(N10097)
         );
  OAI22X1TS U5806 ( .A0(n4716), .A1(n5928), .B0(n4712), .B1(n5960), .Y(N10098)
         );
  OAI22X1TS U5807 ( .A0(n4715), .A1(n5927), .B0(n4712), .B1(n5959), .Y(N10099)
         );
  OAI22X1TS U5808 ( .A0(n4715), .A1(n5926), .B0(n4711), .B1(n5958), .Y(N10100)
         );
  OAI22X1TS U5809 ( .A0(n4715), .A1(n5925), .B0(n4711), .B1(n5957), .Y(N10101)
         );
  OAI22X1TS U5810 ( .A0(n4715), .A1(n5924), .B0(n4712), .B1(n5956), .Y(N10102)
         );
  OAI22X1TS U5811 ( .A0(n4719), .A1(n5923), .B0(n4710), .B1(n5955), .Y(N10103)
         );
  OAI22X1TS U5812 ( .A0(n4724), .A1(n5922), .B0(n4710), .B1(n5954), .Y(N10104)
         );
  OAI22X1TS U5813 ( .A0(n5976), .A1(n5921), .B0(n4709), .B1(n5953), .Y(N10105)
         );
  OAI22X1TS U5814 ( .A0(n5976), .A1(n5920), .B0(n4706), .B1(n5952), .Y(N10106)
         );
  OAI22X1TS U5815 ( .A0(n4722), .A1(n5919), .B0(n4706), .B1(n5951), .Y(N10107)
         );
  OAI22X1TS U5816 ( .A0(n4722), .A1(n5918), .B0(n4706), .B1(n5950), .Y(N10108)
         );
  OAI22X1TS U5817 ( .A0(n4721), .A1(n5917), .B0(n4706), .B1(n5949), .Y(N10109)
         );
  OAI22X1TS U5818 ( .A0(n4723), .A1(n5916), .B0(n4707), .B1(n5948), .Y(N10110)
         );
  OAI22X1TS U5819 ( .A0(n4719), .A1(n5915), .B0(n4707), .B1(n5947), .Y(N10111)
         );
  OAI22X1TS U5820 ( .A0(n4720), .A1(n5914), .B0(n4707), .B1(n5946), .Y(N10112)
         );
  OAI22X1TS U5821 ( .A0(n4724), .A1(n5913), .B0(n4707), .B1(n5945), .Y(N10113)
         );
  OAI22X1TS U5822 ( .A0(n4722), .A1(n5912), .B0(n4708), .B1(n5944), .Y(N10114)
         );
  OAI22X1TS U5823 ( .A0(n4721), .A1(n5911), .B0(n4708), .B1(n5943), .Y(N10115)
         );
  OAI22X1TS U5824 ( .A0(n4722), .A1(n5910), .B0(n4708), .B1(n5942), .Y(N10116)
         );
  OAI22X1TS U5825 ( .A0(n4720), .A1(n5909), .B0(n4708), .B1(n5941), .Y(N10117)
         );
  OAI22X1TS U5826 ( .A0(n4723), .A1(n5908), .B0(n4709), .B1(n5940), .Y(N10118)
         );
  OAI22X1TS U5827 ( .A0(n5676), .A1(n5939), .B0(n5656), .B1(n5971), .Y(N10121)
         );
  OAI22X1TS U5828 ( .A0(n5675), .A1(n5938), .B0(n5656), .B1(n5970), .Y(N10122)
         );
  OAI22X1TS U5829 ( .A0(n5675), .A1(n5937), .B0(n5656), .B1(n5969), .Y(N10123)
         );
  OAI22X1TS U5830 ( .A0(n5675), .A1(n5936), .B0(n5665), .B1(n5968), .Y(N10124)
         );
  OAI22X1TS U5831 ( .A0(n5675), .A1(n5935), .B0(n5665), .B1(n5967), .Y(N10125)
         );
  OAI22X1TS U5832 ( .A0(n5674), .A1(n5934), .B0(n5661), .B1(n5966), .Y(N10126)
         );
  OAI22X1TS U5833 ( .A0(n5674), .A1(n5933), .B0(n1539), .B1(n5965), .Y(N10127)
         );
  OAI22X1TS U5834 ( .A0(n5674), .A1(n5932), .B0(n5664), .B1(n5964), .Y(N10128)
         );
  OAI22X1TS U5835 ( .A0(n5672), .A1(n5931), .B0(n5664), .B1(n5963), .Y(N10129)
         );
  OAI22X1TS U5836 ( .A0(n5674), .A1(n5930), .B0(n5662), .B1(n5962), .Y(N10130)
         );
  OAI22X1TS U5837 ( .A0(n5673), .A1(n5929), .B0(n5667), .B1(n5961), .Y(N10131)
         );
  OAI22X1TS U5838 ( .A0(n5673), .A1(n5928), .B0(n5664), .B1(n5960), .Y(N10132)
         );
  OAI22X1TS U5839 ( .A0(n5673), .A1(n5927), .B0(n5661), .B1(n5959), .Y(N10133)
         );
  OAI22X1TS U5840 ( .A0(n5673), .A1(n5926), .B0(n5665), .B1(n5958), .Y(N10134)
         );
  OAI22X1TS U5841 ( .A0(n5672), .A1(n5925), .B0(n5664), .B1(n5957), .Y(N10135)
         );
  OAI22X1TS U5842 ( .A0(n5672), .A1(n5924), .B0(n5663), .B1(n5956), .Y(N10136)
         );
  OAI22X1TS U5843 ( .A0(n5672), .A1(n5923), .B0(n5663), .B1(n5955), .Y(N10137)
         );
  OAI22X1TS U5844 ( .A0(n5671), .A1(n5922), .B0(n5663), .B1(n5954), .Y(N10138)
         );
  OAI22X1TS U5845 ( .A0(n5671), .A1(n5921), .B0(n5666), .B1(n5953), .Y(N10139)
         );
  OAI22X1TS U5846 ( .A0(n5671), .A1(n5920), .B0(n5660), .B1(n5952), .Y(N10140)
         );
  OAI22X1TS U5847 ( .A0(n5671), .A1(n5919), .B0(n5662), .B1(n5951), .Y(N10141)
         );
  OAI22X1TS U5848 ( .A0(n5670), .A1(n5918), .B0(n5663), .B1(n5950), .Y(N10142)
         );
  OAI22X1TS U5849 ( .A0(n5670), .A1(n5917), .B0(n5667), .B1(n5949), .Y(N10143)
         );
  OAI22X1TS U5850 ( .A0(n5670), .A1(n5916), .B0(n5657), .B1(n5948), .Y(N10144)
         );
  OAI22X1TS U5851 ( .A0(n5670), .A1(n5915), .B0(n5657), .B1(n5947), .Y(N10145)
         );
  OAI22X1TS U5852 ( .A0(n5669), .A1(n5914), .B0(n5657), .B1(n5946), .Y(N10146)
         );
  OAI22X1TS U5853 ( .A0(n5669), .A1(n5913), .B0(n5657), .B1(n5945), .Y(N10147)
         );
  OAI22X1TS U5854 ( .A0(n5669), .A1(n5912), .B0(n5658), .B1(n5944), .Y(N10148)
         );
  OAI22X1TS U5855 ( .A0(n5669), .A1(n5911), .B0(n5658), .B1(n5943), .Y(N10149)
         );
  OAI22X1TS U5856 ( .A0(n5668), .A1(n5910), .B0(n5658), .B1(n5942), .Y(N10150)
         );
  OAI22X1TS U5857 ( .A0(n5668), .A1(n5909), .B0(n5658), .B1(n5941), .Y(N10151)
         );
  OAI22X1TS U5858 ( .A0(n5668), .A1(n5908), .B0(n5659), .B1(n5940), .Y(N10152)
         );
  OAI22X1TS U5859 ( .A0(n5650), .A1(n5939), .B0(n5637), .B1(n5971), .Y(N10155)
         );
  OAI22X1TS U5860 ( .A0(n5649), .A1(n5938), .B0(n5638), .B1(n5970), .Y(N10156)
         );
  OAI22X1TS U5861 ( .A0(n5649), .A1(n5937), .B0(n1548), .B1(n5969), .Y(N10157)
         );
  OAI22X1TS U5862 ( .A0(n5649), .A1(n5936), .B0(n5630), .B1(n5968), .Y(N10158)
         );
  OAI22X1TS U5863 ( .A0(n5649), .A1(n5935), .B0(n5630), .B1(n5967), .Y(N10159)
         );
  OAI22X1TS U5864 ( .A0(n5648), .A1(n5934), .B0(n5630), .B1(n5966), .Y(N10160)
         );
  OAI22X1TS U5865 ( .A0(n5648), .A1(n5933), .B0(n5630), .B1(n5965), .Y(N10161)
         );
  OAI22X1TS U5866 ( .A0(n5648), .A1(n5932), .B0(n5631), .B1(n5964), .Y(N10162)
         );
  OAI22X1TS U5867 ( .A0(n5646), .A1(n5931), .B0(n5631), .B1(n5963), .Y(N10163)
         );
  OAI22X1TS U5868 ( .A0(n5648), .A1(n5930), .B0(n5631), .B1(n5962), .Y(N10164)
         );
  OAI22X1TS U5869 ( .A0(n5647), .A1(n5929), .B0(n5631), .B1(n5961), .Y(N10165)
         );
  OAI22X1TS U5870 ( .A0(n5647), .A1(n5928), .B0(n5632), .B1(n5960), .Y(N10166)
         );
  OAI22X1TS U5871 ( .A0(n5647), .A1(n5927), .B0(n5632), .B1(n5959), .Y(N10167)
         );
  OAI22X1TS U5872 ( .A0(n5647), .A1(n5926), .B0(n5632), .B1(n5958), .Y(N10168)
         );
  OAI22X1TS U5873 ( .A0(n5646), .A1(n5925), .B0(n5632), .B1(n5957), .Y(N10169)
         );
  OAI22X1TS U5874 ( .A0(n5646), .A1(n5924), .B0(n5633), .B1(n5956), .Y(N10170)
         );
  OAI22X1TS U5875 ( .A0(n5646), .A1(n5923), .B0(n5633), .B1(n5955), .Y(N10171)
         );
  OAI22X1TS U5876 ( .A0(n5645), .A1(n5922), .B0(n5633), .B1(n5954), .Y(N10172)
         );
  OAI22X1TS U5877 ( .A0(n5645), .A1(n5921), .B0(n5633), .B1(n5953), .Y(N10173)
         );
  OAI22X1TS U5878 ( .A0(n5645), .A1(n5920), .B0(n5634), .B1(n5952), .Y(N10174)
         );
  OAI22X1TS U5879 ( .A0(n5645), .A1(n5919), .B0(n5634), .B1(n5951), .Y(N10175)
         );
  OAI22X1TS U5880 ( .A0(n5644), .A1(n5918), .B0(n5634), .B1(n5950), .Y(N10176)
         );
  OAI22X1TS U5881 ( .A0(n5644), .A1(n5917), .B0(n5634), .B1(n5949), .Y(N10177)
         );
  OAI22X1TS U5882 ( .A0(n5644), .A1(n5916), .B0(n5635), .B1(n5948), .Y(N10178)
         );
  OAI22X1TS U5883 ( .A0(n5644), .A1(n5915), .B0(n5635), .B1(n5947), .Y(N10179)
         );
  OAI22X1TS U5884 ( .A0(n5643), .A1(n5914), .B0(n5635), .B1(n5946), .Y(N10180)
         );
  OAI22X1TS U5885 ( .A0(n5643), .A1(n5913), .B0(n5635), .B1(n5945), .Y(N10181)
         );
  OAI22X1TS U5886 ( .A0(n5643), .A1(n5912), .B0(n5636), .B1(n5944), .Y(N10182)
         );
  OAI22X1TS U5887 ( .A0(n5643), .A1(n5911), .B0(n5636), .B1(n5943), .Y(N10183)
         );
  OAI22X1TS U5888 ( .A0(n5642), .A1(n5910), .B0(n5636), .B1(n5942), .Y(N10184)
         );
  OAI22X1TS U5889 ( .A0(n5642), .A1(n5909), .B0(n5636), .B1(n5941), .Y(N10185)
         );
  OAI22X1TS U5890 ( .A0(n5642), .A1(n5908), .B0(n5640), .B1(n5940), .Y(N10186)
         );
  OAI22X1TS U5891 ( .A0(n5623), .A1(n5939), .B0(n4725), .B1(n5971), .Y(N10189)
         );
  OAI22X1TS U5892 ( .A0(n5622), .A1(n5938), .B0(n4725), .B1(n5970), .Y(N10190)
         );
  OAI22X1TS U5893 ( .A0(n5622), .A1(n5937), .B0(n4725), .B1(n5969), .Y(N10191)
         );
  OAI22X1TS U5894 ( .A0(n5622), .A1(n5936), .B0(n4733), .B1(n5968), .Y(N10192)
         );
  OAI22X1TS U5895 ( .A0(n5622), .A1(n5935), .B0(n3157), .B1(n5967), .Y(N10193)
         );
  OAI22X1TS U5896 ( .A0(n5621), .A1(n5934), .B0(n4731), .B1(n5966), .Y(N10194)
         );
  OAI22X1TS U5897 ( .A0(n5621), .A1(n5933), .B0(n4732), .B1(n5965), .Y(N10195)
         );
  OAI22X1TS U5898 ( .A0(n5621), .A1(n5932), .B0(n4733), .B1(n5964), .Y(N10196)
         );
  OAI22X1TS U5899 ( .A0(n5619), .A1(n5931), .B0(n4732), .B1(n5963), .Y(N10197)
         );
  OAI22X1TS U5900 ( .A0(n5621), .A1(n5930), .B0(n4734), .B1(n5962), .Y(N10198)
         );
  OAI22X1TS U5901 ( .A0(n5620), .A1(n5929), .B0(n4731), .B1(n5961), .Y(N10199)
         );
  OAI22X1TS U5902 ( .A0(n5620), .A1(n5928), .B0(n4726), .B1(n5960), .Y(N10200)
         );
  OAI22X1TS U5903 ( .A0(n5620), .A1(n5927), .B0(n4726), .B1(n5959), .Y(N10201)
         );
  OAI22X1TS U5904 ( .A0(n5620), .A1(n5926), .B0(n4726), .B1(n5958), .Y(N10202)
         );
  OAI22X1TS U5905 ( .A0(n5619), .A1(n5925), .B0(n4726), .B1(n5957), .Y(N10203)
         );
  OAI22X1TS U5906 ( .A0(n5619), .A1(n5924), .B0(n4727), .B1(n5956), .Y(N10204)
         );
  OAI22X1TS U5907 ( .A0(n5619), .A1(n5923), .B0(n4727), .B1(n5955), .Y(N10205)
         );
  OAI22X1TS U5908 ( .A0(n5618), .A1(n5922), .B0(n4727), .B1(n5954), .Y(N10206)
         );
  OAI22X1TS U5909 ( .A0(n5618), .A1(n5921), .B0(n4727), .B1(n5953), .Y(N10207)
         );
  OAI22X1TS U5910 ( .A0(n5618), .A1(n5920), .B0(n4728), .B1(n5952), .Y(N10208)
         );
  OAI22X1TS U5911 ( .A0(n5618), .A1(n5919), .B0(n4728), .B1(n5951), .Y(N10209)
         );
  OAI22X1TS U5912 ( .A0(n5617), .A1(n5918), .B0(n4728), .B1(n5950), .Y(N10210)
         );
  OAI22X1TS U5913 ( .A0(n5617), .A1(n5917), .B0(n4728), .B1(n5949), .Y(N10211)
         );
  OAI22X1TS U5914 ( .A0(n5617), .A1(n5916), .B0(n4729), .B1(n5948), .Y(N10212)
         );
  OAI22X1TS U5915 ( .A0(n5617), .A1(n5915), .B0(n4729), .B1(n5947), .Y(N10213)
         );
  OAI22X1TS U5916 ( .A0(n5616), .A1(n5914), .B0(n4729), .B1(n5946), .Y(N10214)
         );
  OAI22X1TS U5917 ( .A0(n5616), .A1(n5913), .B0(n4729), .B1(n5945), .Y(N10215)
         );
  OAI22X1TS U5918 ( .A0(n5616), .A1(n5912), .B0(n4730), .B1(n5944), .Y(N10216)
         );
  OAI22X1TS U5919 ( .A0(n5616), .A1(n5911), .B0(n4730), .B1(n5943), .Y(N10217)
         );
  OAI22X1TS U5920 ( .A0(n5615), .A1(n5910), .B0(n4730), .B1(n5942), .Y(N10218)
         );
  OAI22X1TS U5921 ( .A0(n5615), .A1(n5909), .B0(n4730), .B1(n5941), .Y(N10219)
         );
  OAI22X1TS U5922 ( .A0(n5615), .A1(n5908), .B0(n4731), .B1(n5940), .Y(N10220)
         );
  NOR2X1TS U5923 ( .A(n1999), .B(n4601), .Y(n2834) );
  AOI211X1TS U5924 ( .A0(n1757), .A1(n5583), .B0(n4601), .C0(n3708), .Y(n1876)
         );
  OAI21X1TS U5925 ( .A0(n5563), .A1(n1765), .B0(n2235), .Y(n1761) );
  AOI2BB2X1TS U5926 ( .B0(n2238), .B1(n5563), .A0N(n2233), .A1N(n4569), .Y(
        n2237) );
  OAI211X1TS U5927 ( .A0(n5840), .A1(n1770), .B0(n2239), .C0(n1766), .Y(n2238)
         );
  OAI21X1TS U5928 ( .A0(n5564), .A1(n1775), .B0(n5767), .Y(n1771) );
  INVX2TS U5929 ( .A(n2247), .Y(n5767) );
  OAI211X1TS U5930 ( .A0(n5593), .A1(n2248), .B0(n2249), .C0(n2250), .Y(n2247)
         );
  OA21XLTS U5931 ( .A0(n2246), .A1(n4568), .B0(n5693), .Y(n2250) );
  OAI21X1TS U5932 ( .A0(n5564), .A1(n1755), .B0(n5769), .Y(n1750) );
  INVX2TS U5933 ( .A(n2221), .Y(n5769) );
  OAI211X1TS U5934 ( .A0(n5589), .A1(n2222), .B0(n2223), .C0(n2224), .Y(n2221)
         );
  OA21XLTS U5935 ( .A0(n2220), .A1(n4568), .B0(n4697), .Y(n2224) );
  OAI22X1TS U5936 ( .A0(n4823), .A1(n5809), .B0(n5842), .B1(n4834), .Y(n2852)
         );
  OAI22X1TS U5937 ( .A0(n4947), .A1(n5809), .B0(n5842), .B1(n4958), .Y(n2578)
         );
  OAI22X1TS U5938 ( .A0(n5071), .A1(n5809), .B0(n5842), .B1(n5082), .Y(n2299)
         );
  OAI22X1TS U5939 ( .A0(n4885), .A1(n3949), .B0(n4027), .B1(n4895), .Y(n2714)
         );
  OAI22X1TS U5940 ( .A0(n5010), .A1(n5809), .B0(n5842), .B1(n5021), .Y(n2440)
         );
  OAI22X1TS U5941 ( .A0(n4820), .A1(n5821), .B0(n5854), .B1(n4831), .Y(n2900)
         );
  OAI22X1TS U5942 ( .A0(n4944), .A1(n5821), .B0(n5854), .B1(n4955), .Y(n2626)
         );
  OAI22X1TS U5943 ( .A0(n5068), .A1(n5821), .B0(n5854), .B1(n5079), .Y(n2347)
         );
  OAI22X1TS U5944 ( .A0(n4821), .A1(n5820), .B0(n5853), .B1(n4831), .Y(n2896)
         );
  OAI22X1TS U5945 ( .A0(n4945), .A1(n5820), .B0(n5853), .B1(n4955), .Y(n2622)
         );
  OAI22X1TS U5946 ( .A0(n5069), .A1(n5820), .B0(n5853), .B1(n5079), .Y(n2343)
         );
  OAI22X1TS U5947 ( .A0(n4821), .A1(n5819), .B0(n5852), .B1(n4831), .Y(n2892)
         );
  OAI22X1TS U5948 ( .A0(n4945), .A1(n5819), .B0(n5852), .B1(n4955), .Y(n2618)
         );
  OAI22X1TS U5949 ( .A0(n5069), .A1(n5819), .B0(n5852), .B1(n5079), .Y(n2339)
         );
  OAI22X1TS U5950 ( .A0(n4821), .A1(n5818), .B0(n5851), .B1(n4831), .Y(n2888)
         );
  OAI22X1TS U5951 ( .A0(n4945), .A1(n5818), .B0(n5851), .B1(n4955), .Y(n2614)
         );
  OAI22X1TS U5952 ( .A0(n5069), .A1(n5818), .B0(n5851), .B1(n5079), .Y(n2335)
         );
  OAI22X1TS U5953 ( .A0(n4821), .A1(n5817), .B0(n5850), .B1(n4832), .Y(n2884)
         );
  OAI22X1TS U5954 ( .A0(n4945), .A1(n5817), .B0(n5850), .B1(n4956), .Y(n2610)
         );
  OAI22X1TS U5955 ( .A0(n5069), .A1(n5817), .B0(n5850), .B1(n5080), .Y(n2331)
         );
  OAI22X1TS U5956 ( .A0(n4822), .A1(n5816), .B0(n5849), .B1(n4832), .Y(n2880)
         );
  OAI22X1TS U5957 ( .A0(n4946), .A1(n5816), .B0(n5849), .B1(n4956), .Y(n2606)
         );
  OAI22X1TS U5958 ( .A0(n5070), .A1(n5816), .B0(n5849), .B1(n5080), .Y(n2327)
         );
  OAI22X1TS U5959 ( .A0(n4822), .A1(n5815), .B0(n5848), .B1(n4832), .Y(n2876)
         );
  OAI22X1TS U5960 ( .A0(n4946), .A1(n5815), .B0(n5848), .B1(n4956), .Y(n2602)
         );
  OAI22X1TS U5961 ( .A0(n5070), .A1(n5815), .B0(n5848), .B1(n5080), .Y(n2323)
         );
  OAI22X1TS U5962 ( .A0(n4822), .A1(n5814), .B0(n5847), .B1(n4832), .Y(n2872)
         );
  OAI22X1TS U5963 ( .A0(n4946), .A1(n5814), .B0(n5847), .B1(n4956), .Y(n2598)
         );
  OAI22X1TS U5964 ( .A0(n5070), .A1(n5814), .B0(n5847), .B1(n5080), .Y(n2319)
         );
  OAI22X1TS U5965 ( .A0(n4822), .A1(n5813), .B0(n5846), .B1(n4833), .Y(n2868)
         );
  OAI22X1TS U5966 ( .A0(n4946), .A1(n5813), .B0(n5846), .B1(n4957), .Y(n2594)
         );
  OAI22X1TS U5967 ( .A0(n5070), .A1(n5813), .B0(n5846), .B1(n5081), .Y(n2315)
         );
  OAI22X1TS U5968 ( .A0(n4823), .A1(n5812), .B0(n5845), .B1(n4833), .Y(n2864)
         );
  OAI22X1TS U5969 ( .A0(n4947), .A1(n5812), .B0(n5845), .B1(n4957), .Y(n2590)
         );
  OAI22X1TS U5970 ( .A0(n5071), .A1(n5812), .B0(n5845), .B1(n5081), .Y(n2311)
         );
  OAI22X1TS U5971 ( .A0(n4823), .A1(n5811), .B0(n5844), .B1(n4833), .Y(n2860)
         );
  OAI22X1TS U5972 ( .A0(n4947), .A1(n5811), .B0(n5844), .B1(n4957), .Y(n2586)
         );
  OAI22X1TS U5973 ( .A0(n5071), .A1(n5811), .B0(n5844), .B1(n5081), .Y(n2307)
         );
  OAI22X1TS U5974 ( .A0(n4823), .A1(n5810), .B0(n5843), .B1(n4833), .Y(n2856)
         );
  OAI22X1TS U5975 ( .A0(n4947), .A1(n5810), .B0(n5843), .B1(n4957), .Y(n2582)
         );
  OAI22X1TS U5976 ( .A0(n5071), .A1(n5810), .B0(n5843), .B1(n5081), .Y(n2303)
         );
  OAI22X1TS U5977 ( .A0(n4882), .A1(n3925), .B0(n4003), .B1(n4892), .Y(n2762)
         );
  OAI22X1TS U5978 ( .A0(n4883), .A1(n3927), .B0(n4005), .B1(n4892), .Y(n2758)
         );
  OAI22X1TS U5979 ( .A0(n4883), .A1(n3929), .B0(n4007), .B1(n4892), .Y(n2754)
         );
  OAI22X1TS U5980 ( .A0(n4883), .A1(n3931), .B0(n4009), .B1(n4892), .Y(n2750)
         );
  OAI22X1TS U5981 ( .A0(n4883), .A1(n3933), .B0(n4011), .B1(n4893), .Y(n2746)
         );
  OAI22X1TS U5982 ( .A0(n4884), .A1(n3935), .B0(n4013), .B1(n4893), .Y(n2742)
         );
  OAI22X1TS U5983 ( .A0(n4884), .A1(n3937), .B0(n4015), .B1(n4893), .Y(n2738)
         );
  OAI22X1TS U5984 ( .A0(n4884), .A1(n3939), .B0(n4017), .B1(n4893), .Y(n2734)
         );
  OAI22X1TS U5985 ( .A0(n4884), .A1(n3941), .B0(n4019), .B1(n4894), .Y(n2730)
         );
  OAI22X1TS U5986 ( .A0(n4885), .A1(n3943), .B0(n4021), .B1(n4894), .Y(n2726)
         );
  OAI22X1TS U5987 ( .A0(n4885), .A1(n3945), .B0(n4023), .B1(n4894), .Y(n2722)
         );
  OAI22X1TS U5988 ( .A0(n4885), .A1(n3947), .B0(n4025), .B1(n4894), .Y(n2718)
         );
  OAI22X1TS U5989 ( .A0(n5007), .A1(n5821), .B0(n5854), .B1(n5018), .Y(n2488)
         );
  OAI22X1TS U5990 ( .A0(n5008), .A1(n5820), .B0(n5853), .B1(n5018), .Y(n2484)
         );
  OAI22X1TS U5991 ( .A0(n5008), .A1(n5819), .B0(n5852), .B1(n5018), .Y(n2480)
         );
  OAI22X1TS U5992 ( .A0(n5008), .A1(n5818), .B0(n5851), .B1(n5018), .Y(n2476)
         );
  OAI22X1TS U5993 ( .A0(n5008), .A1(n5817), .B0(n5850), .B1(n5019), .Y(n2472)
         );
  OAI22X1TS U5994 ( .A0(n5009), .A1(n5816), .B0(n5849), .B1(n5019), .Y(n2468)
         );
  OAI22X1TS U5995 ( .A0(n5009), .A1(n5815), .B0(n5848), .B1(n5019), .Y(n2464)
         );
  OAI22X1TS U5996 ( .A0(n5009), .A1(n5814), .B0(n5847), .B1(n5019), .Y(n2460)
         );
  OAI22X1TS U5997 ( .A0(n5009), .A1(n5813), .B0(n5846), .B1(n5020), .Y(n2456)
         );
  OAI22X1TS U5998 ( .A0(n5010), .A1(n5812), .B0(n5845), .B1(n5020), .Y(n2452)
         );
  OAI22X1TS U5999 ( .A0(n5010), .A1(n5811), .B0(n5844), .B1(n5020), .Y(n2448)
         );
  OAI22X1TS U6000 ( .A0(n5010), .A1(n5810), .B0(n5843), .B1(n5020), .Y(n2444)
         );
  OAI22X1TS U6001 ( .A0(n4816), .A1(n5839), .B0(n5872), .B1(n4830), .Y(n2973)
         );
  OAI22X1TS U6002 ( .A0(n4940), .A1(n5839), .B0(n5872), .B1(n4949), .Y(n2699)
         );
  OAI22X1TS U6003 ( .A0(n5064), .A1(n5839), .B0(n5872), .B1(n5082), .Y(n2420)
         );
  OAI22X1TS U6004 ( .A0(n4816), .A1(n5838), .B0(n5871), .B1(n4826), .Y(n2968)
         );
  OAI22X1TS U6005 ( .A0(n4940), .A1(n5838), .B0(n5871), .B1(n4949), .Y(n2694)
         );
  OAI22X1TS U6006 ( .A0(n5064), .A1(n5838), .B0(n5871), .B1(n5077), .Y(n2415)
         );
  OAI22X1TS U6007 ( .A0(n4816), .A1(n5837), .B0(n5870), .B1(n4825), .Y(n2964)
         );
  OAI22X1TS U6008 ( .A0(n4940), .A1(n5837), .B0(n5870), .B1(n4950), .Y(n2690)
         );
  OAI22X1TS U6009 ( .A0(n5064), .A1(n5837), .B0(n5870), .B1(n5073), .Y(n2411)
         );
  OAI22X1TS U6010 ( .A0(n4817), .A1(n5836), .B0(n5869), .B1(n4825), .Y(n2960)
         );
  OAI22X1TS U6011 ( .A0(n4941), .A1(n5836), .B0(n5869), .B1(n4950), .Y(n2686)
         );
  OAI22X1TS U6012 ( .A0(n5065), .A1(n5836), .B0(n5869), .B1(n5073), .Y(n2407)
         );
  OAI22X1TS U6013 ( .A0(n4817), .A1(n5835), .B0(n5868), .B1(n4826), .Y(n2956)
         );
  OAI22X1TS U6014 ( .A0(n4941), .A1(n5835), .B0(n5868), .B1(n4951), .Y(n2682)
         );
  OAI22X1TS U6015 ( .A0(n5065), .A1(n5835), .B0(n5868), .B1(n5074), .Y(n2403)
         );
  OAI22X1TS U6016 ( .A0(n4817), .A1(n5834), .B0(n5867), .B1(n4826), .Y(n2952)
         );
  OAI22X1TS U6017 ( .A0(n4941), .A1(n5834), .B0(n5867), .B1(n4951), .Y(n2678)
         );
  OAI22X1TS U6018 ( .A0(n5065), .A1(n5834), .B0(n5867), .B1(n5074), .Y(n2399)
         );
  OAI22X1TS U6019 ( .A0(n4817), .A1(n5833), .B0(n5866), .B1(n4827), .Y(n2948)
         );
  OAI22X1TS U6020 ( .A0(n4941), .A1(n5833), .B0(n5866), .B1(n4952), .Y(n2674)
         );
  OAI22X1TS U6021 ( .A0(n5065), .A1(n5833), .B0(n5866), .B1(n5075), .Y(n2395)
         );
  OAI22X1TS U6022 ( .A0(n4818), .A1(n5832), .B0(n5865), .B1(n4827), .Y(n2944)
         );
  OAI22X1TS U6023 ( .A0(n4942), .A1(n5832), .B0(n5865), .B1(n4952), .Y(n2670)
         );
  OAI22X1TS U6024 ( .A0(n5066), .A1(n5832), .B0(n5865), .B1(n5075), .Y(n2391)
         );
  OAI22X1TS U6025 ( .A0(n4818), .A1(n5831), .B0(n5864), .B1(n4828), .Y(n2940)
         );
  OAI22X1TS U6026 ( .A0(n4942), .A1(n5831), .B0(n5864), .B1(n4953), .Y(n2666)
         );
  OAI22X1TS U6027 ( .A0(n5066), .A1(n5831), .B0(n5864), .B1(n5076), .Y(n2387)
         );
  OAI22X1TS U6028 ( .A0(n4818), .A1(n5830), .B0(n5863), .B1(n4828), .Y(n2936)
         );
  OAI22X1TS U6029 ( .A0(n4942), .A1(n5830), .B0(n5863), .B1(n4953), .Y(n2662)
         );
  OAI22X1TS U6030 ( .A0(n5066), .A1(n5830), .B0(n5863), .B1(n5076), .Y(n2383)
         );
  OAI22X1TS U6031 ( .A0(n4818), .A1(n5829), .B0(n5862), .B1(n4829), .Y(n2932)
         );
  OAI22X1TS U6032 ( .A0(n4942), .A1(n5829), .B0(n5862), .B1(n4961), .Y(n2658)
         );
  OAI22X1TS U6033 ( .A0(n5066), .A1(n5829), .B0(n5862), .B1(n5077), .Y(n2379)
         );
  OAI22X1TS U6034 ( .A0(n4819), .A1(n5828), .B0(n5861), .B1(n4829), .Y(n2928)
         );
  OAI22X1TS U6035 ( .A0(n4943), .A1(n5828), .B0(n5861), .B1(n4949), .Y(n2654)
         );
  OAI22X1TS U6036 ( .A0(n5067), .A1(n5828), .B0(n5861), .B1(n5077), .Y(n2375)
         );
  OAI22X1TS U6037 ( .A0(n4819), .A1(n5827), .B0(n5860), .B1(n4825), .Y(n2924)
         );
  OAI22X1TS U6038 ( .A0(n4943), .A1(n5827), .B0(n5860), .B1(n4958), .Y(n2650)
         );
  OAI22X1TS U6039 ( .A0(n5067), .A1(n5827), .B0(n5860), .B1(n5073), .Y(n2371)
         );
  OAI22X1TS U6040 ( .A0(n4819), .A1(n5826), .B0(n5859), .B1(n4827), .Y(n2920)
         );
  OAI22X1TS U6041 ( .A0(n4943), .A1(n5826), .B0(n5859), .B1(n4958), .Y(n2646)
         );
  OAI22X1TS U6042 ( .A0(n5067), .A1(n5826), .B0(n5859), .B1(n5075), .Y(n2367)
         );
  OAI22X1TS U6043 ( .A0(n4819), .A1(n5825), .B0(n5858), .B1(n4830), .Y(n2916)
         );
  OAI22X1TS U6044 ( .A0(n4943), .A1(n5825), .B0(n5858), .B1(n4954), .Y(n2642)
         );
  OAI22X1TS U6045 ( .A0(n5067), .A1(n5825), .B0(n5858), .B1(n5085), .Y(n2363)
         );
  OAI22X1TS U6046 ( .A0(n4820), .A1(n5824), .B0(n5857), .B1(n4830), .Y(n2912)
         );
  OAI22X1TS U6047 ( .A0(n4944), .A1(n5824), .B0(n5857), .B1(n4954), .Y(n2638)
         );
  OAI22X1TS U6048 ( .A0(n5068), .A1(n5824), .B0(n5857), .B1(n5074), .Y(n2359)
         );
  OAI22X1TS U6049 ( .A0(n4820), .A1(n5823), .B0(n5856), .B1(n4834), .Y(n2908)
         );
  OAI22X1TS U6050 ( .A0(n4944), .A1(n5823), .B0(n5856), .B1(n4954), .Y(n2634)
         );
  OAI22X1TS U6051 ( .A0(n5068), .A1(n5823), .B0(n5856), .B1(n5078), .Y(n2355)
         );
  OAI22X1TS U6052 ( .A0(n4820), .A1(n5822), .B0(n5855), .B1(n4834), .Y(n2904)
         );
  OAI22X1TS U6053 ( .A0(n4944), .A1(n5822), .B0(n5855), .B1(n4953), .Y(n2630)
         );
  OAI22X1TS U6054 ( .A0(n5068), .A1(n5822), .B0(n5855), .B1(n5078), .Y(n2351)
         );
  OAI22X1TS U6055 ( .A0(n4878), .A1(n3889), .B0(n3967), .B1(n4887), .Y(n2835)
         );
  OAI22X1TS U6056 ( .A0(n4878), .A1(n3891), .B0(n3969), .B1(n4887), .Y(n2830)
         );
  OAI22X1TS U6057 ( .A0(n4878), .A1(n3893), .B0(n3971), .B1(n4888), .Y(n2826)
         );
  OAI22X1TS U6058 ( .A0(n4879), .A1(n3895), .B0(n3973), .B1(n4888), .Y(n2822)
         );
  OAI22X1TS U6059 ( .A0(n4879), .A1(n3897), .B0(n3975), .B1(n4889), .Y(n2818)
         );
  OAI22X1TS U6060 ( .A0(n4879), .A1(n3899), .B0(n3977), .B1(n4889), .Y(n2814)
         );
  OAI22X1TS U6061 ( .A0(n4879), .A1(n3901), .B0(n3979), .B1(n4890), .Y(n2810)
         );
  OAI22X1TS U6062 ( .A0(n4880), .A1(n3903), .B0(n3981), .B1(n4890), .Y(n2806)
         );
  OAI22X1TS U6063 ( .A0(n4880), .A1(n3905), .B0(n3983), .B1(n4891), .Y(n2802)
         );
  OAI22X1TS U6064 ( .A0(n4880), .A1(n3907), .B0(n3985), .B1(n4891), .Y(n2798)
         );
  OAI22X1TS U6065 ( .A0(n4880), .A1(n3909), .B0(n3987), .B1(n4887), .Y(n2794)
         );
  OAI22X1TS U6066 ( .A0(n4881), .A1(n3911), .B0(n3989), .B1(n4888), .Y(n2790)
         );
  OAI22X1TS U6067 ( .A0(n4881), .A1(n3913), .B0(n3991), .B1(n4899), .Y(n2786)
         );
  OAI22X1TS U6068 ( .A0(n4881), .A1(n3915), .B0(n3993), .B1(n4889), .Y(n2782)
         );
  OAI22X1TS U6069 ( .A0(n4881), .A1(n3917), .B0(n3995), .B1(n4895), .Y(n2778)
         );
  OAI22X1TS U6070 ( .A0(n4882), .A1(n3919), .B0(n3997), .B1(n4895), .Y(n2774)
         );
  OAI22X1TS U6071 ( .A0(n4882), .A1(n3921), .B0(n3999), .B1(n4890), .Y(n2770)
         );
  OAI22X1TS U6072 ( .A0(n4882), .A1(n3923), .B0(n4001), .B1(n4897), .Y(n2766)
         );
  OAI22X1TS U6073 ( .A0(n5003), .A1(n5839), .B0(n5872), .B1(n5012), .Y(n2561)
         );
  OAI22X1TS U6074 ( .A0(n5003), .A1(n5838), .B0(n5871), .B1(n5012), .Y(n2556)
         );
  OAI22X1TS U6075 ( .A0(n5003), .A1(n5837), .B0(n5870), .B1(n5013), .Y(n2552)
         );
  OAI22X1TS U6076 ( .A0(n5004), .A1(n5836), .B0(n5869), .B1(n5013), .Y(n2548)
         );
  OAI22X1TS U6077 ( .A0(n5004), .A1(n5835), .B0(n5868), .B1(n5014), .Y(n2544)
         );
  OAI22X1TS U6078 ( .A0(n5004), .A1(n5834), .B0(n5867), .B1(n5014), .Y(n2540)
         );
  OAI22X1TS U6079 ( .A0(n5004), .A1(n5833), .B0(n5866), .B1(n5015), .Y(n2536)
         );
  OAI22X1TS U6080 ( .A0(n5005), .A1(n5832), .B0(n5865), .B1(n5015), .Y(n2532)
         );
  OAI22X1TS U6081 ( .A0(n5005), .A1(n5831), .B0(n5864), .B1(n5016), .Y(n2528)
         );
  OAI22X1TS U6082 ( .A0(n5005), .A1(n5830), .B0(n5863), .B1(n5016), .Y(n2524)
         );
  OAI22X1TS U6083 ( .A0(n5005), .A1(n5829), .B0(n5862), .B1(n5002), .Y(n2520)
         );
  OAI22X1TS U6084 ( .A0(n5006), .A1(n5828), .B0(n5861), .B1(n5016), .Y(n2516)
         );
  OAI22X1TS U6085 ( .A0(n5006), .A1(n5827), .B0(n5860), .B1(n5012), .Y(n2512)
         );
  OAI22X1TS U6086 ( .A0(n5006), .A1(n5826), .B0(n5859), .B1(n5013), .Y(n2508)
         );
  OAI22X1TS U6087 ( .A0(n5006), .A1(n5825), .B0(n5858), .B1(n5017), .Y(n2504)
         );
  OAI22X1TS U6088 ( .A0(n5007), .A1(n5824), .B0(n5857), .B1(n5017), .Y(n2500)
         );
  OAI22X1TS U6089 ( .A0(n5007), .A1(n5823), .B0(n5856), .B1(n5023), .Y(n2496)
         );
  OAI22X1TS U6090 ( .A0(n5007), .A1(n5822), .B0(n5855), .B1(n5014), .Y(n2492)
         );
  NAND2X1TS U6091 ( .A(n5805), .B(n3152), .Y(totalAccesses[1]) );
  NAND4X1TS U6092 ( .A(n4561), .B(n4608), .C(n3721), .D(n1824), .Y(n1735) );
  NOR2X1TS U6093 ( .A(n3729), .B(n5561), .Y(n1824) );
  NOR2X1TS U6094 ( .A(n3747), .B(n2131), .Y(n2276) );
  CMPR32X2TS U6095 ( .A(totalAccesses[1]), .B(n5702), .C(
        \add_0_root_sub_0_root_sub_231/carry [1]), .CO(
        \add_0_root_sub_0_root_sub_231/carry [2]), .S(N606) );
  AND2X2TS U6096 ( .A(N615), .B(n3150), .Y(n3644) );
  XOR2X1TS U6097 ( .A(n4595), .B(n4531), .Y(N615) );
  INVX2TS U6098 ( .A(n1529), .Y(n5975) );
  CLKBUFX2TS U6099 ( .A(n1539), .Y(n5666) );
  CLKBUFX2TS U6100 ( .A(n1539), .Y(n5667) );
  CLKBUFX2TS U6101 ( .A(n1548), .Y(n5641) );
  NOR3BX1TS U6102 ( .AN(\r1472/carry[3] ), .B(N6316), .C(n4608), .Y(n2119) );
  NAND4X1TS U6103 ( .A(n5702), .B(n4565), .C(n2253), .D(\r1467/carry[3] ), .Y(
        n1776) );
  NOR2XLTS U6104 ( .A(N6316), .B(n2255), .Y(n2253) );
  OAI22X1TS U6105 ( .A0(n4705), .A1(n3158), .B0(n4719), .B1(n3159), .Y(N10076)
         );
  OAI22X1TS U6106 ( .A0(n5656), .A1(n3158), .B0(n5676), .B1(n3159), .Y(N10077)
         );
  OAI22X1TS U6107 ( .A0(n5641), .A1(n3158), .B0(n5650), .B1(n3159), .Y(N10078)
         );
  OAI22X1TS U6108 ( .A0(n4725), .A1(n3158), .B0(n5623), .B1(n3159), .Y(N10079)
         );
  NOR2X1TS U6109 ( .A(n3743), .B(n5731), .Y(n1555) );
  INVX2TS U6110 ( .A(n4581), .Y(n5976) );
  AND2X2TS U6111 ( .A(n4596), .B(totalAccesses[0]), .Y(n5979) );
  OR3X1TS U6112 ( .A(n4595), .B(N6318), .C(n4608), .Y(n2424) );
  CLKBUFX2TS U6113 ( .A(n3876), .Y(n5744) );
  CLKBUFX2TS U6114 ( .A(n4615), .Y(n5628) );
  CLKBUFX2TS U6115 ( .A(n3876), .Y(n5745) );
  CLKBUFX2TS U6116 ( .A(n4615), .Y(n5629) );
  CLKBUFX2TS U6117 ( .A(n3157), .Y(n4734) );
  AOI211X1TS U6118 ( .A0(n5782), .A1(n4599), .B0(n5790), .C0(n2213), .Y(n2210)
         );
  NOR3X1TS U6119 ( .A(n5708), .B(n4565), .C(n2214), .Y(n2213) );
  AOI211X1TS U6120 ( .A0(n5780), .A1(n3718), .B0(n5788), .C0(n2267), .Y(n2264)
         );
  NOR3X1TS U6121 ( .A(n5707), .B(n3680), .C(n5778), .Y(n2267) );
  CLKBUFX2TS U6122 ( .A(n5655), .Y(n5653) );
  CLKBUFX2TS U6123 ( .A(n5681), .Y(n5680) );
  CLKBUFX2TS U6124 ( .A(n5655), .Y(n5654) );
  CLKBUFX2TS U6125 ( .A(n1748), .Y(n4617) );
  CLKBUFX2TS U6126 ( .A(n5716), .Y(n5710) );
  CLKBUFX2TS U6127 ( .A(n5700), .Y(n5698) );
  NAND4X1TS U6128 ( .A(n5703), .B(n4565), .C(\r1470/carry[3] ), .D(n5785), .Y(
        n1780) );
  CLKBUFX2TS U6129 ( .A(n5717), .Y(n5709) );
  CLKBUFX2TS U6130 ( .A(n5717), .Y(n5707) );
  CLKBUFX2TS U6131 ( .A(n5716), .Y(n5711) );
  CLKBUFX2TS U6132 ( .A(n5701), .Y(n5696) );
  CLKBUFX2TS U6133 ( .A(n5708), .Y(n5712) );
  CLKBUFX2TS U6134 ( .A(n5715), .Y(n5714) );
  CLKBUFX2TS U6135 ( .A(n5700), .Y(n5699) );
  NOR2X1TS U6136 ( .A(n4611), .B(n4593), .Y(n1565) );
  NAND4X1TS U6137 ( .A(n5702), .B(n3680), .C(\r1467/carry[3] ), .D(n5794), .Y(
        n2246) );
  CLKBUFX2TS U6138 ( .A(n5717), .Y(n5708) );
  AND3X2TS U6139 ( .A(\r1470/carry[3] ), .B(n5708), .C(n4564), .Y(n2228) );
  INVX2TS U6140 ( .A(n1783), .Y(n5972) );
  CLKBUFX2TS U6141 ( .A(n880), .Y(n5694) );
  INVX2TS U6142 ( .A(n1740), .Y(n5973) );
  CLKBUFX2TS U6143 ( .A(n5701), .Y(n5697) );
  CLKBUFX2TS U6144 ( .A(n5709), .Y(n5715) );
  AND3X2TS U6145 ( .A(\r1471/carry[3] ), .B(n5712), .C(n4564), .Y(n2227) );
  AND3X2TS U6146 ( .A(\r1472/carry[3] ), .B(n5717), .C(n4565), .Y(n2225) );
  AO21X1TS U6147 ( .A0(n5697), .A1(n4595), .B0(n3806), .Y(n4614) );
  CLKBUFX2TS U6148 ( .A(n5714), .Y(n5713) );
  CLKBUFX2TS U6149 ( .A(n5695), .Y(n5691) );
  CLKBUFX2TS U6150 ( .A(n5695), .Y(n5692) );
  CLKBUFX2TS U6151 ( .A(n5691), .Y(n5693) );
  AOI22XLTS U6152 ( .A0(n4765), .A1(n3968), .B0(n3890), .B1(n4774), .Y(n3107)
         );
  AOI22XLTS U6153 ( .A0(n4765), .A1(n3970), .B0(n3892), .B1(n4781), .Y(n3103)
         );
  AOI22XLTS U6154 ( .A0(n4765), .A1(n3972), .B0(n3894), .B1(n4781), .Y(n3099)
         );
  AOI22XLTS U6155 ( .A0(n4765), .A1(n3974), .B0(n3896), .B1(n4784), .Y(n3095)
         );
  AOI22XLTS U6156 ( .A0(n4766), .A1(n3976), .B0(n3898), .B1(n4784), .Y(n3091)
         );
  AOI22XLTS U6157 ( .A0(n4766), .A1(n3978), .B0(n3900), .B1(n4782), .Y(n3087)
         );
  AOI22XLTS U6158 ( .A0(n4766), .A1(n3980), .B0(n3902), .B1(n4783), .Y(n3083)
         );
  AOI22XLTS U6159 ( .A0(n4766), .A1(n3982), .B0(n3904), .B1(n4784), .Y(n3079)
         );
  AOI22XLTS U6160 ( .A0(n4767), .A1(n3984), .B0(n3906), .B1(n4782), .Y(n3075)
         );
  AOI22XLTS U6161 ( .A0(n4767), .A1(n3986), .B0(n3908), .B1(n4775), .Y(n3071)
         );
  AOI22XLTS U6162 ( .A0(n4767), .A1(n3988), .B0(n3910), .B1(n4775), .Y(n3067)
         );
  AOI22XLTS U6163 ( .A0(n4767), .A1(n3990), .B0(n3912), .B1(n4775), .Y(n3063)
         );
  AOI22XLTS U6164 ( .A0(n4768), .A1(n3992), .B0(n3914), .B1(n4775), .Y(n3059)
         );
  AOI22XLTS U6165 ( .A0(n4768), .A1(n3994), .B0(n3916), .B1(n4776), .Y(n3055)
         );
  AOI22XLTS U6166 ( .A0(n4768), .A1(n3996), .B0(n3918), .B1(n4776), .Y(n3051)
         );
  AOI22XLTS U6167 ( .A0(n4768), .A1(n3998), .B0(n3920), .B1(n4776), .Y(n3047)
         );
  AOI22XLTS U6168 ( .A0(n4769), .A1(n4000), .B0(n3922), .B1(n4776), .Y(n3043)
         );
  AOI22XLTS U6169 ( .A0(n4769), .A1(n4002), .B0(n3924), .B1(n4777), .Y(n3039)
         );
  AOI22XLTS U6170 ( .A0(n4769), .A1(n4004), .B0(n3926), .B1(n4777), .Y(n3035)
         );
  AOI22XLTS U6171 ( .A0(n4769), .A1(n4006), .B0(n3928), .B1(n4777), .Y(n3031)
         );
  AOI22XLTS U6172 ( .A0(n4770), .A1(n4008), .B0(n3930), .B1(n4777), .Y(n3027)
         );
  AOI22XLTS U6173 ( .A0(n4770), .A1(n4010), .B0(n3932), .B1(n4778), .Y(n3023)
         );
  AOI22XLTS U6174 ( .A0(n4770), .A1(n4012), .B0(n3934), .B1(n4778), .Y(n3019)
         );
  AOI22XLTS U6175 ( .A0(n4770), .A1(n4014), .B0(n3936), .B1(n4778), .Y(n3015)
         );
  AOI22XLTS U6176 ( .A0(n4771), .A1(n4016), .B0(n3938), .B1(n4778), .Y(n3011)
         );
  AOI22XLTS U6177 ( .A0(n4771), .A1(n4018), .B0(n3940), .B1(n4779), .Y(n3007)
         );
  AOI22XLTS U6178 ( .A0(n4771), .A1(n4020), .B0(n3942), .B1(n4779), .Y(n3003)
         );
  AOI22XLTS U6179 ( .A0(n4771), .A1(n4022), .B0(n3944), .B1(n4779), .Y(n2999)
         );
  AOI22XLTS U6180 ( .A0(n4772), .A1(n4024), .B0(n3946), .B1(n4779), .Y(n2995)
         );
  AOI22XLTS U6181 ( .A0(n4772), .A1(n4026), .B0(n3948), .B1(n4780), .Y(n2991)
         );
  AOI22XLTS U6182 ( .A0(n4772), .A1(n4028), .B0(n3950), .B1(n4780), .Y(n2987)
         );
  OAI22X1TS U6183 ( .A0(n5875), .A1(n5136), .B0(n5133), .B1(n2982), .Y(n2979)
         );
  AOI22XLTS U6184 ( .A0(n4772), .A1(n4030), .B0(n3952), .B1(n4780), .Y(n2982)
         );
  OAI22X1TS U6185 ( .A0(n2971), .A1(n4847), .B0(n4664), .B1(n1039), .Y(n2970)
         );
  AOI22XLTS U6186 ( .A0(n2973), .A1(n5182), .B0(n5199), .B1(n4291), .Y(n2971)
         );
  OAI22X1TS U6187 ( .A0(n4992), .A1(n1039), .B0(n2695), .B1(n4989), .Y(n3513)
         );
  AOI221XLTS U6188 ( .A0(n5297), .A1(n4158), .B0(n4972), .B1(n4290), .C0(n2696), .Y(n2695) );
  OAI22X1TS U6189 ( .A0(n2697), .A1(n4962), .B0(n5283), .B1(n975), .Y(n2696)
         );
  AOI22XLTS U6190 ( .A0(n2699), .A1(n5260), .B0(n5276), .B1(n4292), .Y(n2697)
         );
  OAI22X1TS U6191 ( .A0(n5116), .A1(n975), .B0(n2416), .B1(n5106), .Y(n3449)
         );
  AOI221XLTS U6192 ( .A0(n5385), .A1(n4159), .B0(n5096), .B1(n4291), .C0(n2417), .Y(n2416) );
  OAI22X1TS U6193 ( .A0(n2418), .A1(n5086), .B0(n1167), .B1(n4679), .Y(n2417)
         );
  AOI22XLTS U6194 ( .A0(n2420), .A1(n5354), .B0(n5370), .B1(n4293), .Y(n2418)
         );
  AOI22XLTS U6195 ( .A0(n2968), .A1(n5182), .B0(n5199), .B1(n4296), .Y(n2967)
         );
  OAI22X1TS U6196 ( .A0(n4992), .A1(n1038), .B0(n2691), .B1(n4991), .Y(n3512)
         );
  AOI221XLTS U6197 ( .A0(n5297), .A1(n4162), .B0(n4972), .B1(n4295), .C0(n2692), .Y(n2691) );
  AOI22XLTS U6198 ( .A0(n2694), .A1(n5260), .B0(n5276), .B1(n4297), .Y(n2693)
         );
  OAI22X1TS U6199 ( .A0(n5116), .A1(n974), .B0(n2412), .B1(n5106), .Y(n3448)
         );
  AOI221XLTS U6200 ( .A0(n5382), .A1(n4163), .B0(n5096), .B1(n4296), .C0(n2413), .Y(n2412) );
  AOI22XLTS U6201 ( .A0(n2415), .A1(n5354), .B0(n5370), .B1(n4298), .Y(n2414)
         );
  OAI22X1TS U6202 ( .A0(n4868), .A1(n1101), .B0(n2961), .B1(n4858), .Y(n3575)
         );
  AOI22XLTS U6203 ( .A0(n2964), .A1(n5182), .B0(n5198), .B1(n4301), .Y(n2963)
         );
  OAI22X1TS U6204 ( .A0(n4992), .A1(n1037), .B0(n2687), .B1(n4991), .Y(n3511)
         );
  AOI221XLTS U6205 ( .A0(n5297), .A1(n4166), .B0(n4972), .B1(n4300), .C0(n2688), .Y(n2687) );
  AOI22XLTS U6206 ( .A0(n2690), .A1(n5260), .B0(n5275), .B1(n4302), .Y(n2689)
         );
  OAI22X1TS U6207 ( .A0(n5116), .A1(n973), .B0(n2408), .B1(n5106), .Y(n3447)
         );
  AOI221XLTS U6208 ( .A0(n5384), .A1(n4167), .B0(n5096), .B1(n4301), .C0(n2409), .Y(n2408) );
  AOI22XLTS U6209 ( .A0(n2411), .A1(n5354), .B0(n5369), .B1(n4303), .Y(n2410)
         );
  OAI22X1TS U6210 ( .A0(n4869), .A1(n1100), .B0(n2957), .B1(n4858), .Y(n3574)
         );
  AOI22XLTS U6211 ( .A0(n2960), .A1(n5182), .B0(n5198), .B1(n4306), .Y(n2959)
         );
  OAI22X1TS U6212 ( .A0(n4993), .A1(n1036), .B0(n2683), .B1(n4990), .Y(n3510)
         );
  AOI221XLTS U6213 ( .A0(n5297), .A1(n4170), .B0(n4972), .B1(n4305), .C0(n2684), .Y(n2683) );
  AOI22XLTS U6214 ( .A0(n2686), .A1(n5260), .B0(n5275), .B1(n4307), .Y(n2685)
         );
  OAI22X1TS U6215 ( .A0(n5117), .A1(n972), .B0(n2404), .B1(n5106), .Y(n3446)
         );
  AOI221XLTS U6216 ( .A0(n5385), .A1(n4171), .B0(n5096), .B1(n4306), .C0(n2405), .Y(n2404) );
  AOI22XLTS U6217 ( .A0(n2407), .A1(n5354), .B0(n5369), .B1(n4308), .Y(n2406)
         );
  OAI22X1TS U6218 ( .A0(n2955), .A1(n4838), .B0(n4669), .B1(n1035), .Y(n2954)
         );
  AOI22XLTS U6219 ( .A0(n2956), .A1(n5181), .B0(n5198), .B1(n4311), .Y(n2955)
         );
  OAI22X1TS U6220 ( .A0(n4993), .A1(n1035), .B0(n2679), .B1(n4982), .Y(n3509)
         );
  AOI221XLTS U6221 ( .A0(n5306), .A1(n4174), .B0(n4973), .B1(n4310), .C0(n2680), .Y(n2679) );
  OAI22X1TS U6222 ( .A0(n2681), .A1(n4963), .B0(n5290), .B1(n971), .Y(n2680)
         );
  AOI22XLTS U6223 ( .A0(n2682), .A1(n5259), .B0(n5275), .B1(n4312), .Y(n2681)
         );
  OAI22X1TS U6224 ( .A0(n5117), .A1(n971), .B0(n2400), .B1(n5115), .Y(n3445)
         );
  AOI221XLTS U6225 ( .A0(n5386), .A1(n4175), .B0(n5097), .B1(n4311), .C0(n2401), .Y(n2400) );
  OAI22X1TS U6226 ( .A0(n2402), .A1(n5087), .B0(n1163), .B1(n4688), .Y(n2401)
         );
  AOI22XLTS U6227 ( .A0(n2403), .A1(n5353), .B0(n5369), .B1(n4313), .Y(n2402)
         );
  OAI22X1TS U6228 ( .A0(n4869), .A1(n1098), .B0(n2949), .B1(n4865), .Y(n3572)
         );
  AOI221XLTS U6229 ( .A0(n2009), .A1(n4180), .B0(n4849), .B1(n4318), .C0(n2950), .Y(n2949) );
  AOI22XLTS U6230 ( .A0(n2952), .A1(n5181), .B0(n5198), .B1(n4316), .Y(n2951)
         );
  OAI22X1TS U6231 ( .A0(n4993), .A1(n1034), .B0(n2675), .B1(n4982), .Y(n3508)
         );
  AOI221XLTS U6232 ( .A0(n5308), .A1(n4178), .B0(n4973), .B1(n4315), .C0(n2676), .Y(n2675) );
  AOI22XLTS U6233 ( .A0(n2678), .A1(n5259), .B0(n5275), .B1(n4317), .Y(n2677)
         );
  OAI22X1TS U6234 ( .A0(n5117), .A1(n970), .B0(n2396), .B1(n5113), .Y(n3444)
         );
  AOI221XLTS U6235 ( .A0(n1831), .A1(n4179), .B0(n5097), .B1(n4316), .C0(n2397), .Y(n2396) );
  AOI22XLTS U6236 ( .A0(n2399), .A1(n5353), .B0(n5369), .B1(n4318), .Y(n2398)
         );
  OAI22X1TS U6237 ( .A0(n4869), .A1(n1097), .B0(n2945), .B1(n4867), .Y(n3571)
         );
  AOI221XLTS U6238 ( .A0(n5212), .A1(n4184), .B0(n4849), .B1(n4323), .C0(n2946), .Y(n2945) );
  AOI22XLTS U6239 ( .A0(n2948), .A1(n5181), .B0(n5197), .B1(n4321), .Y(n2947)
         );
  OAI22X1TS U6240 ( .A0(n4993), .A1(n1033), .B0(n2671), .B1(n4982), .Y(n3507)
         );
  AOI221XLTS U6241 ( .A0(n1920), .A1(n4182), .B0(n4973), .B1(n4320), .C0(n2672), .Y(n2671) );
  AOI22XLTS U6242 ( .A0(n2674), .A1(n5259), .B0(n5274), .B1(n4322), .Y(n2673)
         );
  OAI22X1TS U6243 ( .A0(n5117), .A1(n969), .B0(n2392), .B1(n5115), .Y(n3443)
         );
  AOI221XLTS U6244 ( .A0(n5384), .A1(n4183), .B0(n5097), .B1(n4321), .C0(n2393), .Y(n2392) );
  AOI22XLTS U6245 ( .A0(n2395), .A1(n5353), .B0(n5368), .B1(n4323), .Y(n2394)
         );
  OAI22X1TS U6246 ( .A0(n4870), .A1(n1096), .B0(n2941), .B1(n4865), .Y(n3570)
         );
  AOI221XLTS U6247 ( .A0(n5213), .A1(n4188), .B0(n4849), .B1(n4328), .C0(n2942), .Y(n2941) );
  AOI22XLTS U6248 ( .A0(n2944), .A1(n5181), .B0(n5197), .B1(n4326), .Y(n2943)
         );
  OAI22X1TS U6249 ( .A0(n4994), .A1(n1032), .B0(n2667), .B1(n4982), .Y(n3506)
         );
  AOI221XLTS U6250 ( .A0(n1920), .A1(n4186), .B0(n4973), .B1(n4325), .C0(n2668), .Y(n2667) );
  AOI22XLTS U6251 ( .A0(n2670), .A1(n5259), .B0(n5274), .B1(n4327), .Y(n2669)
         );
  OAI22X1TS U6252 ( .A0(n5118), .A1(n968), .B0(n2388), .B1(n5113), .Y(n3442)
         );
  AOI221XLTS U6253 ( .A0(n1831), .A1(n4187), .B0(n5097), .B1(n4326), .C0(n2389), .Y(n2388) );
  AOI22XLTS U6254 ( .A0(n2391), .A1(n5353), .B0(n5368), .B1(n4328), .Y(n2390)
         );
  OAI22X1TS U6255 ( .A0(n4870), .A1(n1095), .B0(n2937), .B1(n4859), .Y(n3569)
         );
  AOI221XLTS U6256 ( .A0(n5210), .A1(n4192), .B0(n4856), .B1(n4333), .C0(n2938), .Y(n2937) );
  OAI22X1TS U6257 ( .A0(n2939), .A1(n4839), .B0(n4668), .B1(n1031), .Y(n2938)
         );
  AOI22XLTS U6258 ( .A0(n2940), .A1(n5180), .B0(n5190), .B1(n4331), .Y(n2939)
         );
  OAI22X1TS U6259 ( .A0(n4994), .A1(n1031), .B0(n2663), .B1(n4983), .Y(n3505)
         );
  AOI221XLTS U6260 ( .A0(n5305), .A1(n4190), .B0(n4974), .B1(n4330), .C0(n2664), .Y(n2663) );
  OAI22X1TS U6261 ( .A0(n2665), .A1(n4964), .B0(n5289), .B1(n967), .Y(n2664)
         );
  AOI22XLTS U6262 ( .A0(n2666), .A1(n5258), .B0(n5265), .B1(n4332), .Y(n2665)
         );
  OAI22X1TS U6263 ( .A0(n5118), .A1(n967), .B0(n2384), .B1(n5107), .Y(n3441)
         );
  AOI221XLTS U6264 ( .A0(n5383), .A1(n4191), .B0(n5104), .B1(n4331), .C0(n2385), .Y(n2384) );
  OAI22X1TS U6265 ( .A0(n2386), .A1(n5092), .B0(n1159), .B1(n4685), .Y(n2385)
         );
  AOI22XLTS U6266 ( .A0(n2387), .A1(n5352), .B0(n5359), .B1(n4333), .Y(n2386)
         );
  OAI22X1TS U6267 ( .A0(n4870), .A1(n1094), .B0(n2933), .B1(n4859), .Y(n3568)
         );
  AOI221XLTS U6268 ( .A0(n5210), .A1(n4196), .B0(n4856), .B1(n4338), .C0(n2934), .Y(n2933) );
  AOI22XLTS U6269 ( .A0(n2936), .A1(n5179), .B0(n5190), .B1(n4336), .Y(n2935)
         );
  OAI22X1TS U6270 ( .A0(n4994), .A1(n1030), .B0(n2659), .B1(n4983), .Y(n3504)
         );
  AOI221XLTS U6271 ( .A0(n5302), .A1(n4194), .B0(n4974), .B1(n4335), .C0(n2660), .Y(n2659) );
  AOI22XLTS U6272 ( .A0(n2662), .A1(n5257), .B0(n5265), .B1(n4337), .Y(n2661)
         );
  OAI22X1TS U6273 ( .A0(n5118), .A1(n966), .B0(n2380), .B1(n5107), .Y(n3440)
         );
  AOI221XLTS U6274 ( .A0(n5386), .A1(n4195), .B0(n5104), .B1(n4336), .C0(n2381), .Y(n2380) );
  AOI22XLTS U6275 ( .A0(n2383), .A1(n5351), .B0(n5359), .B1(n4338), .Y(n2382)
         );
  OAI22X1TS U6276 ( .A0(n4870), .A1(n1093), .B0(n2929), .B1(n4859), .Y(n3567)
         );
  AOI221XLTS U6277 ( .A0(n5214), .A1(n4200), .B0(n4854), .B1(n4343), .C0(n2930), .Y(n2929) );
  AOI22XLTS U6278 ( .A0(n2932), .A1(n5180), .B0(n5191), .B1(n4341), .Y(n2931)
         );
  OAI22X1TS U6279 ( .A0(n4994), .A1(n1029), .B0(n2655), .B1(n4983), .Y(n3503)
         );
  AOI221XLTS U6280 ( .A0(n5308), .A1(n4198), .B0(n4974), .B1(n4340), .C0(n2656), .Y(n2655) );
  AOI22XLTS U6281 ( .A0(n2658), .A1(n5258), .B0(n5266), .B1(n4342), .Y(n2657)
         );
  OAI22X1TS U6282 ( .A0(n5118), .A1(n965), .B0(n2376), .B1(n5107), .Y(n3439)
         );
  AOI221XLTS U6283 ( .A0(n5383), .A1(n4199), .B0(n5102), .B1(n4341), .C0(n2377), .Y(n2376) );
  AOI22XLTS U6284 ( .A0(n2379), .A1(n5352), .B0(n5360), .B1(n4343), .Y(n2378)
         );
  OAI22X1TS U6285 ( .A0(n4875), .A1(n1092), .B0(n2925), .B1(n4859), .Y(n3566)
         );
  AOI221XLTS U6286 ( .A0(n5212), .A1(n4204), .B0(n4854), .B1(n4348), .C0(n2926), .Y(n2925) );
  AOI22XLTS U6287 ( .A0(n2928), .A1(n5180), .B0(n5191), .B1(n4346), .Y(n2927)
         );
  OAI22X1TS U6288 ( .A0(n4995), .A1(n1028), .B0(n2651), .B1(n4983), .Y(n3502)
         );
  AOI221XLTS U6289 ( .A0(n5306), .A1(n4202), .B0(n4974), .B1(n4345), .C0(n2652), .Y(n2651) );
  AOI22XLTS U6290 ( .A0(n2654), .A1(n5258), .B0(n5266), .B1(n4347), .Y(n2653)
         );
  OAI22X1TS U6291 ( .A0(n5119), .A1(n964), .B0(n2372), .B1(n5107), .Y(n3438)
         );
  AOI221XLTS U6292 ( .A0(n5385), .A1(n4203), .B0(n5102), .B1(n4346), .C0(n2373), .Y(n2372) );
  AOI22XLTS U6293 ( .A0(n2375), .A1(n5352), .B0(n5360), .B1(n4348), .Y(n2374)
         );
  OAI22X1TS U6294 ( .A0(n4877), .A1(n1091), .B0(n2921), .B1(n4860), .Y(n3565)
         );
  AOI221XLTS U6295 ( .A0(n5203), .A1(n4208), .B0(n4856), .B1(n4353), .C0(n2922), .Y(n2921) );
  OAI22X1TS U6296 ( .A0(n2923), .A1(n4840), .B0(n4667), .B1(n1027), .Y(n2922)
         );
  AOI22XLTS U6297 ( .A0(n2924), .A1(n5180), .B0(n5192), .B1(n4351), .Y(n2923)
         );
  OAI22X1TS U6298 ( .A0(n4995), .A1(n1027), .B0(n2647), .B1(n4984), .Y(n3501)
         );
  AOI221XLTS U6299 ( .A0(n5305), .A1(n4206), .B0(n4975), .B1(n4350), .C0(n2648), .Y(n2647) );
  OAI22X1TS U6300 ( .A0(n2649), .A1(n4965), .B0(n5288), .B1(n963), .Y(n2648)
         );
  AOI22XLTS U6301 ( .A0(n2650), .A1(n5258), .B0(n5267), .B1(n4352), .Y(n2649)
         );
  OAI22X1TS U6302 ( .A0(n5119), .A1(n963), .B0(n2368), .B1(n5108), .Y(n3437)
         );
  AOI221XLTS U6303 ( .A0(n5375), .A1(n4207), .B0(n5104), .B1(n4351), .C0(n2369), .Y(n2368) );
  OAI22X1TS U6304 ( .A0(n2370), .A1(n5093), .B0(n1155), .B1(n4684), .Y(n2369)
         );
  AOI22XLTS U6305 ( .A0(n2371), .A1(n5352), .B0(n5361), .B1(n4353), .Y(n2370)
         );
  AOI221XLTS U6306 ( .A0(n5203), .A1(n4212), .B0(n4856), .B1(n4358), .C0(n2918), .Y(n2917) );
  AOI22XLTS U6307 ( .A0(n2920), .A1(n5179), .B0(n5192), .B1(n4356), .Y(n2919)
         );
  OAI22X1TS U6308 ( .A0(n4995), .A1(n1026), .B0(n2643), .B1(n4984), .Y(n3500)
         );
  AOI221XLTS U6309 ( .A0(n5305), .A1(n4210), .B0(n4975), .B1(n4355), .C0(n2644), .Y(n2643) );
  AOI22XLTS U6310 ( .A0(n2646), .A1(n5257), .B0(n5267), .B1(n4357), .Y(n2645)
         );
  OAI22X1TS U6311 ( .A0(n5119), .A1(n962), .B0(n2364), .B1(n5108), .Y(n3436)
         );
  AOI221XLTS U6312 ( .A0(n5375), .A1(n4211), .B0(n5104), .B1(n4356), .C0(n2365), .Y(n2364) );
  AOI22XLTS U6313 ( .A0(n2367), .A1(n5351), .B0(n5361), .B1(n4358), .Y(n2366)
         );
  OAI22X1TS U6314 ( .A0(n4877), .A1(n1089), .B0(n2913), .B1(n4860), .Y(n3563)
         );
  AOI221XLTS U6315 ( .A0(n5203), .A1(n4216), .B0(n4857), .B1(n4363), .C0(n2914), .Y(n2913) );
  AOI22XLTS U6316 ( .A0(n2916), .A1(n5179), .B0(n5193), .B1(n4361), .Y(n2915)
         );
  OAI22X1TS U6317 ( .A0(n4995), .A1(n1025), .B0(n2639), .B1(n4984), .Y(n3499)
         );
  AOI221XLTS U6318 ( .A0(n5306), .A1(n4214), .B0(n4975), .B1(n4360), .C0(n2640), .Y(n2639) );
  AOI22XLTS U6319 ( .A0(n2642), .A1(n5257), .B0(n5268), .B1(n4362), .Y(n2641)
         );
  OAI22X1TS U6320 ( .A0(n5119), .A1(n961), .B0(n2360), .B1(n5108), .Y(n3435)
         );
  AOI221XLTS U6321 ( .A0(n5375), .A1(n4215), .B0(n5105), .B1(n4361), .C0(n2361), .Y(n2360) );
  AOI22XLTS U6322 ( .A0(n2363), .A1(n5351), .B0(n5362), .B1(n4363), .Y(n2362)
         );
  OAI22X1TS U6323 ( .A0(n4876), .A1(n1088), .B0(n2909), .B1(n4860), .Y(n3562)
         );
  AOI221XLTS U6324 ( .A0(n5203), .A1(n4220), .B0(n4855), .B1(n4368), .C0(n2910), .Y(n2909) );
  AOI22XLTS U6325 ( .A0(n2912), .A1(n5179), .B0(n5193), .B1(n4366), .Y(n2911)
         );
  OAI22X1TS U6326 ( .A0(n4999), .A1(n1024), .B0(n2635), .B1(n4984), .Y(n3498)
         );
  AOI221XLTS U6327 ( .A0(n5305), .A1(n4218), .B0(n4975), .B1(n4365), .C0(n2636), .Y(n2635) );
  AOI22XLTS U6328 ( .A0(n2638), .A1(n5257), .B0(n5268), .B1(n4367), .Y(n2637)
         );
  OAI22X1TS U6329 ( .A0(n5123), .A1(n960), .B0(n2356), .B1(n5108), .Y(n3434)
         );
  AOI221XLTS U6330 ( .A0(n5375), .A1(n4219), .B0(n5103), .B1(n4366), .C0(n2357), .Y(n2356) );
  AOI22XLTS U6331 ( .A0(n2359), .A1(n5351), .B0(n5362), .B1(n4368), .Y(n2358)
         );
  OAI22X1TS U6332 ( .A0(n4875), .A1(n1087), .B0(n2905), .B1(n4861), .Y(n3561)
         );
  AOI221XLTS U6333 ( .A0(n5204), .A1(n4224), .B0(n4850), .B1(n4373), .C0(n2906), .Y(n2905) );
  OAI22X1TS U6334 ( .A0(n2907), .A1(n4841), .B0(n4666), .B1(n1023), .Y(n2906)
         );
  AOI22XLTS U6335 ( .A0(n2908), .A1(n5185), .B0(n5194), .B1(n4371), .Y(n2907)
         );
  OAI22X1TS U6336 ( .A0(n5001), .A1(n1023), .B0(n2631), .B1(n4985), .Y(n3497)
         );
  AOI221XLTS U6337 ( .A0(n5304), .A1(n4222), .B0(n4976), .B1(n4370), .C0(n2632), .Y(n2631) );
  OAI22X1TS U6338 ( .A0(n2633), .A1(n4969), .B0(n5287), .B1(n959), .Y(n2632)
         );
  AOI22XLTS U6339 ( .A0(n2634), .A1(n5256), .B0(n5269), .B1(n4372), .Y(n2633)
         );
  OAI22X1TS U6340 ( .A0(n5125), .A1(n959), .B0(n2352), .B1(n5109), .Y(n3433)
         );
  AOI221XLTS U6341 ( .A0(n5376), .A1(n4223), .B0(n5098), .B1(n4371), .C0(n2353), .Y(n2352) );
  OAI22X1TS U6342 ( .A0(n2354), .A1(n5088), .B0(n1151), .B1(n4683), .Y(n2353)
         );
  AOI22XLTS U6343 ( .A0(n2355), .A1(n5357), .B0(n5363), .B1(n4373), .Y(n2354)
         );
  AOI22XLTS U6344 ( .A0(n2904), .A1(n5185), .B0(n5199), .B1(n4376), .Y(n2903)
         );
  OAI22X1TS U6345 ( .A0(n2566), .A1(n1022), .B0(n2627), .B1(n4985), .Y(n3496)
         );
  AOI221XLTS U6346 ( .A0(n5304), .A1(n4226), .B0(n4976), .B1(n4375), .C0(n2628), .Y(n2627) );
  AOI22XLTS U6347 ( .A0(n2630), .A1(n5256), .B0(n5269), .B1(n4377), .Y(n2629)
         );
  OAI22X1TS U6348 ( .A0(n2287), .A1(n958), .B0(n2348), .B1(n5109), .Y(n3432)
         );
  AOI221XLTS U6349 ( .A0(n5376), .A1(n4227), .B0(n5098), .B1(n4376), .C0(n2349), .Y(n2348) );
  AOI22XLTS U6350 ( .A0(n2351), .A1(n5357), .B0(n5363), .B1(n4378), .Y(n2350)
         );
  OAI22X1TS U6351 ( .A0(n4874), .A1(n1085), .B0(n2897), .B1(n4861), .Y(n3559)
         );
  AOI221XLTS U6352 ( .A0(n5204), .A1(n4232), .B0(n4850), .B1(n4383), .C0(n2898), .Y(n2897) );
  AOI22XLTS U6353 ( .A0(n2900), .A1(n2012), .B0(n5191), .B1(n4381), .Y(n2899)
         );
  OAI22X1TS U6354 ( .A0(n5001), .A1(n1021), .B0(n2623), .B1(n4985), .Y(n3495)
         );
  AOI221XLTS U6355 ( .A0(n5307), .A1(n4230), .B0(n4976), .B1(n4380), .C0(n2624), .Y(n2623) );
  AOI22XLTS U6356 ( .A0(n2626), .A1(n5256), .B0(n5270), .B1(n4382), .Y(n2625)
         );
  OAI22X1TS U6357 ( .A0(n5125), .A1(n957), .B0(n2344), .B1(n5109), .Y(n3431)
         );
  AOI221XLTS U6358 ( .A0(n5376), .A1(n4231), .B0(n5098), .B1(n4381), .C0(n2345), .Y(n2344) );
  AOI22XLTS U6359 ( .A0(n2347), .A1(n1834), .B0(n5364), .B1(n4383), .Y(n2346)
         );
  OAI22X1TS U6360 ( .A0(n4871), .A1(n1084), .B0(n2893), .B1(n4861), .Y(n3558)
         );
  AOI221XLTS U6361 ( .A0(n5204), .A1(n4236), .B0(n4850), .B1(n4388), .C0(n2894), .Y(n2893) );
  AOI22XLTS U6362 ( .A0(n2896), .A1(n2012), .B0(n5189), .B1(n4386), .Y(n2895)
         );
  OAI22X1TS U6363 ( .A0(n5000), .A1(n1020), .B0(n2619), .B1(n4985), .Y(n3494)
         );
  AOI221XLTS U6364 ( .A0(n5302), .A1(n4234), .B0(n4976), .B1(n4385), .C0(n2620), .Y(n2619) );
  AOI22XLTS U6365 ( .A0(n2622), .A1(n5256), .B0(n5270), .B1(n4387), .Y(n2621)
         );
  OAI22X1TS U6366 ( .A0(n5124), .A1(n956), .B0(n2340), .B1(n5109), .Y(n3430)
         );
  AOI221XLTS U6367 ( .A0(n5376), .A1(n4235), .B0(n5098), .B1(n4386), .C0(n2341), .Y(n2340) );
  AOI22XLTS U6368 ( .A0(n2343), .A1(n1834), .B0(n5364), .B1(n4388), .Y(n2342)
         );
  OAI22X1TS U6369 ( .A0(n4871), .A1(n1083), .B0(n2889), .B1(n4862), .Y(n3557)
         );
  AOI221XLTS U6370 ( .A0(n5205), .A1(n4240), .B0(n4851), .B1(n4393), .C0(n2890), .Y(n2889) );
  OAI22X1TS U6371 ( .A0(n2891), .A1(n4842), .B0(n4665), .B1(n1019), .Y(n2890)
         );
  AOI22XLTS U6372 ( .A0(n2892), .A1(n5178), .B0(n5194), .B1(n4391), .Y(n2891)
         );
  OAI22X1TS U6373 ( .A0(n4998), .A1(n1019), .B0(n2615), .B1(n4986), .Y(n3493)
         );
  AOI221XLTS U6374 ( .A0(n5303), .A1(n4238), .B0(n4979), .B1(n4390), .C0(n2616), .Y(n2615) );
  OAI22X1TS U6375 ( .A0(n2617), .A1(n4966), .B0(n5286), .B1(n955), .Y(n2616)
         );
  AOI22XLTS U6376 ( .A0(n2618), .A1(n5255), .B0(n5271), .B1(n4392), .Y(n2617)
         );
  OAI22X1TS U6377 ( .A0(n5122), .A1(n955), .B0(n2336), .B1(n5110), .Y(n3429)
         );
  AOI221XLTS U6378 ( .A0(n5377), .A1(n4239), .B0(n5099), .B1(n4391), .C0(n2337), .Y(n2336) );
  OAI22X1TS U6379 ( .A0(n2338), .A1(n5089), .B0(n1147), .B1(n4682), .Y(n2337)
         );
  AOI22XLTS U6380 ( .A0(n2339), .A1(n5350), .B0(n5365), .B1(n4393), .Y(n2338)
         );
  OAI22X1TS U6381 ( .A0(n4871), .A1(n1082), .B0(n2885), .B1(n4862), .Y(n3556)
         );
  AOI221XLTS U6382 ( .A0(n5205), .A1(n4244), .B0(n4851), .B1(n4398), .C0(n2886), .Y(n2885) );
  AOI22XLTS U6383 ( .A0(n2888), .A1(n5178), .B0(n5194), .B1(n4396), .Y(n2887)
         );
  OAI22X1TS U6384 ( .A0(n4998), .A1(n1018), .B0(n2611), .B1(n4986), .Y(n3492)
         );
  AOI221XLTS U6385 ( .A0(n5304), .A1(n4242), .B0(n4979), .B1(n4395), .C0(n2612), .Y(n2611) );
  AOI22XLTS U6386 ( .A0(n2614), .A1(n5255), .B0(n5271), .B1(n4397), .Y(n2613)
         );
  OAI22X1TS U6387 ( .A0(n5122), .A1(n954), .B0(n2332), .B1(n5110), .Y(n3428)
         );
  AOI221XLTS U6388 ( .A0(n5377), .A1(n4243), .B0(n5099), .B1(n4396), .C0(n2333), .Y(n2332) );
  AOI22XLTS U6389 ( .A0(n2335), .A1(n5350), .B0(n5365), .B1(n4398), .Y(n2334)
         );
  OAI22X1TS U6390 ( .A0(n4871), .A1(n1081), .B0(n2881), .B1(n4862), .Y(n3555)
         );
  AOI221XLTS U6391 ( .A0(n5205), .A1(n4248), .B0(n4851), .B1(n4403), .C0(n2882), .Y(n2881) );
  AOI22XLTS U6392 ( .A0(n2884), .A1(n5178), .B0(n5195), .B1(n4401), .Y(n2883)
         );
  OAI22X1TS U6393 ( .A0(n4998), .A1(n1017), .B0(n2607), .B1(n4986), .Y(n3491)
         );
  AOI221XLTS U6394 ( .A0(n5303), .A1(n4246), .B0(n4979), .B1(n4400), .C0(n2608), .Y(n2607) );
  AOI22XLTS U6395 ( .A0(n2610), .A1(n5255), .B0(n5272), .B1(n4402), .Y(n2609)
         );
  OAI22X1TS U6396 ( .A0(n5122), .A1(n953), .B0(n2328), .B1(n5110), .Y(n3427)
         );
  AOI221XLTS U6397 ( .A0(n5377), .A1(n4247), .B0(n5099), .B1(n4401), .C0(n2329), .Y(n2328) );
  AOI22XLTS U6398 ( .A0(n2331), .A1(n5350), .B0(n5366), .B1(n4403), .Y(n2330)
         );
  OAI22X1TS U6399 ( .A0(n4872), .A1(n1080), .B0(n2877), .B1(n4862), .Y(n3554)
         );
  AOI221XLTS U6400 ( .A0(n5205), .A1(n4252), .B0(n4851), .B1(n4408), .C0(n2878), .Y(n2877) );
  AOI22XLTS U6401 ( .A0(n2880), .A1(n5178), .B0(n5195), .B1(n4406), .Y(n2879)
         );
  OAI22X1TS U6402 ( .A0(n4996), .A1(n1016), .B0(n2603), .B1(n4986), .Y(n3490)
         );
  AOI221XLTS U6403 ( .A0(n5304), .A1(n4250), .B0(n4981), .B1(n4405), .C0(n2604), .Y(n2603) );
  AOI22XLTS U6404 ( .A0(n2606), .A1(n5255), .B0(n5272), .B1(n4407), .Y(n2605)
         );
  OAI22X1TS U6405 ( .A0(n5120), .A1(n952), .B0(n2324), .B1(n5110), .Y(n3426)
         );
  AOI221XLTS U6406 ( .A0(n5377), .A1(n4251), .B0(n5099), .B1(n4406), .C0(n2325), .Y(n2324) );
  AOI22XLTS U6407 ( .A0(n2327), .A1(n5350), .B0(n5366), .B1(n4408), .Y(n2326)
         );
  OAI22X1TS U6408 ( .A0(n4872), .A1(n1079), .B0(n2873), .B1(n4863), .Y(n3553)
         );
  AOI221XLTS U6409 ( .A0(n5206), .A1(n4256), .B0(n4852), .B1(n4413), .C0(n2874), .Y(n2873) );
  OAI22X1TS U6410 ( .A0(n2875), .A1(n4843), .B0(n5972), .B1(n1015), .Y(n2874)
         );
  AOI22XLTS U6411 ( .A0(n2876), .A1(n5177), .B0(n5195), .B1(n4411), .Y(n2875)
         );
  OAI22X1TS U6412 ( .A0(n4996), .A1(n1015), .B0(n2599), .B1(n4987), .Y(n3489)
         );
  AOI221XLTS U6413 ( .A0(n5298), .A1(n4254), .B0(n4977), .B1(n4410), .C0(n2600), .Y(n2599) );
  OAI22X1TS U6414 ( .A0(n2601), .A1(n4967), .B0(n5285), .B1(n951), .Y(n2600)
         );
  AOI22XLTS U6415 ( .A0(n2602), .A1(n5254), .B0(n5272), .B1(n4412), .Y(n2601)
         );
  OAI22X1TS U6416 ( .A0(n5120), .A1(n951), .B0(n2320), .B1(n5111), .Y(n3425)
         );
  AOI221XLTS U6417 ( .A0(n5378), .A1(n4255), .B0(n5100), .B1(n4411), .C0(n2321), .Y(n2320) );
  OAI22X1TS U6418 ( .A0(n2322), .A1(n5090), .B0(n1143), .B1(n4681), .Y(n2321)
         );
  AOI22XLTS U6419 ( .A0(n2323), .A1(n5349), .B0(n5366), .B1(n4413), .Y(n2322)
         );
  OAI22X1TS U6420 ( .A0(n4872), .A1(n1078), .B0(n2869), .B1(n4863), .Y(n3552)
         );
  AOI221XLTS U6421 ( .A0(n5206), .A1(n4260), .B0(n4852), .B1(n4418), .C0(n2870), .Y(n2869) );
  AOI22XLTS U6422 ( .A0(n2872), .A1(n5177), .B0(n5195), .B1(n4416), .Y(n2871)
         );
  OAI22X1TS U6423 ( .A0(n4996), .A1(n1014), .B0(n2595), .B1(n4987), .Y(n3488)
         );
  AOI221XLTS U6424 ( .A0(n5298), .A1(n4258), .B0(n4977), .B1(n4415), .C0(n2596), .Y(n2595) );
  AOI22XLTS U6425 ( .A0(n2598), .A1(n5254), .B0(n5272), .B1(n4417), .Y(n2597)
         );
  OAI22X1TS U6426 ( .A0(n5120), .A1(n950), .B0(n2316), .B1(n5111), .Y(n3424)
         );
  AOI221XLTS U6427 ( .A0(n5378), .A1(n4259), .B0(n5100), .B1(n4416), .C0(n2317), .Y(n2316) );
  AOI22XLTS U6428 ( .A0(n2319), .A1(n5349), .B0(n5366), .B1(n4418), .Y(n2318)
         );
  OAI22X1TS U6429 ( .A0(n4872), .A1(n1077), .B0(n2865), .B1(n4863), .Y(n3551)
         );
  AOI221XLTS U6430 ( .A0(n5206), .A1(n4264), .B0(n4852), .B1(n4423), .C0(n2866), .Y(n2865) );
  AOI22XLTS U6431 ( .A0(n2868), .A1(n5177), .B0(n5196), .B1(n4421), .Y(n2867)
         );
  OAI22X1TS U6432 ( .A0(n4996), .A1(n1013), .B0(n2591), .B1(n4987), .Y(n3487)
         );
  AOI221XLTS U6433 ( .A0(n5298), .A1(n4262), .B0(n4977), .B1(n4420), .C0(n2592), .Y(n2591) );
  AOI22XLTS U6434 ( .A0(n2594), .A1(n5254), .B0(n5273), .B1(n4422), .Y(n2593)
         );
  OAI22X1TS U6435 ( .A0(n5120), .A1(n949), .B0(n2312), .B1(n5111), .Y(n3423)
         );
  AOI221XLTS U6436 ( .A0(n5378), .A1(n4263), .B0(n5100), .B1(n4421), .C0(n2313), .Y(n2312) );
  AOI22XLTS U6437 ( .A0(n2315), .A1(n5349), .B0(n5367), .B1(n4423), .Y(n2314)
         );
  OAI22X1TS U6438 ( .A0(n4873), .A1(n1076), .B0(n2861), .B1(n4863), .Y(n3550)
         );
  AOI221XLTS U6439 ( .A0(n5206), .A1(n4268), .B0(n4852), .B1(n4428), .C0(n2862), .Y(n2861) );
  AOI22XLTS U6440 ( .A0(n2864), .A1(n5177), .B0(n5196), .B1(n4426), .Y(n2863)
         );
  OAI22X1TS U6441 ( .A0(n4997), .A1(n1012), .B0(n2587), .B1(n4987), .Y(n3486)
         );
  AOI221XLTS U6442 ( .A0(n5298), .A1(n4266), .B0(n4977), .B1(n4425), .C0(n2588), .Y(n2587) );
  AOI22XLTS U6443 ( .A0(n2590), .A1(n5254), .B0(n5273), .B1(n4427), .Y(n2589)
         );
  OAI22X1TS U6444 ( .A0(n5121), .A1(n948), .B0(n2308), .B1(n5111), .Y(n3422)
         );
  AOI221XLTS U6445 ( .A0(n5378), .A1(n4267), .B0(n5100), .B1(n4426), .C0(n2309), .Y(n2308) );
  AOI22XLTS U6446 ( .A0(n2311), .A1(n5349), .B0(n5367), .B1(n4428), .Y(n2310)
         );
  OAI22X1TS U6447 ( .A0(n2859), .A1(n4844), .B0(n4670), .B1(n1011), .Y(n2858)
         );
  AOI22XLTS U6448 ( .A0(n2860), .A1(n5176), .B0(n5196), .B1(n4431), .Y(n2859)
         );
  OAI22X1TS U6449 ( .A0(n4997), .A1(n1011), .B0(n2583), .B1(n4988), .Y(n3485)
         );
  AOI221XLTS U6450 ( .A0(n5299), .A1(n4270), .B0(n4978), .B1(n4430), .C0(n2584), .Y(n2583) );
  OAI22X1TS U6451 ( .A0(n2585), .A1(n4968), .B0(n5284), .B1(n947), .Y(n2584)
         );
  AOI22XLTS U6452 ( .A0(n2586), .A1(n5263), .B0(n5273), .B1(n4432), .Y(n2585)
         );
  OAI22X1TS U6453 ( .A0(n5121), .A1(n947), .B0(n2304), .B1(n5112), .Y(n3421)
         );
  AOI221XLTS U6454 ( .A0(n5379), .A1(n4271), .B0(n5101), .B1(n4431), .C0(n2305), .Y(n2304) );
  OAI22X1TS U6455 ( .A0(n2306), .A1(n5091), .B0(n1139), .B1(n4680), .Y(n2305)
         );
  AOI22XLTS U6456 ( .A0(n2307), .A1(n5348), .B0(n5367), .B1(n4433), .Y(n2306)
         );
  OAI22X1TS U6457 ( .A0(n4873), .A1(n1074), .B0(n2853), .B1(n4864), .Y(n3548)
         );
  AOI221XLTS U6458 ( .A0(n5207), .A1(n4276), .B0(n4853), .B1(n4438), .C0(n2854), .Y(n2853) );
  AOI22XLTS U6459 ( .A0(n2856), .A1(n5176), .B0(n5196), .B1(n4436), .Y(n2855)
         );
  OAI22X1TS U6460 ( .A0(n4997), .A1(n1010), .B0(n2579), .B1(n4988), .Y(n3484)
         );
  AOI221XLTS U6461 ( .A0(n5299), .A1(n4274), .B0(n4978), .B1(n4435), .C0(n2580), .Y(n2579) );
  AOI22XLTS U6462 ( .A0(n2582), .A1(n1924), .B0(n5273), .B1(n4437), .Y(n2581)
         );
  OAI22X1TS U6463 ( .A0(n5121), .A1(n946), .B0(n2300), .B1(n5112), .Y(n3420)
         );
  AOI221XLTS U6464 ( .A0(n5379), .A1(n4275), .B0(n5101), .B1(n4436), .C0(n2301), .Y(n2300) );
  AOI22XLTS U6465 ( .A0(n2303), .A1(n5348), .B0(n5367), .B1(n4438), .Y(n2302)
         );
  OAI22X1TS U6466 ( .A0(n4873), .A1(n1073), .B0(n2849), .B1(n4864), .Y(n3547)
         );
  AOI221XLTS U6467 ( .A0(n5207), .A1(n4280), .B0(n4853), .B1(n4443), .C0(n2850), .Y(n2849) );
  AOI22XLTS U6468 ( .A0(n2852), .A1(n5176), .B0(n5197), .B1(n4441), .Y(n2851)
         );
  OAI22X1TS U6469 ( .A0(n4997), .A1(n1009), .B0(n2575), .B1(n4988), .Y(n3483)
         );
  AOI221XLTS U6470 ( .A0(n5299), .A1(n4278), .B0(n4978), .B1(n4440), .C0(n2576), .Y(n2575) );
  AOI22XLTS U6471 ( .A0(n2578), .A1(n1924), .B0(n5274), .B1(n4442), .Y(n2577)
         );
  OAI22X1TS U6472 ( .A0(n5121), .A1(n945), .B0(n2296), .B1(n5112), .Y(n3419)
         );
  AOI221XLTS U6473 ( .A0(n5379), .A1(n4279), .B0(n5101), .B1(n4441), .C0(n2297), .Y(n2296) );
  AOI22XLTS U6474 ( .A0(n2299), .A1(n5348), .B0(n5368), .B1(n4443), .Y(n2298)
         );
  OAI22X1TS U6475 ( .A0(n4876), .A1(n1072), .B0(n2841), .B1(n4864), .Y(n3546)
         );
  AOI221XLTS U6476 ( .A0(n5207), .A1(n4284), .B0(n4853), .B1(n4448), .C0(n2844), .Y(n2841) );
  OAI22X1TS U6477 ( .A0(n5000), .A1(n1008), .B0(n2567), .B1(n4988), .Y(n3482)
         );
  AOI221XLTS U6478 ( .A0(n5299), .A1(n4282), .B0(n4978), .B1(n4445), .C0(n2570), .Y(n2567) );
  OAI22X1TS U6479 ( .A0(n5124), .A1(n944), .B0(n2288), .B1(n5112), .Y(n3418)
         );
  AOI221XLTS U6480 ( .A0(n5379), .A1(n4283), .B0(n5101), .B1(n4446), .C0(n2291), .Y(n2288) );
  AOI221XLTS U6481 ( .A0(n5242), .A1(n4158), .B0(n4910), .B1(n4293), .C0(n2832), .Y(n2831) );
  OAI22X1TS U6482 ( .A0(n2833), .A1(n4900), .B0(n5690), .B1(n1007), .Y(n2832)
         );
  AOI22XLTS U6483 ( .A0(n2835), .A1(n5221), .B0(n5237), .B1(n4291), .Y(n2833)
         );
  AOI221XLTS U6484 ( .A0(n5242), .A1(n4162), .B0(n4910), .B1(n4298), .C0(n2828), .Y(n2827) );
  OAI22X1TS U6485 ( .A0(n2829), .A1(n4900), .B0(n5690), .B1(n1006), .Y(n2828)
         );
  AOI22XLTS U6486 ( .A0(n2830), .A1(n5221), .B0(n5237), .B1(n4296), .Y(n2829)
         );
  AOI221XLTS U6487 ( .A0(n5242), .A1(n4166), .B0(n4910), .B1(n4303), .C0(n2824), .Y(n2823) );
  OAI22X1TS U6488 ( .A0(n2825), .A1(n4900), .B0(n5689), .B1(n1005), .Y(n2824)
         );
  AOI22XLTS U6489 ( .A0(n2826), .A1(n5221), .B0(n5236), .B1(n4301), .Y(n2825)
         );
  AOI221XLTS U6490 ( .A0(n5242), .A1(n4170), .B0(n4910), .B1(n4308), .C0(n2820), .Y(n2819) );
  OAI22X1TS U6491 ( .A0(n2821), .A1(n4900), .B0(n5688), .B1(n1004), .Y(n2820)
         );
  AOI22XLTS U6492 ( .A0(n2822), .A1(n5221), .B0(n5236), .B1(n4306), .Y(n2821)
         );
  AOI221XLTS U6493 ( .A0(n5243), .A1(n4174), .B0(n4911), .B1(n4313), .C0(n2816), .Y(n2815) );
  OAI22X1TS U6494 ( .A0(n2817), .A1(n4901), .B0(n5689), .B1(n1003), .Y(n2816)
         );
  AOI22XLTS U6495 ( .A0(n2818), .A1(n5220), .B0(n5236), .B1(n4311), .Y(n2817)
         );
  AOI221XLTS U6496 ( .A0(n5243), .A1(n4178), .B0(n4911), .B1(n4318), .C0(n2812), .Y(n2811) );
  OAI22X1TS U6497 ( .A0(n2813), .A1(n4901), .B0(n5689), .B1(n1002), .Y(n2812)
         );
  AOI22XLTS U6498 ( .A0(n2814), .A1(n5220), .B0(n5236), .B1(n4316), .Y(n2813)
         );
  AOI221XLTS U6499 ( .A0(n5243), .A1(n4182), .B0(n4911), .B1(n4323), .C0(n2808), .Y(n2807) );
  OAI22X1TS U6500 ( .A0(n2809), .A1(n4901), .B0(n5689), .B1(n1001), .Y(n2808)
         );
  AOI22XLTS U6501 ( .A0(n2810), .A1(n5220), .B0(n5235), .B1(n4321), .Y(n2809)
         );
  AOI221XLTS U6502 ( .A0(n5243), .A1(n4186), .B0(n4911), .B1(n4328), .C0(n2804), .Y(n2803) );
  OAI22X1TS U6503 ( .A0(n2805), .A1(n4901), .B0(n5688), .B1(n1000), .Y(n2804)
         );
  AOI22XLTS U6504 ( .A0(n2806), .A1(n5220), .B0(n5235), .B1(n4326), .Y(n2805)
         );
  AOI221XLTS U6505 ( .A0(n5244), .A1(n4190), .B0(n4912), .B1(n4333), .C0(n2800), .Y(n2799) );
  OAI22X1TS U6506 ( .A0(n2801), .A1(n4908), .B0(n5685), .B1(n999), .Y(n2800)
         );
  AOI22XLTS U6507 ( .A0(n2802), .A1(n5219), .B0(n5226), .B1(n4331), .Y(n2801)
         );
  AOI221XLTS U6508 ( .A0(n5244), .A1(n4194), .B0(n4912), .B1(n4338), .C0(n2796), .Y(n2795) );
  OAI22X1TS U6509 ( .A0(n2797), .A1(n4909), .B0(n5688), .B1(n998), .Y(n2796)
         );
  AOI22XLTS U6510 ( .A0(n2798), .A1(n5218), .B0(n5226), .B1(n4336), .Y(n2797)
         );
  AOI221XLTS U6511 ( .A0(n5244), .A1(n4198), .B0(n4912), .B1(n4343), .C0(n2792), .Y(n2791) );
  OAI22X1TS U6512 ( .A0(n2793), .A1(n4908), .B0(n5688), .B1(n997), .Y(n2792)
         );
  AOI22XLTS U6513 ( .A0(n2794), .A1(n5219), .B0(n5227), .B1(n4341), .Y(n2793)
         );
  AOI221XLTS U6514 ( .A0(n5244), .A1(n4202), .B0(n4912), .B1(n4348), .C0(n2788), .Y(n2787) );
  OAI22X1TS U6515 ( .A0(n2789), .A1(n4907), .B0(n5687), .B1(n996), .Y(n2788)
         );
  AOI22XLTS U6516 ( .A0(n2790), .A1(n5219), .B0(n5227), .B1(n4346), .Y(n2789)
         );
  AOI221XLTS U6517 ( .A0(n5245), .A1(n4206), .B0(n4913), .B1(n4353), .C0(n2784), .Y(n2783) );
  OAI22X1TS U6518 ( .A0(n2785), .A1(n4902), .B0(n5687), .B1(n995), .Y(n2784)
         );
  AOI22XLTS U6519 ( .A0(n2786), .A1(n5219), .B0(n5228), .B1(n4351), .Y(n2785)
         );
  AOI221XLTS U6520 ( .A0(n5245), .A1(n4210), .B0(n4913), .B1(n4358), .C0(n2780), .Y(n2779) );
  OAI22X1TS U6521 ( .A0(n2781), .A1(n4902), .B0(n5687), .B1(n994), .Y(n2780)
         );
  AOI22XLTS U6522 ( .A0(n2782), .A1(n5218), .B0(n5228), .B1(n4356), .Y(n2781)
         );
  AOI221XLTS U6523 ( .A0(n5245), .A1(n4214), .B0(n4913), .B1(n4363), .C0(n2776), .Y(n2775) );
  OAI22X1TS U6524 ( .A0(n2777), .A1(n4902), .B0(n5687), .B1(n993), .Y(n2776)
         );
  AOI22XLTS U6525 ( .A0(n2778), .A1(n5218), .B0(n5229), .B1(n4361), .Y(n2777)
         );
  AOI221XLTS U6526 ( .A0(n5245), .A1(n4218), .B0(n4913), .B1(n4368), .C0(n2772), .Y(n2771) );
  OAI22X1TS U6527 ( .A0(n2773), .A1(n4902), .B0(n5686), .B1(n992), .Y(n2772)
         );
  AOI22XLTS U6528 ( .A0(n2774), .A1(n5218), .B0(n5229), .B1(n4366), .Y(n2773)
         );
  AOI221XLTS U6529 ( .A0(n5246), .A1(n4222), .B0(n4917), .B1(n4373), .C0(n2768), .Y(n2767) );
  OAI22X1TS U6530 ( .A0(n2769), .A1(n4903), .B0(n5686), .B1(n991), .Y(n2768)
         );
  AOI22XLTS U6531 ( .A0(n2770), .A1(n5224), .B0(n5230), .B1(n4371), .Y(n2769)
         );
  AOI221XLTS U6532 ( .A0(n5246), .A1(n4226), .B0(n4919), .B1(n4378), .C0(n2764), .Y(n2763) );
  OAI22X1TS U6533 ( .A0(n2765), .A1(n4903), .B0(n5686), .B1(n990), .Y(n2764)
         );
  AOI22XLTS U6534 ( .A0(n2766), .A1(n5224), .B0(n5230), .B1(n4376), .Y(n2765)
         );
  AOI221XLTS U6535 ( .A0(n5246), .A1(n4230), .B0(n4919), .B1(n4383), .C0(n2760), .Y(n2759) );
  OAI22X1TS U6536 ( .A0(n2761), .A1(n4903), .B0(n5686), .B1(n989), .Y(n2760)
         );
  AOI22XLTS U6537 ( .A0(n2762), .A1(n1968), .B0(n5231), .B1(n4381), .Y(n2761)
         );
  AOI221XLTS U6538 ( .A0(n5246), .A1(n4234), .B0(n4918), .B1(n4388), .C0(n2756), .Y(n2755) );
  OAI22X1TS U6539 ( .A0(n2757), .A1(n4903), .B0(n5685), .B1(n988), .Y(n2756)
         );
  AOI22XLTS U6540 ( .A0(n2758), .A1(n1968), .B0(n5231), .B1(n4386), .Y(n2757)
         );
  AOI221XLTS U6541 ( .A0(n5247), .A1(n4238), .B0(n4914), .B1(n4393), .C0(n2752), .Y(n2751) );
  OAI22X1TS U6542 ( .A0(n2753), .A1(n4904), .B0(n5685), .B1(n987), .Y(n2752)
         );
  AOI22XLTS U6543 ( .A0(n2754), .A1(n5217), .B0(n5232), .B1(n4391), .Y(n2753)
         );
  AOI221XLTS U6544 ( .A0(n5247), .A1(n4242), .B0(n4914), .B1(n4398), .C0(n2748), .Y(n2747) );
  OAI22X1TS U6545 ( .A0(n2749), .A1(n4904), .B0(n5685), .B1(n986), .Y(n2748)
         );
  AOI22XLTS U6546 ( .A0(n2750), .A1(n5217), .B0(n5232), .B1(n4396), .Y(n2749)
         );
  AOI221XLTS U6547 ( .A0(n5247), .A1(n4246), .B0(n4914), .B1(n4403), .C0(n2744), .Y(n2743) );
  OAI22X1TS U6548 ( .A0(n2745), .A1(n4904), .B0(n5684), .B1(n985), .Y(n2744)
         );
  AOI22XLTS U6549 ( .A0(n2746), .A1(n5217), .B0(n5233), .B1(n4401), .Y(n2745)
         );
  AOI221XLTS U6550 ( .A0(n5247), .A1(n4250), .B0(n4914), .B1(n4408), .C0(n2740), .Y(n2739) );
  OAI22X1TS U6551 ( .A0(n2741), .A1(n4904), .B0(n5684), .B1(n984), .Y(n2740)
         );
  AOI22XLTS U6552 ( .A0(n2742), .A1(n5217), .B0(n5233), .B1(n4406), .Y(n2741)
         );
  AOI221XLTS U6553 ( .A0(n5253), .A1(n4254), .B0(n4915), .B1(n4413), .C0(n2736), .Y(n2735) );
  OAI22X1TS U6554 ( .A0(n2737), .A1(n4905), .B0(n5684), .B1(n983), .Y(n2736)
         );
  AOI22XLTS U6555 ( .A0(n2738), .A1(n5216), .B0(n5233), .B1(n4411), .Y(n2737)
         );
  AOI221XLTS U6556 ( .A0(n5249), .A1(n4258), .B0(n4915), .B1(n4418), .C0(n2732), .Y(n2731) );
  OAI22X1TS U6557 ( .A0(n2733), .A1(n4905), .B0(n5684), .B1(n982), .Y(n2732)
         );
  AOI22XLTS U6558 ( .A0(n2734), .A1(n5216), .B0(n5233), .B1(n4416), .Y(n2733)
         );
  AOI221XLTS U6559 ( .A0(n5251), .A1(n4262), .B0(n4915), .B1(n4423), .C0(n2728), .Y(n2727) );
  OAI22X1TS U6560 ( .A0(n2729), .A1(n4905), .B0(n5692), .B1(n981), .Y(n2728)
         );
  AOI22XLTS U6561 ( .A0(n2730), .A1(n5216), .B0(n5234), .B1(n4421), .Y(n2729)
         );
  AOI221XLTS U6562 ( .A0(n5252), .A1(n4266), .B0(n4915), .B1(n4428), .C0(n2724), .Y(n2723) );
  OAI22X1TS U6563 ( .A0(n2725), .A1(n4905), .B0(n880), .B1(n980), .Y(n2724) );
  AOI22XLTS U6564 ( .A0(n2726), .A1(n5216), .B0(n5234), .B1(n4426), .Y(n2725)
         );
  AOI221XLTS U6565 ( .A0(n5248), .A1(n4270), .B0(n4916), .B1(n4433), .C0(n2720), .Y(n2719) );
  OAI22X1TS U6566 ( .A0(n2721), .A1(n4906), .B0(n880), .B1(n979), .Y(n2720) );
  AOI22XLTS U6567 ( .A0(n2722), .A1(n5215), .B0(n5234), .B1(n4431), .Y(n2721)
         );
  AOI221XLTS U6568 ( .A0(n5248), .A1(n4274), .B0(n4916), .B1(n4438), .C0(n2716), .Y(n2715) );
  OAI22X1TS U6569 ( .A0(n2717), .A1(n4906), .B0(n5694), .B1(n978), .Y(n2716)
         );
  AOI22XLTS U6570 ( .A0(n2718), .A1(n5215), .B0(n5234), .B1(n4436), .Y(n2717)
         );
  AOI221XLTS U6571 ( .A0(n5248), .A1(n4278), .B0(n4916), .B1(n4443), .C0(n2712), .Y(n2711) );
  OAI22X1TS U6572 ( .A0(n2713), .A1(n4906), .B0(n5692), .B1(n977), .Y(n2712)
         );
  AOI22XLTS U6573 ( .A0(n2714), .A1(n5215), .B0(n5235), .B1(n4441), .Y(n2713)
         );
  AOI221XLTS U6574 ( .A0(n5248), .A1(n4282), .B0(n4916), .B1(n4448), .C0(n2706), .Y(n2703) );
  OAI22X1TS U6575 ( .A0(n2707), .A1(n4906), .B0(n5693), .B1(n976), .Y(n2706)
         );
  AOI221XLTS U6576 ( .A0(n5336), .A1(n4160), .B0(n5034), .B1(n4292), .C0(n2558), .Y(n2557) );
  OAI22X1TS U6577 ( .A0(n2559), .A1(n5024), .B0(n4700), .B1(n943), .Y(n2558)
         );
  AOI22XLTS U6578 ( .A0(n2561), .A1(n5315), .B0(n5331), .B1(n4290), .Y(n2559)
         );
  AOI221XLTS U6579 ( .A0(n5336), .A1(n4164), .B0(n5034), .B1(n4297), .C0(n2554), .Y(n2553) );
  OAI22X1TS U6580 ( .A0(n2555), .A1(n5024), .B0(n4695), .B1(n942), .Y(n2554)
         );
  AOI22XLTS U6581 ( .A0(n2556), .A1(n5315), .B0(n5331), .B1(n4295), .Y(n2555)
         );
  AOI221XLTS U6582 ( .A0(n5336), .A1(n4168), .B0(n5034), .B1(n4302), .C0(n2550), .Y(n2549) );
  OAI22X1TS U6583 ( .A0(n2551), .A1(n5024), .B0(n4697), .B1(n941), .Y(n2550)
         );
  AOI22XLTS U6584 ( .A0(n2552), .A1(n5315), .B0(n5330), .B1(n4300), .Y(n2551)
         );
  AOI221XLTS U6585 ( .A0(n5336), .A1(n4172), .B0(n5034), .B1(n4307), .C0(n2546), .Y(n2545) );
  OAI22X1TS U6586 ( .A0(n2547), .A1(n5024), .B0(n4697), .B1(n940), .Y(n2546)
         );
  AOI22XLTS U6587 ( .A0(n2548), .A1(n5315), .B0(n5330), .B1(n4305), .Y(n2547)
         );
  AOI221XLTS U6588 ( .A0(n5337), .A1(n4176), .B0(n5035), .B1(n4312), .C0(n2542), .Y(n2541) );
  OAI22X1TS U6589 ( .A0(n2543), .A1(n5025), .B0(n4696), .B1(n939), .Y(n2542)
         );
  AOI22XLTS U6590 ( .A0(n2544), .A1(n5314), .B0(n5330), .B1(n4310), .Y(n2543)
         );
  AOI221XLTS U6591 ( .A0(n5337), .A1(n4180), .B0(n5035), .B1(n4317), .C0(n2538), .Y(n2537) );
  OAI22X1TS U6592 ( .A0(n2539), .A1(n5025), .B0(n4695), .B1(n938), .Y(n2538)
         );
  AOI22XLTS U6593 ( .A0(n2540), .A1(n5314), .B0(n5330), .B1(n4315), .Y(n2539)
         );
  AOI221XLTS U6594 ( .A0(n5337), .A1(n4184), .B0(n5035), .B1(n4322), .C0(n2534), .Y(n2533) );
  OAI22X1TS U6595 ( .A0(n2535), .A1(n5025), .B0(n4696), .B1(n937), .Y(n2534)
         );
  AOI22XLTS U6596 ( .A0(n2536), .A1(n5314), .B0(n5329), .B1(n4320), .Y(n2535)
         );
  AOI221XLTS U6597 ( .A0(n5337), .A1(n4188), .B0(n5035), .B1(n4327), .C0(n2530), .Y(n2529) );
  OAI22X1TS U6598 ( .A0(n2531), .A1(n5025), .B0(n4696), .B1(n936), .Y(n2530)
         );
  AOI22XLTS U6599 ( .A0(n2532), .A1(n5314), .B0(n5329), .B1(n4325), .Y(n2531)
         );
  AOI221XLTS U6600 ( .A0(n5346), .A1(n4192), .B0(n5036), .B1(n4332), .C0(n2526), .Y(n2525) );
  OAI22X1TS U6601 ( .A0(n2527), .A1(n5026), .B0(n4696), .B1(n935), .Y(n2526)
         );
  AOI22XLTS U6602 ( .A0(n2528), .A1(n5313), .B0(n5320), .B1(n4330), .Y(n2527)
         );
  AOI221XLTS U6603 ( .A0(n5347), .A1(n4196), .B0(n5036), .B1(n4337), .C0(n2522), .Y(n2521) );
  OAI22X1TS U6604 ( .A0(n2523), .A1(n5026), .B0(n4692), .B1(n934), .Y(n2522)
         );
  AOI22XLTS U6605 ( .A0(n2524), .A1(n5312), .B0(n5320), .B1(n4335), .Y(n2523)
         );
  AOI221XLTS U6606 ( .A0(n5345), .A1(n4200), .B0(n5036), .B1(n4342), .C0(n2518), .Y(n2517) );
  OAI22X1TS U6607 ( .A0(n2519), .A1(n5026), .B0(n4695), .B1(n933), .Y(n2518)
         );
  AOI22XLTS U6608 ( .A0(n2520), .A1(n5313), .B0(n5321), .B1(n4340), .Y(n2519)
         );
  AOI221XLTS U6609 ( .A0(n5345), .A1(n4204), .B0(n5036), .B1(n4347), .C0(n2514), .Y(n2513) );
  OAI22X1TS U6610 ( .A0(n2515), .A1(n5026), .B0(n4695), .B1(n932), .Y(n2514)
         );
  AOI22XLTS U6611 ( .A0(n2516), .A1(n5313), .B0(n5321), .B1(n4345), .Y(n2515)
         );
  AOI221XLTS U6612 ( .A0(n5338), .A1(n4208), .B0(n5037), .B1(n4352), .C0(n2510), .Y(n2509) );
  OAI22X1TS U6613 ( .A0(n2511), .A1(n5027), .B0(n4694), .B1(n931), .Y(n2510)
         );
  AOI22XLTS U6614 ( .A0(n2512), .A1(n5313), .B0(n5322), .B1(n4350), .Y(n2511)
         );
  AOI221XLTS U6615 ( .A0(n5338), .A1(n4212), .B0(n5037), .B1(n4357), .C0(n2506), .Y(n2505) );
  OAI22X1TS U6616 ( .A0(n2507), .A1(n5027), .B0(n4694), .B1(n930), .Y(n2506)
         );
  AOI22XLTS U6617 ( .A0(n2508), .A1(n5312), .B0(n5322), .B1(n4355), .Y(n2507)
         );
  AOI221XLTS U6618 ( .A0(n5338), .A1(n4216), .B0(n5037), .B1(n4362), .C0(n2502), .Y(n2501) );
  OAI22X1TS U6619 ( .A0(n2503), .A1(n5027), .B0(n4694), .B1(n929), .Y(n2502)
         );
  AOI22XLTS U6620 ( .A0(n2504), .A1(n5312), .B0(n5323), .B1(n4360), .Y(n2503)
         );
  AOI221XLTS U6621 ( .A0(n5338), .A1(n4220), .B0(n5037), .B1(n4367), .C0(n2498), .Y(n2497) );
  OAI22X1TS U6622 ( .A0(n2499), .A1(n5027), .B0(n4694), .B1(n928), .Y(n2498)
         );
  AOI22XLTS U6623 ( .A0(n2500), .A1(n5312), .B0(n5323), .B1(n4365), .Y(n2499)
         );
  AOI221XLTS U6624 ( .A0(n5339), .A1(n4224), .B0(n5038), .B1(n4372), .C0(n2494), .Y(n2493) );
  OAI22X1TS U6625 ( .A0(n2495), .A1(n5028), .B0(n4693), .B1(n927), .Y(n2494)
         );
  AOI22XLTS U6626 ( .A0(n2496), .A1(n5311), .B0(n5324), .B1(n4370), .Y(n2495)
         );
  AOI221XLTS U6627 ( .A0(n5339), .A1(n4228), .B0(n5038), .B1(n4377), .C0(n2490), .Y(n2489) );
  OAI22X1TS U6628 ( .A0(n2491), .A1(n5028), .B0(n4693), .B1(n926), .Y(n2490)
         );
  AOI22XLTS U6629 ( .A0(n2492), .A1(n5311), .B0(n5324), .B1(n4375), .Y(n2491)
         );
  AOI221XLTS U6630 ( .A0(n5339), .A1(n4232), .B0(n5038), .B1(n4382), .C0(n2486), .Y(n2485) );
  OAI22X1TS U6631 ( .A0(n2487), .A1(n5028), .B0(n4693), .B1(n925), .Y(n2486)
         );
  AOI22XLTS U6632 ( .A0(n2488), .A1(n5311), .B0(n5325), .B1(n4380), .Y(n2487)
         );
  AOI221XLTS U6633 ( .A0(n5339), .A1(n4236), .B0(n5038), .B1(n4387), .C0(n2482), .Y(n2481) );
  OAI22X1TS U6634 ( .A0(n2483), .A1(n5028), .B0(n4693), .B1(n924), .Y(n2482)
         );
  AOI22XLTS U6635 ( .A0(n2484), .A1(n5311), .B0(n5325), .B1(n4385), .Y(n2483)
         );
  AOI221XLTS U6636 ( .A0(n5340), .A1(n4240), .B0(n5041), .B1(n4392), .C0(n2478), .Y(n2477) );
  OAI22X1TS U6637 ( .A0(n2479), .A1(n5029), .B0(n4692), .B1(n923), .Y(n2478)
         );
  AOI22XLTS U6638 ( .A0(n2480), .A1(n5310), .B0(n5326), .B1(n4390), .Y(n2479)
         );
  AOI221XLTS U6639 ( .A0(n5340), .A1(n4244), .B0(n5041), .B1(n4397), .C0(n2474), .Y(n2473) );
  OAI22X1TS U6640 ( .A0(n2475), .A1(n5029), .B0(n4692), .B1(n922), .Y(n2474)
         );
  AOI22XLTS U6641 ( .A0(n2476), .A1(n5310), .B0(n5326), .B1(n4395), .Y(n2475)
         );
  AOI221XLTS U6642 ( .A0(n5340), .A1(n4248), .B0(n5041), .B1(n4402), .C0(n2470), .Y(n2469) );
  OAI22X1TS U6643 ( .A0(n2471), .A1(n5029), .B0(n4692), .B1(n921), .Y(n2470)
         );
  AOI22XLTS U6644 ( .A0(n2472), .A1(n5310), .B0(n5327), .B1(n4400), .Y(n2471)
         );
  AOI221XLTS U6645 ( .A0(n5340), .A1(n4252), .B0(n5043), .B1(n4407), .C0(n2466), .Y(n2465) );
  OAI22X1TS U6646 ( .A0(n2467), .A1(n5029), .B0(n4701), .B1(n920), .Y(n2466)
         );
  AOI22XLTS U6647 ( .A0(n2468), .A1(n5310), .B0(n5327), .B1(n4405), .Y(n2467)
         );
  AOI221XLTS U6648 ( .A0(n5341), .A1(n4256), .B0(n5039), .B1(n4412), .C0(n2462), .Y(n2461) );
  OAI22X1TS U6649 ( .A0(n2463), .A1(n5031), .B0(n4702), .B1(n919), .Y(n2462)
         );
  AOI22XLTS U6650 ( .A0(n2464), .A1(n5309), .B0(n5327), .B1(n4410), .Y(n2463)
         );
  AOI221XLTS U6651 ( .A0(n5341), .A1(n4260), .B0(n5039), .B1(n4417), .C0(n2458), .Y(n2457) );
  OAI22X1TS U6652 ( .A0(n2459), .A1(n5032), .B0(n4702), .B1(n918), .Y(n2458)
         );
  AOI22XLTS U6653 ( .A0(n2460), .A1(n5309), .B0(n5327), .B1(n4415), .Y(n2459)
         );
  AOI221XLTS U6654 ( .A0(n5341), .A1(n4264), .B0(n5039), .B1(n4422), .C0(n2454), .Y(n2453) );
  OAI22X1TS U6655 ( .A0(n2455), .A1(n5031), .B0(n4702), .B1(n917), .Y(n2454)
         );
  AOI22XLTS U6656 ( .A0(n2456), .A1(n5309), .B0(n5328), .B1(n4420), .Y(n2455)
         );
  AOI221XLTS U6657 ( .A0(n5341), .A1(n4268), .B0(n5039), .B1(n4427), .C0(n2450), .Y(n2449) );
  OAI22X1TS U6658 ( .A0(n2451), .A1(n5033), .B0(n4701), .B1(n916), .Y(n2450)
         );
  AOI22XLTS U6659 ( .A0(n2452), .A1(n5309), .B0(n5328), .B1(n4425), .Y(n2451)
         );
  AOI221XLTS U6660 ( .A0(n5342), .A1(n4272), .B0(n5040), .B1(n4432), .C0(n2446), .Y(n2445) );
  OAI22X1TS U6661 ( .A0(n2447), .A1(n5030), .B0(n4698), .B1(n915), .Y(n2446)
         );
  AOI22XLTS U6662 ( .A0(n2448), .A1(n5318), .B0(n5328), .B1(n4430), .Y(n2447)
         );
  AOI221XLTS U6663 ( .A0(n5342), .A1(n4276), .B0(n5040), .B1(n4437), .C0(n2442), .Y(n2441) );
  OAI22X1TS U6664 ( .A0(n2443), .A1(n5030), .B0(n4703), .B1(n914), .Y(n2442)
         );
  AOI22XLTS U6665 ( .A0(n2444), .A1(n1879), .B0(n5328), .B1(n4435), .Y(n2443)
         );
  AOI221XLTS U6666 ( .A0(n5342), .A1(n4280), .B0(n5040), .B1(n4442), .C0(n2438), .Y(n2437) );
  OAI22X1TS U6667 ( .A0(n2439), .A1(n5030), .B0(n4703), .B1(n913), .Y(n2438)
         );
  AOI22XLTS U6668 ( .A0(n2440), .A1(n1879), .B0(n5329), .B1(n4440), .Y(n2439)
         );
  AOI221XLTS U6669 ( .A0(n5342), .A1(n4284), .B0(n5040), .B1(n4447), .C0(n2432), .Y(n2429) );
  OAI22X1TS U6670 ( .A0(n2433), .A1(n5030), .B0(n4701), .B1(n912), .Y(n2432)
         );
  OAI22X1TS U6671 ( .A0(n1284), .A1(n1588), .B0(n1589), .B1(n1590), .Y(n3191)
         );
  AOI222XLTS U6672 ( .A0(n4061), .A1(n5570), .B0(n4060), .B1(n3865), .C0(n4622), .C1(n4032), .Y(n1589) );
  OAI22X1TS U6673 ( .A0(n1283), .A1(n1588), .B0(n1592), .B1(n1590), .Y(n3192)
         );
  AOI222XLTS U6674 ( .A0(n4064), .A1(n5572), .B0(n4063), .B1(n3864), .C0(n4622), .C1(n4034), .Y(n1592) );
  OAI22X1TS U6675 ( .A0(n1282), .A1(n4533), .B0(n1593), .B1(n1590), .Y(n3193)
         );
  AOI222XLTS U6676 ( .A0(n4067), .A1(n5573), .B0(n4066), .B1(n3866), .C0(n4623), .C1(n4036), .Y(n1593) );
  OAI22X1TS U6677 ( .A0(n1281), .A1(n4533), .B0(n1594), .B1(n4524), .Y(n3194)
         );
  AOI222XLTS U6678 ( .A0(n4070), .A1(n5574), .B0(n4069), .B1(n3863), .C0(n4622), .C1(n4038), .Y(n1594) );
  OAI22X1TS U6679 ( .A0(n1280), .A1(n4533), .B0(n1595), .B1(n4524), .Y(n3195)
         );
  AOI222XLTS U6680 ( .A0(n4073), .A1(n5571), .B0(n4072), .B1(n3865), .C0(n4623), .C1(n4040), .Y(n1595) );
  OAI22X1TS U6681 ( .A0(n1279), .A1(n4533), .B0(n1596), .B1(n4524), .Y(n3196)
         );
  AOI222XLTS U6682 ( .A0(n4076), .A1(n5572), .B0(n4075), .B1(n3866), .C0(n4623), .C1(n4042), .Y(n1596) );
  OAI22X1TS U6683 ( .A0(n4517), .A1(n1224), .B0(n2039), .B1(n4574), .Y(n3325)
         );
  AOI221XLTS U6684 ( .A0(n3759), .A1(n2040), .B0(n5208), .B1(n4126), .C0(n2041), .Y(n2039) );
  OAI22X1TS U6685 ( .A0(n3833), .A1(n5183), .B0(n5189), .B1(n2042), .Y(n2040)
         );
  OAI22X1TS U6686 ( .A0(n4672), .A1(n1208), .B0(n3778), .B1(n3832), .Y(n2041)
         );
  OAI22X1TS U6687 ( .A0(n4529), .A1(n1208), .B0(n1951), .B1(n4556), .Y(n3309)
         );
  AOI221XLTS U6688 ( .A0(n3757), .A1(n1952), .B0(n5300), .B1(n4128), .C0(n1953), .Y(n1951) );
  OAI22X1TS U6689 ( .A0(n3834), .A1(n5261), .B0(n5276), .B1(n1954), .Y(n1952)
         );
  OAI22X1TS U6690 ( .A0(n5282), .A1(n1192), .B0(n3780), .B1(n3833), .Y(n1953)
         );
  OAI22X1TS U6691 ( .A0(n4515), .A1(n1192), .B0(n1861), .B1(n4572), .Y(n3293)
         );
  AOI221XLTS U6692 ( .A0(n3761), .A1(n1862), .B0(n5380), .B1(n4126), .C0(n1863), .Y(n1861) );
  OAI22X1TS U6693 ( .A0(n3833), .A1(n5355), .B0(n5364), .B1(n1864), .Y(n1862)
         );
  OAI22X1TS U6694 ( .A0(n1240), .A1(n4587), .B0(n2100), .B1(n4554), .Y(n3341)
         );
  AOI222XLTS U6695 ( .A0(\addressToWriteBuffer[2][0] ), .A1(n5571), .B0(n4044), 
        .B1(n3865), .C0(n4127), .C1(n4625), .Y(n2100) );
  OAI22X1TS U6696 ( .A0(n4518), .A1(n1223), .B0(n2035), .B1(n4574), .Y(n3324)
         );
  AOI221XLTS U6697 ( .A0(n3760), .A1(n2036), .B0(n5208), .B1(n4130), .C0(n2037), .Y(n2035) );
  OAI22X1TS U6698 ( .A0(n3837), .A1(n5183), .B0(n5189), .B1(n2038), .Y(n2036)
         );
  OAI22X1TS U6699 ( .A0(n4674), .A1(n1207), .B0(n3779), .B1(n3836), .Y(n2037)
         );
  OAI22X1TS U6700 ( .A0(n4528), .A1(n1207), .B0(n1947), .B1(n4556), .Y(n3308)
         );
  AOI221XLTS U6701 ( .A0(n3758), .A1(n1948), .B0(n5300), .B1(n4132), .C0(n1949), .Y(n1947) );
  OAI22X1TS U6702 ( .A0(n3838), .A1(n5261), .B0(n5276), .B1(n1950), .Y(n1948)
         );
  OAI22X1TS U6703 ( .A0(n5282), .A1(n1191), .B0(n3781), .B1(n3837), .Y(n1949)
         );
  OAI22X1TS U6704 ( .A0(n4516), .A1(n1191), .B0(n1857), .B1(n4572), .Y(n3292)
         );
  AOI221XLTS U6705 ( .A0(n3762), .A1(n1858), .B0(n5380), .B1(n4130), .C0(n1859), .Y(n1857) );
  OAI22X1TS U6706 ( .A0(n3837), .A1(n5355), .B0(n5370), .B1(n1860), .Y(n1858)
         );
  OAI22X1TS U6707 ( .A0(n1239), .A1(n4586), .B0(n2099), .B1(n4554), .Y(n3340)
         );
  AOI222XLTS U6708 ( .A0(\addressToWriteBuffer[2][1] ), .A1(n5573), .B0(n4046), 
        .B1(n3866), .C0(n4131), .C1(n4625), .Y(n2099) );
  OAI22X1TS U6709 ( .A0(n4518), .A1(n1222), .B0(n2031), .B1(n4574), .Y(n3323)
         );
  AOI221XLTS U6710 ( .A0(n3759), .A1(n2032), .B0(n5208), .B1(n4134), .C0(n2033), .Y(n2031) );
  OAI22X1TS U6711 ( .A0(n3841), .A1(n5183), .B0(n5188), .B1(n2034), .Y(n2032)
         );
  OAI22X1TS U6712 ( .A0(n4672), .A1(n1206), .B0(n3777), .B1(n3840), .Y(n2033)
         );
  OAI22X1TS U6713 ( .A0(n4529), .A1(n1206), .B0(n1943), .B1(n4556), .Y(n3307)
         );
  AOI221XLTS U6714 ( .A0(n3757), .A1(n1944), .B0(n5300), .B1(n4136), .C0(n1945), .Y(n1943) );
  OAI22X1TS U6715 ( .A0(n3842), .A1(n5261), .B0(n5264), .B1(n1946), .Y(n1944)
         );
  OAI22X1TS U6716 ( .A0(n5282), .A1(n1190), .B0(n3782), .B1(n3841), .Y(n1945)
         );
  OAI22X1TS U6717 ( .A0(n4516), .A1(n1190), .B0(n1853), .B1(n4572), .Y(n3291)
         );
  AOI221XLTS U6718 ( .A0(n3761), .A1(n1854), .B0(n5380), .B1(n4134), .C0(n1855), .Y(n1853) );
  OAI22X1TS U6719 ( .A0(n3841), .A1(n5355), .B0(n5358), .B1(n1856), .Y(n1854)
         );
  OAI22X1TS U6720 ( .A0(n1238), .A1(n4587), .B0(n2098), .B1(n4554), .Y(n3339)
         );
  AOI222XLTS U6721 ( .A0(\addressToWriteBuffer[2][2] ), .A1(n5573), .B0(n4048), 
        .B1(n3863), .C0(n4135), .C1(n4625), .Y(n2098) );
  OAI22X1TS U6722 ( .A0(n4517), .A1(n1221), .B0(n2027), .B1(n4574), .Y(n3322)
         );
  AOI221XLTS U6723 ( .A0(n3760), .A1(n2028), .B0(n5208), .B1(n4138), .C0(n2029), .Y(n2027) );
  OAI22X1TS U6724 ( .A0(n3845), .A1(n5184), .B0(n5187), .B1(n2030), .Y(n2028)
         );
  OAI22X1TS U6725 ( .A0(n4673), .A1(n1205), .B0(n3778), .B1(n3844), .Y(n2029)
         );
  OAI22X1TS U6726 ( .A0(n4528), .A1(n1205), .B0(n1939), .B1(n4556), .Y(n3306)
         );
  AOI221XLTS U6727 ( .A0(n3758), .A1(n1940), .B0(n5300), .B1(n4140), .C0(n1941), .Y(n1939) );
  OAI22X1TS U6728 ( .A0(n3846), .A1(n5262), .B0(n5271), .B1(n1942), .Y(n1940)
         );
  OAI22X1TS U6729 ( .A0(n5282), .A1(n1189), .B0(n3780), .B1(n3845), .Y(n1941)
         );
  OAI22X1TS U6730 ( .A0(n4515), .A1(n1189), .B0(n1849), .B1(n4572), .Y(n3290)
         );
  AOI221XLTS U6731 ( .A0(n3762), .A1(n1850), .B0(n5380), .B1(n4138), .C0(n1851), .Y(n1849) );
  OAI22X1TS U6732 ( .A0(n3845), .A1(n5356), .B0(n5370), .B1(n1852), .Y(n1850)
         );
  OAI22X1TS U6733 ( .A0(n1237), .A1(n4586), .B0(n2097), .B1(n4554), .Y(n3338)
         );
  AOI222XLTS U6734 ( .A0(\addressToWriteBuffer[2][3] ), .A1(n5573), .B0(n4050), 
        .B1(n3864), .C0(n4139), .C1(n4625), .Y(n2097) );
  OAI22X1TS U6735 ( .A0(n4518), .A1(n1220), .B0(n2023), .B1(n4575), .Y(n3321)
         );
  AOI221XLTS U6736 ( .A0(n3759), .A1(n2024), .B0(n5209), .B1(n4142), .C0(n2025), .Y(n2023) );
  OAI22X1TS U6737 ( .A0(n3849), .A1(n5184), .B0(n5187), .B1(n2026), .Y(n2024)
         );
  OAI22X1TS U6738 ( .A0(n4663), .A1(n1204), .B0(n3779), .B1(n3848), .Y(n2025)
         );
  OAI22X1TS U6739 ( .A0(n4529), .A1(n1204), .B0(n1935), .B1(n4557), .Y(n3305)
         );
  AOI221XLTS U6740 ( .A0(n3757), .A1(n1936), .B0(n5301), .B1(n4144), .C0(n1937), .Y(n1935) );
  OAI22X1TS U6741 ( .A0(n3850), .A1(n5262), .B0(n5271), .B1(n1938), .Y(n1936)
         );
  OAI22X1TS U6742 ( .A0(n5281), .A1(n1188), .B0(n3781), .B1(n3849), .Y(n1937)
         );
  OAI22X1TS U6743 ( .A0(n4516), .A1(n1188), .B0(n1845), .B1(n4573), .Y(n3289)
         );
  AOI221XLTS U6744 ( .A0(n3761), .A1(n1846), .B0(n5381), .B1(n4142), .C0(n1847), .Y(n1845) );
  OAI22X1TS U6745 ( .A0(n3849), .A1(n5356), .B0(n5363), .B1(n1848), .Y(n1846)
         );
  OAI22X1TS U6746 ( .A0(n1236), .A1(n4587), .B0(n2096), .B1(n4555), .Y(n3337)
         );
  AOI222XLTS U6747 ( .A0(\addressToWriteBuffer[2][4] ), .A1(n5574), .B0(n4052), 
        .B1(n3865), .C0(n4143), .C1(n4624), .Y(n2096) );
  OAI22X1TS U6748 ( .A0(n4517), .A1(n1219), .B0(n2019), .B1(n4575), .Y(n3320)
         );
  AOI221XLTS U6749 ( .A0(n3760), .A1(n2020), .B0(n5209), .B1(n4146), .C0(n2021), .Y(n2019) );
  OAI22X1TS U6750 ( .A0(n4663), .A1(n1203), .B0(n3777), .B1(n3852), .Y(n2021)
         );
  OAI22X1TS U6751 ( .A0(n4528), .A1(n1203), .B0(n1931), .B1(n4557), .Y(n3304)
         );
  AOI221XLTS U6752 ( .A0(n3758), .A1(n1932), .B0(n5301), .B1(n4148), .C0(n1933), .Y(n1931) );
  OAI22X1TS U6753 ( .A0(n5281), .A1(n1187), .B0(n3782), .B1(n3853), .Y(n1933)
         );
  OAI22X1TS U6754 ( .A0(n4515), .A1(n1187), .B0(n1841), .B1(n4573), .Y(n3288)
         );
  AOI221XLTS U6755 ( .A0(n3762), .A1(n1842), .B0(n5381), .B1(n4146), .C0(n1843), .Y(n1841) );
  OAI22X1TS U6756 ( .A0(n1235), .A1(n4586), .B0(n2095), .B1(n4555), .Y(n3336)
         );
  AOI222XLTS U6757 ( .A0(\addressToWriteBuffer[2][5] ), .A1(n5571), .B0(n4054), 
        .B1(n3866), .C0(n4147), .C1(n4624), .Y(n2095) );
  OAI22X1TS U6758 ( .A0(n4517), .A1(n1218), .B0(n2015), .B1(n4575), .Y(n3319)
         );
  AOI221XLTS U6759 ( .A0(n3759), .A1(n2016), .B0(n5209), .B1(n4150), .C0(n2017), .Y(n2015) );
  OAI22X1TS U6760 ( .A0(n4663), .A1(n1202), .B0(n3778), .B1(n3856), .Y(n2017)
         );
  OAI22X1TS U6761 ( .A0(n4529), .A1(n1202), .B0(n1927), .B1(n4557), .Y(n3303)
         );
  AOI221XLTS U6762 ( .A0(n3757), .A1(n1928), .B0(n5301), .B1(n4152), .C0(n1929), .Y(n1927) );
  OAI22X1TS U6763 ( .A0(n5281), .A1(n1186), .B0(n3780), .B1(n3857), .Y(n1929)
         );
  OAI22X1TS U6764 ( .A0(n4515), .A1(n1186), .B0(n1837), .B1(n4573), .Y(n3287)
         );
  AOI221XLTS U6765 ( .A0(n3761), .A1(n1838), .B0(n5381), .B1(n4150), .C0(n1839), .Y(n1837) );
  OAI22X1TS U6766 ( .A0(n1234), .A1(n4587), .B0(n2094), .B1(n4555), .Y(n3335)
         );
  AOI222XLTS U6767 ( .A0(\addressToWriteBuffer[2][6] ), .A1(n5572), .B0(n4056), 
        .B1(n3863), .C0(n4151), .C1(n4624), .Y(n2094) );
  OAI22X1TS U6768 ( .A0(n4518), .A1(n1217), .B0(n2005), .B1(n4575), .Y(n3318)
         );
  AOI221XLTS U6769 ( .A0(n3760), .A1(n2008), .B0(n5209), .B1(n4154), .C0(n2010), .Y(n2005) );
  OAI22X1TS U6770 ( .A0(n3861), .A1(n5183), .B0(n5188), .B1(n2013), .Y(n2008)
         );
  OAI22X1TS U6771 ( .A0(n4664), .A1(n1201), .B0(n3779), .B1(n3860), .Y(n2010)
         );
  OAI22X1TS U6772 ( .A0(n4528), .A1(n1201), .B0(n1916), .B1(n4557), .Y(n3302)
         );
  AOI221XLTS U6773 ( .A0(n3758), .A1(n1919), .B0(n5301), .B1(n4156), .C0(n1921), .Y(n1916) );
  OAI22X1TS U6774 ( .A0(n3862), .A1(n5261), .B0(n5264), .B1(n1925), .Y(n1919)
         );
  OAI22X1TS U6775 ( .A0(n5283), .A1(n1185), .B0(n3781), .B1(n3861), .Y(n1921)
         );
  OAI22X1TS U6776 ( .A0(n4516), .A1(n1185), .B0(n1827), .B1(n4573), .Y(n3286)
         );
  AOI221XLTS U6777 ( .A0(n3762), .A1(n1830), .B0(n5381), .B1(n4154), .C0(n1832), .Y(n1827) );
  OAI22X1TS U6778 ( .A0(n3861), .A1(n5355), .B0(n5358), .B1(n1835), .Y(n1830)
         );
  OAI22X1TS U6779 ( .A0(n1233), .A1(n4586), .B0(n2092), .B1(n4555), .Y(n3334)
         );
  AOI222XLTS U6780 ( .A0(\addressToWriteBuffer[2][7] ), .A1(n5571), .B0(n4058), 
        .B1(n3864), .C0(n4155), .C1(n4624), .Y(n2092) );
  OAI22X1TS U6781 ( .A0(n1232), .A1(n4522), .B0(n2081), .B1(n4541), .Y(n3333)
         );
  AOI221XLTS U6782 ( .A0(n5169), .A1(n4128), .B0(n5155), .B1(n2082), .C0(n2083), .Y(n2081) );
  OAI22X1TS U6783 ( .A0(n3832), .A1(n5136), .B0(n5134), .B1(n2084), .Y(n2082)
         );
  OAI22X1TS U6784 ( .A0(n5401), .A1(n1216), .B0(n3810), .B1(n3834), .Y(n2083)
         );
  OAI22X1TS U6785 ( .A0(n1231), .A1(n4521), .B0(n2077), .B1(n4541), .Y(n3332)
         );
  AOI221XLTS U6786 ( .A0(n5169), .A1(n4132), .B0(n5155), .B1(n2078), .C0(n2079), .Y(n2077) );
  OAI22X1TS U6787 ( .A0(n3836), .A1(n5136), .B0(n5134), .B1(n2080), .Y(n2078)
         );
  OAI22X1TS U6788 ( .A0(n5400), .A1(n1215), .B0(n3811), .B1(n3838), .Y(n2079)
         );
  OAI22X1TS U6789 ( .A0(n1230), .A1(n4522), .B0(n2073), .B1(n4541), .Y(n3331)
         );
  AOI221XLTS U6790 ( .A0(n5169), .A1(n4136), .B0(n5155), .B1(n2074), .C0(n2075), .Y(n2073) );
  OAI22X1TS U6791 ( .A0(n3840), .A1(n5138), .B0(n5134), .B1(n2076), .Y(n2074)
         );
  OAI22X1TS U6792 ( .A0(n5400), .A1(n1214), .B0(n3811), .B1(n3842), .Y(n2075)
         );
  OAI22X1TS U6793 ( .A0(n1229), .A1(n4521), .B0(n2069), .B1(n4541), .Y(n3330)
         );
  AOI221XLTS U6794 ( .A0(n5169), .A1(n4140), .B0(n5155), .B1(n2070), .C0(n2071), .Y(n2069) );
  OAI22X1TS U6795 ( .A0(n3844), .A1(n5141), .B0(n5134), .B1(n2072), .Y(n2070)
         );
  OAI22X1TS U6796 ( .A0(n5400), .A1(n1213), .B0(n3810), .B1(n3846), .Y(n2071)
         );
  OAI22X1TS U6797 ( .A0(n1228), .A1(n4522), .B0(n2065), .B1(n4542), .Y(n3329)
         );
  AOI221XLTS U6798 ( .A0(n5170), .A1(n4144), .B0(n5156), .B1(n2066), .C0(n2067), .Y(n2065) );
  OAI22X1TS U6799 ( .A0(n3848), .A1(n5142), .B0(n5135), .B1(n2068), .Y(n2066)
         );
  OAI22X1TS U6800 ( .A0(n5404), .A1(n1212), .B0(n3811), .B1(n3850), .Y(n2067)
         );
  OAI22X1TS U6801 ( .A0(n1227), .A1(n4521), .B0(n2061), .B1(n4542), .Y(n3328)
         );
  AOI221XLTS U6802 ( .A0(n5170), .A1(n4148), .B0(n5156), .B1(n2062), .C0(n2063), .Y(n2061) );
  OAI22X1TS U6803 ( .A0(n3852), .A1(n5151), .B0(n5135), .B1(n2064), .Y(n2062)
         );
  OAI22X1TS U6804 ( .A0(n5399), .A1(n1211), .B0(n3810), .B1(n3854), .Y(n2063)
         );
  OAI22X1TS U6805 ( .A0(n1226), .A1(n4522), .B0(n2057), .B1(n4542), .Y(n3327)
         );
  AOI221XLTS U6806 ( .A0(n5170), .A1(n4152), .B0(n5156), .B1(n2058), .C0(n2059), .Y(n2057) );
  OAI22X1TS U6807 ( .A0(n3856), .A1(n5151), .B0(n5135), .B1(n2060), .Y(n2058)
         );
  OAI22X1TS U6808 ( .A0(n5399), .A1(n1210), .B0(n3811), .B1(n3858), .Y(n2059)
         );
  OAI22X1TS U6809 ( .A0(n1225), .A1(n4521), .B0(n2048), .B1(n4542), .Y(n3326)
         );
  AOI221XLTS U6810 ( .A0(n5170), .A1(n4156), .B0(n5156), .B1(n2052), .C0(n2053), .Y(n2048) );
  OAI22X1TS U6811 ( .A0(n3860), .A1(n5143), .B0(n5135), .B1(n2055), .Y(n2052)
         );
  OAI22X1TS U6812 ( .A0(n5399), .A1(n1209), .B0(n3660), .B1(n3862), .Y(n2053)
         );
  AOI221XLTS U6813 ( .A0(n3765), .A1(n1996), .B0(n5253), .B1(n4127), .C0(n1997), .Y(n1995) );
  OAI22X1TS U6814 ( .A0(n3834), .A1(n5222), .B0(n5237), .B1(n1998), .Y(n1996)
         );
  OAI22X1TS U6815 ( .A0(n5691), .A1(n1200), .B0(n3787), .B1(n4043), .Y(n1997)
         );
  AOI221XLTS U6816 ( .A0(n3766), .A1(n1992), .B0(n5250), .B1(n4131), .C0(n1993), .Y(n1991) );
  OAI22X1TS U6817 ( .A0(n3838), .A1(n5222), .B0(n5237), .B1(n1994), .Y(n1992)
         );
  OAI22X1TS U6818 ( .A0(n5683), .A1(n1199), .B0(n3788), .B1(n4045), .Y(n1993)
         );
  AOI221XLTS U6819 ( .A0(n3765), .A1(n1988), .B0(n5250), .B1(n4135), .C0(n1989), .Y(n1987) );
  OAI22X1TS U6820 ( .A0(n3842), .A1(n5222), .B0(n5230), .B1(n1990), .Y(n1988)
         );
  OAI22X1TS U6821 ( .A0(n5683), .A1(n1198), .B0(n3786), .B1(n4047), .Y(n1989)
         );
  AOI221XLTS U6822 ( .A0(n3766), .A1(n1984), .B0(n5253), .B1(n4139), .C0(n1985), .Y(n1983) );
  OAI22X1TS U6823 ( .A0(n3846), .A1(n5223), .B0(n5232), .B1(n1986), .Y(n1984)
         );
  OAI22X1TS U6824 ( .A0(n5683), .A1(n1197), .B0(n3787), .B1(n4049), .Y(n1985)
         );
  AOI221XLTS U6825 ( .A0(n3765), .A1(n1980), .B0(n1965), .B1(n4143), .C0(n1981), .Y(n1979) );
  OAI22X1TS U6826 ( .A0(n3850), .A1(n5223), .B0(n5241), .B1(n1982), .Y(n1980)
         );
  OAI22X1TS U6827 ( .A0(n5683), .A1(n1196), .B0(n3788), .B1(n4051), .Y(n1981)
         );
  AOI221XLTS U6828 ( .A0(n3766), .A1(n1976), .B0(n1965), .B1(n4147), .C0(n1977), .Y(n1975) );
  OAI22X1TS U6829 ( .A0(n3854), .A1(n5223), .B0(n5225), .B1(n1978), .Y(n1976)
         );
  OAI22X1TS U6830 ( .A0(n5682), .A1(n1195), .B0(n3786), .B1(n3853), .Y(n1977)
         );
  AOI221XLTS U6831 ( .A0(n3765), .A1(n1972), .B0(n5249), .B1(n4151), .C0(n1973), .Y(n1971) );
  OAI22X1TS U6832 ( .A0(n3858), .A1(n5223), .B0(n5225), .B1(n1974), .Y(n1972)
         );
  OAI22X1TS U6833 ( .A0(n5682), .A1(n1194), .B0(n3787), .B1(n3857), .Y(n1973)
         );
  AOI221XLTS U6834 ( .A0(n3766), .A1(n1964), .B0(n5251), .B1(n4155), .C0(n1966), .Y(n1961) );
  OAI22X1TS U6835 ( .A0(n3862), .A1(n5222), .B0(n5229), .B1(n1969), .Y(n1964)
         );
  OAI22X1TS U6836 ( .A0(n5695), .A1(n1193), .B0(n3788), .B1(n4057), .Y(n1966)
         );
  OAI22X1TS U6837 ( .A0(n4513), .A1(n1200), .B0(n1906), .B1(n4552), .Y(n3301)
         );
  AOI221XLTS U6838 ( .A0(n3767), .A1(n1907), .B0(n5344), .B1(n4127), .C0(n1908), .Y(n1906) );
  OAI22X1TS U6839 ( .A0(n3834), .A1(n5316), .B0(n5331), .B1(n1909), .Y(n1907)
         );
  OAI22X1TS U6840 ( .A0(n4701), .A1(n1184), .B0(n3789), .B1(n3833), .Y(n1908)
         );
  OAI22X1TS U6841 ( .A0(n4514), .A1(n1199), .B0(n1902), .B1(n4552), .Y(n3300)
         );
  AOI221XLTS U6842 ( .A0(n3768), .A1(n1903), .B0(n5344), .B1(n4131), .C0(n1904), .Y(n1902) );
  OAI22X1TS U6843 ( .A0(n3838), .A1(n5316), .B0(n5324), .B1(n1905), .Y(n1903)
         );
  OAI22X1TS U6844 ( .A0(n4699), .A1(n1183), .B0(n3790), .B1(n3837), .Y(n1904)
         );
  OAI22X1TS U6845 ( .A0(n4513), .A1(n1198), .B0(n1898), .B1(n4552), .Y(n3299)
         );
  AOI221XLTS U6846 ( .A0(n3767), .A1(n1899), .B0(n5347), .B1(n4135), .C0(n1900), .Y(n1898) );
  OAI22X1TS U6847 ( .A0(n3842), .A1(n5316), .B0(n5326), .B1(n1901), .Y(n1899)
         );
  OAI22X1TS U6848 ( .A0(n4700), .A1(n1182), .B0(n3791), .B1(n3841), .Y(n1900)
         );
  OAI22X1TS U6849 ( .A0(n4513), .A1(n1197), .B0(n1894), .B1(n4552), .Y(n3298)
         );
  AOI221XLTS U6850 ( .A0(n3768), .A1(n1895), .B0(n5346), .B1(n4139), .C0(n1896), .Y(n1894) );
  OAI22X1TS U6851 ( .A0(n3846), .A1(n5317), .B0(n5319), .B1(n1897), .Y(n1895)
         );
  OAI22X1TS U6852 ( .A0(n4704), .A1(n1181), .B0(n3789), .B1(n3845), .Y(n1896)
         );
  OAI22X1TS U6853 ( .A0(n4514), .A1(n1196), .B0(n1890), .B1(n4553), .Y(n3297)
         );
  AOI221XLTS U6854 ( .A0(n3767), .A1(n1891), .B0(n5343), .B1(n4143), .C0(n1892), .Y(n1890) );
  OAI22X1TS U6855 ( .A0(n3850), .A1(n5317), .B0(n5319), .B1(n1893), .Y(n1891)
         );
  OAI22X1TS U6856 ( .A0(n4698), .A1(n1180), .B0(n3790), .B1(n3849), .Y(n1892)
         );
  OAI22X1TS U6857 ( .A0(n1871), .A1(n1195), .B0(n1886), .B1(n4553), .Y(n3296)
         );
  AOI221XLTS U6858 ( .A0(n3768), .A1(n1887), .B0(n5343), .B1(n4147), .C0(n1888), .Y(n1886) );
  OAI22X1TS U6859 ( .A0(n4691), .A1(n1179), .B0(n3791), .B1(n3854), .Y(n1888)
         );
  OAI22X1TS U6860 ( .A0(n4513), .A1(n1194), .B0(n1882), .B1(n4553), .Y(n3295)
         );
  AOI221XLTS U6861 ( .A0(n3767), .A1(n1883), .B0(n5343), .B1(n4151), .C0(n1884), .Y(n1882) );
  OAI22X1TS U6862 ( .A0(n4691), .A1(n1178), .B0(n3789), .B1(n3858), .Y(n1884)
         );
  OAI22X1TS U6863 ( .A0(n4514), .A1(n1193), .B0(n1872), .B1(n4553), .Y(n3294)
         );
  AOI221XLTS U6864 ( .A0(n3768), .A1(n1875), .B0(n5343), .B1(n4155), .C0(n1877), .Y(n1872) );
  OAI22X1TS U6865 ( .A0(n3862), .A1(n5316), .B0(n5331), .B1(n1880), .Y(n1875)
         );
  OAI22X1TS U6866 ( .A0(n4699), .A1(n1177), .B0(n3790), .B1(n3861), .Y(n1877)
         );
  OAI22X1TS U6867 ( .A0(n1167), .A1(n4762), .B0(n3148), .B1(n4745), .Y(n3641)
         );
  AOI222XLTS U6868 ( .A0(\dataToWriteBuffer[2][0] ), .A1(n5572), .B0(n4735), 
        .B1(n4292), .C0(n4159), .C1(n4631), .Y(n3148) );
  OAI22X1TS U6869 ( .A0(n1166), .A1(n4762), .B0(n3147), .B1(n4745), .Y(n3640)
         );
  AOI222XLTS U6870 ( .A0(\dataToWriteBuffer[2][1] ), .A1(n5578), .B0(n4735), 
        .B1(n4297), .C0(n4163), .C1(n4623), .Y(n3147) );
  OAI22X1TS U6871 ( .A0(n1165), .A1(n4762), .B0(n3146), .B1(n4745), .Y(n3639)
         );
  AOI222XLTS U6872 ( .A0(\dataToWriteBuffer[2][2] ), .A1(n5582), .B0(n4735), 
        .B1(n4302), .C0(n4167), .C1(n4636), .Y(n3146) );
  OAI22X1TS U6873 ( .A0(n1164), .A1(n4763), .B0(n3145), .B1(n4745), .Y(n3638)
         );
  AOI222XLTS U6874 ( .A0(\dataToWriteBuffer[2][3] ), .A1(n5582), .B0(n4735), 
        .B1(n4307), .C0(n4171), .C1(n4634), .Y(n3145) );
  OAI22X1TS U6875 ( .A0(n1163), .A1(n3114), .B0(n3144), .B1(n4746), .Y(n3637)
         );
  AOI222XLTS U6876 ( .A0(\dataToWriteBuffer[2][4] ), .A1(n5581), .B0(n4736), 
        .B1(n4312), .C0(n4175), .C1(n4632), .Y(n3144) );
  OAI22X1TS U6877 ( .A0(n1162), .A1(n3114), .B0(n3143), .B1(n4746), .Y(n3636)
         );
  AOI222XLTS U6878 ( .A0(\dataToWriteBuffer[2][5] ), .A1(n5581), .B0(n4736), 
        .B1(n4317), .C0(n4179), .C1(n4636), .Y(n3143) );
  OAI22X1TS U6879 ( .A0(n1161), .A1(n4761), .B0(n3142), .B1(n4746), .Y(n3635)
         );
  AOI222XLTS U6880 ( .A0(\dataToWriteBuffer[2][6] ), .A1(n5581), .B0(n4736), 
        .B1(n4322), .C0(n4183), .C1(n4633), .Y(n3142) );
  OAI22X1TS U6881 ( .A0(n1160), .A1(n4760), .B0(n3141), .B1(n4746), .Y(n3634)
         );
  AOI222XLTS U6882 ( .A0(\dataToWriteBuffer[2][7] ), .A1(n5581), .B0(n4736), 
        .B1(n4327), .C0(n4187), .C1(n4633), .Y(n3141) );
  OAI22X1TS U6883 ( .A0(n1159), .A1(n4760), .B0(n3140), .B1(n4747), .Y(n3633)
         );
  AOI222XLTS U6884 ( .A0(\dataToWriteBuffer[2][8] ), .A1(n5580), .B0(n4737), 
        .B1(n4332), .C0(n4191), .C1(n4635), .Y(n3140) );
  OAI22X1TS U6885 ( .A0(n1158), .A1(n4764), .B0(n3139), .B1(n4747), .Y(n3632)
         );
  AOI222XLTS U6886 ( .A0(\dataToWriteBuffer[2][9] ), .A1(n5579), .B0(n4737), 
        .B1(n4337), .C0(n4195), .C1(n4632), .Y(n3139) );
  OAI22X1TS U6887 ( .A0(n1157), .A1(n4763), .B0(n3138), .B1(n4747), .Y(n3631)
         );
  AOI222XLTS U6888 ( .A0(\dataToWriteBuffer[2][10] ), .A1(n5580), .B0(n4737), 
        .B1(n4342), .C0(n4199), .C1(n4629), .Y(n3138) );
  OAI22X1TS U6889 ( .A0(n1156), .A1(n4755), .B0(n3137), .B1(n4747), .Y(n3630)
         );
  AOI222XLTS U6890 ( .A0(\dataToWriteBuffer[2][11] ), .A1(n5580), .B0(n4737), 
        .B1(n4347), .C0(n4203), .C1(n4629), .Y(n3137) );
  OAI22X1TS U6891 ( .A0(n1155), .A1(n4755), .B0(n3136), .B1(n4748), .Y(n3629)
         );
  AOI222XLTS U6892 ( .A0(\dataToWriteBuffer[2][12] ), .A1(n5579), .B0(n4738), 
        .B1(n4352), .C0(n4207), .C1(n4629), .Y(n3136) );
  OAI22X1TS U6893 ( .A0(n1154), .A1(n4755), .B0(n3135), .B1(n4748), .Y(n3628)
         );
  AOI222XLTS U6894 ( .A0(\dataToWriteBuffer[2][13] ), .A1(n5580), .B0(n4738), 
        .B1(n4357), .C0(n4211), .C1(n4629), .Y(n3135) );
  OAI22X1TS U6895 ( .A0(n1153), .A1(n4755), .B0(n3134), .B1(n4748), .Y(n3627)
         );
  AOI222XLTS U6896 ( .A0(\dataToWriteBuffer[2][14] ), .A1(n5579), .B0(n4738), 
        .B1(n4362), .C0(n4215), .C1(n4628), .Y(n3134) );
  OAI22X1TS U6897 ( .A0(n1152), .A1(n4756), .B0(n3133), .B1(n4748), .Y(n3626)
         );
  AOI222XLTS U6898 ( .A0(\dataToWriteBuffer[2][15] ), .A1(n5578), .B0(n4738), 
        .B1(n4367), .C0(n4219), .C1(n4628), .Y(n3133) );
  OAI22X1TS U6899 ( .A0(n1151), .A1(n4756), .B0(n3132), .B1(n4749), .Y(n3625)
         );
  AOI222XLTS U6900 ( .A0(\dataToWriteBuffer[2][16] ), .A1(n5579), .B0(n4739), 
        .B1(n4372), .C0(n4223), .C1(n4628), .Y(n3132) );
  OAI22X1TS U6901 ( .A0(n1150), .A1(n4756), .B0(n3131), .B1(n4749), .Y(n3624)
         );
  AOI222XLTS U6902 ( .A0(\dataToWriteBuffer[2][17] ), .A1(n5577), .B0(n4739), 
        .B1(n4377), .C0(n4227), .C1(n4628), .Y(n3131) );
  OAI22X1TS U6903 ( .A0(n1149), .A1(n4756), .B0(n3130), .B1(n4749), .Y(n3623)
         );
  AOI222XLTS U6904 ( .A0(\dataToWriteBuffer[2][18] ), .A1(n5575), .B0(n4739), 
        .B1(n4382), .C0(n4231), .C1(n4631), .Y(n3130) );
  OAI22X1TS U6905 ( .A0(n1148), .A1(n4757), .B0(n3129), .B1(n4749), .Y(n3622)
         );
  AOI222XLTS U6906 ( .A0(\dataToWriteBuffer[2][19] ), .A1(n5578), .B0(n4739), 
        .B1(n4387), .C0(n4235), .C1(n4630), .Y(n3129) );
  OAI22X1TS U6907 ( .A0(n1147), .A1(n4757), .B0(n3128), .B1(n4752), .Y(n3621)
         );
  AOI222XLTS U6908 ( .A0(\dataToWriteBuffer[2][20] ), .A1(n5578), .B0(n4742), 
        .B1(n4392), .C0(n4239), .C1(n4634), .Y(n3128) );
  OAI22X1TS U6909 ( .A0(n1146), .A1(n4757), .B0(n3127), .B1(n4753), .Y(n3620)
         );
  AOI222XLTS U6910 ( .A0(\dataToWriteBuffer[2][21] ), .A1(n5577), .B0(n4744), 
        .B1(n4397), .C0(n4243), .C1(n5760), .Y(n3127) );
  OAI22X1TS U6911 ( .A0(n1145), .A1(n4757), .B0(n3126), .B1(n4752), .Y(n3619)
         );
  AOI222XLTS U6912 ( .A0(\dataToWriteBuffer[2][22] ), .A1(n5577), .B0(n4743), 
        .B1(n4402), .C0(n4247), .C1(n4631), .Y(n3126) );
  OAI22X1TS U6913 ( .A0(n1144), .A1(n4758), .B0(n3125), .B1(n4753), .Y(n3618)
         );
  AOI222XLTS U6914 ( .A0(\dataToWriteBuffer[2][23] ), .A1(n5575), .B0(n4742), 
        .B1(n4407), .C0(n4251), .C1(n4630), .Y(n3125) );
  OAI22X1TS U6915 ( .A0(n1143), .A1(n4758), .B0(n3124), .B1(n4750), .Y(n3617)
         );
  AOI222XLTS U6916 ( .A0(\dataToWriteBuffer[2][24] ), .A1(n5576), .B0(n4740), 
        .B1(n4412), .C0(n4255), .C1(n4631), .Y(n3124) );
  OAI22X1TS U6917 ( .A0(n1142), .A1(n4758), .B0(n3123), .B1(n4750), .Y(n3616)
         );
  AOI222XLTS U6918 ( .A0(\dataToWriteBuffer[2][25] ), .A1(n5577), .B0(n4740), 
        .B1(n4417), .C0(n4259), .C1(n4627), .Y(n3123) );
  OAI22X1TS U6919 ( .A0(n1141), .A1(n4758), .B0(n3122), .B1(n4750), .Y(n3615)
         );
  AOI222XLTS U6920 ( .A0(\dataToWriteBuffer[2][26] ), .A1(n5576), .B0(n4740), 
        .B1(n4422), .C0(n4263), .C1(n4627), .Y(n3122) );
  OAI22X1TS U6921 ( .A0(n1140), .A1(n4759), .B0(n3121), .B1(n4750), .Y(n3614)
         );
  AOI222XLTS U6922 ( .A0(\dataToWriteBuffer[2][27] ), .A1(n5576), .B0(n4740), 
        .B1(n4427), .C0(n4267), .C1(n4627), .Y(n3121) );
  OAI22X1TS U6923 ( .A0(n1139), .A1(n4759), .B0(n3120), .B1(n4751), .Y(n3613)
         );
  AOI222XLTS U6924 ( .A0(\dataToWriteBuffer[2][28] ), .A1(n5576), .B0(n4741), 
        .B1(n4432), .C0(n4271), .C1(n4627), .Y(n3120) );
  OAI22X1TS U6925 ( .A0(n1138), .A1(n4759), .B0(n3119), .B1(n4751), .Y(n3612)
         );
  AOI222XLTS U6926 ( .A0(\dataToWriteBuffer[2][29] ), .A1(n5575), .B0(n4741), 
        .B1(n4437), .C0(n4275), .C1(n4626), .Y(n3119) );
  OAI22X1TS U6927 ( .A0(n1137), .A1(n4759), .B0(n3118), .B1(n4751), .Y(n3611)
         );
  AOI222XLTS U6928 ( .A0(\dataToWriteBuffer[2][30] ), .A1(n5575), .B0(n4741), 
        .B1(n4442), .C0(n4279), .C1(n4626), .Y(n3118) );
  OAI22X1TS U6929 ( .A0(n1136), .A1(n4760), .B0(n3115), .B1(n4751), .Y(n3610)
         );
  AOI222XLTS U6930 ( .A0(\dataToWriteBuffer[2][31] ), .A1(n5574), .B0(n4741), 
        .B1(n4447), .C0(n4283), .C1(n4626), .Y(n3115) );
  AOI221XLTS U6931 ( .A0(n5173), .A1(n4159), .B0(n5152), .B1(n3105), .C0(n3106), .Y(n3104) );
  OAI22X1TS U6932 ( .A0(n5399), .A1(n1071), .B0(n5906), .B1(n4786), .Y(n3106)
         );
  OAI22X1TS U6933 ( .A0(n5906), .A1(n5147), .B0(n5126), .B1(n3107), .Y(n3105)
         );
  AOI221XLTS U6934 ( .A0(n5174), .A1(n4163), .B0(n5152), .B1(n3101), .C0(n3102), .Y(n3100) );
  OAI22X1TS U6935 ( .A0(n5407), .A1(n1070), .B0(n5905), .B1(n4786), .Y(n3102)
         );
  OAI22X1TS U6936 ( .A0(n5905), .A1(n5147), .B0(n5126), .B1(n3103), .Y(n3101)
         );
  AOI221XLTS U6937 ( .A0(n5175), .A1(n4167), .B0(n5152), .B1(n3097), .C0(n3098), .Y(n3096) );
  OAI22X1TS U6938 ( .A0(n5409), .A1(n1069), .B0(n5904), .B1(n4786), .Y(n3098)
         );
  OAI22X1TS U6939 ( .A0(n5904), .A1(n5147), .B0(n5126), .B1(n3099), .Y(n3097)
         );
  AOI221XLTS U6940 ( .A0(n5174), .A1(n4171), .B0(n5152), .B1(n3093), .C0(n3094), .Y(n3092) );
  OAI22X1TS U6941 ( .A0(n5408), .A1(n1068), .B0(n5903), .B1(n4786), .Y(n3094)
         );
  OAI22X1TS U6942 ( .A0(n5903), .A1(n5147), .B0(n5126), .B1(n3095), .Y(n3093)
         );
  AOI221XLTS U6943 ( .A0(n5171), .A1(n4175), .B0(n5161), .B1(n3089), .C0(n3090), .Y(n3088) );
  OAI22X1TS U6944 ( .A0(n5407), .A1(n1067), .B0(n5902), .B1(n4787), .Y(n3090)
         );
  OAI22X1TS U6945 ( .A0(n5902), .A1(n5146), .B0(n5127), .B1(n3091), .Y(n3089)
         );
  AOI221XLTS U6946 ( .A0(n2050), .A1(n4179), .B0(n5157), .B1(n3085), .C0(n3086), .Y(n3084) );
  OAI22X1TS U6947 ( .A0(n5408), .A1(n1066), .B0(n5901), .B1(n4787), .Y(n3086)
         );
  OAI22X1TS U6948 ( .A0(n5901), .A1(n5146), .B0(n5127), .B1(n3087), .Y(n3085)
         );
  AOI221XLTS U6949 ( .A0(n5173), .A1(n4183), .B0(n2051), .B1(n3081), .C0(n3082), .Y(n3080) );
  OAI22X1TS U6950 ( .A0(n5408), .A1(n1065), .B0(n5900), .B1(n4787), .Y(n3082)
         );
  OAI22X1TS U6951 ( .A0(n5900), .A1(n5146), .B0(n5127), .B1(n3083), .Y(n3081)
         );
  AOI221XLTS U6952 ( .A0(n5171), .A1(n4187), .B0(n5157), .B1(n3077), .C0(n3078), .Y(n3076) );
  OAI22X1TS U6953 ( .A0(n5408), .A1(n1064), .B0(n5899), .B1(n4787), .Y(n3078)
         );
  OAI22X1TS U6954 ( .A0(n5899), .A1(n5146), .B0(n5127), .B1(n3079), .Y(n3077)
         );
  AOI221XLTS U6955 ( .A0(n5172), .A1(n4191), .B0(n5160), .B1(n3073), .C0(n3074), .Y(n3072) );
  OAI22X1TS U6956 ( .A0(n5407), .A1(n1063), .B0(n5898), .B1(n4788), .Y(n3074)
         );
  OAI22X1TS U6957 ( .A0(n5898), .A1(n5145), .B0(n5128), .B1(n3075), .Y(n3073)
         );
  AOI221XLTS U6958 ( .A0(n5175), .A1(n4195), .B0(n5163), .B1(n3069), .C0(n3070), .Y(n3068) );
  OAI22X1TS U6959 ( .A0(n5407), .A1(n1062), .B0(n5897), .B1(n4788), .Y(n3070)
         );
  OAI22X1TS U6960 ( .A0(n5897), .A1(n5145), .B0(n5128), .B1(n3071), .Y(n3069)
         );
  AOI221XLTS U6961 ( .A0(n5172), .A1(n4199), .B0(n5163), .B1(n3065), .C0(n3066), .Y(n3064) );
  OAI22X1TS U6962 ( .A0(n5406), .A1(n1061), .B0(n5896), .B1(n4788), .Y(n3066)
         );
  OAI22X1TS U6963 ( .A0(n5896), .A1(n5145), .B0(n5128), .B1(n3067), .Y(n3065)
         );
  AOI221XLTS U6964 ( .A0(n2050), .A1(n4203), .B0(n2051), .B1(n3061), .C0(n3062), .Y(n3060) );
  OAI22X1TS U6965 ( .A0(n5406), .A1(n1060), .B0(n5895), .B1(n4788), .Y(n3062)
         );
  OAI22X1TS U6966 ( .A0(n5895), .A1(n5145), .B0(n5128), .B1(n3063), .Y(n3061)
         );
  AOI221XLTS U6967 ( .A0(n5164), .A1(n4207), .B0(n5160), .B1(n3057), .C0(n3058), .Y(n3056) );
  OAI22X1TS U6968 ( .A0(n5406), .A1(n1059), .B0(n5894), .B1(n4789), .Y(n3058)
         );
  OAI22X1TS U6969 ( .A0(n5894), .A1(n5144), .B0(n5129), .B1(n3059), .Y(n3057)
         );
  AOI221XLTS U6970 ( .A0(n5164), .A1(n4211), .B0(n5160), .B1(n3053), .C0(n3054), .Y(n3052) );
  OAI22X1TS U6971 ( .A0(n5406), .A1(n1058), .B0(n5893), .B1(n4789), .Y(n3054)
         );
  OAI22X1TS U6972 ( .A0(n5893), .A1(n5144), .B0(n5129), .B1(n3055), .Y(n3053)
         );
  AOI221XLTS U6973 ( .A0(n5164), .A1(n4215), .B0(n5160), .B1(n3049), .C0(n3050), .Y(n3048) );
  OAI22X1TS U6974 ( .A0(n5405), .A1(n1057), .B0(n5892), .B1(n4789), .Y(n3050)
         );
  OAI22X1TS U6975 ( .A0(n5892), .A1(n5144), .B0(n5129), .B1(n3051), .Y(n3049)
         );
  AOI221XLTS U6976 ( .A0(n5164), .A1(n4219), .B0(n5161), .B1(n3045), .C0(n3046), .Y(n3044) );
  OAI22X1TS U6977 ( .A0(n5405), .A1(n1056), .B0(n5891), .B1(n4789), .Y(n3046)
         );
  OAI22X1TS U6978 ( .A0(n5891), .A1(n5144), .B0(n5129), .B1(n3047), .Y(n3045)
         );
  AOI221XLTS U6979 ( .A0(n5165), .A1(n4223), .B0(n5159), .B1(n3041), .C0(n3042), .Y(n3040) );
  OAI22X1TS U6980 ( .A0(n5405), .A1(n1055), .B0(n5890), .B1(n4794), .Y(n3042)
         );
  OAI22X1TS U6981 ( .A0(n5890), .A1(n5143), .B0(n5130), .B1(n3043), .Y(n3041)
         );
  AOI221XLTS U6982 ( .A0(n5165), .A1(n4227), .B0(n5159), .B1(n3037), .C0(n3038), .Y(n3036) );
  OAI22X1TS U6983 ( .A0(n5405), .A1(n1054), .B0(n5889), .B1(n4795), .Y(n3038)
         );
  OAI22X1TS U6984 ( .A0(n5889), .A1(n5143), .B0(n5130), .B1(n3039), .Y(n3037)
         );
  AOI221XLTS U6985 ( .A0(n5165), .A1(n4231), .B0(n5162), .B1(n3033), .C0(n3034), .Y(n3032) );
  OAI22X1TS U6986 ( .A0(n5404), .A1(n1053), .B0(n5888), .B1(n4794), .Y(n3034)
         );
  OAI22X1TS U6987 ( .A0(n5888), .A1(n5143), .B0(n5130), .B1(n3035), .Y(n3033)
         );
  AOI221XLTS U6988 ( .A0(n5165), .A1(n4235), .B0(n5161), .B1(n3029), .C0(n3030), .Y(n3028) );
  OAI22X1TS U6989 ( .A0(n5404), .A1(n1052), .B0(n5887), .B1(n4793), .Y(n3030)
         );
  OAI22X1TS U6990 ( .A0(n5887), .A1(n5142), .B0(n5130), .B1(n3031), .Y(n3029)
         );
  AOI221XLTS U6991 ( .A0(n5166), .A1(n4239), .B0(n5158), .B1(n3025), .C0(n3026), .Y(n3024) );
  OAI22X1TS U6992 ( .A0(n5404), .A1(n1051), .B0(n5886), .B1(n4790), .Y(n3026)
         );
  OAI22X1TS U6993 ( .A0(n5886), .A1(n5142), .B0(n5131), .B1(n3027), .Y(n3025)
         );
  AOI221XLTS U6994 ( .A0(n5166), .A1(n4243), .B0(n5159), .B1(n3021), .C0(n3022), .Y(n3020) );
  OAI22X1TS U6995 ( .A0(n5403), .A1(n1050), .B0(n5885), .B1(n4790), .Y(n3022)
         );
  OAI22X1TS U6996 ( .A0(n5885), .A1(n5141), .B0(n5131), .B1(n3023), .Y(n3021)
         );
  AOI221XLTS U6997 ( .A0(n5166), .A1(n4247), .B0(n5158), .B1(n3017), .C0(n3018), .Y(n3016) );
  OAI22X1TS U6998 ( .A0(n5403), .A1(n1049), .B0(n5884), .B1(n4790), .Y(n3018)
         );
  OAI22X1TS U6999 ( .A0(n5884), .A1(n5141), .B0(n5131), .B1(n3019), .Y(n3017)
         );
  AOI221XLTS U7000 ( .A0(n5166), .A1(n4251), .B0(n5159), .B1(n3013), .C0(n3014), .Y(n3012) );
  OAI22X1TS U7001 ( .A0(n5403), .A1(n1048), .B0(n5883), .B1(n4790), .Y(n3014)
         );
  OAI22X1TS U7002 ( .A0(n5883), .A1(n5140), .B0(n5131), .B1(n3015), .Y(n3013)
         );
  AOI221XLTS U7003 ( .A0(n5167), .A1(n4255), .B0(n5153), .B1(n3009), .C0(n3010), .Y(n3008) );
  OAI22X1TS U7004 ( .A0(n5403), .A1(n1047), .B0(n5882), .B1(n4791), .Y(n3010)
         );
  OAI22X1TS U7005 ( .A0(n5882), .A1(n5140), .B0(n5132), .B1(n3011), .Y(n3009)
         );
  AOI221XLTS U7006 ( .A0(n5167), .A1(n4259), .B0(n5153), .B1(n3005), .C0(n3006), .Y(n3004) );
  OAI22X1TS U7007 ( .A0(n5402), .A1(n1046), .B0(n5881), .B1(n4791), .Y(n3006)
         );
  OAI22X1TS U7008 ( .A0(n5881), .A1(n5139), .B0(n5132), .B1(n3007), .Y(n3005)
         );
  AOI221XLTS U7009 ( .A0(n5167), .A1(n4263), .B0(n5153), .B1(n3001), .C0(n3002), .Y(n3000) );
  OAI22X1TS U7010 ( .A0(n5402), .A1(n1045), .B0(n5880), .B1(n4791), .Y(n3002)
         );
  OAI22X1TS U7011 ( .A0(n5880), .A1(n5139), .B0(n5132), .B1(n3003), .Y(n3001)
         );
  AOI221XLTS U7012 ( .A0(n5167), .A1(n4267), .B0(n5153), .B1(n2997), .C0(n2998), .Y(n2996) );
  OAI22X1TS U7013 ( .A0(n5402), .A1(n1044), .B0(n5879), .B1(n4791), .Y(n2998)
         );
  OAI22X1TS U7014 ( .A0(n5879), .A1(n5138), .B0(n5132), .B1(n2999), .Y(n2997)
         );
  AOI221XLTS U7015 ( .A0(n5168), .A1(n4271), .B0(n5154), .B1(n2993), .C0(n2994), .Y(n2992) );
  OAI22X1TS U7016 ( .A0(n5402), .A1(n1043), .B0(n5878), .B1(n4792), .Y(n2994)
         );
  OAI22X1TS U7017 ( .A0(n5878), .A1(n5138), .B0(n5133), .B1(n2995), .Y(n2993)
         );
  AOI221XLTS U7018 ( .A0(n5168), .A1(n4275), .B0(n5154), .B1(n2989), .C0(n2990), .Y(n2988) );
  OAI22X1TS U7019 ( .A0(n5401), .A1(n1042), .B0(n5877), .B1(n4792), .Y(n2990)
         );
  OAI22X1TS U7020 ( .A0(n5877), .A1(n5137), .B0(n5133), .B1(n2991), .Y(n2989)
         );
  AOI221XLTS U7021 ( .A0(n5168), .A1(n4279), .B0(n5154), .B1(n2985), .C0(n2986), .Y(n2984) );
  OAI22X1TS U7022 ( .A0(n5401), .A1(n1041), .B0(n5876), .B1(n4792), .Y(n2986)
         );
  OAI22X1TS U7023 ( .A0(n5876), .A1(n5137), .B0(n5133), .B1(n2987), .Y(n2985)
         );
  AOI221XLTS U7024 ( .A0(n5168), .A1(n4283), .B0(n5154), .B1(n2979), .C0(n2980), .Y(n2977) );
  OAI22X1TS U7025 ( .A0(n5401), .A1(n1040), .B0(n5875), .B1(n4792), .Y(n2980)
         );
  OAI32X1TS U7026 ( .A0(n5751), .A1(n5732), .A2(n2229), .B0(n1761), .B1(n1170), 
        .Y(n3381) );
  INVX2TS U7027 ( .A(n1761), .Y(n5751) );
  AOI221XLTS U7028 ( .A0(n4288), .A1(n1764), .B0(isWrite[6]), .B1(n5294), .C0(
        n2230), .Y(n2229) );
  OAI32X1TS U7029 ( .A0(n5293), .A1(n2231), .A2(n2232), .B0(n3782), .B1(n3807), 
        .Y(n2230) );
  OAI222X1TS U7030 ( .A0(n3832), .A1(n5391), .B0(n4125), .B1(n4638), .C0(n5417), .C1(n1184), .Y(n3285) );
  OAI222X1TS U7031 ( .A0(n3836), .A1(n5391), .B0(n4129), .B1(n4638), .C0(n5417), .C1(n1183), .Y(n3284) );
  OAI222X1TS U7032 ( .A0(n3840), .A1(n5391), .B0(n4133), .B1(n4638), .C0(n5416), .C1(n1182), .Y(n3283) );
  OAI222X1TS U7033 ( .A0(n3844), .A1(n5391), .B0(n4137), .B1(n4637), .C0(n5416), .C1(n1181), .Y(n3282) );
  OAI222X1TS U7034 ( .A0(n3848), .A1(n5392), .B0(n4141), .B1(n4637), .C0(n5416), .C1(n1180), .Y(n3281) );
  OAI222X1TS U7035 ( .A0(n3852), .A1(n5392), .B0(n4145), .B1(n4637), .C0(n5416), .C1(n1179), .Y(n3280) );
  OAI222X1TS U7036 ( .A0(n3856), .A1(n5392), .B0(n4149), .B1(n4637), .C0(n5415), .C1(n1178), .Y(n3279) );
  OAI222X1TS U7037 ( .A0(n3860), .A1(n5392), .B0(n4153), .B1(n4648), .C0(n5417), .C1(n1177), .Y(n3278) );
  OAI222XLTS U7038 ( .A0(n5906), .A1(n5396), .B0(n4157), .B1(n4648), .C0(n5415), .C1(n943), .Y(n3417) );
  OAI222XLTS U7039 ( .A0(n5905), .A1(n5393), .B0(n4161), .B1(n4644), .C0(n1737), .C1(n942), .Y(n3416) );
  OAI222XLTS U7040 ( .A0(n5904), .A1(n1825), .B0(n4165), .B1(n4644), .C0(n1737), .C1(n941), .Y(n3415) );
  OAI222XLTS U7041 ( .A0(n5903), .A1(n5396), .B0(n4169), .B1(n4643), .C0(n5424), .C1(n940), .Y(n3414) );
  OAI222XLTS U7042 ( .A0(n5902), .A1(n5396), .B0(n4173), .B1(n4643), .C0(n5424), .C1(n939), .Y(n3413) );
  OAI222XLTS U7043 ( .A0(n5901), .A1(n5393), .B0(n4177), .B1(n4643), .C0(n5424), .C1(n938), .Y(n3412) );
  OAI222XLTS U7044 ( .A0(n5900), .A1(n5396), .B0(n4181), .B1(n4643), .C0(n5424), .C1(n937), .Y(n3411) );
  OAI222XLTS U7045 ( .A0(n5899), .A1(n1825), .B0(n4185), .B1(n4642), .C0(n5423), .C1(n936), .Y(n3410) );
  OAI222XLTS U7046 ( .A0(n5898), .A1(n5395), .B0(n4189), .B1(n4642), .C0(n5423), .C1(n935), .Y(n3409) );
  OAI222XLTS U7047 ( .A0(n5897), .A1(n5395), .B0(n4193), .B1(n4642), .C0(n5423), .C1(n934), .Y(n3408) );
  OAI222XLTS U7048 ( .A0(n5896), .A1(n5395), .B0(n4197), .B1(n4642), .C0(n5423), .C1(n933), .Y(n3407) );
  OAI222XLTS U7049 ( .A0(n5895), .A1(n5397), .B0(n4201), .B1(n4641), .C0(n5422), .C1(n932), .Y(n3406) );
  OAI222XLTS U7050 ( .A0(n5894), .A1(n5394), .B0(n4205), .B1(n4641), .C0(n5422), .C1(n931), .Y(n3405) );
  OAI222XLTS U7051 ( .A0(n5893), .A1(n5395), .B0(n4209), .B1(n4641), .C0(n5422), .C1(n930), .Y(n3404) );
  OAI222XLTS U7052 ( .A0(n5892), .A1(n5398), .B0(n4213), .B1(n4641), .C0(n5422), .C1(n929), .Y(n3403) );
  OAI222XLTS U7053 ( .A0(n5891), .A1(n5398), .B0(n4217), .B1(n4640), .C0(n5421), .C1(n928), .Y(n3402) );
  OAI222XLTS U7054 ( .A0(n5890), .A1(n5387), .B0(n4221), .B1(n4640), .C0(n5421), .C1(n927), .Y(n3401) );
  OAI222XLTS U7055 ( .A0(n5889), .A1(n5387), .B0(n4225), .B1(n4640), .C0(n5421), .C1(n926), .Y(n3400) );
  OAI222XLTS U7056 ( .A0(n5888), .A1(n5387), .B0(n4229), .B1(n4640), .C0(n5421), .C1(n925), .Y(n3399) );
  OAI222XLTS U7057 ( .A0(n5887), .A1(n5387), .B0(n4233), .B1(n4639), .C0(n5420), .C1(n924), .Y(n3398) );
  OAI222XLTS U7058 ( .A0(n5886), .A1(n5388), .B0(n4237), .B1(n4639), .C0(n5420), .C1(n923), .Y(n3397) );
  OAI222XLTS U7059 ( .A0(n5885), .A1(n5388), .B0(n4241), .B1(n4639), .C0(n5420), .C1(n922), .Y(n3396) );
  OAI222XLTS U7060 ( .A0(n5884), .A1(n5388), .B0(n4245), .B1(n4648), .C0(n5419), .C1(n921), .Y(n3395) );
  OAI222XLTS U7061 ( .A0(n5883), .A1(n5388), .B0(n4249), .B1(n4646), .C0(n5419), .C1(n920), .Y(n3394) );
  OAI222XLTS U7062 ( .A0(n5882), .A1(n5389), .B0(n4253), .B1(n4649), .C0(n5419), .C1(n919), .Y(n3393) );
  OAI222XLTS U7063 ( .A0(n5881), .A1(n5389), .B0(n4257), .B1(n5771), .C0(n5419), .C1(n918), .Y(n3392) );
  OAI222XLTS U7064 ( .A0(n5880), .A1(n5389), .B0(n4261), .B1(n4644), .C0(n5418), .C1(n917), .Y(n3391) );
  OAI222XLTS U7065 ( .A0(n5879), .A1(n5389), .B0(n4265), .B1(n4647), .C0(n5418), .C1(n916), .Y(n3390) );
  OAI222XLTS U7066 ( .A0(n5878), .A1(n5390), .B0(n4269), .B1(n4644), .C0(n5418), .C1(n915), .Y(n3389) );
  OAI222XLTS U7067 ( .A0(n5877), .A1(n5390), .B0(n4273), .B1(n5771), .C0(n5418), .C1(n914), .Y(n3388) );
  OAI222XLTS U7068 ( .A0(n5876), .A1(n5390), .B0(n4277), .B1(n4638), .C0(n5420), .C1(n913), .Y(n3387) );
  OAI222XLTS U7069 ( .A0(n5875), .A1(n5390), .B0(n4281), .B1(n4639), .C0(n5417), .C1(n912), .Y(n3386) );
  OAI32X1TS U7070 ( .A0(n5748), .A1(n5738), .A2(n2104), .B0(n1176), .B1(n2105), 
        .Y(n3343) );
  INVX2TS U7071 ( .A(n2105), .Y(n5748) );
  OAI211X1TS U7072 ( .A0(n5582), .A1(n3726), .B0(n5727), .C0(n2115), .Y(n2105)
         );
  AOI222XLTS U7073 ( .A0(n3966), .A1(n2106), .B0(n3863), .B1(n3686), .C0(n2107), .C1(n2108), .Y(n2104) );
  OAI32X1TS U7074 ( .A0(n5749), .A1(n5728), .A2(n2257), .B0(n1781), .B1(n1172), 
        .Y(n3383) );
  INVX2TS U7075 ( .A(n1781), .Y(n5749) );
  AOI221XLTS U7076 ( .A0(n4286), .A1(n1785), .B0(isWrite[4]), .B1(n4543), .C0(
        n2258), .Y(n2257) );
  OAI32XLTS U7077 ( .A0(n2259), .A1(n4543), .A2(n2260), .B0(n3777), .B1(n3808), 
        .Y(n2258) );
  OAI32X1TS U7078 ( .A0(n5752), .A1(n5731), .A2(n2201), .B0(n1738), .B1(n1168), 
        .Y(n3379) );
  INVX2TS U7079 ( .A(n1738), .Y(n5752) );
  AOI221XLTS U7080 ( .A0(n4288), .A1(n1742), .B0(isWrite[0]), .B1(n4534), .C0(
        n2202), .Y(n2201) );
  OAI32X1TS U7081 ( .A0(n2203), .A1(n4534), .A2(n2204), .B0(n3785), .B1(n3808), 
        .Y(n2202) );
  OAI32X1TS U7082 ( .A0(n5756), .A1(n5734), .A2(n2241), .B0(n1771), .B1(n1171), 
        .Y(n3382) );
  INVX2TS U7083 ( .A(n1771), .Y(n5756) );
  AOI221XLTS U7084 ( .A0(n4287), .A1(n1774), .B0(isWrite[5]), .B1(n5699), .C0(
        n2242), .Y(n2241) );
  OAI32X1TS U7085 ( .A0(n2243), .A1(n5699), .A2(n2244), .B0(n3786), .B1(n3807), 
        .Y(n2242) );
  OAI32X1TS U7086 ( .A0(n5757), .A1(n5733), .A2(n2215), .B0(n1750), .B1(n1169), 
        .Y(n3380) );
  INVX2TS U7087 ( .A(n1750), .Y(n5757) );
  AOI221XLTS U7088 ( .A0(n4287), .A1(n1754), .B0(isWrite[7]), .B1(n3805), .C0(
        n2216), .Y(n2215) );
  OAI32X1TS U7089 ( .A0(n2091), .A1(n5730), .A2(n2279), .B0(n1174), .B1(n4585), 
        .Y(n3385) );
  AOI222XLTS U7090 ( .A0(isWrite[2]), .A1(n5574), .B0(n3771), .B1(n3864), .C0(
        n4286), .C1(n4626), .Y(n2279) );
  AOI22XLTS U7091 ( .A0(n2847), .A1(n5176), .B0(n5197), .B1(n4446), .Y(n2845)
         );
  OAI22X1TS U7092 ( .A0(n4824), .A1(n5808), .B0(n5841), .B1(n4834), .Y(n2847)
         );
  INVX2TS U7093 ( .A(n4828), .Y(n4824) );
  AOI22XLTS U7094 ( .A0(n2573), .A1(n5263), .B0(n5274), .B1(n4447), .Y(n2571)
         );
  OAI22X1TS U7095 ( .A0(n4948), .A1(n5808), .B0(n5841), .B1(n4958), .Y(n2573)
         );
  INVX2TS U7096 ( .A(n4949), .Y(n4948) );
  AOI22XLTS U7097 ( .A0(n2294), .A1(n5348), .B0(n5368), .B1(n4448), .Y(n2292)
         );
  OAI22X1TS U7098 ( .A0(n5072), .A1(n5808), .B0(n5841), .B1(n5082), .Y(n2294)
         );
  INVX2TS U7099 ( .A(n5082), .Y(n5072) );
  AOI22XLTS U7100 ( .A0(n2709), .A1(n5215), .B0(n5235), .B1(n4446), .Y(n2707)
         );
  OAI22X1TS U7101 ( .A0(n4886), .A1(n3951), .B0(n4029), .B1(n4895), .Y(n2709)
         );
  INVX2TS U7102 ( .A(n4887), .Y(n4886) );
  AOI22XLTS U7103 ( .A0(n2435), .A1(n5318), .B0(n5329), .B1(n4445), .Y(n2433)
         );
  OAI22X1TS U7104 ( .A0(n5011), .A1(n5808), .B0(n5841), .B1(n5015), .Y(n2435)
         );
  INVX2TS U7105 ( .A(n5012), .Y(n5011) );
  AOI22XLTS U7106 ( .A0(n3812), .A1(n4103), .B0(n4079), .B1(n3793), .Y(n1909)
         );
  AOI22XLTS U7107 ( .A0(n3813), .A1(n4106), .B0(n4082), .B1(n3794), .Y(n1905)
         );
  AOI22XLTS U7108 ( .A0(n3667), .A1(n4109), .B0(n4085), .B1(n3792), .Y(n1901)
         );
  AOI22XLTS U7109 ( .A0(n3812), .A1(n4112), .B0(n4088), .B1(n3793), .Y(n1897)
         );
  AOI22XLTS U7110 ( .A0(n3813), .A1(n4115), .B0(n4091), .B1(n3794), .Y(n1893)
         );
  AOI22XLTS U7111 ( .A0(n3813), .A1(n4118), .B0(n4094), .B1(n3793), .Y(n1889)
         );
  AOI22XLTS U7112 ( .A0(n3813), .A1(n4121), .B0(n4097), .B1(n3794), .Y(n1885)
         );
  AOI22XLTS U7113 ( .A0(n3812), .A1(n4124), .B0(n4100), .B1(n3792), .Y(n1880)
         );
  AOI22XLTS U7114 ( .A0(n3814), .A1(n4103), .B0(n4079), .B1(n3796), .Y(n1864)
         );
  AOI22XLTS U7115 ( .A0(n3815), .A1(n4106), .B0(n4082), .B1(n3797), .Y(n1860)
         );
  AOI22XLTS U7116 ( .A0(n3815), .A1(n4109), .B0(n4085), .B1(n3795), .Y(n1856)
         );
  AOI22XLTS U7117 ( .A0(n3814), .A1(n4112), .B0(n4088), .B1(n3796), .Y(n1852)
         );
  AOI22XLTS U7118 ( .A0(n3815), .A1(n4115), .B0(n4091), .B1(n3797), .Y(n1848)
         );
  AOI22XLTS U7119 ( .A0(n3814), .A1(n4117), .B0(n4093), .B1(n3796), .Y(n1844)
         );
  AOI22XLTS U7120 ( .A0(n3815), .A1(n4120), .B0(n4096), .B1(n3797), .Y(n1840)
         );
  AOI22XLTS U7121 ( .A0(n3814), .A1(n4124), .B0(n4100), .B1(n3795), .Y(n1835)
         );
  AOI22XLTS U7122 ( .A0(n3773), .A1(n4102), .B0(n4078), .B1(n3823), .Y(n2084)
         );
  AOI22XLTS U7123 ( .A0(n3774), .A1(n4105), .B0(n4081), .B1(n3824), .Y(n2080)
         );
  AOI22XLTS U7124 ( .A0(n3773), .A1(n4108), .B0(n4084), .B1(n3822), .Y(n2076)
         );
  AOI22XLTS U7125 ( .A0(n3774), .A1(n4111), .B0(n4087), .B1(n3823), .Y(n2072)
         );
  AOI22XLTS U7126 ( .A0(n3773), .A1(n4114), .B0(n4090), .B1(n3824), .Y(n2068)
         );
  AOI22XLTS U7127 ( .A0(n3773), .A1(n4117), .B0(n4093), .B1(n3824), .Y(n2064)
         );
  AOI22XLTS U7128 ( .A0(n3774), .A1(n4120), .B0(n4096), .B1(n3822), .Y(n2060)
         );
  AOI22XLTS U7129 ( .A0(n3774), .A1(n4123), .B0(n4099), .B1(n3822), .Y(n2055)
         );
  AOI22XLTS U7130 ( .A0(n3775), .A1(n4102), .B0(n4078), .B1(n3830), .Y(n1954)
         );
  AOI22XLTS U7131 ( .A0(n3776), .A1(n4105), .B0(n4081), .B1(n1926), .Y(n1950)
         );
  AOI22XLTS U7132 ( .A0(n3775), .A1(n4108), .B0(n4084), .B1(n3829), .Y(n1946)
         );
  AOI22XLTS U7133 ( .A0(n3776), .A1(n4111), .B0(n4087), .B1(n3830), .Y(n1942)
         );
  AOI22XLTS U7134 ( .A0(n3775), .A1(n4114), .B0(n4090), .B1(n1926), .Y(n1938)
         );
  AOI22XLTS U7135 ( .A0(n3776), .A1(n4118), .B0(n4094), .B1(n3830), .Y(n1934)
         );
  AOI22XLTS U7136 ( .A0(n3775), .A1(n4121), .B0(n4097), .B1(n1926), .Y(n1930)
         );
  AOI22XLTS U7137 ( .A0(n3776), .A1(n4123), .B0(n4099), .B1(n3829), .Y(n1925)
         );
  AOI221XLTS U7138 ( .A0(n4286), .A1(n1797), .B0(isWrite[3]), .B1(n4611), .C0(
        n2269), .Y(n2268) );
  OAI22X1TS U7139 ( .A0(n1278), .A1(n4620), .B0(n1619), .B1(n1620), .Y(n3203)
         );
  AOI222XLTS U7140 ( .A0(n4032), .A1(n1621), .B0(n3739), .B1(n1622), .C0(n4061), .C1(n3755), .Y(n1619) );
  OAI2BB2XLTS U7141 ( .B0(n3870), .B1(n1624), .A0N(n4060), .A1N(n3871), .Y(
        n1622) );
  AOI22XLTS U7142 ( .A0(n3821), .A1(n3954), .B0(n3878), .B1(n3827), .Y(n1624)
         );
  AOI222XLTS U7143 ( .A0(n4034), .A1(n3747), .B0(n3740), .B1(n1627), .C0(n4063), .C1(n3756), .Y(n1626) );
  OAI2BB2XLTS U7144 ( .B0(n3868), .B1(n1628), .A0N(n4063), .A1N(n3869), .Y(
        n1627) );
  AOI22XLTS U7145 ( .A0(n3820), .A1(n3956), .B0(n3880), .B1(n3825), .Y(n1628)
         );
  AOI222XLTS U7146 ( .A0(n4036), .A1(n1621), .B0(n3739), .B1(n1630), .C0(n4066), .C1(n3755), .Y(n1629) );
  OAI2BB2XLTS U7147 ( .B0(n3869), .B1(n1631), .A0N(n4066), .A1N(n3870), .Y(
        n1630) );
  AOI22XLTS U7148 ( .A0(n3821), .A1(n3958), .B0(n3882), .B1(n3826), .Y(n1631)
         );
  AOI222XLTS U7149 ( .A0(n4038), .A1(n3747), .B0(n3740), .B1(n1633), .C0(n4069), .C1(n3756), .Y(n1632) );
  OAI2BB2XLTS U7150 ( .B0(n3870), .B1(n1634), .A0N(n4069), .A1N(n3871), .Y(
        n1633) );
  AOI22XLTS U7151 ( .A0(n3820), .A1(n3960), .B0(n3884), .B1(n3827), .Y(n1634)
         );
  AOI222XLTS U7152 ( .A0(n4040), .A1(n1621), .B0(n3739), .B1(n1636), .C0(n4072), .C1(n3755), .Y(n1635) );
  OAI2BB2XLTS U7153 ( .B0(n3871), .B1(n1637), .A0N(n4072), .A1N(n3868), .Y(
        n1636) );
  AOI22XLTS U7154 ( .A0(n3820), .A1(n3962), .B0(n3886), .B1(n3825), .Y(n1637)
         );
  AOI222XLTS U7155 ( .A0(n4042), .A1(n3747), .B0(n3740), .B1(n1639), .C0(n4075), .C1(n3756), .Y(n1638) );
  OAI2BB2XLTS U7156 ( .B0(n3868), .B1(n1640), .A0N(n4075), .A1N(n3869), .Y(
        n1639) );
  AOI22XLTS U7157 ( .A0(n3821), .A1(n3964), .B0(n3888), .B1(n3826), .Y(n1640)
         );
  NOR2X1TS U7158 ( .A(n1797), .B(n1801), .Y(n1800) );
  OAI32X1TS U7159 ( .A0(n3825), .A1(n3871), .A2(n5974), .B0(n5409), .B1(n1258), 
        .Y(n1801) );
  OAI22X1TS U7160 ( .A0(n1781), .A1(n1260), .B0(n5737), .B1(n1789), .Y(n3263)
         );
  AOI211XLTS U7161 ( .A0(n4543), .A1(\requesterPortBuffer[4][0] ), .B0(n1785), 
        .C0(n1790), .Y(n1789) );
  NOR4XLTS U7162 ( .A(n3717), .B(n5788), .C(n1788), .D(n1791), .Y(n1790) );
  OAI22X1TS U7163 ( .A0(n1738), .A1(n1252), .B0(n5735), .B1(n1746), .Y(n3255)
         );
  AOI211XLTS U7164 ( .A0(n4534), .A1(\requesterPortBuffer[0][0] ), .B0(n1742), 
        .C0(n1747), .Y(n1746) );
  NOR4XLTS U7165 ( .A(n4617), .B(n5790), .C(n1745), .D(n1749), .Y(n1747) );
  OAI22X1TS U7166 ( .A0(n1781), .A1(n1259), .B0(n5737), .B1(n1782), .Y(n3262)
         );
  AOI211XLTS U7167 ( .A0(n4543), .A1(\requesterPortBuffer[4][1] ), .B0(n1784), 
        .C0(n1785), .Y(n1782) );
  OAI22X1TS U7168 ( .A0(n5562), .A1(n1786), .B0(n1787), .B1(n1788), .Y(n1784)
         );
  OAI22X1TS U7169 ( .A0(n1761), .A1(n1255), .B0(n5736), .B1(n1762), .Y(n3258)
         );
  AOI211X1TS U7170 ( .A0(\requesterPortBuffer[6][1] ), .A1(n4614), .B0(n1763), 
        .C0(n1764), .Y(n1762) );
  OAI22X1TS U7171 ( .A0(n5562), .A1(n1765), .B0(n1766), .B1(n1767), .Y(n1763)
         );
  OAI22X1TS U7172 ( .A0(n1738), .A1(n1251), .B0(n5735), .B1(n1739), .Y(n3254)
         );
  AOI211XLTS U7173 ( .A0(n4534), .A1(\requesterPortBuffer[0][1] ), .B0(n1741), 
        .C0(n1742), .Y(n1739) );
  OAI22X1TS U7174 ( .A0(n5561), .A1(n1743), .B0(n1744), .B1(n1745), .Y(n1741)
         );
  AOI211X1TS U7175 ( .A0(n5754), .A1(n5594), .B0(n1796), .C0(n1797), .Y(n1795)
         );
  OAI22X1TS U7176 ( .A0(n5400), .A1(n1257), .B0(n5974), .B1(n1799), .Y(n1796)
         );
  OAI22X1TS U7177 ( .A0(n1771), .A1(n1258), .B0(n5737), .B1(n1778), .Y(n3261)
         );
  AOI211X1TS U7178 ( .A0(\requesterPortBuffer[5][0] ), .A1(n5700), .B0(n1774), 
        .C0(n1779), .Y(n1778) );
  NOR4XLTS U7179 ( .A(n4547), .B(n5791), .C(n1777), .D(n1780), .Y(n1779) );
  OAI22X1TS U7180 ( .A0(n1771), .A1(n1257), .B0(n5736), .B1(n1772), .Y(n3260)
         );
  AOI211X1TS U7181 ( .A0(\requesterPortBuffer[5][1] ), .A1(n5701), .B0(n1773), 
        .C0(n1774), .Y(n1772) );
  OAI22X1TS U7182 ( .A0(n5562), .A1(n1775), .B0(n1776), .B1(n1777), .Y(n1773)
         );
  OAI22X1TS U7183 ( .A0(n1750), .A1(n1254), .B0(n5735), .B1(n1758), .Y(n3257)
         );
  AOI211X1TS U7184 ( .A0(n1752), .A1(\requesterPortBuffer[7][0] ), .B0(n1754), 
        .C0(n1759), .Y(n1758) );
  NOR4XLTS U7185 ( .A(n3717), .B(n5787), .C(n1757), .D(n1760), .Y(n1759) );
  OAI22X1TS U7186 ( .A0(n1750), .A1(n1253), .B0(n5738), .B1(n1751), .Y(n3256)
         );
  AOI211X1TS U7187 ( .A0(n3806), .A1(\requesterPortBuffer[7][1] ), .B0(n1753), 
        .C0(n1754), .Y(n1751) );
  OAI22X1TS U7188 ( .A0(n5562), .A1(n1755), .B0(n1756), .B1(n1757), .Y(n1753)
         );
  OAI2BB2XLTS U7189 ( .B0(n5427), .B1(n2198), .A0N(n5426), .A1N(isWrite[7]), 
        .Y(n3378) );
  AOI22XLTS U7190 ( .A0(n3772), .A1(n2199), .B0(n4287), .B1(n2200), .Y(n2198)
         );
  OAI2BB2XLTS U7191 ( .B0(n5734), .B1(n1804), .A0N(\requesterPortBuffer[0][0] ), .A1N(n1802), .Y(n3269) );
  AOI21X1TS U7192 ( .A0(\requesterPortBuffer[2][0] ), .A1(n5564), .B0(n4622), 
        .Y(n1804) );
  AOI21X1TS U7193 ( .A0(n2116), .A1(n5565), .B0(n2106), .Y(n2115) );
  OAI21X1TS U7194 ( .A0(n4547), .A1(n2113), .B0(n2118), .Y(n2116) );
  AOI32X1TS U7195 ( .A0(n4621), .A1(n5714), .A2(n2119), .B0(n2111), .B1(n4591), 
        .Y(n2118) );
  OAI22X1TS U7196 ( .A0(n1761), .A1(n1256), .B0(n5736), .B1(n1768), .Y(n3259)
         );
  AOI211X1TS U7197 ( .A0(\requesterPortBuffer[6][0] ), .A1(n4614), .B0(n1764), 
        .C0(n1769), .Y(n1768) );
  NOR4XLTS U7198 ( .A(n4547), .B(n5789), .C(n1767), .D(n1770), .Y(n1769) );
  AO22X1TS U7199 ( .A0(\requesterPortBuffer[0][1] ), .A1(n1802), .B0(n5726), 
        .B1(n1803), .Y(n3268) );
  OAI221XLTS U7200 ( .A0(n1259), .A1(n5594), .B0(n3726), .B1(n5585), .C0(n1598), .Y(n1803) );
  OAI2BB1X1TS U7201 ( .A0N(n5425), .A1N(\requesterPortBuffer[7][0] ), .B0(
        n4647), .Y(n3253) );
  OAI32X1TS U7202 ( .A0(n2124), .A1(n5730), .A2(n2125), .B0(n1175), .B1(n5753), 
        .Y(n3345) );
  INVX2TS U7203 ( .A(n2124), .Y(n5753) );
  AOI222XLTS U7204 ( .A0(n3966), .A1(n2126), .B0(n3686), .B1(n3756), .C0(n2127), .C1(n2128), .Y(n2125) );
  OAI221XLTS U7205 ( .A0(n4550), .A1(n1736), .B0(n5415), .B1(n1250), .C0(n4646), .Y(n3252) );
  OAI211X1TS U7206 ( .A0(n5492), .A1(n4077), .B0(n1805), .C0(n1806), .Y(n3270)
         );
  AOI22XLTS U7207 ( .A0(\addressToWriteBuffer[0][0] ), .A1(n5442), .B0(n5430), 
        .B1(n4044), .Y(n1805) );
  AOI222XLTS U7208 ( .A0(cacheAddressIn_A[0]), .A1(n5606), .B0(n5485), .B1(
        n4102), .C0(n5476), .C1(n4126), .Y(n1806) );
  OAI211X1TS U7209 ( .A0(n5492), .A1(n4080), .B0(n1807), .C0(n1808), .Y(n3271)
         );
  AOI22XLTS U7210 ( .A0(\addressToWriteBuffer[0][1] ), .A1(n5442), .B0(n5430), 
        .B1(n4046), .Y(n1807) );
  AOI222XLTS U7211 ( .A0(cacheAddressIn_A[1]), .A1(n5606), .B0(n5485), .B1(
        n4105), .C0(n5477), .C1(n4130), .Y(n1808) );
  OAI211X1TS U7212 ( .A0(n5492), .A1(n4083), .B0(n1809), .C0(n1810), .Y(n3272)
         );
  AOI22XLTS U7213 ( .A0(\addressToWriteBuffer[0][2] ), .A1(n5442), .B0(n5430), 
        .B1(n4048), .Y(n1809) );
  AOI222XLTS U7214 ( .A0(cacheAddressIn_A[2]), .A1(n5606), .B0(n5485), .B1(
        n4108), .C0(n1667), .C1(n4134), .Y(n1810) );
  OAI211X1TS U7215 ( .A0(n5492), .A1(n4086), .B0(n1811), .C0(n1812), .Y(n3273)
         );
  AOI22XLTS U7216 ( .A0(\addressToWriteBuffer[0][3] ), .A1(n5442), .B0(n5430), 
        .B1(n4050), .Y(n1811) );
  AOI222XLTS U7217 ( .A0(cacheAddressIn_A[3]), .A1(n5606), .B0(n5485), .B1(
        n4111), .C0(n1667), .C1(n4138), .Y(n1812) );
  OAI211X1TS U7218 ( .A0(n5491), .A1(n4089), .B0(n1813), .C0(n1814), .Y(n3274)
         );
  AOI22XLTS U7219 ( .A0(\addressToWriteBuffer[0][4] ), .A1(n5441), .B0(n5429), 
        .B1(n4052), .Y(n1813) );
  AOI222XLTS U7220 ( .A0(cacheAddressIn_A[4]), .A1(n5607), .B0(n5486), .B1(
        n4114), .C0(n5476), .C1(n4142), .Y(n1814) );
  OAI211X1TS U7221 ( .A0(n5491), .A1(n4092), .B0(n1815), .C0(n1816), .Y(n3275)
         );
  AOI22XLTS U7222 ( .A0(\addressToWriteBuffer[0][5] ), .A1(n5441), .B0(n5429), 
        .B1(n4054), .Y(n1815) );
  AOI222XLTS U7223 ( .A0(cacheAddressIn_A[5]), .A1(n5607), .B0(n5486), .B1(
        n4117), .C0(n5476), .C1(n4146), .Y(n1816) );
  OAI211X1TS U7224 ( .A0(n5491), .A1(n4095), .B0(n1817), .C0(n1818), .Y(n3276)
         );
  AOI22XLTS U7225 ( .A0(\addressToWriteBuffer[0][6] ), .A1(n5441), .B0(n5429), 
        .B1(n4056), .Y(n1817) );
  AOI222XLTS U7226 ( .A0(cacheAddressIn_A[6]), .A1(n5607), .B0(n5486), .B1(
        n4120), .C0(n5476), .C1(n4150), .Y(n1818) );
  OAI211X1TS U7227 ( .A0(n5491), .A1(n4098), .B0(n1819), .C0(n1820), .Y(n3277)
         );
  AOI22XLTS U7228 ( .A0(\addressToWriteBuffer[0][7] ), .A1(n5441), .B0(n5429), 
        .B1(n4058), .Y(n1819) );
  AOI222XLTS U7229 ( .A0(cacheAddressIn_A[7]), .A1(n5613), .B0(n5486), .B1(
        n4123), .C0(n5478), .C1(n4154), .Y(n1820) );
  OAI211X1TS U7230 ( .A0(n5501), .A1(n3889), .B0(n1664), .C0(n1665), .Y(n3218)
         );
  AOI22XLTS U7231 ( .A0(\dataToWriteBuffer[0][0] ), .A1(n5450), .B0(n4291), 
        .B1(n5435), .Y(n1664) );
  AOI222XLTS U7232 ( .A0(cacheDataIn_A[0]), .A1(n5612), .B0(n3968), .B1(n5487), 
        .C0(n4158), .C1(n5471), .Y(n1665) );
  OAI211X1TS U7233 ( .A0(n5501), .A1(n3891), .B0(n1670), .C0(n1671), .Y(n3219)
         );
  AOI22XLTS U7234 ( .A0(\dataToWriteBuffer[0][1] ), .A1(n5450), .B0(n4296), 
        .B1(n5435), .Y(n1670) );
  AOI222XLTS U7235 ( .A0(cacheDataIn_A[1]), .A1(n5608), .B0(n3970), .B1(n5487), 
        .C0(n4162), .C1(n5471), .Y(n1671) );
  OAI211X1TS U7236 ( .A0(n5500), .A1(n3893), .B0(n1672), .C0(n1673), .Y(n3220)
         );
  AOI22XLTS U7237 ( .A0(\dataToWriteBuffer[0][2] ), .A1(n5450), .B0(n4301), 
        .B1(n5435), .Y(n1672) );
  AOI222XLTS U7238 ( .A0(cacheDataIn_A[2]), .A1(n5610), .B0(n3972), .B1(n5490), 
        .C0(n4166), .C1(n5471), .Y(n1673) );
  OAI211X1TS U7239 ( .A0(n5499), .A1(n3895), .B0(n1674), .C0(n1675), .Y(n3221)
         );
  AOI22XLTS U7240 ( .A0(\dataToWriteBuffer[0][3] ), .A1(n5450), .B0(n4306), 
        .B1(n5435), .Y(n1674) );
  AOI222XLTS U7241 ( .A0(cacheDataIn_A[3]), .A1(n5609), .B0(n3974), .B1(n1666), 
        .C0(n4170), .C1(n5471), .Y(n1675) );
  OAI211X1TS U7242 ( .A0(n5498), .A1(n3897), .B0(n1676), .C0(n1677), .Y(n3222)
         );
  AOI22XLTS U7243 ( .A0(\dataToWriteBuffer[0][4] ), .A1(n5449), .B0(n4311), 
        .B1(n5434), .Y(n1676) );
  AOI222XLTS U7244 ( .A0(cacheDataIn_A[4]), .A1(n5608), .B0(n3976), .B1(n5479), 
        .C0(n4174), .C1(n5470), .Y(n1677) );
  OAI211X1TS U7245 ( .A0(n5498), .A1(n3899), .B0(n1678), .C0(n1679), .Y(n3223)
         );
  AOI22XLTS U7246 ( .A0(\dataToWriteBuffer[0][5] ), .A1(n5449), .B0(n4316), 
        .B1(n5434), .Y(n1678) );
  AOI222XLTS U7247 ( .A0(cacheDataIn_A[5]), .A1(n5610), .B0(n3978), .B1(n5479), 
        .C0(n4178), .C1(n5470), .Y(n1679) );
  OAI211X1TS U7248 ( .A0(n5498), .A1(n3901), .B0(n1680), .C0(n1681), .Y(n3224)
         );
  AOI22XLTS U7249 ( .A0(\dataToWriteBuffer[0][6] ), .A1(n5449), .B0(n4321), 
        .B1(n5434), .Y(n1680) );
  AOI222XLTS U7250 ( .A0(cacheDataIn_A[6]), .A1(n5609), .B0(n3980), .B1(n5479), 
        .C0(n4182), .C1(n5470), .Y(n1681) );
  OAI211X1TS U7251 ( .A0(n5498), .A1(n3903), .B0(n1682), .C0(n1683), .Y(n3225)
         );
  AOI22XLTS U7252 ( .A0(\dataToWriteBuffer[0][7] ), .A1(n5449), .B0(n4326), 
        .B1(n5434), .Y(n1682) );
  AOI222XLTS U7253 ( .A0(cacheDataIn_A[7]), .A1(n5612), .B0(n3982), .B1(n5479), 
        .C0(n4186), .C1(n5470), .Y(n1683) );
  OAI211X1TS U7254 ( .A0(n5497), .A1(n3905), .B0(n1684), .C0(n1685), .Y(n3226)
         );
  AOI22XLTS U7255 ( .A0(\dataToWriteBuffer[0][8] ), .A1(n5448), .B0(n4331), 
        .B1(n5433), .Y(n1684) );
  AOI222XLTS U7256 ( .A0(cacheDataIn_A[8]), .A1(n5602), .B0(n3984), .B1(n5480), 
        .C0(n4190), .C1(n5469), .Y(n1685) );
  OAI211X1TS U7257 ( .A0(n5497), .A1(n3907), .B0(n1686), .C0(n1687), .Y(n3227)
         );
  AOI22XLTS U7258 ( .A0(\dataToWriteBuffer[0][9] ), .A1(n5448), .B0(n4336), 
        .B1(n5433), .Y(n1686) );
  AOI222XLTS U7259 ( .A0(cacheDataIn_A[9]), .A1(n5611), .B0(n3986), .B1(n5480), 
        .C0(n4194), .C1(n5469), .Y(n1687) );
  OAI211X1TS U7260 ( .A0(n5497), .A1(n3909), .B0(n1688), .C0(n1689), .Y(n3228)
         );
  AOI22XLTS U7261 ( .A0(\dataToWriteBuffer[0][10] ), .A1(n5448), .B0(n4341), 
        .B1(n5433), .Y(n1688) );
  AOI222XLTS U7262 ( .A0(cacheDataIn_A[10]), .A1(n5611), .B0(n3988), .B1(n5480), .C0(n4198), .C1(n5469), .Y(n1689) );
  OAI211X1TS U7263 ( .A0(n5497), .A1(n3911), .B0(n1690), .C0(n1691), .Y(n3229)
         );
  AOI22XLTS U7264 ( .A0(\dataToWriteBuffer[0][11] ), .A1(n5448), .B0(n4346), 
        .B1(n5433), .Y(n1690) );
  AOI222XLTS U7265 ( .A0(cacheDataIn_A[11]), .A1(n5612), .B0(n3990), .B1(n5480), .C0(n4202), .C1(n5469), .Y(n1691) );
  OAI211X1TS U7266 ( .A0(n5496), .A1(n3913), .B0(n1692), .C0(n1693), .Y(n3230)
         );
  AOI22XLTS U7267 ( .A0(\dataToWriteBuffer[0][12] ), .A1(n5447), .B0(n4351), 
        .B1(n5432), .Y(n1692) );
  AOI222XLTS U7268 ( .A0(cacheDataIn_A[12]), .A1(n5612), .B0(n3992), .B1(n5481), .C0(n4206), .C1(n5468), .Y(n1693) );
  OAI211X1TS U7269 ( .A0(n5496), .A1(n3915), .B0(n1694), .C0(n1695), .Y(n3231)
         );
  AOI22XLTS U7270 ( .A0(\dataToWriteBuffer[0][13] ), .A1(n5447), .B0(n4356), 
        .B1(n5432), .Y(n1694) );
  AOI222XLTS U7271 ( .A0(cacheDataIn_A[13]), .A1(n5611), .B0(n3994), .B1(n5481), .C0(n4210), .C1(n5468), .Y(n1695) );
  OAI211X1TS U7272 ( .A0(n5496), .A1(n3917), .B0(n1696), .C0(n1697), .Y(n3232)
         );
  AOI22XLTS U7273 ( .A0(\dataToWriteBuffer[0][14] ), .A1(n5447), .B0(n4361), 
        .B1(n5432), .Y(n1696) );
  AOI222XLTS U7274 ( .A0(cacheDataIn_A[14]), .A1(n5607), .B0(n3996), .B1(n5481), .C0(n4214), .C1(n5468), .Y(n1697) );
  OAI211X1TS U7275 ( .A0(n5496), .A1(n3919), .B0(n1698), .C0(n1699), .Y(n3233)
         );
  AOI22XLTS U7276 ( .A0(\dataToWriteBuffer[0][15] ), .A1(n5447), .B0(n4366), 
        .B1(n5432), .Y(n1698) );
  AOI222XLTS U7277 ( .A0(cacheDataIn_A[15]), .A1(n5611), .B0(n3998), .B1(n5481), .C0(n4218), .C1(n5468), .Y(n1699) );
  OAI211X1TS U7278 ( .A0(n5502), .A1(n3921), .B0(n1700), .C0(n1701), .Y(n3234)
         );
  AOI22XLTS U7279 ( .A0(\dataToWriteBuffer[0][16] ), .A1(n5446), .B0(n4371), 
        .B1(n5439), .Y(n1700) );
  AOI222XLTS U7280 ( .A0(cacheDataIn_A[16]), .A1(n5614), .B0(n4000), .B1(n5482), .C0(n4222), .C1(n5467), .Y(n1701) );
  OAI211X1TS U7281 ( .A0(n5500), .A1(n3923), .B0(n1702), .C0(n1703), .Y(n3235)
         );
  AOI22XLTS U7282 ( .A0(\dataToWriteBuffer[0][17] ), .A1(n5446), .B0(n4376), 
        .B1(n1669), .Y(n1702) );
  AOI222XLTS U7283 ( .A0(cacheDataIn_A[17]), .A1(n5602), .B0(n4002), .B1(n5482), .C0(n4226), .C1(n5467), .Y(n1703) );
  OAI211X1TS U7284 ( .A0(n5502), .A1(n3925), .B0(n1704), .C0(n1705), .Y(n3236)
         );
  AOI22XLTS U7285 ( .A0(\dataToWriteBuffer[0][18] ), .A1(n5446), .B0(n4381), 
        .B1(n1669), .Y(n1704) );
  AOI222XLTS U7286 ( .A0(cacheDataIn_A[18]), .A1(n5602), .B0(n4004), .B1(n5482), .C0(n4230), .C1(n5467), .Y(n1705) );
  OAI211X1TS U7287 ( .A0(n5502), .A1(n3927), .B0(n1706), .C0(n1707), .Y(n3237)
         );
  AOI22XLTS U7288 ( .A0(\dataToWriteBuffer[0][19] ), .A1(n5446), .B0(n4386), 
        .B1(n5438), .Y(n1706) );
  AOI222XLTS U7289 ( .A0(cacheDataIn_A[19]), .A1(n5602), .B0(n4006), .B1(n5482), .C0(n4234), .C1(n5467), .Y(n1707) );
  OAI211X1TS U7290 ( .A0(n5495), .A1(n3929), .B0(n1708), .C0(n1709), .Y(n3238)
         );
  AOI22XLTS U7291 ( .A0(\dataToWriteBuffer[0][20] ), .A1(n5445), .B0(n4391), 
        .B1(n5439), .Y(n1708) );
  AOI222XLTS U7292 ( .A0(cacheDataIn_A[20]), .A1(n5603), .B0(n4008), .B1(n5483), .C0(n4238), .C1(n5474), .Y(n1709) );
  OAI211X1TS U7293 ( .A0(n5495), .A1(n3931), .B0(n1710), .C0(n1711), .Y(n3239)
         );
  AOI22XLTS U7294 ( .A0(\dataToWriteBuffer[0][21] ), .A1(n5445), .B0(n4396), 
        .B1(n5436), .Y(n1710) );
  AOI222XLTS U7295 ( .A0(cacheDataIn_A[21]), .A1(n5603), .B0(n4010), .B1(n5483), .C0(n4242), .C1(n5474), .Y(n1711) );
  OAI211X1TS U7296 ( .A0(n5495), .A1(n3933), .B0(n1712), .C0(n1713), .Y(n3240)
         );
  AOI22XLTS U7297 ( .A0(\dataToWriteBuffer[0][22] ), .A1(n5445), .B0(n4401), 
        .B1(n5438), .Y(n1712) );
  AOI222XLTS U7298 ( .A0(cacheDataIn_A[22]), .A1(n5603), .B0(n4012), .B1(n5483), .C0(n4246), .C1(n5472), .Y(n1713) );
  OAI211X1TS U7299 ( .A0(n5495), .A1(n3935), .B0(n1714), .C0(n1715), .Y(n3241)
         );
  AOI22XLTS U7300 ( .A0(\dataToWriteBuffer[0][23] ), .A1(n5445), .B0(n4406), 
        .B1(n5437), .Y(n1714) );
  AOI222XLTS U7301 ( .A0(cacheDataIn_A[23]), .A1(n5603), .B0(n4014), .B1(n5483), .C0(n4250), .C1(n5473), .Y(n1715) );
  OAI211X1TS U7302 ( .A0(n5494), .A1(n3937), .B0(n1716), .C0(n1717), .Y(n3242)
         );
  AOI22XLTS U7303 ( .A0(\dataToWriteBuffer[0][24] ), .A1(n5444), .B0(n4411), 
        .B1(n5440), .Y(n1716) );
  AOI222XLTS U7304 ( .A0(cacheDataIn_A[24]), .A1(n5604), .B0(n4016), .B1(n5488), .C0(n4254), .C1(n5475), .Y(n1717) );
  OAI211X1TS U7305 ( .A0(n5494), .A1(n3939), .B0(n1718), .C0(n1719), .Y(n3243)
         );
  AOI22XLTS U7306 ( .A0(\dataToWriteBuffer[0][25] ), .A1(n5444), .B0(n4416), 
        .B1(n5436), .Y(n1718) );
  AOI222XLTS U7307 ( .A0(cacheDataIn_A[25]), .A1(n5604), .B0(n4018), .B1(n5488), .C0(n4258), .C1(n5475), .Y(n1719) );
  OAI211X1TS U7308 ( .A0(n5494), .A1(n3941), .B0(n1720), .C0(n1721), .Y(n3244)
         );
  AOI22XLTS U7309 ( .A0(\dataToWriteBuffer[0][26] ), .A1(n5444), .B0(n4421), 
        .B1(n5440), .Y(n1720) );
  AOI222XLTS U7310 ( .A0(cacheDataIn_A[26]), .A1(n5604), .B0(n4020), .B1(n5489), .C0(n4262), .C1(n5472), .Y(n1721) );
  OAI211X1TS U7311 ( .A0(n5494), .A1(n3943), .B0(n1722), .C0(n1723), .Y(n3245)
         );
  AOI22XLTS U7312 ( .A0(\dataToWriteBuffer[0][27] ), .A1(n5444), .B0(n4426), 
        .B1(n5437), .Y(n1722) );
  AOI222XLTS U7313 ( .A0(cacheDataIn_A[27]), .A1(n5604), .B0(n4022), .B1(n5489), .C0(n4266), .C1(n5473), .Y(n1723) );
  OAI211X1TS U7314 ( .A0(n5493), .A1(n3945), .B0(n1724), .C0(n1725), .Y(n3246)
         );
  AOI22XLTS U7315 ( .A0(\dataToWriteBuffer[0][28] ), .A1(n5443), .B0(n4431), 
        .B1(n5431), .Y(n1724) );
  AOI222XLTS U7316 ( .A0(cacheDataIn_A[28]), .A1(n5605), .B0(n4024), .B1(n5484), .C0(n4270), .C1(n5478), .Y(n1725) );
  OAI211X1TS U7317 ( .A0(n5493), .A1(n3947), .B0(n1726), .C0(n1727), .Y(n3247)
         );
  AOI22XLTS U7318 ( .A0(\dataToWriteBuffer[0][29] ), .A1(n5443), .B0(n4436), 
        .B1(n5431), .Y(n1726) );
  AOI222XLTS U7319 ( .A0(cacheDataIn_A[29]), .A1(n5605), .B0(n4026), .B1(n5484), .C0(n4274), .C1(n5475), .Y(n1727) );
  OAI211X1TS U7320 ( .A0(n5493), .A1(n3949), .B0(n1728), .C0(n1729), .Y(n3248)
         );
  AOI22XLTS U7321 ( .A0(\dataToWriteBuffer[0][30] ), .A1(n5443), .B0(n4441), 
        .B1(n5431), .Y(n1728) );
  AOI222XLTS U7322 ( .A0(cacheDataIn_A[30]), .A1(n5605), .B0(n4028), .B1(n5484), .C0(n4278), .C1(n5475), .Y(n1729) );
  OAI211X1TS U7323 ( .A0(n5493), .A1(n3951), .B0(n1730), .C0(n1731), .Y(n3249)
         );
  AOI22XLTS U7324 ( .A0(\dataToWriteBuffer[0][31] ), .A1(n5443), .B0(n4446), 
        .B1(n5431), .Y(n1730) );
  AOI222XLTS U7325 ( .A0(cacheDataIn_A[31]), .A1(n5605), .B0(n4030), .B1(n5484), .C0(n4282), .C1(n5474), .Y(n1731) );
  INVX2TS U7326 ( .A(n1547), .Y(n5655) );
  NAND2BX1TS U7327 ( .AN(n3645), .B(n3693), .Y(n1547) );
  NOR2XLTS U7328 ( .A(n4286), .B(n3966), .Y(n2421) );
  AOI22XLTS U7329 ( .A0(n3818), .A1(n4103), .B0(n4079), .B1(n3802), .Y(n1998)
         );
  AOI22XLTS U7330 ( .A0(n3819), .A1(n4106), .B0(n4082), .B1(n3803), .Y(n1994)
         );
  AOI22XLTS U7331 ( .A0(n3819), .A1(n4109), .B0(n4085), .B1(n3801), .Y(n1990)
         );
  AOI22XLTS U7332 ( .A0(n3818), .A1(n4112), .B0(n4088), .B1(n3802), .Y(n1986)
         );
  AOI22XLTS U7333 ( .A0(n3819), .A1(n4115), .B0(n4091), .B1(n3803), .Y(n1982)
         );
  AOI22XLTS U7334 ( .A0(n3818), .A1(n4117), .B0(n4093), .B1(n3802), .Y(n1978)
         );
  AOI22XLTS U7335 ( .A0(n3819), .A1(n4120), .B0(n4096), .B1(n3803), .Y(n1974)
         );
  AOI22XLTS U7336 ( .A0(n3818), .A1(n4124), .B0(n4100), .B1(n3801), .Y(n1969)
         );
  AOI22XLTS U7337 ( .A0(n3816), .A1(n4102), .B0(n4078), .B1(n3799), .Y(n2042)
         );
  AOI22XLTS U7338 ( .A0(n3817), .A1(n4105), .B0(n4081), .B1(n3800), .Y(n2038)
         );
  AOI22XLTS U7339 ( .A0(n3817), .A1(n4108), .B0(n4084), .B1(n3798), .Y(n2034)
         );
  AOI22XLTS U7340 ( .A0(n3816), .A1(n4111), .B0(n4087), .B1(n3799), .Y(n2030)
         );
  AOI22XLTS U7341 ( .A0(n3817), .A1(n4114), .B0(n4090), .B1(n3800), .Y(n2026)
         );
  AOI22XLTS U7342 ( .A0(n3816), .A1(n4118), .B0(n4094), .B1(n3799), .Y(n2022)
         );
  AOI22XLTS U7343 ( .A0(n3817), .A1(n4121), .B0(n4097), .B1(n3800), .Y(n2018)
         );
  AOI22XLTS U7344 ( .A0(n3816), .A1(n4123), .B0(n4099), .B1(n3798), .Y(n2013)
         );
  NAND3X1TS U7345 ( .A(n5668), .B(n1241), .C(prevRequesterPort_B[0]), .Y(n1539) );
  NAND3X1TS U7346 ( .A(n5642), .B(n1243), .C(n4523), .Y(n1548) );
  INVX2TS U7347 ( .A(n1538), .Y(n5681) );
  NAND2BX1TS U7348 ( .AN(n3646), .B(n3694), .Y(n1538) );
  OAI221XLTS U7349 ( .A0(n4576), .A1(n4031), .B0(n5797), .B1(n1272), .C0(n1582), .Y(n3190) );
  AOI222XLTS U7350 ( .A0(\requesterAddressBuffer[0][0] ), .A1(n3769), .B0(
        n3733), .B1(n1583), .C0(n4061), .C1(n3737), .Y(n1582) );
  AO22XLTS U7351 ( .A0(n4532), .A1(n3954), .B0(n4561), .B1(n3878), .Y(n1583)
         );
  OAI221XLTS U7352 ( .A0(n4576), .A1(n4033), .B0(n5797), .B1(n1271), .C0(n1580), .Y(n3189) );
  AOI222XLTS U7353 ( .A0(\requesterAddressBuffer[0][1] ), .A1(n3770), .B0(
        n3734), .B1(n1581), .C0(n4064), .C1(n3738), .Y(n1580) );
  AO22XLTS U7354 ( .A0(n5801), .A1(n3956), .B0(n4562), .B1(n3880), .Y(n1581)
         );
  OAI221XLTS U7355 ( .A0(n4576), .A1(n4035), .B0(n4540), .B1(n1270), .C0(n1578), .Y(n3188) );
  AOI222XLTS U7356 ( .A0(\requesterAddressBuffer[0][2] ), .A1(n3769), .B0(
        n3733), .B1(n1579), .C0(n4067), .C1(n3737), .Y(n1578) );
  AO22XLTS U7357 ( .A0(n4606), .A1(n3958), .B0(n4563), .B1(n3882), .Y(n1579)
         );
  OAI221XLTS U7358 ( .A0(n4576), .A1(n4037), .B0(n4540), .B1(n1269), .C0(n1576), .Y(n3187) );
  AOI222XLTS U7359 ( .A0(\requesterAddressBuffer[0][3] ), .A1(n3770), .B0(
        n3734), .B1(n1577), .C0(n4070), .C1(n3738), .Y(n1576) );
  AO22XLTS U7360 ( .A0(n4606), .A1(n3960), .B0(n4562), .B1(n3884), .Y(n1577)
         );
  OAI221XLTS U7361 ( .A0(n4577), .A1(n4039), .B0(n4540), .B1(n1268), .C0(n1574), .Y(n3186) );
  AOI222XLTS U7362 ( .A0(\requesterAddressBuffer[0][4] ), .A1(n3769), .B0(
        n3733), .B1(n1575), .C0(n4073), .C1(n3737), .Y(n1574) );
  AO22XLTS U7363 ( .A0(n4606), .A1(n3962), .B0(n4563), .B1(n3886), .Y(n1575)
         );
  OAI221XLTS U7364 ( .A0(n4577), .A1(n4041), .B0(n4540), .B1(n1267), .C0(n1568), .Y(n3185) );
  AOI222XLTS U7365 ( .A0(\requesterAddressBuffer[0][5] ), .A1(n3770), .B0(
        n3734), .B1(n1571), .C0(n4076), .C1(n3738), .Y(n1568) );
  AO22XLTS U7366 ( .A0(n4606), .A1(n3964), .B0(n4563), .B1(n3888), .Y(n1571)
         );
  OAI221XLTS U7367 ( .A0(n4558), .A1(n1278), .B0(n4584), .B1(n1249), .C0(n1614), .Y(n3202) );
  AOI22XLTS U7368 ( .A0(n3735), .A1(n1615), .B0(n3751), .B1(n4032), .Y(n1614)
         );
  AO22XLTS U7369 ( .A0(n4060), .A1(n5539), .B0(n5541), .B1(n3954), .Y(n1615)
         );
  INVX2TS U7370 ( .A(n5540), .Y(n5539) );
  OAI221XLTS U7371 ( .A0(n4558), .A1(n1277), .B0(n4583), .B1(n1248), .C0(n1612), .Y(n3201) );
  AOI22XLTS U7372 ( .A0(n3736), .A1(n1613), .B0(n1604), .B1(n4034), .Y(n1612)
         );
  AO22XLTS U7373 ( .A0(n4064), .A1(n5538), .B0(n5542), .B1(n3956), .Y(n1613)
         );
  OAI221XLTS U7374 ( .A0(n4558), .A1(n1276), .B0(n4584), .B1(n1247), .C0(n1610), .Y(n3200) );
  AOI22XLTS U7375 ( .A0(n3735), .A1(n1611), .B0(n3751), .B1(n4036), .Y(n1610)
         );
  AO22XLTS U7376 ( .A0(n4067), .A1(n5538), .B0(n5543), .B1(n3958), .Y(n1611)
         );
  OAI221XLTS U7377 ( .A0(n4559), .A1(n1275), .B0(n4583), .B1(n1246), .C0(n1608), .Y(n3199) );
  AOI22XLTS U7378 ( .A0(n3736), .A1(n1609), .B0(n1604), .B1(n4038), .Y(n1608)
         );
  AO22XLTS U7379 ( .A0(n4070), .A1(n5538), .B0(n5544), .B1(n3960), .Y(n1609)
         );
  OAI221XLTS U7380 ( .A0(n4559), .A1(n1274), .B0(n4584), .B1(n1245), .C0(n1606), .Y(n3198) );
  AOI22XLTS U7381 ( .A0(n3735), .A1(n1607), .B0(n3751), .B1(n4040), .Y(n1606)
         );
  AO22XLTS U7382 ( .A0(n4073), .A1(n5538), .B0(n5545), .B1(n3962), .Y(n1607)
         );
  OAI221XLTS U7383 ( .A0(n4559), .A1(n1273), .B0(n4583), .B1(n1244), .C0(n1601), .Y(n3197) );
  AOI22XLTS U7384 ( .A0(n3736), .A1(n1603), .B0(n1604), .B1(n4042), .Y(n1601)
         );
  AO22XLTS U7385 ( .A0(n4076), .A1(n5537), .B0(n5546), .B1(n3964), .Y(n1603)
         );
  OAI221XLTS U7386 ( .A0(n5457), .A1(n1232), .B0(n1642), .B1(n5519), .C0(n1644), .Y(n3209) );
  AOI22XLTS U7387 ( .A0(n4103), .A1(n5541), .B0(n4044), .B1(n5528), .Y(n1642)
         );
  AOI22XLTS U7388 ( .A0(n4128), .A1(n5513), .B0(cacheAddressIn_B[0]), .B1(
        n4657), .Y(n1644) );
  OAI221XLTS U7389 ( .A0(n5451), .A1(n1231), .B0(n1646), .B1(n5519), .C0(n1647), .Y(n3210) );
  AOI22XLTS U7390 ( .A0(n4106), .A1(n5541), .B0(n4046), .B1(n5528), .Y(n1646)
         );
  AOI22XLTS U7391 ( .A0(n4132), .A1(n5513), .B0(cacheAddressIn_B[1]), .B1(
        n4650), .Y(n1647) );
  OAI221XLTS U7392 ( .A0(n5451), .A1(n1230), .B0(n1648), .B1(n5519), .C0(n1649), .Y(n3211) );
  AOI22XLTS U7393 ( .A0(n4109), .A1(n5542), .B0(n4048), .B1(n5528), .Y(n1648)
         );
  AOI22XLTS U7394 ( .A0(n4136), .A1(n5512), .B0(cacheAddressIn_B[2]), .B1(
        n4650), .Y(n1649) );
  OAI221XLTS U7395 ( .A0(n5452), .A1(n1229), .B0(n1650), .B1(n5519), .C0(n1651), .Y(n3212) );
  AOI22XLTS U7396 ( .A0(n4112), .A1(n5542), .B0(n4050), .B1(n5528), .Y(n1650)
         );
  AOI22XLTS U7397 ( .A0(n4140), .A1(n5512), .B0(cacheAddressIn_B[3]), .B1(
        n4651), .Y(n1651) );
  OAI221XLTS U7398 ( .A0(n5452), .A1(n1228), .B0(n1652), .B1(n5518), .C0(n1653), .Y(n3213) );
  AOI22XLTS U7399 ( .A0(n4115), .A1(n5543), .B0(n4052), .B1(n5529), .Y(n1652)
         );
  AOI22XLTS U7400 ( .A0(n4144), .A1(n5510), .B0(cacheAddressIn_B[4]), .B1(
        n4651), .Y(n1653) );
  OAI221XLTS U7401 ( .A0(n5452), .A1(n1227), .B0(n1654), .B1(n5518), .C0(n1655), .Y(n3214) );
  AOI22XLTS U7402 ( .A0(n4118), .A1(n5543), .B0(n4054), .B1(n5529), .Y(n1654)
         );
  AOI22XLTS U7403 ( .A0(n4148), .A1(n5510), .B0(cacheAddressIn_B[5]), .B1(
        n4651), .Y(n1655) );
  OAI221XLTS U7404 ( .A0(n5453), .A1(n1226), .B0(n1656), .B1(n5518), .C0(n1657), .Y(n3215) );
  AOI22XLTS U7405 ( .A0(n4121), .A1(n5544), .B0(n4056), .B1(n5532), .Y(n1656)
         );
  AOI22XLTS U7406 ( .A0(n4152), .A1(n5510), .B0(cacheAddressIn_B[6]), .B1(
        n4651), .Y(n1657) );
  OAI221XLTS U7407 ( .A0(n5453), .A1(n1225), .B0(n1658), .B1(n5518), .C0(n1659), .Y(n3216) );
  AOI22XLTS U7408 ( .A0(n4124), .A1(n5544), .B0(n4058), .B1(n5529), .Y(n1658)
         );
  AOI22XLTS U7409 ( .A0(n4156), .A1(n5510), .B0(cacheAddressIn_B[7]), .B1(
        n4652), .Y(n1659) );
  OAI221XLTS U7410 ( .A0(n5453), .A1(n1135), .B0(n2133), .B1(n5517), .C0(n2134), .Y(n3346) );
  AOI22XLTS U7411 ( .A0(n3968), .A1(n5545), .B0(n4290), .B1(n5529), .Y(n2133)
         );
  AOI22XLTS U7412 ( .A0(n4160), .A1(n5509), .B0(cacheDataIn_B[0]), .B1(n4652), 
        .Y(n2134) );
  OAI221XLTS U7413 ( .A0(n5454), .A1(n1134), .B0(n2135), .B1(n5517), .C0(n2136), .Y(n3347) );
  AOI22XLTS U7414 ( .A0(n3970), .A1(n5545), .B0(n4295), .B1(n5530), .Y(n2135)
         );
  AOI22XLTS U7415 ( .A0(n4164), .A1(n5509), .B0(cacheDataIn_B[1]), .B1(n4652), 
        .Y(n2136) );
  OAI221XLTS U7416 ( .A0(n5454), .A1(n1133), .B0(n2137), .B1(n5517), .C0(n2138), .Y(n3348) );
  AOI22XLTS U7417 ( .A0(n3972), .A1(n5546), .B0(n4300), .B1(n5530), .Y(n2137)
         );
  AOI22XLTS U7418 ( .A0(n4168), .A1(n5509), .B0(cacheDataIn_B[2]), .B1(n4652), 
        .Y(n2138) );
  OAI221XLTS U7419 ( .A0(n5454), .A1(n1132), .B0(n2139), .B1(n5517), .C0(n2140), .Y(n3349) );
  AOI22XLTS U7420 ( .A0(n3974), .A1(n5546), .B0(n4305), .B1(n5530), .Y(n2139)
         );
  AOI22XLTS U7421 ( .A0(n4172), .A1(n5509), .B0(cacheDataIn_B[3]), .B1(n4653), 
        .Y(n2140) );
  OAI221XLTS U7422 ( .A0(n5455), .A1(n1131), .B0(n2141), .B1(n5516), .C0(n2142), .Y(n3350) );
  AOI22XLTS U7423 ( .A0(n3976), .A1(n5547), .B0(n4310), .B1(n5530), .Y(n2141)
         );
  AOI22XLTS U7424 ( .A0(n4176), .A1(n5508), .B0(cacheDataIn_B[4]), .B1(n4653), 
        .Y(n2142) );
  OAI221XLTS U7425 ( .A0(n5455), .A1(n1130), .B0(n2143), .B1(n5516), .C0(n2144), .Y(n3351) );
  AOI22XLTS U7426 ( .A0(n3978), .A1(n5547), .B0(n4315), .B1(n5531), .Y(n2143)
         );
  AOI22XLTS U7427 ( .A0(n4180), .A1(n5508), .B0(cacheDataIn_B[5]), .B1(n4653), 
        .Y(n2144) );
  OAI221XLTS U7428 ( .A0(n5455), .A1(n1129), .B0(n2145), .B1(n5516), .C0(n2146), .Y(n3352) );
  AOI22XLTS U7429 ( .A0(n3980), .A1(n5548), .B0(n4320), .B1(n5531), .Y(n2145)
         );
  AOI22XLTS U7430 ( .A0(n4184), .A1(n5508), .B0(cacheDataIn_B[6]), .B1(n4653), 
        .Y(n2146) );
  OAI221XLTS U7431 ( .A0(n5456), .A1(n1128), .B0(n2147), .B1(n5516), .C0(n2148), .Y(n3353) );
  AOI22XLTS U7432 ( .A0(n3982), .A1(n5548), .B0(n4325), .B1(n5531), .Y(n2147)
         );
  AOI22XLTS U7433 ( .A0(n4188), .A1(n5508), .B0(cacheDataIn_B[7]), .B1(n4654), 
        .Y(n2148) );
  OAI221XLTS U7434 ( .A0(n5456), .A1(n1127), .B0(n2149), .B1(n5515), .C0(n2150), .Y(n3354) );
  AOI22XLTS U7435 ( .A0(n3984), .A1(n5557), .B0(n4330), .B1(n5531), .Y(n2149)
         );
  AOI22XLTS U7436 ( .A0(n4192), .A1(n5511), .B0(cacheDataIn_B[8]), .B1(n4654), 
        .Y(n2150) );
  OAI221XLTS U7437 ( .A0(n5456), .A1(n1126), .B0(n2151), .B1(n5515), .C0(n2152), .Y(n3355) );
  AOI22XLTS U7438 ( .A0(n3986), .A1(n5557), .B0(n4335), .B1(n5532), .Y(n2151)
         );
  AOI22XLTS U7439 ( .A0(n4196), .A1(n5514), .B0(cacheDataIn_B[9]), .B1(n4654), 
        .Y(n2152) );
  OAI221XLTS U7440 ( .A0(n5457), .A1(n1125), .B0(n2153), .B1(n5515), .C0(n2154), .Y(n3356) );
  AOI22XLTS U7441 ( .A0(n3988), .A1(n5558), .B0(n4340), .B1(n5532), .Y(n2153)
         );
  AOI22XLTS U7442 ( .A0(n4200), .A1(n5514), .B0(cacheDataIn_B[10]), .B1(n4654), 
        .Y(n2154) );
  OAI221XLTS U7443 ( .A0(n5457), .A1(n1124), .B0(n2155), .B1(n5515), .C0(n2156), .Y(n3357) );
  AOI22XLTS U7444 ( .A0(n3990), .A1(n5548), .B0(n4345), .B1(n5532), .Y(n2155)
         );
  AOI22XLTS U7445 ( .A0(n4204), .A1(n5514), .B0(cacheDataIn_B[11]), .B1(n5798), 
        .Y(n2156) );
  OAI221XLTS U7446 ( .A0(n5458), .A1(n1123), .B0(n2157), .B1(n5521), .C0(n2158), .Y(n3358) );
  AOI22XLTS U7447 ( .A0(n3992), .A1(n5558), .B0(n4350), .B1(n5533), .Y(n2157)
         );
  AOI22XLTS U7448 ( .A0(n4208), .A1(n5507), .B0(cacheDataIn_B[12]), .B1(n4660), 
        .Y(n2158) );
  OAI221XLTS U7449 ( .A0(n5458), .A1(n1122), .B0(n2159), .B1(n5522), .C0(n2160), .Y(n3359) );
  AOI22XLTS U7450 ( .A0(n3994), .A1(n5556), .B0(n4355), .B1(n5533), .Y(n2159)
         );
  AOI22XLTS U7451 ( .A0(n4212), .A1(n5507), .B0(cacheDataIn_B[13]), .B1(n4660), 
        .Y(n2160) );
  OAI221XLTS U7452 ( .A0(n5458), .A1(n1121), .B0(n2161), .B1(n1643), .C0(n2162), .Y(n3360) );
  AOI22XLTS U7453 ( .A0(n3996), .A1(n5556), .B0(n4360), .B1(n5533), .Y(n2161)
         );
  AOI22XLTS U7454 ( .A0(n4216), .A1(n5507), .B0(cacheDataIn_B[14]), .B1(n4657), 
        .Y(n2162) );
  OAI221XLTS U7455 ( .A0(n5459), .A1(n1120), .B0(n2163), .B1(n1643), .C0(n2164), .Y(n3361) );
  AOI22XLTS U7456 ( .A0(n3998), .A1(n5549), .B0(n4365), .B1(n5533), .Y(n2163)
         );
  AOI22XLTS U7457 ( .A0(n4220), .A1(n5507), .B0(cacheDataIn_B[15]), .B1(n4662), 
        .Y(n2164) );
  OAI221XLTS U7458 ( .A0(n5459), .A1(n1119), .B0(n2165), .B1(n5523), .C0(n2166), .Y(n3362) );
  AOI22XLTS U7459 ( .A0(n4000), .A1(n5549), .B0(n4370), .B1(n5534), .Y(n2165)
         );
  AOI22XLTS U7460 ( .A0(n4224), .A1(n5506), .B0(cacheDataIn_B[16]), .B1(n4661), 
        .Y(n2166) );
  OAI221XLTS U7461 ( .A0(n5459), .A1(n1118), .B0(n2167), .B1(n5523), .C0(n2168), .Y(n3363) );
  AOI22XLTS U7462 ( .A0(n4002), .A1(n5549), .B0(n4375), .B1(n5534), .Y(n2167)
         );
  AOI22XLTS U7463 ( .A0(n4228), .A1(n5506), .B0(cacheDataIn_B[17]), .B1(n5798), 
        .Y(n2168) );
  OAI221XLTS U7464 ( .A0(n5460), .A1(n1117), .B0(n2169), .B1(n5522), .C0(n2170), .Y(n3364) );
  AOI22XLTS U7465 ( .A0(n4004), .A1(n5549), .B0(n4380), .B1(n5534), .Y(n2169)
         );
  AOI22XLTS U7466 ( .A0(n4232), .A1(n5506), .B0(cacheDataIn_B[18]), .B1(n4662), 
        .Y(n2170) );
  OAI221XLTS U7467 ( .A0(n5460), .A1(n1116), .B0(n2171), .B1(n5520), .C0(n2172), .Y(n3365) );
  AOI22XLTS U7468 ( .A0(n4006), .A1(n5550), .B0(n4385), .B1(n5534), .Y(n2171)
         );
  AOI22XLTS U7469 ( .A0(n4236), .A1(n5506), .B0(cacheDataIn_B[19]), .B1(n4657), 
        .Y(n2172) );
  OAI221XLTS U7470 ( .A0(n5460), .A1(n1115), .B0(n2173), .B1(n5523), .C0(n2174), .Y(n3366) );
  AOI22XLTS U7471 ( .A0(n4008), .A1(n5550), .B0(n4390), .B1(n5535), .Y(n2173)
         );
  AOI22XLTS U7472 ( .A0(n4240), .A1(n5505), .B0(cacheDataIn_B[20]), .B1(n4662), 
        .Y(n2174) );
  OAI221XLTS U7473 ( .A0(n5461), .A1(n1114), .B0(n2175), .B1(n5523), .C0(n2176), .Y(n3367) );
  AOI22XLTS U7474 ( .A0(n4010), .A1(n5550), .B0(n4395), .B1(n5535), .Y(n2175)
         );
  AOI22XLTS U7475 ( .A0(n4244), .A1(n5505), .B0(cacheDataIn_B[21]), .B1(n4659), 
        .Y(n2176) );
  OAI221XLTS U7476 ( .A0(n5461), .A1(n1113), .B0(n2177), .B1(n5520), .C0(n2178), .Y(n3368) );
  AOI22XLTS U7477 ( .A0(n4012), .A1(n5551), .B0(n4400), .B1(n5535), .Y(n2177)
         );
  AOI22XLTS U7478 ( .A0(n4248), .A1(n5505), .B0(cacheDataIn_B[22]), .B1(n4656), 
        .Y(n2178) );
  OAI221XLTS U7479 ( .A0(n5462), .A1(n1112), .B0(n2179), .B1(n5521), .C0(n2180), .Y(n3369) );
  AOI22XLTS U7480 ( .A0(n4014), .A1(n5550), .B0(n4405), .B1(n5535), .Y(n2179)
         );
  AOI22XLTS U7481 ( .A0(n4252), .A1(n5505), .B0(cacheDataIn_B[23]), .B1(n4656), 
        .Y(n2180) );
  OAI221XLTS U7482 ( .A0(n5462), .A1(n1111), .B0(n2181), .B1(n5524), .C0(n2182), .Y(n3370) );
  AOI22XLTS U7483 ( .A0(n4016), .A1(n4613), .B0(n4410), .B1(n5536), .Y(n2181)
         );
  AOI22XLTS U7484 ( .A0(n4256), .A1(n5504), .B0(cacheDataIn_B[24]), .B1(n4659), 
        .Y(n2182) );
  OAI221XLTS U7485 ( .A0(n5462), .A1(n1110), .B0(n2183), .B1(n5524), .C0(n2184), .Y(n3371) );
  AOI22XLTS U7486 ( .A0(n4018), .A1(n5551), .B0(n4415), .B1(n5536), .Y(n2183)
         );
  AOI22XLTS U7487 ( .A0(n4260), .A1(n5504), .B0(cacheDataIn_B[25]), .B1(n4655), 
        .Y(n2184) );
  OAI221XLTS U7488 ( .A0(n5461), .A1(n1109), .B0(n2185), .B1(n5525), .C0(n2186), .Y(n3372) );
  AOI22XLTS U7489 ( .A0(n4020), .A1(n5552), .B0(n4420), .B1(n5536), .Y(n2185)
         );
  AOI22XLTS U7490 ( .A0(n4264), .A1(n5504), .B0(cacheDataIn_B[26]), .B1(n4658), 
        .Y(n2186) );
  OAI221XLTS U7491 ( .A0(n5462), .A1(n1108), .B0(n2187), .B1(n5522), .C0(n2188), .Y(n3373) );
  AOI22XLTS U7492 ( .A0(n4022), .A1(n5551), .B0(n4425), .B1(n5536), .Y(n2187)
         );
  AOI22XLTS U7493 ( .A0(n4268), .A1(n5504), .B0(cacheDataIn_B[27]), .B1(n4655), 
        .Y(n2188) );
  OAI221XLTS U7494 ( .A0(n5463), .A1(n1107), .B0(n2189), .B1(n5526), .C0(n2190), .Y(n3374) );
  AOI22XLTS U7495 ( .A0(n4024), .A1(n5552), .B0(n4430), .B1(n5537), .Y(n2189)
         );
  AOI22XLTS U7496 ( .A0(n4272), .A1(n5503), .B0(cacheDataIn_B[28]), .B1(n4655), 
        .Y(n2190) );
  OAI221XLTS U7497 ( .A0(n5463), .A1(n1106), .B0(n2191), .B1(n5524), .C0(n2192), .Y(n3375) );
  AOI22XLTS U7498 ( .A0(n4026), .A1(n5552), .B0(n4435), .B1(n5537), .Y(n2191)
         );
  AOI22XLTS U7499 ( .A0(n4276), .A1(n5503), .B0(cacheDataIn_B[29]), .B1(n4656), 
        .Y(n2192) );
  OAI221XLTS U7500 ( .A0(n5461), .A1(n1105), .B0(n2193), .B1(n5524), .C0(n2194), .Y(n3376) );
  AOI22XLTS U7501 ( .A0(n4028), .A1(n5551), .B0(n4440), .B1(n5537), .Y(n2193)
         );
  AOI22XLTS U7502 ( .A0(n4280), .A1(n5503), .B0(cacheDataIn_B[30]), .B1(n4655), 
        .Y(n2194) );
  OAI221XLTS U7503 ( .A0(n5451), .A1(n1104), .B0(n2195), .B1(n5526), .C0(n2196), .Y(n3377) );
  AOI22XLTS U7504 ( .A0(n4030), .A1(n5540), .B0(n4445), .B1(n5527), .Y(n2195)
         );
  AOI22XLTS U7505 ( .A0(n4284), .A1(n5503), .B0(cacheDataIn_B[31]), .B1(n4650), 
        .Y(n2196) );
  OAI22XLTS U7506 ( .A0(n4288), .A1(n5802), .B0(n3730), .B1(n2102), .Y(n1566)
         );
  AOI22X1TS U7507 ( .A0(n2103), .A1(n3704), .B0(n3720), .B1(n3807), .Y(n2102)
         );
  OAI22XLTS U7508 ( .A0(n3692), .A1(n4562), .B0(n4532), .B1(n3684), .Y(n2103)
         );
  AOI22XLTS U7509 ( .A0(n2273), .A1(n1799), .B0(n3870), .B1(n3772), .Y(n2270)
         );
  OAI22X1TS U7510 ( .A0(n3821), .A1(n3741), .B0(n3827), .B1(n3753), .Y(n2273)
         );
  OAI22X1TS U7511 ( .A0(n1799), .A1(n5873), .B0(n3869), .B1(n2129), .Y(n2128)
         );
  AOI22XLTS U7512 ( .A0(n3688), .A1(n3654), .B0(n3826), .B1(n3682), .Y(n2129)
         );
  AOI22XLTS U7513 ( .A0(n3772), .A1(n5789), .B0(n2234), .B1(n1766), .Y(n2231)
         );
  OAI221XLTS U7514 ( .A0(n1770), .A1(n3753), .B0(n5781), .B1(n3741), .C0(n3716), .Y(n2234) );
  INVX2TS U7515 ( .A(n1770), .Y(n5781) );
  AOI22XLTS U7516 ( .A0(n3771), .A1(n5790), .B0(n2206), .B1(n1744), .Y(n2204)
         );
  OAI221XLTS U7517 ( .A0(n1749), .A1(n3752), .B0(n5782), .B1(n3683), .C0(n3715), .Y(n2206) );
  AOI22XLTS U7518 ( .A0(n3772), .A1(n5787), .B0(n2219), .B1(n1756), .Y(n2218)
         );
  OAI221XLTS U7519 ( .A0(n1760), .A1(n3753), .B0(n5779), .B1(n3741), .C0(n3716), .Y(n2219) );
  AOI22XLTS U7520 ( .A0(n3771), .A1(n5788), .B0(n2261), .B1(n1787), .Y(n2260)
         );
  OAI221XLTS U7521 ( .A0(n1791), .A1(n3752), .B0(n5780), .B1(n3683), .C0(n3715), .Y(n2261) );
  AOI22XLTS U7522 ( .A0(n3771), .A1(n5791), .B0(n2245), .B1(n1776), .Y(n2244)
         );
  OAI221XLTS U7523 ( .A0(n1780), .A1(n3752), .B0(n5784), .B1(n3741), .C0(n3715), .Y(n2245) );
  AOI211X1TS U7524 ( .A0(n1241), .A1(n4520), .B0(n5678), .C0(n5739), .Y(n1536)
         );
  AOI211X1TS U7525 ( .A0(n1243), .A1(n4523), .B0(n5652), .C0(n5740), .Y(n1545)
         );
  OAI211X1TS U7526 ( .A0(n4563), .A1(n1586), .B0(n4577), .C0(n1732), .Y(n3250)
         );
  AOI22X1TS U7527 ( .A0(\requesterPortBuffer[0][0] ), .A1(n3770), .B0(n3694), 
        .B1(n1733), .Y(n1732) );
  OAI211X1TS U7528 ( .A0(n3721), .A1(n1586), .B0(n4577), .C0(n1734), .Y(n3251)
         );
  AOI22X1TS U7529 ( .A0(\requesterPortBuffer[0][1] ), .A1(n3769), .B0(n3646), 
        .B1(n1733), .Y(n1734) );
  AOI211X1TS U7530 ( .A0(n1241), .A1(n1243), .B0(n4580), .C0(n5740), .Y(n1528)
         );
  AND2X2TS U7531 ( .A(n3646), .B(n3694), .Y(n4615) );
  NAND3X1TS U7532 ( .A(n4520), .B(n5615), .C(prevRequesterPort_B[1]), .Y(n3157) );
  OAI2BB2XLTS U7533 ( .B0(n5734), .B1(n1527), .A0N(
        requesterAddressOut_NORTH[0]), .A1N(n1528), .Y(n3160) );
  AOI22X1TS U7534 ( .A0(prevRequesterAddress_B[0]), .A1(n1529), .B0(
        prevRequesterAddress_A[0]), .B1(n4581), .Y(n1527) );
  OAI2BB2XLTS U7535 ( .B0(n5737), .B1(n1531), .A0N(
        requesterAddressOut_NORTH[1]), .A1N(n1528), .Y(n3161) );
  AOI22X1TS U7536 ( .A0(prevRequesterAddress_B[1]), .A1(n1529), .B0(
        prevRequesterAddress_A[1]), .B1(n4580), .Y(n1531) );
  OAI2BB2XLTS U7537 ( .B0(n5732), .B1(n1532), .A0N(
        requesterAddressOut_NORTH[2]), .A1N(n1528), .Y(n3162) );
  AOI22X1TS U7538 ( .A0(prevRequesterAddress_B[2]), .A1(n1529), .B0(
        prevRequesterAddress_A[2]), .B1(n4581), .Y(n1532) );
  OAI2BB2XLTS U7539 ( .B0(n5736), .B1(n1533), .A0N(
        requesterAddressOut_NORTH[3]), .A1N(n4537), .Y(n3163) );
  AOI22X1TS U7540 ( .A0(prevRequesterAddress_B[3]), .A1(n4551), .B0(
        prevRequesterAddress_A[3]), .B1(n4580), .Y(n1533) );
  OAI2BB2XLTS U7541 ( .B0(n5729), .B1(n1534), .A0N(
        requesterAddressOut_NORTH[4]), .A1N(n4537), .Y(n3164) );
  AOI22X1TS U7542 ( .A0(prevRequesterAddress_B[4]), .A1(n4551), .B0(
        prevRequesterAddress_A[4]), .B1(n4581), .Y(n1534) );
  OAI2BB2XLTS U7543 ( .B0(n5734), .B1(n1535), .A0N(
        requesterAddressOut_NORTH[5]), .A1N(n4537), .Y(n3165) );
  AOI22X1TS U7544 ( .A0(prevRequesterAddress_B[5]), .A1(n4551), .B0(
        prevRequesterAddress_A[5]), .B1(n4580), .Y(n1535) );
  NAND3BX1TS U7545 ( .AN(n2214), .B(n3873), .C(n5709), .Y(n2239) );
  OAI2BB2XLTS U7546 ( .B0(n1563), .B1(n1564), .A0N(memWrite_A), .A1N(n5613), 
        .Y(n3184) );
  AOI221X1TS U7547 ( .A0(n5582), .A1(n1174), .B0(n5594), .B1(n1566), .C0(n5732), .Y(n1564) );
  OA22XLTS U7548 ( .A0(n3727), .A1(n2123), .B0(n4287), .B1(n5805), .Y(n1662)
         );
  AOI22X1TS U7549 ( .A0(n5540), .A1(n3752), .B0(n5527), .B1(n3808), .Y(n2123)
         );
  AOI21X1TS U7550 ( .A0(n5784), .A1(n4599), .B0(n2252), .Y(n2248) );
  OAI31X1TS U7551 ( .A0(n5713), .A1(n5778), .A2(n4621), .B0(n1776), .Y(n2252)
         );
  OAI211X1TS U7552 ( .A0(n1616), .A1(n5807), .B0(n3750), .C0(n1793), .Y(n3265)
         );
  OA22X1TS U7553 ( .A0(n1243), .A1(n4583), .B0(n1262), .B1(n4558), .Y(n1793)
         );
  NAND2X1TS U7554 ( .A(n5718), .B(n2277), .Y(n2131) );
  OAI31X1TS U7555 ( .A0(n2278), .A1(n3868), .A2(n3820), .B0(n5585), .Y(n2277)
         );
  NOR3X1TS U7556 ( .A(n3874), .B(n5703), .C(n5778), .Y(n2278) );
  AO22X1TS U7557 ( .A0(requesterAddressOut_SOUTH[0]), .A1(n1536), .B0(n1537), 
        .B1(n5726), .Y(n3166) );
  OAI22X1TS U7558 ( .A0(n1272), .A1(n5676), .B0(n1249), .B1(n5660), .Y(n1537)
         );
  AO22X1TS U7559 ( .A0(requesterAddressOut_SOUTH[1]), .A1(n1536), .B0(n1540), 
        .B1(n5726), .Y(n3167) );
  OAI22X1TS U7560 ( .A0(n1271), .A1(n5677), .B0(n1248), .B1(n5660), .Y(n1540)
         );
  AO22X1TS U7561 ( .A0(requesterAddressOut_SOUTH[2]), .A1(n1536), .B0(n1541), 
        .B1(n5725), .Y(n3168) );
  OAI22X1TS U7562 ( .A0(n1270), .A1(n5677), .B0(n1247), .B1(n5660), .Y(n1541)
         );
  AO22X1TS U7563 ( .A0(requesterAddressOut_SOUTH[3]), .A1(n4571), .B0(n1542), 
        .B1(n5726), .Y(n3169) );
  OAI22X1TS U7564 ( .A0(n1269), .A1(n5677), .B0(n1246), .B1(n5659), .Y(n1542)
         );
  AO22X1TS U7565 ( .A0(requesterAddressOut_SOUTH[4]), .A1(n4571), .B0(n1543), 
        .B1(n5725), .Y(n3170) );
  OAI22X1TS U7566 ( .A0(n1268), .A1(n5677), .B0(n1245), .B1(n5659), .Y(n1543)
         );
  AO22X1TS U7567 ( .A0(requesterAddressOut_SOUTH[5]), .A1(n4571), .B0(n1544), 
        .B1(n5725), .Y(n3171) );
  OAI22X1TS U7568 ( .A0(n1267), .A1(n5676), .B0(n1244), .B1(n5659), .Y(n1544)
         );
  AO22X1TS U7569 ( .A0(requesterAddressOut_EAST[0]), .A1(n1545), .B0(n1546), 
        .B1(n5727), .Y(n3172) );
  OAI22X1TS U7570 ( .A0(n1272), .A1(n5650), .B0(n1249), .B1(n5637), .Y(n1546)
         );
  AO22X1TS U7571 ( .A0(requesterAddressOut_EAST[1]), .A1(n1545), .B0(n1549), 
        .B1(n5725), .Y(n3173) );
  OAI22X1TS U7572 ( .A0(n1271), .A1(n5651), .B0(n1248), .B1(n5637), .Y(n1549)
         );
  AO22X1TS U7573 ( .A0(requesterAddressOut_EAST[2]), .A1(n1545), .B0(n1550), 
        .B1(n5727), .Y(n3174) );
  OAI22X1TS U7574 ( .A0(n1270), .A1(n5651), .B0(n1247), .B1(n5637), .Y(n1550)
         );
  AO22X1TS U7575 ( .A0(requesterAddressOut_EAST[3]), .A1(n4530), .B0(n1551), 
        .B1(n3875), .Y(n3175) );
  OAI22X1TS U7576 ( .A0(n1269), .A1(n5651), .B0(n1246), .B1(n5639), .Y(n1551)
         );
  AO22X1TS U7577 ( .A0(requesterAddressOut_EAST[4]), .A1(n4530), .B0(n1552), 
        .B1(n5724), .Y(n3176) );
  OAI22X1TS U7578 ( .A0(n1268), .A1(n5651), .B0(n1245), .B1(n5640), .Y(n1552)
         );
  AO22X1TS U7579 ( .A0(requesterAddressOut_EAST[5]), .A1(n4530), .B0(n1553), 
        .B1(n3875), .Y(n3177) );
  OAI22X1TS U7580 ( .A0(n1267), .A1(n5650), .B0(n1244), .B1(n5639), .Y(n1553)
         );
  AO22X1TS U7581 ( .A0(requesterAddressOut_WEST[0]), .A1(n1554), .B0(n1555), 
        .B1(n1556), .Y(n3178) );
  OAI22X1TS U7582 ( .A0(n1272), .A1(n5623), .B0(n5627), .B1(n1249), .Y(n1556)
         );
  AO22X1TS U7583 ( .A0(requesterAddressOut_WEST[1]), .A1(n3743), .B0(n1555), 
        .B1(n1558), .Y(n3179) );
  OAI22X1TS U7584 ( .A0(n1271), .A1(n5624), .B0(n5627), .B1(n1248), .Y(n1558)
         );
  AO22X1TS U7585 ( .A0(requesterAddressOut_WEST[2]), .A1(n1554), .B0(n1555), 
        .B1(n1559), .Y(n3180) );
  OAI22X1TS U7586 ( .A0(n1270), .A1(n5624), .B0(n5626), .B1(n1247), .Y(n1559)
         );
  AO22X1TS U7587 ( .A0(requesterAddressOut_WEST[3]), .A1(n3743), .B0(n4570), 
        .B1(n1560), .Y(n3181) );
  OAI22X1TS U7588 ( .A0(n1269), .A1(n5624), .B0(n5627), .B1(n1246), .Y(n1560)
         );
  AO22X1TS U7589 ( .A0(requesterAddressOut_WEST[4]), .A1(n1554), .B0(n4570), 
        .B1(n1561), .Y(n3182) );
  OAI22X1TS U7590 ( .A0(n1268), .A1(n5624), .B0(n5626), .B1(n1245), .Y(n1561)
         );
  AO22X1TS U7591 ( .A0(requesterAddressOut_WEST[5]), .A1(n3743), .B0(n4570), 
        .B1(n1562), .Y(n3183) );
  OAI22X1TS U7592 ( .A0(n1267), .A1(n5623), .B0(n5626), .B1(n1244), .Y(n1562)
         );
  AO22X1TS U7593 ( .A0(memWrite_B), .A1(n4656), .B0(n1660), .B1(n1661), .Y(
        n3217) );
  OAI221XLTS U7594 ( .A0(n1662), .A1(n5583), .B0(isWrite[1]), .B1(n5594), .C0(
        n5727), .Y(n1660) );
  OAI32X1TS U7595 ( .A0(n4550), .A1(n5800), .A2(n2101), .B0(n5463), .B1(n1176), 
        .Y(n3342) );
  INVX2TS U7596 ( .A(n1566), .Y(n5800) );
  OAI32X1TS U7597 ( .A0(n2122), .A1(n1662), .A2(n2101), .B0(n5463), .B1(n1175), 
        .Y(n3344) );
  OAI21X1TS U7598 ( .A0(n4525), .A1(n5806), .B0(n4538), .Y(n2122) );
  INVX2TS U7599 ( .A(totalAccesses[0]), .Y(n5806) );
  AOI211X1TS U7600 ( .A0(n5779), .A1(n4597), .B0(n5787), .C0(n2226), .Y(n2222)
         );
  NOR3X1TS U7601 ( .A(n2214), .B(n5703), .C(n3874), .Y(n2226) );
  OAI211X1TS U7602 ( .A0(n4559), .A1(n1261), .B0(n3750), .C0(n1792), .Y(n3264)
         );
  OA22X1TS U7603 ( .A0(n5540), .A1(n1616), .B0(n1241), .B1(n4584), .Y(n1792)
         );
  NAND2X1TS U7604 ( .A(prevMemRead_B), .B(n5721), .Y(n3158) );
  NAND2X1TS U7605 ( .A(prevMemRead_A), .B(n5722), .Y(n3159) );
  OAI2BB2XLTS U7606 ( .B0(n5873), .B1(n2110), .A0N(n4616), .A1N(n2110), .Y(
        n2108) );
  NAND2X1TS U7607 ( .A(n2111), .B(n4590), .Y(n2110) );
  CLKBUFX2TS U7608 ( .A(N651), .Y(n5700) );
  INVXLTS U7609 ( .A(n3686), .Y(n5873) );
  CLKBUFX2TS U7610 ( .A(N650), .Y(n5716) );
  CLKBUFX2TS U7611 ( .A(N651), .Y(n5701) );
  INVXLTS U7612 ( .A(n4290), .Y(n5906) );
  INVXLTS U7613 ( .A(n4295), .Y(n5905) );
  INVXLTS U7614 ( .A(n4300), .Y(n5904) );
  INVXLTS U7615 ( .A(n4305), .Y(n5903) );
  INVXLTS U7616 ( .A(n4310), .Y(n5902) );
  INVXLTS U7617 ( .A(n4315), .Y(n5901) );
  INVXLTS U7618 ( .A(n4320), .Y(n5900) );
  INVXLTS U7619 ( .A(n4325), .Y(n5899) );
  INVXLTS U7620 ( .A(n4330), .Y(n5898) );
  INVXLTS U7621 ( .A(n4335), .Y(n5897) );
  INVXLTS U7622 ( .A(n4340), .Y(n5896) );
  INVXLTS U7623 ( .A(n4345), .Y(n5895) );
  INVXLTS U7624 ( .A(n4350), .Y(n5894) );
  INVXLTS U7625 ( .A(n4355), .Y(n5893) );
  INVXLTS U7626 ( .A(n4360), .Y(n5892) );
  INVXLTS U7627 ( .A(n4365), .Y(n5891) );
  INVXLTS U7628 ( .A(n4370), .Y(n5890) );
  INVXLTS U7629 ( .A(n4375), .Y(n5889) );
  INVXLTS U7630 ( .A(n4380), .Y(n5888) );
  INVXLTS U7631 ( .A(n4385), .Y(n5887) );
  INVXLTS U7632 ( .A(n4390), .Y(n5886) );
  INVXLTS U7633 ( .A(n4395), .Y(n5885) );
  INVXLTS U7634 ( .A(n4400), .Y(n5884) );
  INVXLTS U7635 ( .A(n4405), .Y(n5883) );
  INVXLTS U7636 ( .A(n4410), .Y(n5882) );
  INVXLTS U7637 ( .A(n4415), .Y(n5881) );
  INVXLTS U7638 ( .A(n4420), .Y(n5880) );
  INVXLTS U7639 ( .A(n4425), .Y(n5879) );
  INVXLTS U7640 ( .A(n4430), .Y(n5878) );
  INVXLTS U7641 ( .A(n4435), .Y(n5877) );
  INVXLTS U7642 ( .A(n4440), .Y(n5876) );
  INVXLTS U7643 ( .A(n4445), .Y(n5875) );
  CLKBUFX2TS U7644 ( .A(N650), .Y(n5717) );
  CLKBUFX2TS U7645 ( .A(n880), .Y(n5695) );
  XOR2X1TS U7646 ( .A(N6701), .B(\add_0_root_sub_278_I2/carry [4]), .Y(N6622)
         );
  AND2X1TS U7647 ( .A(\add_0_root_sub_278_I2/carry [3]), .B(N6701), .Y(
        \add_0_root_sub_278_I2/carry [4]) );
  XOR2X1TS U7648 ( .A(N6701), .B(\add_0_root_sub_278_I2/carry [3]), .Y(N6621)
         );
  AND2X1TS U7649 ( .A(\add_0_root_sub_278_I2/carry [2]), .B(
        \add_0_root_sub_278_I2/B[2] ), .Y(\add_0_root_sub_278_I2/carry [3]) );
  XOR2X1TS U7650 ( .A(n4578), .B(\add_0_root_sub_278_I2/carry [2]), .Y(N6620)
         );
  AND2X1TS U7651 ( .A(\add_0_root_sub_278_I2/carry [1]), .B(n5706), .Y(
        \add_0_root_sub_278_I2/carry [2]) );
  XOR2X1TS U7652 ( .A(n5705), .B(\add_0_root_sub_278_I2/carry [1]), .Y(N6619)
         );
  AND2X1TS U7653 ( .A(n4546), .B(n4594), .Y(\add_0_root_sub_278_I2/carry [1])
         );
  XOR2X1TS U7654 ( .A(n4594), .B(n4546), .Y(N6618) );
  OR2X1TS U7655 ( .A(n5700), .B(n5715), .Y(\r1472/carry[3] ) );
  XNOR2X1TS U7656 ( .A(n5712), .B(n5697), .Y(N8209) );
  OR2X1TS U7657 ( .A(N651), .B(n5715), .Y(\r1467/carry[3] ) );
  XNOR2X1TS U7658 ( .A(n5712), .B(n5698), .Y(N6316) );
  OR2X1TS U7659 ( .A(n5698), .B(n5715), .Y(\r1471/carry[3] ) );
  OR2X1TS U7660 ( .A(N651), .B(n5714), .Y(\r1470/carry[3] ) );
  XNOR2X1TS U7661 ( .A(n5710), .B(n5699), .Y(N6699) );
  XOR2X1TS U7662 ( .A(N6318), .B(\add_0_root_sub_277_I2/carry [4]), .Y(N6375)
         );
  AND2X1TS U7663 ( .A(\add_0_root_sub_277_I2/carry [3]), .B(n4612), .Y(
        \add_0_root_sub_277_I2/carry [4]) );
  XOR2X1TS U7664 ( .A(N6318), .B(\add_0_root_sub_277_I2/carry [3]), .Y(N6374)
         );
  AND2X1TS U7665 ( .A(\add_0_root_sub_277_I2/carry [2]), .B(
        \add_0_root_sub_278_I2/B[2] ), .Y(\add_0_root_sub_277_I2/carry [3]) );
  XOR2X1TS U7666 ( .A(\add_0_root_sub_278_I2/B[2] ), .B(
        \add_0_root_sub_277_I2/carry [2]), .Y(N6373) );
  AND2X1TS U7667 ( .A(\add_0_root_sub_277_I2/carry [1]), .B(n5706), .Y(
        \add_0_root_sub_277_I2/carry [2]) );
  XOR2X1TS U7668 ( .A(n5704), .B(\add_0_root_sub_277_I2/carry [1]), .Y(N6372)
         );
  AND2X1TS U7669 ( .A(n4546), .B(n4593), .Y(\add_0_root_sub_277_I2/carry [1])
         );
  XOR2X1TS U7670 ( .A(n4594), .B(n4607), .Y(N6371) );
  XNOR2X1TS U7671 ( .A(n5710), .B(n5698), .Y(\add_0_root_sub_278_I2/B[2] ) );
  XOR2X1TS U7672 ( .A(n5807), .B(\add_0_root_r1459/carry [3]), .Y(
        \add_0_root_r1459/SUM[3] ) );
  AND2X1TS U7673 ( .A(n4593), .B(\add_0_root_r1459/B[0] ), .Y(
        \add_0_root_r1459/carry [1]) );
  XOR2X1TS U7674 ( .A(\add_0_root_r1459/B[0] ), .B(n4595), .Y(
        \add_0_root_r1459/SUM[0] ) );
  XOR2X1TS U7675 ( .A(n4548), .B(\add_0_root_r1463/carry [4]), .Y(
        \add_0_root_r1463/SUM[4] ) );
  AND2X1TS U7676 ( .A(\add_0_root_r1463/carry [3]), .B(\add_0_root_r1463/B[4] ), .Y(\add_0_root_r1463/carry [4]) );
  XOR2X1TS U7677 ( .A(n4548), .B(\add_0_root_r1463/carry [3]), .Y(
        \add_0_root_r1463/SUM[3] ) );
  XOR2X1TS U7678 ( .A(n4612), .B(\add_0_root_sub_0_root_sub_231/carry [4]), 
        .Y(N609) );
  AND2X1TS U7679 ( .A(\add_0_root_sub_0_root_sub_231/carry [3]), .B(n4612), 
        .Y(\add_0_root_sub_0_root_sub_231/carry [4]) );
  XOR2X1TS U7680 ( .A(n4612), .B(\add_0_root_sub_0_root_sub_231/carry [3]), 
        .Y(N608) );
  XNOR2X1TS U7681 ( .A(n5712), .B(n5698), .Y(
        \add_0_root_sub_0_root_sub_231/B[2] ) );
  AND2X1TS U7682 ( .A(totalAccesses[0]), .B(n4596), .Y(
        \add_0_root_sub_0_root_sub_231/carry [1]) );
  XOR2X1TS U7683 ( .A(n4594), .B(totalAccesses[0]), .Y(N605) );
  NAND3X1TS U7684 ( .A(N606), .B(N605), .C(N607), .Y(n5746) );
  NOR3BX1TS U7685 ( .AN(n5746), .B(N609), .C(N608), .Y(N610) );
endmodule

