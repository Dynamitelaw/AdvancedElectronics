##
## LEF for PtnCells ;
## created by Encounter v14.23-s044_1 on Wed Feb 27 22:15:21 2019
##

VERSION 5.5 ;

NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO lfsr1
  CLASS BLOCK ;
  SIZE 67.0000 BY 52.0000 ;
  FOREIGN lfsr1 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.86 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.682 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.7016 LAYER M3  ;
    ANTENNAMAXAREACAR 5.59473 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 20.969 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.0470146 LAYER VL  ;
    PORT
      LAYER M3 ;
        RECT 0.0000 10.9000 0.6000 11.1000 ;
    END
  END clk
  PIN resetn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.98 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.866 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.9648 LAYER M3  ;
    ANTENNAMAXAREACAR 19.492 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 75.3915 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.968523 LAYER VL  ;
    PORT
      LAYER M3 ;
        RECT 0.0000 14.9000 0.6000 15.1000 ;
    END
  END resetn
  PIN lfsr_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.12 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.644 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 2.44 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.176 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2552 LAYER M3  ;
    ANTENNAMAXAREACAR 3.40913 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 12.9484 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.358423 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 52.4000 0.0000 52.6000 0.6000 ;
    END
  END lfsr_out[27]
  PIN lfsr_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.14 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.018 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 2.4 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.176 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0896 LAYER M3  ;
    ANTENNAMAXAREACAR 6.06375 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 26.2548 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 50.9000 0.0000 51.1000 0.6000 ;
    END
  END lfsr_out[26]
  PIN lfsr_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.14 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.018 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 0.54 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.146 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0896 LAYER M3  ;
    ANTENNAMAXAREACAR 3.0443 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 12.5133 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.731155 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 49.4000 0.0000 49.6000 0.6000 ;
    END
  END lfsr_out[25]
  PIN lfsr_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.7 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.39 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 3.4 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.728 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0896 LAYER M3  ;
    ANTENNAMAXAREACAR 12.5371 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 50.0702 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 47.9000 0.0000 48.1000 0.6000 ;
    END
  END lfsr_out[24]
  PIN lfsr_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.7 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.538 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1136 LAYER M2  ;
    ANTENNAMAXAREACAR 5.91662 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 22.4156 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAMAXCUTCAR 0.526116 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 1.48 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.624 LAYER M3  ;
    ANTENNAGATEAREA 1.1712 LAYER M3  ;
    ANTENNAMAXAREACAR 7.18029 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 27.2175 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 46.4000 0.0000 46.6000 0.6000 ;
    END
  END lfsr_out[23]
  PIN lfsr_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.94 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.278 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2  ;
    ANTENNAMAXAREACAR 87.5417 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 324.882 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAMAXCUTCAR 1.38889 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 1.96 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.4 LAYER M3  ;
    ANTENNAGATEAREA 1.0896 LAYER M3  ;
    ANTENNAMAXAREACAR 89.3405 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 331.673 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 44.9000 0.0000 45.1000 0.6000 ;
    END
  END lfsr_out[22]
  PIN lfsr_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.37 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 3.98 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.022 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0896 LAYER M3  ;
    ANTENNAMAXAREACAR 10.2916 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 41.8978 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 43.4000 0.0000 43.6000 0.6000 ;
    END
  END lfsr_out[21]
  PIN lfsr_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.258 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 3.32 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.58 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0896 LAYER M3  ;
    ANTENNAMAXAREACAR 6.9081 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 29.3789 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 41.9000 0.0000 42.1000 0.6000 ;
    END
  END lfsr_out[20]
  PIN lfsr_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.48 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.176 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 2.04 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.696 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0896 LAYER M3  ;
    ANTENNAMAXAREACAR 15.4556 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 60.8687 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 40.4000 0.0000 40.6000 0.6000 ;
    END
  END lfsr_out[19]
  PIN lfsr_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.14 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.218 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 0.68 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.664 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0896 LAYER M3  ;
    ANTENNAMAXAREACAR 4.12726 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 16.5203 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.731155 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 38.9000 0.0000 39.1000 0.6000 ;
    END
  END lfsr_out[18]
  PIN lfsr_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.06 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.322 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 0.62 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.442 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0896 LAYER M3  ;
    ANTENNAMAXAREACAR 3.0443 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 12.5133 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.731155 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 37.4000 0.0000 37.6000 0.6000 ;
    END
  END lfsr_out[17]
  PIN lfsr_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.25 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 3.48 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.172 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2288 LAYER M3  ;
    ANTENNAMAXAREACAR 6.26179 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 24.5231 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.767866 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 35.9000 0.0000 36.1000 0.6000 ;
    END
  END lfsr_out[16]
  PIN lfsr_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.64 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.868 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 LAYER M2  ;
    ANTENNAMAXAREACAR 99.6944 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 369.847 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAMAXCUTCAR 1.38889 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 1 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.848 LAYER M3  ;
    ANTENNAGATEAREA 1.0896 LAYER M3  ;
    ANTENNAMAXAREACAR 100.612 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 373.379 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 34.4000 0.0000 34.6000 0.6000 ;
    END
  END lfsr_out[15]
  PIN lfsr_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.94 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.978 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 0.6 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.368 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0896 LAYER M3  ;
    ANTENNAMAXAREACAR 3.02594 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 12.4454 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.731155 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 32.9000 0.0000 33.1000 0.6000 ;
    END
  END lfsr_out[14]
  PIN lfsr_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.37 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 2.06 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.77 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0896 LAYER M3  ;
    ANTENNAMAXAREACAR 9.65223 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 36.9627 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.731155 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 31.4000 0.0000 31.6000 0.6000 ;
    END
  END lfsr_out[13]
  PIN lfsr_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.86 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.882 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 0.32 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.332 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0896 LAYER M3  ;
    ANTENNAMAXAREACAR 6.14635 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 23.9909 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.731155 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 29.9000 0.0000 30.1000 0.6000 ;
    END
  END lfsr_out[12]
  PIN lfsr_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.66 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.842 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 1.38 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.254 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0896 LAYER M3  ;
    ANTENNAMAXAREACAR 5.02668 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 19.984 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.731155 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 28.4000 0.0000 28.6000 0.6000 ;
    END
  END lfsr_out[11]
  PIN lfsr_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.46 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.802 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 0.68 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.664 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0896 LAYER M3  ;
    ANTENNAMAXAREACAR 3.31963 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 13.5321 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.731155 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 26.9000 0.0000 27.1000 0.6000 ;
    END
  END lfsr_out[10]
  PIN lfsr_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.74 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.138 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 0.62 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.442 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0896 LAYER M3  ;
    ANTENNAMAXAREACAR 4.14562 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 16.5882 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.731155 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 25.4000 0.0000 25.6000 0.6000 ;
    END
  END lfsr_out[9]
  PIN lfsr_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.94 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.178 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 1.44 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.476 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0896 LAYER M3  ;
    ANTENNAMAXAREACAR 4.2374 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 16.9278 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.731155 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 23.9000 0.0000 24.1000 0.6000 ;
    END
  END lfsr_out[8]
  PIN lfsr_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.88 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0896 LAYER M2  ;
    ANTENNAMAXAREACAR 3.98042 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 15.7053 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 22.4000 0.0000 22.6000 0.6000 ;
    END
  END lfsr_out[7]
  PIN lfsr_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.33 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 1.96 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.4 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0896 LAYER M3  ;
    ANTENNAMAXAREACAR 5.44885 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 21.4102 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.731155 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 20.9000 0.0000 21.1000 0.6000 ;
    END
  END lfsr_out[6]
  PIN lfsr_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.72 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.764 LAYER M2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0896 LAYER M2  ;
    ANTENNAMAXAREACAR 5.19187 LAYER M2  ;
    ANTENNAMAXSIDEAREACAR 20.1877 LAYER M2  ;
    ANTENNAMAXCUTCAR 0.694444 LAYER V2  ;
    PORT
      LAYER M2 ;
        RECT 19.4000 0.0000 19.6000 0.6000 ;
    END
  END lfsr_out[5]
  PIN lfsr_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.74 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.738 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 1.52 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.772 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0896 LAYER M3  ;
    ANTENNAMAXAREACAR 6.58688 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 25.6209 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.731155 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 17.9000 0.0000 18.1000 0.6000 ;
    END
  END lfsr_out[4]
  PIN lfsr_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.02 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.874 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 0.54 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.146 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0896 LAYER M3  ;
    ANTENNAMAXAREACAR 3.33798 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 13.6 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.731155 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 16.4000 0.0000 16.6000 0.6000 ;
    END
  END lfsr_out[3]
  PIN lfsr_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.69 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 0.84 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.256 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0896 LAYER M3  ;
    ANTENNAMAXAREACAR 4.49437 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 17.8786 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.731155 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 14.9000 0.0000 15.1000 0.6000 ;
    END
  END lfsr_out[2]
  PIN lfsr_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.06 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.722 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 1.14 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.366 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0896 LAYER M3  ;
    ANTENNAMAXAREACAR 4.32917 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 17.2674 LAYER M3  ;
    ANTENNAMAXCUTCAR 0.731155 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 13.4000 0.0000 13.6000 0.6000 ;
    END
  END lfsr_out[1]
  PIN lfsr_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.26 LAYER M2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.362 LAYER M2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER V2  ;
    ANTENNAPARTIALMETALAREA 6.84 LAYER M3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.604 LAYER M3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2288 LAYER M3  ;
    ANTENNAMAXAREACAR 19.9572 LAYER M3  ;
    ANTENNAMAXSIDEAREACAR 75.3883 LAYER M3  ;
    ANTENNAMAXCUTCAR 1.38889 LAYER VL  ;
    PORT
      LAYER M2 ;
        RECT 11.9000 0.0000 12.1000 0.6000 ;
    END
  END lfsr_out[0]
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 67.0000 52.0000 ;
    LAYER M2 ;
      RECT 0.0000 2.5200 67.0000 52.0000 ;
      RECT 54.5200 0.0000 67.0000 2.5200 ;
      RECT 0.0000 0.0000 9.9800 2.5200 ;
    LAYER M3 ;
      RECT 0.0000 17.0200 67.0000 52.0000 ;
      RECT 2.5200 8.9800 67.0000 17.0200 ;
      RECT 0.0000 0.0000 67.0000 8.9800 ;
    LAYER MQ ;
      RECT 0.0000 0.0000 67.0000 52.0000 ;
  END
END lfsr1

END LIBRARY
