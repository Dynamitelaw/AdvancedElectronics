
//`include "../rtl/CacheMem.v"

module cacheBank ( clk, reset, cacheDataIn_A, cacheAddressIn_A, memWrite_A, 
        cacheDataOut_A, portA_writtenTo, cacheDataIn_B, cacheAddressIn_B, 
        memWrite_B, cacheDataOut_B, portB_writtenTo );
  input [31:0] cacheDataIn_A;
  input [7:0] cacheAddressIn_A;
  output [31:0] cacheDataOut_A;
  input [31:0] cacheDataIn_B;
  input [7:0] cacheAddressIn_B;
  output [31:0] cacheDataOut_B;
  input clk, reset, memWrite_A, memWrite_B;
  output portA_writtenTo, portB_writtenTo;

CacheMem Memory( .QA(cacheDataOut_A), .QB(cacheDataOut_B), .CLKA(clk), .CENA(reset), .WENA(memWrite_A), .AA(cacheAddressIn_A), .DA(cacheDataIn_A), .CLKB(clk), .CENB(reset), .WENB(memWrite_B), .AB(cacheAddressIn_B), .DB(cacheDataIn_B));

endmodule



module incomingPortHandler_0 ( clk, reset, localRouterAddress, 
        destinationAddressIn, requesterAddressIn, readIn, writeIn, 
        outputPortSelect, memRead, memWrite );
  input [5:0] localRouterAddress;
  input [13:0] destinationAddressIn;
  input [5:0] requesterAddressIn;
  output [3:0] outputPortSelect;
  input clk, reset, readIn, writeIn;
  output memRead, memWrite;
  wire   n44, n42, n45, n43, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32;

  DFFQX1TS memWrite_reg ( .D(n30), .CK(clk), .Q(memWrite) );
  DFFQX1TS memRead_reg ( .D(n31), .CK(clk), .Q(memRead) );
  DFFHQX4TS \outputPortSelect_reg[3]  ( .D(n45), .CK(clk), .Q(
        outputPortSelect[3]) );
  DFFHQX1TS \outputPortSelect_reg[2]  ( .D(n44), .CK(clk), .Q(
        outputPortSelect[2]) );
  DFFHQX1TS \outputPortSelect_reg[1]  ( .D(n43), .CK(clk), .Q(
        outputPortSelect[1]) );
  DFFHQX1TS \outputPortSelect_reg[0]  ( .D(n42), .CK(clk), .Q(
        outputPortSelect[0]) );
  INVXLTS U1 ( .A(localRouterAddress[2]), .Y(n5) );
  INVXLTS U2 ( .A(localRouterAddress[1]), .Y(n6) );
  INVXLTS U3 ( .A(localRouterAddress[3]), .Y(n3) );
  INVXLTS U4 ( .A(destinationAddressIn[12]), .Y(n7) );
  OAI22XLTS U5 ( .A0(destinationAddressIn[10]), .A1(n5), .B0(n15), .B1(n4), 
        .Y(n13) );
  OAI21XLTS U6 ( .A0(localRouterAddress[4]), .A1(n7), .B0(n29), .Y(n20) );
  CLKBUFX2TS U7 ( .A(reset), .Y(n32) );
  NAND4BBX1TS U8 ( .AN(n17), .BN(n18), .C(n12), .D(n19), .Y(n14) );
  NOR2X1TS U9 ( .A(n20), .B(n21), .Y(n19) );
  OR2X2TS U10 ( .A(n32), .B(n10), .Y(n21) );
  NOR2BX1TS U11 ( .AN(n13), .B(n14), .Y(n45) );
  NOR2X1TS U12 ( .A(n14), .B(n13), .Y(n44) );
  NAND2BX1TS U13 ( .AN(n26), .B(n27), .Y(n18) );
  XOR2X1TS U14 ( .A(n8), .B(n3), .Y(n17) );
  INVX2TS U15 ( .A(n20), .Y(n2) );
  INVX2TS U16 ( .A(n12), .Y(n1) );
  AOI211X1TS U17 ( .A0(n2), .A1(n25), .B0(n21), .C0(n26), .Y(n43) );
  NAND3XLTS U18 ( .A(n27), .B(n3), .C(destinationAddressIn[11]), .Y(n25) );
  AOI22XLTS U19 ( .A0(n6), .A1(destinationAddressIn[9]), .B0(n5), .B1(
        destinationAddressIn[10]), .Y(n16) );
  NAND4X1TS U20 ( .A(n2), .B(n16), .C(n22), .D(n23), .Y(n12) );
  XNOR2XLTS U21 ( .A(destinationAddressIn[8]), .B(localRouterAddress[0]), .Y(
        n22) );
  NOR3X1TS U22 ( .A(n24), .B(n18), .C(n17), .Y(n23) );
  OAI22XLTS U23 ( .A0(destinationAddressIn[9]), .A1(n6), .B0(
        destinationAddressIn[10]), .B1(n5), .Y(n24) );
  NOR2XLTS U24 ( .A(readIn), .B(writeIn), .Y(n10) );
  NOR2BXLTS U25 ( .AN(localRouterAddress[5]), .B(destinationAddressIn[13]), 
        .Y(n26) );
  NAND2XLTS U26 ( .A(localRouterAddress[4]), .B(n7), .Y(n27) );
  NAND2BXLTS U27 ( .AN(localRouterAddress[5]), .B(destinationAddressIn[13]), 
        .Y(n29) );
  OA21XLTS U28 ( .A0(n6), .A1(destinationAddressIn[9]), .B0(
        destinationAddressIn[8]), .Y(n15) );
  INVX2TS U29 ( .A(n16), .Y(n4) );
  NOR2X1TS U30 ( .A(n28), .B(n21), .Y(n42) );
  AOI32XLTS U31 ( .A0(localRouterAddress[3]), .A1(n8), .A2(n2), .B0(n18), .B1(
        n29), .Y(n28) );
  NOR2X1TS U32 ( .A(n32), .B(n11), .Y(n31) );
  AOI22XLTS U33 ( .A0(memRead), .A1(n10), .B0(readIn), .B1(n1), .Y(n11) );
  NOR2X1TS U34 ( .A(n32), .B(n9), .Y(n30) );
  AOI22XLTS U35 ( .A0(memWrite), .A1(n10), .B0(writeIn), .B1(n1), .Y(n9) );
  INVXLTS U36 ( .A(destinationAddressIn[11]), .Y(n8) );
endmodule


module incomingPortHandler_3 ( clk, reset, localRouterAddress, 
        destinationAddressIn, requesterAddressIn, readIn, writeIn, 
        outputPortSelect, memRead, memWrite );
  input [5:0] localRouterAddress;
  input [13:0] destinationAddressIn;
  input [5:0] requesterAddressIn;
  output [3:0] outputPortSelect;
  input clk, reset, readIn, writeIn;
  output memRead, memWrite;
  wire   n44, n42, n43, n45, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32;

  DFFHQX1TS memWrite_reg ( .D(n30), .CK(clk), .Q(memWrite) );
  DFFHQX1TS memRead_reg ( .D(n31), .CK(clk), .Q(memRead) );
  DFFHQX4TS \outputPortSelect_reg[3]  ( .D(n45), .CK(clk), .Q(
        outputPortSelect[3]) );
  DFFHQX4TS \outputPortSelect_reg[1]  ( .D(n43), .CK(clk), .Q(
        outputPortSelect[1]) );
  DFFHQX1TS \outputPortSelect_reg[0]  ( .D(n42), .CK(clk), .Q(
        outputPortSelect[0]) );
  DFFHQX1TS \outputPortSelect_reg[2]  ( .D(n44), .CK(clk), .Q(
        outputPortSelect[2]) );
  INVXLTS U1 ( .A(localRouterAddress[2]), .Y(n5) );
  INVXLTS U2 ( .A(localRouterAddress[1]), .Y(n6) );
  INVXLTS U3 ( .A(localRouterAddress[3]), .Y(n3) );
  INVXLTS U4 ( .A(destinationAddressIn[12]), .Y(n7) );
  OAI22XLTS U5 ( .A0(destinationAddressIn[10]), .A1(n5), .B0(n15), .B1(n4), 
        .Y(n13) );
  OAI21XLTS U6 ( .A0(localRouterAddress[4]), .A1(n7), .B0(n29), .Y(n20) );
  CLKBUFX2TS U7 ( .A(reset), .Y(n32) );
  NAND4BBX1TS U8 ( .AN(n17), .BN(n18), .C(n12), .D(n19), .Y(n14) );
  NOR2X1TS U9 ( .A(n20), .B(n21), .Y(n19) );
  OR2X2TS U10 ( .A(n32), .B(n10), .Y(n21) );
  NOR2BX1TS U11 ( .AN(n13), .B(n14), .Y(n45) );
  NOR2X1TS U12 ( .A(n14), .B(n13), .Y(n44) );
  NAND2BX1TS U13 ( .AN(n26), .B(n27), .Y(n18) );
  XOR2X1TS U14 ( .A(n8), .B(n3), .Y(n17) );
  INVX2TS U15 ( .A(n20), .Y(n2) );
  INVX2TS U16 ( .A(n12), .Y(n1) );
  AOI211X1TS U17 ( .A0(n2), .A1(n25), .B0(n21), .C0(n26), .Y(n43) );
  NAND3XLTS U18 ( .A(n27), .B(n3), .C(destinationAddressIn[11]), .Y(n25) );
  AOI22XLTS U19 ( .A0(n6), .A1(destinationAddressIn[9]), .B0(n5), .B1(
        destinationAddressIn[10]), .Y(n16) );
  NAND4X1TS U20 ( .A(n2), .B(n16), .C(n22), .D(n23), .Y(n12) );
  XNOR2XLTS U21 ( .A(destinationAddressIn[8]), .B(localRouterAddress[0]), .Y(
        n22) );
  NOR3X1TS U22 ( .A(n24), .B(n18), .C(n17), .Y(n23) );
  OAI22XLTS U23 ( .A0(destinationAddressIn[9]), .A1(n6), .B0(
        destinationAddressIn[10]), .B1(n5), .Y(n24) );
  NOR2XLTS U24 ( .A(readIn), .B(writeIn), .Y(n10) );
  NOR2BXLTS U25 ( .AN(localRouterAddress[5]), .B(destinationAddressIn[13]), 
        .Y(n26) );
  NAND2XLTS U26 ( .A(localRouterAddress[4]), .B(n7), .Y(n27) );
  NAND2BXLTS U27 ( .AN(localRouterAddress[5]), .B(destinationAddressIn[13]), 
        .Y(n29) );
  OA21XLTS U28 ( .A0(n6), .A1(destinationAddressIn[9]), .B0(
        destinationAddressIn[8]), .Y(n15) );
  INVX2TS U29 ( .A(n16), .Y(n4) );
  NOR2X1TS U30 ( .A(n28), .B(n21), .Y(n42) );
  AOI32XLTS U31 ( .A0(localRouterAddress[3]), .A1(n8), .A2(n2), .B0(n18), .B1(
        n29), .Y(n28) );
  NOR2X1TS U32 ( .A(n32), .B(n11), .Y(n31) );
  AOI22XLTS U33 ( .A0(memRead), .A1(n10), .B0(readIn), .B1(n1), .Y(n11) );
  NOR2X1TS U34 ( .A(n32), .B(n9), .Y(n30) );
  AOI22XLTS U35 ( .A0(memWrite), .A1(n10), .B0(writeIn), .B1(n1), .Y(n9) );
  INVXLTS U36 ( .A(destinationAddressIn[11]), .Y(n8) );
endmodule


module incomingPortHandler_2 ( clk, reset, localRouterAddress, 
        destinationAddressIn, requesterAddressIn, readIn, writeIn, 
        outputPortSelect, memRead, memWrite );
  input [5:0] localRouterAddress;
  input [13:0] destinationAddressIn;
  input [5:0] requesterAddressIn;
  output [3:0] outputPortSelect;
  input clk, reset, readIn, writeIn;
  output memRead, memWrite;
  wire   n42, n43, n44, n45, n69, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32;
  assign memWrite = n69;

  DFFHQX1TS \outputPortSelect_reg[2]  ( .D(n44), .CK(clk), .Q(
        outputPortSelect[2]) );
  DFFHQX1TS \outputPortSelect_reg[3]  ( .D(n45), .CK(clk), .Q(
        outputPortSelect[3]) );
  DFFHQX1TS \outputPortSelect_reg[1]  ( .D(n43), .CK(clk), .Q(
        outputPortSelect[1]) );
  DFFQX1TS memRead_reg ( .D(n30), .CK(clk), .Q(memRead) );
  DFFQX4TS memWrite_reg ( .D(n31), .CK(clk), .Q(n69) );
  DFFHQX1TS \outputPortSelect_reg[0]  ( .D(n42), .CK(clk), .Q(
        outputPortSelect[0]) );
  INVXLTS U1 ( .A(localRouterAddress[2]), .Y(n5) );
  INVXLTS U2 ( .A(localRouterAddress[1]), .Y(n6) );
  INVXLTS U3 ( .A(localRouterAddress[3]), .Y(n3) );
  INVXLTS U4 ( .A(destinationAddressIn[12]), .Y(n7) );
  OAI22XLTS U5 ( .A0(destinationAddressIn[10]), .A1(n5), .B0(n15), .B1(n4), 
        .Y(n13) );
  OAI21XLTS U6 ( .A0(localRouterAddress[4]), .A1(n7), .B0(n29), .Y(n20) );
  CLKBUFX2TS U7 ( .A(reset), .Y(n32) );
  NAND4BBX1TS U8 ( .AN(n17), .BN(n18), .C(n12), .D(n19), .Y(n14) );
  NOR2X1TS U9 ( .A(n20), .B(n21), .Y(n19) );
  OR2X2TS U10 ( .A(n32), .B(n10), .Y(n21) );
  NOR2BX1TS U11 ( .AN(n13), .B(n14), .Y(n45) );
  NOR2X1TS U12 ( .A(n14), .B(n13), .Y(n44) );
  NAND2BX1TS U13 ( .AN(n26), .B(n27), .Y(n18) );
  XOR2X1TS U14 ( .A(n8), .B(n3), .Y(n17) );
  INVX2TS U15 ( .A(n20), .Y(n2) );
  INVX2TS U16 ( .A(n12), .Y(n1) );
  AOI211X1TS U17 ( .A0(n2), .A1(n25), .B0(n21), .C0(n26), .Y(n43) );
  NAND3XLTS U18 ( .A(n27), .B(n3), .C(destinationAddressIn[11]), .Y(n25) );
  AOI22XLTS U19 ( .A0(n6), .A1(destinationAddressIn[9]), .B0(n5), .B1(
        destinationAddressIn[10]), .Y(n16) );
  NAND4X1TS U20 ( .A(n2), .B(n16), .C(n22), .D(n23), .Y(n12) );
  XNOR2XLTS U21 ( .A(destinationAddressIn[8]), .B(localRouterAddress[0]), .Y(
        n22) );
  NOR3X1TS U22 ( .A(n24), .B(n18), .C(n17), .Y(n23) );
  OAI22XLTS U23 ( .A0(destinationAddressIn[9]), .A1(n6), .B0(
        destinationAddressIn[10]), .B1(n5), .Y(n24) );
  NOR2XLTS U24 ( .A(readIn), .B(writeIn), .Y(n10) );
  NOR2BXLTS U25 ( .AN(localRouterAddress[5]), .B(destinationAddressIn[13]), 
        .Y(n26) );
  NAND2XLTS U26 ( .A(localRouterAddress[4]), .B(n7), .Y(n27) );
  NAND2BXLTS U27 ( .AN(localRouterAddress[5]), .B(destinationAddressIn[13]), 
        .Y(n29) );
  OA21XLTS U28 ( .A0(n6), .A1(destinationAddressIn[9]), .B0(
        destinationAddressIn[8]), .Y(n15) );
  INVX2TS U29 ( .A(n16), .Y(n4) );
  NOR2X1TS U30 ( .A(n28), .B(n21), .Y(n42) );
  AOI32XLTS U31 ( .A0(localRouterAddress[3]), .A1(n8), .A2(n2), .B0(n18), .B1(
        n29), .Y(n28) );
  NOR2X1TS U32 ( .A(n32), .B(n11), .Y(n31) );
  AOI22XLTS U33 ( .A0(n69), .A1(n10), .B0(writeIn), .B1(n1), .Y(n11) );
  NOR2X1TS U34 ( .A(n32), .B(n9), .Y(n30) );
  AOI22XLTS U35 ( .A0(memRead), .A1(n10), .B0(readIn), .B1(n1), .Y(n9) );
  INVXLTS U36 ( .A(destinationAddressIn[11]), .Y(n8) );
endmodule


module incomingPortHandler_1 ( clk, reset, localRouterAddress, 
        destinationAddressIn, requesterAddressIn, readIn, writeIn, 
        outputPortSelect, memRead, memWrite );
  input [5:0] localRouterAddress;
  input [13:0] destinationAddressIn;
  input [5:0] requesterAddressIn;
  output [3:0] outputPortSelect;
  input clk, reset, readIn, writeIn;
  output memRead, memWrite;
  wire   n70, n43, n45, n44, n42, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32;

  DFFQX1TS memWrite_reg ( .D(n31), .CK(clk), .Q(n70) );
  DFFQX1TS memRead_reg ( .D(n30), .CK(clk), .Q(memRead) );
  DFFQX1TS \outputPortSelect_reg[0]  ( .D(n42), .CK(clk), .Q(
        outputPortSelect[0]) );
  DFFQX1TS \outputPortSelect_reg[3]  ( .D(n45), .CK(clk), .Q(
        outputPortSelect[3]) );
  DFFQX1TS \outputPortSelect_reg[2]  ( .D(n44), .CK(clk), .Q(
        outputPortSelect[2]) );
  DFFQX1TS \outputPortSelect_reg[1]  ( .D(n43), .CK(clk), .Q(
        outputPortSelect[1]) );
  INVXLTS U1 ( .A(n70), .Y(n32) );
  INVXLTS U2 ( .A(n32), .Y(memWrite) );
  INVXLTS U3 ( .A(localRouterAddress[2]), .Y(n5) );
  INVXLTS U4 ( .A(localRouterAddress[1]), .Y(n6) );
  INVXLTS U5 ( .A(localRouterAddress[3]), .Y(n3) );
  INVXLTS U6 ( .A(destinationAddressIn[12]), .Y(n7) );
  OAI22XLTS U7 ( .A0(destinationAddressIn[10]), .A1(n5), .B0(n15), .B1(n4), 
        .Y(n13) );
  OAI21XLTS U8 ( .A0(localRouterAddress[4]), .A1(n7), .B0(n29), .Y(n20) );
  NAND4BBX1TS U9 ( .AN(n17), .BN(n18), .C(n12), .D(n19), .Y(n14) );
  NOR2X1TS U10 ( .A(n20), .B(n21), .Y(n19) );
  OR2X2TS U11 ( .A(reset), .B(n10), .Y(n21) );
  NOR2BX1TS U12 ( .AN(n13), .B(n14), .Y(n45) );
  NOR2X1TS U13 ( .A(n14), .B(n13), .Y(n44) );
  NAND2BX1TS U14 ( .AN(n26), .B(n27), .Y(n18) );
  XOR2X1TS U15 ( .A(n8), .B(n3), .Y(n17) );
  INVX2TS U16 ( .A(n20), .Y(n2) );
  INVX2TS U17 ( .A(n12), .Y(n1) );
  AOI211X1TS U18 ( .A0(n2), .A1(n25), .B0(n21), .C0(n26), .Y(n43) );
  NAND3XLTS U19 ( .A(n27), .B(n3), .C(destinationAddressIn[11]), .Y(n25) );
  AOI22XLTS U20 ( .A0(n6), .A1(destinationAddressIn[9]), .B0(n5), .B1(
        destinationAddressIn[10]), .Y(n16) );
  NAND4X1TS U21 ( .A(n2), .B(n16), .C(n22), .D(n23), .Y(n12) );
  XNOR2XLTS U22 ( .A(destinationAddressIn[8]), .B(localRouterAddress[0]), .Y(
        n22) );
  NOR3X1TS U23 ( .A(n24), .B(n18), .C(n17), .Y(n23) );
  OAI22XLTS U24 ( .A0(destinationAddressIn[9]), .A1(n6), .B0(
        destinationAddressIn[10]), .B1(n5), .Y(n24) );
  NOR2XLTS U25 ( .A(readIn), .B(writeIn), .Y(n10) );
  NOR2BXLTS U26 ( .AN(localRouterAddress[5]), .B(destinationAddressIn[13]), 
        .Y(n26) );
  NAND2XLTS U27 ( .A(localRouterAddress[4]), .B(n7), .Y(n27) );
  NAND2BXLTS U28 ( .AN(localRouterAddress[5]), .B(destinationAddressIn[13]), 
        .Y(n29) );
  OA21XLTS U29 ( .A0(n6), .A1(destinationAddressIn[9]), .B0(
        destinationAddressIn[8]), .Y(n15) );
  INVX2TS U30 ( .A(n16), .Y(n4) );
  NOR2X1TS U31 ( .A(n28), .B(n21), .Y(n42) );
  AOI32XLTS U32 ( .A0(localRouterAddress[3]), .A1(n8), .A2(n2), .B0(n18), .B1(
        n29), .Y(n28) );
  NOR2X1TS U33 ( .A(reset), .B(n11), .Y(n31) );
  AOI22XLTS U34 ( .A0(n70), .A1(n10), .B0(writeIn), .B1(n1), .Y(n11) );
  NOR2X1TS U35 ( .A(reset), .B(n9), .Y(n30) );
  AOI22XLTS U36 ( .A0(memRead), .A1(n10), .B0(readIn), .B1(n1), .Y(n9) );
  INVXLTS U37 ( .A(destinationAddressIn[11]), .Y(n8) );
endmodule


module cacheAccessArbiter ( clk, reset, cacheAddressIn_NORTH, 
        requesterAddressIn_NORTH, memRead_NORTH, memWrite_NORTH, dataIn_NORTH, 
        readReady_NORTH, requesterAddressOut_NORTH, cacheDataOut_NORTH, 
        cacheAddressIn_SOUTH, requesterAddressIn_SOUTH, memRead_SOUTH, 
        memWrite_SOUTH, dataIn_SOUTH, readReady_SOUTH, 
        requesterAddressOut_SOUTH, cacheDataOut_SOUTH, cacheAddressIn_EAST, 
        requesterAddressIn_EAST, memRead_EAST, memWrite_EAST, dataIn_EAST, 
        readReady_EAST, requesterAddressOut_EAST, cacheDataOut_EAST, 
        cacheAddressIn_WEST, requesterAddressIn_WEST, memRead_WEST, 
        memWrite_WEST, dataIn_WEST, readReady_WEST, requesterAddressOut_WEST, 
        cacheDataOut_WEST, cacheDataIn_A, cacheAddressIn_A, cacheDataOut_A, 
        memWrite_A, cacheDataIn_B, cacheAddressIn_B, cacheDataOut_B, 
        memWrite_B );
  input [7:0] cacheAddressIn_NORTH;
  input [5:0] requesterAddressIn_NORTH;
  input [31:0] dataIn_NORTH;
  output [5:0] requesterAddressOut_NORTH;
  output [31:0] cacheDataOut_NORTH;
  input [7:0] cacheAddressIn_SOUTH;
  input [5:0] requesterAddressIn_SOUTH;
  input [31:0] dataIn_SOUTH;
  output [5:0] requesterAddressOut_SOUTH;
  output [31:0] cacheDataOut_SOUTH;
  input [7:0] cacheAddressIn_EAST;
  input [5:0] requesterAddressIn_EAST;
  input [31:0] dataIn_EAST;
  output [5:0] requesterAddressOut_EAST;
  output [31:0] cacheDataOut_EAST;
  input [7:0] cacheAddressIn_WEST;
  input [5:0] requesterAddressIn_WEST;
  input [31:0] dataIn_WEST;
  output [5:0] requesterAddressOut_WEST;
  output [31:0] cacheDataOut_WEST;
  output [31:0] cacheDataIn_A;
  output [7:0] cacheAddressIn_A;
  input [31:0] cacheDataOut_A;
  output [31:0] cacheDataIn_B;
  output [7:0] cacheAddressIn_B;
  input [31:0] cacheDataOut_B;
  input clk, reset, memRead_NORTH, memWrite_NORTH, memRead_SOUTH,
         memWrite_SOUTH, memRead_EAST, memWrite_EAST, memRead_WEST,
         memWrite_WEST;
  output readReady_NORTH, readReady_SOUTH, readReady_EAST, readReady_WEST,
         memWrite_A, memWrite_B;
  wire   \requesterPortBuffer[4][0] , \requesterPortBuffer[6][0] ,
         \requesterPortBuffer[2][0] , n3253, n3252, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, \requesterPortBuffer[0][0] , n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3345, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3208, n3207, n3206, n3205, n3204, n3203, n3268,
         \requesterPortBuffer[0][1] , n3343, n45, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3310, n79, n3311, n78, n3312, n77, n3313,
         n76, n3314, n75, n3315, n74, n3316, n73, n3317, n72, n3286, n3302,
         n62, n3287, n3303, n60, n3288, n3304, n58, n3289, n3305, n56, n3290,
         n3306, n54, n3291, n3307, n52, n3292, n3308, n50, n3293, n3309, n48,
         n3514, n1922, n3515, n1921, n3516, n1920, n3517, n1919, n3518, n1918,
         n3519, n1917, n3520, n1916, n3521, n1915, n3522, n1914, n3523, n1913,
         n3524, n1912, n3525, n1911, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3266, n47, n3267, n46, n3643, n910,
         n3642, n880, n3344, n3197, n3198, n3199, n3200, n3201, n3202, n3185,
         n3186, n3187, n3188, n3189, n3190, n3265, \prevRequesterPort_B[0] ,
         n3264, n3277, n1974, n3276, n1973, n3275, n1972, n3274, n1971, n3273,
         n1970, n3272, n1969, n3271, n1968, n3270, n1967, n3249, n2006, n3248,
         n2005, n3247, n2004, n3246, n2003, n3245, n2002, n3244, n2001, n3243,
         n2000, n3242, n1999, n3241, n1998, n3240, n1997, n3239, n1996, n3238,
         n1995, n3237, n1994, n3236, n1993, n3235, n1992, n3234, n1991, n3233,
         n1990, n3232, n1989, n3231, n1988, n3230, n1987, n3229, n1986, n3228,
         n1985, n3227, n1984, n3226, n1983, n3225, n1982, n3224, n1981, n3223,
         n1980, n3222, n1979, n3221, n1978, n3220, n1977, n3219, n1976, n3218,
         n1975, n3184, n2095, n3217, n2097, n3377, n2092, n3376, n2090, n3375,
         n2088, n3374, n2086, n3373, n2084, n3372, n2082, n3371, n2080, n3370,
         n2078, n3369, n2076, n3368, n2074, n3367, n2072, n3366, n2070, n3365,
         n2068, n3364, n2066, n3363, n2064, n3362, n2062, n3361, n2060, n3360,
         n2058, n3359, n2056, n3358, n2054, n3357, n2052, n3356, n2050, n3355,
         n2048, n3354, n2046, n3353, n2044, n3352, n2042, n3351, n2040, n3350,
         n2038, n3349, n2036, n3348, n2034, n3347, n2032, n3346, n2030, n3216,
         n2028, n3215, n2026, n3214, n2024, n3213, n2022, n3212, n2020, n3211,
         n2018, n3210, n2016, n3209, n2014, N10040, N10030, N10020, N10010,
         n3165, n3164, n3163, n3162, n3161, n3160, n3177, n3176, n3175, n3174,
         n3173, n3172, n3171, n3170, n3169, n3168, n3167, n3166, n3183, n3182,
         n3181, n3180, n3179, n3178, N10216, N10215, N10214, N10213, N10212,
         N10211, N10210, N10209, N10208, N10207, N10206, N10205, N10204,
         N10203, N10202, N10201, N10200, N10199, N10198, N10197, N10196,
         N10195, N10194, N10193, N10192, N10191, N10190, N10189, N10188,
         N10187, N10186, N10185, N10182, N10181, N10180, N10179, N10178,
         N10177, N10176, N10175, N10174, N10173, N10172, N10171, N10170,
         N10169, N10168, N10167, N10166, N10165, N10164, N10163, N10162,
         N10161, N10160, N10159, N10158, N10157, N10156, N10155, N10154,
         N10153, N10152, N10151, N10148, N10147, N10146, N10145, N10144,
         N10143, N10142, N10141, N10140, N10139, N10138, N10137, N10136,
         N10135, N10134, N10133, N10132, N10131, N10130, N10129, N10128,
         N10127, N10126, N10125, N10124, N10123, N10122, N10121, N10120,
         N10119, N10118, N10117, N10114, N10113, N10112, N10111, N10110,
         N10109, N10108, N10107, N10106, N10105, N10104, N10103, N10102,
         N10101, N10100, N10099, N10098, N10097, N10096, N10095, N10094,
         N10093, N10092, N10091, N10090, N10089, N10088, N10087, N10086,
         N10085, N10084, N10083, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         \requesterAddressBuffer[0][5] , \requesterAddressBuffer[0][4] ,
         \requesterAddressBuffer[0][2] , \requesterAddressBuffer[0][3] ,
         \requesterAddressBuffer[0][1] , \requesterAddressBuffer[0][0] , n3610,
         n783, n3617, n790, n3620, n793, n3625, n720, n3629, n724, n3633, n728,
         n3637, n732, n3641, n736, n3611, n784, n3612, n785, n3613, n786,
         n3614, n787, n3615, n788, n3616, n789, n3618, n791, n3619, n792,
         n3621, n716, n3622, n717, n3623, n718, n3624, n719, n3626, n721,
         n3627, n722, n3628, n723, n3630, n725, n3631, n726, n3632, n727,
         n3634, n729, n3635, n730, n3636, n731, n3638, n733, n3639, n734,
         n3640, n735, n3378, n3379, n3381, n3383, n3385, n3341, n782, n3251,
         n3250, n740, n3335, n776, n3337, n778, n3339, n780, n3340, n781,
         n3334, n775, n3336, n777, n3338, n779, n3384, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3644, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n737,
         n738, n739, n742, n743, n748, n754, n755, n756, n757, n758, n759,
         n770, n771, n773, n774, n794, n795, n796, n797, n798, n800, n801,
         n802, n803, n805, n808, n809, n810, n811, n812, n813, n814, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n957, n958, n960, n961, n962, n963, n964, n965, n966, n975,
         n976, n977, n1024, n1025, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n2007,
         n2008, n2009, n2010, n2011, n2012, n2013, n2015, n2017, n2019, n2021,
         n2023, n2025, n2027, n2029, n2031, n2033, n2035, n2037, n2039, n2041,
         n2043, n2045, n2047, n2049, n2051, n2053, n2055, n2057, n2059, n2061,
         n2063, n2065, n2067, n2069, n2071, n2073, n2075, n2077, n2079, n2081,
         n2083, n2089, n2091, n2093, n2094, n2096, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n49, n51, n53, n55, n57, n59, n61,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n683, n684, n685, n686, n687, n688, n689, n690,
         n741, n744, n745, n746, n747, n749, n750, n751, n752, n753, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n772, n799,
         n804, n806, n807, n815, n816, n831, n935, n955, n956, n959, n967,
         n968, n969, n970, n971, n972, n973, n974, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1136, n1137, n1263, n1377, n1489, n1500, n1599, n1607,
         n1681, n1739, n1752, n1767, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1965, n1966, n2085, n2087, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506;
  wire   [5:0] prevRequesterAddress_B;
  wire   [5:0] prevRequesterAddress_A;

  DFFNSRX2TS \cacheAddressIn_A_reg[7]  ( .D(n3277), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_A[7]), .QN(n1974) );
  DFFNSRX2TS \cacheAddressIn_A_reg[6]  ( .D(n3276), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_A[6]), .QN(n1973) );
  DFFNSRX2TS \cacheAddressIn_A_reg[5]  ( .D(n3275), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_A[5]), .QN(n1972) );
  DFFNSRX2TS \cacheAddressIn_A_reg[4]  ( .D(n3274), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_A[4]), .QN(n1971) );
  DFFNSRX2TS \cacheAddressIn_A_reg[3]  ( .D(n3273), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_A[3]), .QN(n1970) );
  DFFNSRX2TS \cacheAddressIn_A_reg[2]  ( .D(n3272), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_A[2]), .QN(n1969) );
  DFFNSRX2TS \cacheAddressIn_A_reg[1]  ( .D(n3271), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_A[1]), .QN(n1968) );
  DFFNSRX2TS \cacheAddressIn_A_reg[0]  ( .D(n3270), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_A[0]), .QN(n1967) );
  DFFNSRX2TS \cacheDataIn_A_reg[31]  ( .D(n3249), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[31]), .QN(n2006) );
  DFFNSRX2TS \cacheDataIn_A_reg[30]  ( .D(n3248), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[30]), .QN(n2005) );
  DFFNSRX2TS \cacheDataIn_A_reg[29]  ( .D(n3247), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[29]), .QN(n2004) );
  DFFNSRX2TS \cacheDataIn_A_reg[28]  ( .D(n3246), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[28]), .QN(n2003) );
  DFFNSRX2TS \cacheDataIn_A_reg[27]  ( .D(n3245), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[27]), .QN(n2002) );
  DFFNSRX2TS \cacheDataIn_A_reg[26]  ( .D(n3244), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[26]), .QN(n2001) );
  DFFNSRX2TS \cacheDataIn_A_reg[25]  ( .D(n3243), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[25]), .QN(n2000) );
  DFFNSRX2TS \cacheDataIn_A_reg[24]  ( .D(n3242), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[24]), .QN(n1999) );
  DFFNSRX2TS \cacheDataIn_A_reg[23]  ( .D(n3241), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[23]), .QN(n1998) );
  DFFNSRX2TS \cacheDataIn_A_reg[22]  ( .D(n3240), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[22]), .QN(n1997) );
  DFFNSRX2TS \cacheDataIn_A_reg[21]  ( .D(n3239), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[21]), .QN(n1996) );
  DFFNSRX2TS \cacheDataIn_A_reg[20]  ( .D(n3238), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[20]), .QN(n1995) );
  DFFNSRX2TS \cacheDataIn_A_reg[19]  ( .D(n3237), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[19]), .QN(n1994) );
  DFFNSRX2TS \cacheDataIn_A_reg[18]  ( .D(n3236), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[18]), .QN(n1993) );
  DFFNSRX2TS \cacheDataIn_A_reg[17]  ( .D(n3235), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[17]), .QN(n1992) );
  DFFNSRX2TS \cacheDataIn_A_reg[16]  ( .D(n3234), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[16]), .QN(n1991) );
  DFFNSRX2TS \cacheDataIn_A_reg[15]  ( .D(n3233), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[15]), .QN(n1990) );
  DFFNSRX2TS \cacheDataIn_A_reg[14]  ( .D(n3232), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[14]), .QN(n1989) );
  DFFNSRX2TS \cacheDataIn_A_reg[13]  ( .D(n3231), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[13]), .QN(n1988) );
  DFFNSRX2TS \cacheDataIn_A_reg[12]  ( .D(n3230), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[12]), .QN(n1987) );
  DFFNSRX2TS \cacheDataIn_A_reg[11]  ( .D(n3229), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[11]), .QN(n1986) );
  DFFNSRX2TS \cacheDataIn_A_reg[10]  ( .D(n3228), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[10]), .QN(n1985) );
  DFFNSRX2TS \cacheDataIn_A_reg[9]  ( .D(n3227), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[9]), .QN(n1984) );
  DFFNSRX2TS \cacheDataIn_A_reg[8]  ( .D(n3226), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[8]), .QN(n1983) );
  DFFNSRX2TS \cacheDataIn_A_reg[7]  ( .D(n3225), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[7]), .QN(n1982) );
  DFFNSRX2TS \cacheDataIn_A_reg[6]  ( .D(n3224), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[6]), .QN(n1981) );
  DFFNSRX2TS \cacheDataIn_A_reg[5]  ( .D(n3223), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[5]), .QN(n1980) );
  DFFNSRX2TS \cacheDataIn_A_reg[4]  ( .D(n3222), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[4]), .QN(n1979) );
  DFFNSRX2TS \cacheDataIn_A_reg[3]  ( .D(n3221), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[3]), .QN(n1978) );
  DFFNSRX2TS \cacheDataIn_A_reg[2]  ( .D(n3220), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[2]), .QN(n1977) );
  DFFNSRX2TS \cacheDataIn_A_reg[1]  ( .D(n3219), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[1]), .QN(n1976) );
  DFFNSRX2TS \cacheDataIn_A_reg[0]  ( .D(n3218), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_A[0]), .QN(n1975) );
  DFFNSRX2TS \cacheDataIn_B_reg[31]  ( .D(n3377), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[31]), .QN(n2092) );
  DFFNSRX2TS \cacheDataIn_B_reg[30]  ( .D(n3376), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[30]), .QN(n2090) );
  DFFNSRX2TS \cacheDataIn_B_reg[29]  ( .D(n3375), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[29]), .QN(n2088) );
  DFFNSRX2TS \cacheDataIn_B_reg[28]  ( .D(n3374), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[28]), .QN(n2086) );
  DFFNSRX2TS \cacheDataIn_B_reg[27]  ( .D(n3373), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[27]), .QN(n2084) );
  DFFNSRX2TS \cacheDataIn_B_reg[26]  ( .D(n3372), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[26]), .QN(n2082) );
  DFFNSRX2TS \cacheDataIn_B_reg[25]  ( .D(n3371), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[25]), .QN(n2080) );
  DFFNSRX2TS \cacheDataIn_B_reg[24]  ( .D(n3370), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[24]), .QN(n2078) );
  DFFNSRX2TS \cacheDataIn_B_reg[23]  ( .D(n3369), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[23]), .QN(n2076) );
  DFFNSRX2TS \cacheDataIn_B_reg[22]  ( .D(n3368), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[22]), .QN(n2074) );
  DFFNSRX2TS \cacheDataIn_B_reg[21]  ( .D(n3367), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[21]), .QN(n2072) );
  DFFNSRX2TS \cacheDataIn_B_reg[20]  ( .D(n3366), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[20]), .QN(n2070) );
  DFFNSRX2TS \cacheDataIn_B_reg[19]  ( .D(n3365), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[19]), .QN(n2068) );
  DFFNSRX2TS \cacheDataIn_B_reg[18]  ( .D(n3364), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[18]), .QN(n2066) );
  DFFNSRX2TS \cacheDataIn_B_reg[17]  ( .D(n3363), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[17]), .QN(n2064) );
  DFFNSRX2TS \cacheDataIn_B_reg[16]  ( .D(n3362), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[16]), .QN(n2062) );
  DFFNSRX2TS \cacheDataIn_B_reg[15]  ( .D(n3361), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[15]), .QN(n2060) );
  DFFNSRX2TS \cacheDataIn_B_reg[14]  ( .D(n3360), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[14]), .QN(n2058) );
  DFFNSRX2TS \cacheDataIn_B_reg[13]  ( .D(n3359), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[13]), .QN(n2056) );
  DFFNSRX2TS \cacheDataIn_B_reg[12]  ( .D(n3358), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[12]), .QN(n2054) );
  DFFNSRX2TS \cacheDataIn_B_reg[11]  ( .D(n3357), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[11]), .QN(n2052) );
  DFFNSRX2TS \cacheDataIn_B_reg[10]  ( .D(n3356), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[10]), .QN(n2050) );
  DFFNSRX2TS \cacheDataIn_B_reg[9]  ( .D(n3355), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[9]), .QN(n2048) );
  DFFNSRX2TS \cacheDataIn_B_reg[8]  ( .D(n3354), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[8]), .QN(n2046) );
  DFFNSRX2TS \cacheDataIn_B_reg[7]  ( .D(n3353), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[7]), .QN(n2044) );
  DFFNSRX2TS \cacheDataIn_B_reg[6]  ( .D(n3352), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[6]), .QN(n2042) );
  DFFNSRX2TS \cacheDataIn_B_reg[5]  ( .D(n3351), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[5]), .QN(n2040) );
  DFFNSRX2TS \cacheDataIn_B_reg[4]  ( .D(n3350), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[4]), .QN(n2038) );
  DFFNSRX2TS \cacheDataIn_B_reg[3]  ( .D(n3349), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[3]), .QN(n2036) );
  DFFNSRX2TS \cacheDataIn_B_reg[2]  ( .D(n3348), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[2]), .QN(n2034) );
  DFFNSRX2TS \cacheDataIn_B_reg[1]  ( .D(n3347), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[1]), .QN(n2032) );
  DFFNSRX2TS \cacheDataIn_B_reg[0]  ( .D(n3346), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheDataIn_B[0]), .QN(n2030) );
  DFFNSRX2TS \cacheAddressIn_B_reg[7]  ( .D(n3216), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_B[7]), .QN(n2028) );
  DFFNSRX2TS \cacheAddressIn_B_reg[6]  ( .D(n3215), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_B[6]), .QN(n2026) );
  DFFNSRX2TS \cacheAddressIn_B_reg[5]  ( .D(n3214), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_B[5]), .QN(n2024) );
  DFFNSRX2TS \cacheAddressIn_B_reg[4]  ( .D(n3213), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_B[4]), .QN(n2022) );
  DFFNSRX2TS \cacheAddressIn_B_reg[3]  ( .D(n3212), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_B[3]), .QN(n2020) );
  DFFNSRX2TS \cacheAddressIn_B_reg[2]  ( .D(n3211), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_B[2]), .QN(n2018) );
  DFFNSRX2TS \cacheAddressIn_B_reg[1]  ( .D(n3210), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_B[1]), .QN(n2016) );
  DFFNSRX2TS \cacheAddressIn_B_reg[0]  ( .D(n3209), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(cacheAddressIn_B[0]), .QN(n2014) );
  DFFNSRX2TS memWrite_A_reg ( .D(n3184), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        memWrite_A), .QN(n2095) );
  DFFNSRX2TS memWrite_B_reg ( .D(n3217), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        memWrite_B), .QN(n2097) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][31]  ( .D(n3450), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1880) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][30]  ( .D(n3451), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1879) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][29]  ( .D(n3452), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1878) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][28]  ( .D(n3453), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1877) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][27]  ( .D(n3454), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1876) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][26]  ( .D(n3455), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1875) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][25]  ( .D(n3456), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1874) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][24]  ( .D(n3457), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1873) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][23]  ( .D(n3458), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1872) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][22]  ( .D(n3459), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1871) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][21]  ( .D(n3460), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1870) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][20]  ( .D(n3461), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1869) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][19]  ( .D(n3462), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1868) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][18]  ( .D(n3463), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1867) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][17]  ( .D(n3464), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1866) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][16]  ( .D(n3465), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1865) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][15]  ( .D(n3466), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1864) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][14]  ( .D(n3467), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1863) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][13]  ( .D(n3468), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1862) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][12]  ( .D(n3469), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1861) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][11]  ( .D(n3470), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1860) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][10]  ( .D(n3471), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1859) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][9]  ( .D(n3472), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1858) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][8]  ( .D(n3473), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1857) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][7]  ( .D(n3474), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1856) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][6]  ( .D(n3475), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1855) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][5]  ( .D(n3476), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1854) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][4]  ( .D(n3477), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1853) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][3]  ( .D(n3478), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1852) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][2]  ( .D(n3479), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1851) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][1]  ( .D(n3480), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1850) );
  DFFNSRX2TS \dataToWriteBuffer_reg[5][0]  ( .D(n3481), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1849) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][31]  ( .D(n3418), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1848) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][30]  ( .D(n3419), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1847) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][29]  ( .D(n3420), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1846) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][28]  ( .D(n3421), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1845) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][27]  ( .D(n3422), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1843) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][26]  ( .D(n3423), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1842) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][25]  ( .D(n3424), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1841) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][24]  ( .D(n3425), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1840) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][23]  ( .D(n3426), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1838) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][22]  ( .D(n3427), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1837) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][21]  ( .D(n3428), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1836) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][20]  ( .D(n3429), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1835) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][19]  ( .D(n3430), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1833) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][18]  ( .D(n3431), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1832) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][17]  ( .D(n3432), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1831) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][16]  ( .D(n3433), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1830) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][3]  ( .D(n3446), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1813) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][2]  ( .D(n3447), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1812) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][1]  ( .D(n3448), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1811) );
  DFFNSRX2TS \dataToWriteBuffer_reg[6][0]  ( .D(n3449), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1810) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][31]  ( .D(n3482), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1808) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][30]  ( .D(n3483), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1807) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][29]  ( .D(n3484), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1806) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][28]  ( .D(n3485), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1844) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][27]  ( .D(n3486), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1805) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][26]  ( .D(n3487), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1804) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][25]  ( .D(n3488), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1803) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][24]  ( .D(n3489), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1839) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][23]  ( .D(n3490), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1802) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][22]  ( .D(n3491), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1801) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][21]  ( .D(n3492), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1800) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][20]  ( .D(n3493), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1834) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][19]  ( .D(n3494), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1799) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][18]  ( .D(n3495), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1798) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][17]  ( .D(n3496), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1797) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][16]  ( .D(n3497), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1829) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][15]  ( .D(n3498), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1796) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][14]  ( .D(n3499), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1795) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][13]  ( .D(n3500), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1794) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][12]  ( .D(n3501), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1824) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][11]  ( .D(n3502), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1793) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][10]  ( .D(n3503), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1792) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][9]  ( .D(n3504), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1791) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][8]  ( .D(n3505), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1819) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][7]  ( .D(n3506), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1790) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][6]  ( .D(n3507), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1789) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][5]  ( .D(n3508), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1788) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][4]  ( .D(n3509), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1814) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][3]  ( .D(n3510), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1787) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][2]  ( .D(n3511), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1786) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][1]  ( .D(n3512), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1785) );
  DFFNSRX2TS \dataToWriteBuffer_reg[4][0]  ( .D(n3513), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1809) );
  DFFNSRX2TS \addressToWriteBuffer_reg[4][7]  ( .D(n3302), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n62) );
  DFFNSRX2TS \addressToWriteBuffer_reg[4][6]  ( .D(n3303), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n60) );
  DFFNSRX2TS \addressToWriteBuffer_reg[4][5]  ( .D(n3304), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n58) );
  DFFNSRX2TS \addressToWriteBuffer_reg[4][4]  ( .D(n3305), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n56) );
  DFFNSRX2TS \addressToWriteBuffer_reg[4][3]  ( .D(n3306), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n54) );
  DFFNSRX2TS \addressToWriteBuffer_reg[4][2]  ( .D(n3307), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n52) );
  DFFNSRX2TS \addressToWriteBuffer_reg[4][1]  ( .D(n3308), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n50) );
  DFFNSRX2TS \addressToWriteBuffer_reg[4][0]  ( .D(n3309), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n48) );
  DFFNSRX2TS \addressToWriteBuffer_reg[5][7]  ( .D(n3294), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n675) );
  DFFNSRX2TS \addressToWriteBuffer_reg[5][6]  ( .D(n3295), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n676) );
  DFFNSRX2TS \addressToWriteBuffer_reg[5][5]  ( .D(n3296), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n677) );
  DFFNSRX2TS \addressToWriteBuffer_reg[5][4]  ( .D(n3297), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n678) );
  DFFNSRX2TS \addressToWriteBuffer_reg[5][3]  ( .D(n3298), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n679) );
  DFFNSRX2TS \addressToWriteBuffer_reg[5][2]  ( .D(n3299), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n680) );
  DFFNSRX2TS \addressToWriteBuffer_reg[5][1]  ( .D(n3300), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n681) );
  DFFNSRX2TS \addressToWriteBuffer_reg[5][0]  ( .D(n3301), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n682) );
  DFFNSRX2TS \addressToWriteBuffer_reg[6][7]  ( .D(n3286), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n691) );
  DFFNSRX2TS \addressToWriteBuffer_reg[6][6]  ( .D(n3287), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n692) );
  DFFNSRX2TS \addressToWriteBuffer_reg[6][5]  ( .D(n3288), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n693) );
  DFFNSRX2TS \addressToWriteBuffer_reg[6][4]  ( .D(n3289), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n694) );
  DFFNSRX2TS \addressToWriteBuffer_reg[6][3]  ( .D(n3290), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n695) );
  DFFNSRX2TS \addressToWriteBuffer_reg[6][2]  ( .D(n3291), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n696) );
  DFFNSRX2TS \addressToWriteBuffer_reg[6][1]  ( .D(n3292), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n697) );
  DFFNSRX2TS \addressToWriteBuffer_reg[6][0]  ( .D(n3293), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n698) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][19]  ( .D(n3526), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n699) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][18]  ( .D(n3527), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n700) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][17]  ( .D(n3528), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n701) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][16]  ( .D(n3529), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n702) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][15]  ( .D(n3530), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n703) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][14]  ( .D(n3531), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n704) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][13]  ( .D(n3532), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n705) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][12]  ( .D(n3533), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n706) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][11]  ( .D(n3534), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n707) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][10]  ( .D(n3535), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n708) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][9]  ( .D(n3536), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n709) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][8]  ( .D(n3537), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n710) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][7]  ( .D(n3538), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n711) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][6]  ( .D(n3539), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n712) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][5]  ( .D(n3540), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n713) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][4]  ( .D(n3541), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n714) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][3]  ( .D(n3542), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n715) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][2]  ( .D(n3543), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n737) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][1]  ( .D(n3544), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n738) );
  DFFNSRX2TS \dataToWriteBuffer_reg[3][0]  ( .D(n3545), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n739) );
  DFFNSRX2TS \addressToWriteBuffer_reg[3][7]  ( .D(n3310), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n24), .QN(n79) );
  DFFNSRX2TS \addressToWriteBuffer_reg[3][6]  ( .D(n3311), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n23), .QN(n78) );
  DFFNSRX2TS \addressToWriteBuffer_reg[3][5]  ( .D(n3312), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n22), .QN(n77) );
  DFFNSRX2TS \addressToWriteBuffer_reg[3][4]  ( .D(n3313), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n21), .QN(n76) );
  DFFNSRX2TS \addressToWriteBuffer_reg[3][3]  ( .D(n3314), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n20), .QN(n75) );
  DFFNSRX2TS \addressToWriteBuffer_reg[3][2]  ( .D(n3315), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n19), .QN(n74) );
  DFFNSRX2TS \addressToWriteBuffer_reg[3][1]  ( .D(n3316), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n18), .QN(n73) );
  DFFNSRX2TS \addressToWriteBuffer_reg[3][0]  ( .D(n3317), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n17), .QN(n72) );
  DFFNSRX2TS \nextEmptyBuffer_reg[1]  ( .D(n3643), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n347), .QN(n910) );
  DFFNSRX2TS \nextEmptyBuffer_reg[0]  ( .D(n3644), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n5), .QN(n1) );
  DFFNSRX2TS \prevRequesterPort_B_reg[0]  ( .D(n3265), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\prevRequesterPort_B[0] ), .QN(n348) );
  EDFFX2TS \readReady_Concatenated_reg[2]  ( .D(N10030), .E(n2497), .CK(clk), 
        .Q(readReady_EAST) );
  EDFFX2TS \readReady_Concatenated_reg[0]  ( .D(N10010), .E(n2495), .CK(clk), 
        .Q(readReady_NORTH) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[2][5]  ( .D(n3177), .CK(clk), 
        .Q(requesterAddressOut_EAST[5]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[2][4]  ( .D(n3176), .CK(clk), 
        .Q(requesterAddressOut_EAST[4]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[2][3]  ( .D(n3175), .CK(clk), 
        .Q(requesterAddressOut_EAST[3]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[2][2]  ( .D(n3174), .CK(clk), 
        .Q(requesterAddressOut_EAST[2]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[2][1]  ( .D(n3173), .CK(clk), 
        .Q(requesterAddressOut_EAST[1]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[2][0]  ( .D(n3172), .CK(clk), 
        .Q(requesterAddressOut_EAST[0]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[1][5]  ( .D(n3171), .CK(clk), 
        .Q(requesterAddressOut_SOUTH[5]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[1][4]  ( .D(n3170), .CK(clk), 
        .Q(requesterAddressOut_SOUTH[4]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[1][3]  ( .D(n3169), .CK(clk), 
        .Q(requesterAddressOut_SOUTH[3]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[1][2]  ( .D(n3168), .CK(clk), 
        .Q(requesterAddressOut_SOUTH[2]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[1][1]  ( .D(n3167), .CK(clk), 
        .Q(requesterAddressOut_SOUTH[1]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[1][0]  ( .D(n3166), .CK(clk), 
        .Q(requesterAddressOut_SOUTH[0]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[3][5]  ( .D(n3183), .CK(clk), 
        .Q(requesterAddressOut_WEST[5]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[3][4]  ( .D(n3182), .CK(clk), 
        .Q(requesterAddressOut_WEST[4]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[3][3]  ( .D(n3181), .CK(clk), 
        .Q(requesterAddressOut_WEST[3]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[3][2]  ( .D(n3180), .CK(clk), 
        .Q(requesterAddressOut_WEST[2]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[3][1]  ( .D(n3179), .CK(clk), 
        .Q(requesterAddressOut_WEST[1]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[3][0]  ( .D(n3178), .CK(clk), 
        .Q(requesterAddressOut_WEST[0]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[0][5]  ( .D(n3165), .CK(clk), 
        .Q(requesterAddressOut_NORTH[5]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[0][4]  ( .D(n3164), .CK(clk), 
        .Q(requesterAddressOut_NORTH[4]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[0][3]  ( .D(n3163), .CK(clk), 
        .Q(requesterAddressOut_NORTH[3]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[0][2]  ( .D(n3162), .CK(clk), 
        .Q(requesterAddressOut_NORTH[2]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[0][1]  ( .D(n3161), .CK(clk), 
        .Q(requesterAddressOut_NORTH[1]) );
  DFFQX1TS \requesterAddressOut_Concatenated_reg[0][0]  ( .D(n3160), .CK(clk), 
        .Q(requesterAddressOut_NORTH[0]) );
  TLATXLTS \dataOut_Concatenated_reg[2][31]  ( .G(clk), .D(N10182), .Q(
        cacheDataOut_EAST[31]) );
  TLATXLTS \dataOut_Concatenated_reg[2][30]  ( .G(clk), .D(N10181), .Q(
        cacheDataOut_EAST[30]) );
  TLATXLTS \dataOut_Concatenated_reg[2][29]  ( .G(clk), .D(N10180), .Q(
        cacheDataOut_EAST[29]) );
  TLATXLTS \dataOut_Concatenated_reg[2][28]  ( .G(clk), .D(N10179), .Q(
        cacheDataOut_EAST[28]) );
  TLATXLTS \dataOut_Concatenated_reg[2][27]  ( .G(clk), .D(N10178), .Q(
        cacheDataOut_EAST[27]) );
  TLATXLTS \dataOut_Concatenated_reg[2][26]  ( .G(clk), .D(N10177), .Q(
        cacheDataOut_EAST[26]) );
  TLATXLTS \dataOut_Concatenated_reg[2][25]  ( .G(clk), .D(N10176), .Q(
        cacheDataOut_EAST[25]) );
  TLATXLTS \dataOut_Concatenated_reg[2][24]  ( .G(clk), .D(N10175), .Q(
        cacheDataOut_EAST[24]) );
  TLATXLTS \dataOut_Concatenated_reg[2][23]  ( .G(clk), .D(N10174), .Q(
        cacheDataOut_EAST[23]) );
  TLATXLTS \dataOut_Concatenated_reg[2][22]  ( .G(clk), .D(N10173), .Q(
        cacheDataOut_EAST[22]) );
  TLATXLTS \dataOut_Concatenated_reg[2][21]  ( .G(clk), .D(N10172), .Q(
        cacheDataOut_EAST[21]) );
  TLATXLTS \dataOut_Concatenated_reg[2][20]  ( .G(clk), .D(N10171), .Q(
        cacheDataOut_EAST[20]) );
  TLATXLTS \dataOut_Concatenated_reg[2][19]  ( .G(clk), .D(N10170), .Q(
        cacheDataOut_EAST[19]) );
  TLATXLTS \dataOut_Concatenated_reg[2][18]  ( .G(clk), .D(N10169), .Q(
        cacheDataOut_EAST[18]) );
  TLATXLTS \dataOut_Concatenated_reg[2][17]  ( .G(clk), .D(N10168), .Q(
        cacheDataOut_EAST[17]) );
  TLATXLTS \dataOut_Concatenated_reg[2][16]  ( .G(clk), .D(N10167), .Q(
        cacheDataOut_EAST[16]) );
  TLATXLTS \dataOut_Concatenated_reg[2][15]  ( .G(clk), .D(N10166), .Q(
        cacheDataOut_EAST[15]) );
  TLATXLTS \dataOut_Concatenated_reg[2][14]  ( .G(clk), .D(N10165), .Q(
        cacheDataOut_EAST[14]) );
  TLATXLTS \dataOut_Concatenated_reg[2][13]  ( .G(clk), .D(N10164), .Q(
        cacheDataOut_EAST[13]) );
  TLATXLTS \dataOut_Concatenated_reg[2][12]  ( .G(clk), .D(N10163), .Q(
        cacheDataOut_EAST[12]) );
  TLATXLTS \dataOut_Concatenated_reg[2][11]  ( .G(clk), .D(N10162), .Q(
        cacheDataOut_EAST[11]) );
  TLATXLTS \dataOut_Concatenated_reg[2][10]  ( .G(clk), .D(N10161), .Q(
        cacheDataOut_EAST[10]) );
  TLATXLTS \dataOut_Concatenated_reg[2][9]  ( .G(clk), .D(N10160), .Q(
        cacheDataOut_EAST[9]) );
  TLATXLTS \dataOut_Concatenated_reg[2][8]  ( .G(clk), .D(N10159), .Q(
        cacheDataOut_EAST[8]) );
  TLATXLTS \dataOut_Concatenated_reg[2][7]  ( .G(clk), .D(N10158), .Q(
        cacheDataOut_EAST[7]) );
  TLATXLTS \dataOut_Concatenated_reg[2][6]  ( .G(clk), .D(N10157), .Q(
        cacheDataOut_EAST[6]) );
  TLATXLTS \dataOut_Concatenated_reg[2][5]  ( .G(clk), .D(N10156), .Q(
        cacheDataOut_EAST[5]) );
  TLATXLTS \dataOut_Concatenated_reg[2][4]  ( .G(clk), .D(N10155), .Q(
        cacheDataOut_EAST[4]) );
  TLATXLTS \dataOut_Concatenated_reg[2][3]  ( .G(clk), .D(N10154), .Q(
        cacheDataOut_EAST[3]) );
  TLATXLTS \dataOut_Concatenated_reg[2][2]  ( .G(clk), .D(N10153), .Q(
        cacheDataOut_EAST[2]) );
  TLATXLTS \dataOut_Concatenated_reg[2][1]  ( .G(clk), .D(N10152), .Q(
        cacheDataOut_EAST[1]) );
  TLATXLTS \dataOut_Concatenated_reg[2][0]  ( .G(clk), .D(N10151), .Q(
        cacheDataOut_EAST[0]) );
  TLATXLTS \dataOut_Concatenated_reg[1][31]  ( .G(clk), .D(N10148), .Q(
        cacheDataOut_SOUTH[31]) );
  TLATXLTS \dataOut_Concatenated_reg[1][30]  ( .G(clk), .D(N10147), .Q(
        cacheDataOut_SOUTH[30]) );
  TLATXLTS \dataOut_Concatenated_reg[1][29]  ( .G(clk), .D(N10146), .Q(
        cacheDataOut_SOUTH[29]) );
  TLATXLTS \dataOut_Concatenated_reg[1][28]  ( .G(clk), .D(N10145), .Q(
        cacheDataOut_SOUTH[28]) );
  TLATXLTS \dataOut_Concatenated_reg[1][27]  ( .G(clk), .D(N10144), .Q(
        cacheDataOut_SOUTH[27]) );
  TLATXLTS \dataOut_Concatenated_reg[1][26]  ( .G(clk), .D(N10143), .Q(
        cacheDataOut_SOUTH[26]) );
  TLATXLTS \dataOut_Concatenated_reg[1][25]  ( .G(clk), .D(N10142), .Q(
        cacheDataOut_SOUTH[25]) );
  TLATXLTS \dataOut_Concatenated_reg[1][24]  ( .G(clk), .D(N10141), .Q(
        cacheDataOut_SOUTH[24]) );
  TLATXLTS \dataOut_Concatenated_reg[1][23]  ( .G(clk), .D(N10140), .Q(
        cacheDataOut_SOUTH[23]) );
  TLATXLTS \dataOut_Concatenated_reg[1][22]  ( .G(clk), .D(N10139), .Q(
        cacheDataOut_SOUTH[22]) );
  TLATXLTS \dataOut_Concatenated_reg[1][21]  ( .G(clk), .D(N10138), .Q(
        cacheDataOut_SOUTH[21]) );
  TLATXLTS \dataOut_Concatenated_reg[1][20]  ( .G(clk), .D(N10137), .Q(
        cacheDataOut_SOUTH[20]) );
  TLATXLTS \dataOut_Concatenated_reg[1][19]  ( .G(clk), .D(N10136), .Q(
        cacheDataOut_SOUTH[19]) );
  TLATXLTS \dataOut_Concatenated_reg[1][18]  ( .G(clk), .D(N10135), .Q(
        cacheDataOut_SOUTH[18]) );
  TLATXLTS \dataOut_Concatenated_reg[1][17]  ( .G(clk), .D(N10134), .Q(
        cacheDataOut_SOUTH[17]) );
  TLATXLTS \dataOut_Concatenated_reg[1][16]  ( .G(clk), .D(N10133), .Q(
        cacheDataOut_SOUTH[16]) );
  TLATXLTS \dataOut_Concatenated_reg[1][15]  ( .G(clk), .D(N10132), .Q(
        cacheDataOut_SOUTH[15]) );
  TLATXLTS \dataOut_Concatenated_reg[1][14]  ( .G(clk), .D(N10131), .Q(
        cacheDataOut_SOUTH[14]) );
  TLATXLTS \dataOut_Concatenated_reg[1][13]  ( .G(clk), .D(N10130), .Q(
        cacheDataOut_SOUTH[13]) );
  TLATXLTS \dataOut_Concatenated_reg[1][12]  ( .G(clk), .D(N10129), .Q(
        cacheDataOut_SOUTH[12]) );
  TLATXLTS \dataOut_Concatenated_reg[1][11]  ( .G(clk), .D(N10128), .Q(
        cacheDataOut_SOUTH[11]) );
  TLATXLTS \dataOut_Concatenated_reg[1][10]  ( .G(clk), .D(N10127), .Q(
        cacheDataOut_SOUTH[10]) );
  TLATXLTS \dataOut_Concatenated_reg[1][9]  ( .G(clk), .D(N10126), .Q(
        cacheDataOut_SOUTH[9]) );
  TLATXLTS \dataOut_Concatenated_reg[1][8]  ( .G(clk), .D(N10125), .Q(
        cacheDataOut_SOUTH[8]) );
  TLATXLTS \dataOut_Concatenated_reg[1][7]  ( .G(clk), .D(N10124), .Q(
        cacheDataOut_SOUTH[7]) );
  TLATXLTS \dataOut_Concatenated_reg[1][6]  ( .G(clk), .D(N10123), .Q(
        cacheDataOut_SOUTH[6]) );
  TLATXLTS \dataOut_Concatenated_reg[1][5]  ( .G(clk), .D(N10122), .Q(
        cacheDataOut_SOUTH[5]) );
  TLATXLTS \dataOut_Concatenated_reg[1][4]  ( .G(clk), .D(N10121), .Q(
        cacheDataOut_SOUTH[4]) );
  TLATXLTS \dataOut_Concatenated_reg[1][3]  ( .G(clk), .D(N10120), .Q(
        cacheDataOut_SOUTH[3]) );
  TLATXLTS \dataOut_Concatenated_reg[1][2]  ( .G(clk), .D(N10119), .Q(
        cacheDataOut_SOUTH[2]) );
  TLATXLTS \dataOut_Concatenated_reg[1][1]  ( .G(clk), .D(N10118), .Q(
        cacheDataOut_SOUTH[1]) );
  TLATXLTS \dataOut_Concatenated_reg[1][0]  ( .G(clk), .D(N10117), .Q(
        cacheDataOut_SOUTH[0]) );
  TLATXLTS \dataOut_Concatenated_reg[3][31]  ( .G(clk), .D(N10216), .Q(
        cacheDataOut_WEST[31]) );
  TLATXLTS \dataOut_Concatenated_reg[3][30]  ( .G(clk), .D(N10215), .Q(
        cacheDataOut_WEST[30]) );
  TLATXLTS \dataOut_Concatenated_reg[3][29]  ( .G(clk), .D(N10214), .Q(
        cacheDataOut_WEST[29]) );
  TLATXLTS \dataOut_Concatenated_reg[3][28]  ( .G(clk), .D(N10213), .Q(
        cacheDataOut_WEST[28]) );
  TLATXLTS \dataOut_Concatenated_reg[3][27]  ( .G(clk), .D(N10212), .Q(
        cacheDataOut_WEST[27]) );
  TLATXLTS \dataOut_Concatenated_reg[3][26]  ( .G(clk), .D(N10211), .Q(
        cacheDataOut_WEST[26]) );
  TLATXLTS \dataOut_Concatenated_reg[3][25]  ( .G(clk), .D(N10210), .Q(
        cacheDataOut_WEST[25]) );
  TLATXLTS \dataOut_Concatenated_reg[3][24]  ( .G(clk), .D(N10209), .Q(
        cacheDataOut_WEST[24]) );
  TLATXLTS \dataOut_Concatenated_reg[3][23]  ( .G(clk), .D(N10208), .Q(
        cacheDataOut_WEST[23]) );
  TLATXLTS \dataOut_Concatenated_reg[3][22]  ( .G(clk), .D(N10207), .Q(
        cacheDataOut_WEST[22]) );
  TLATXLTS \dataOut_Concatenated_reg[3][21]  ( .G(clk), .D(N10206), .Q(
        cacheDataOut_WEST[21]) );
  TLATXLTS \dataOut_Concatenated_reg[3][20]  ( .G(clk), .D(N10205), .Q(
        cacheDataOut_WEST[20]) );
  TLATXLTS \dataOut_Concatenated_reg[3][19]  ( .G(clk), .D(N10204), .Q(
        cacheDataOut_WEST[19]) );
  TLATXLTS \dataOut_Concatenated_reg[3][18]  ( .G(clk), .D(N10203), .Q(
        cacheDataOut_WEST[18]) );
  TLATXLTS \dataOut_Concatenated_reg[3][17]  ( .G(clk), .D(N10202), .Q(
        cacheDataOut_WEST[17]) );
  TLATXLTS \dataOut_Concatenated_reg[3][16]  ( .G(clk), .D(N10201), .Q(
        cacheDataOut_WEST[16]) );
  TLATXLTS \dataOut_Concatenated_reg[3][15]  ( .G(clk), .D(N10200), .Q(
        cacheDataOut_WEST[15]) );
  TLATXLTS \dataOut_Concatenated_reg[3][14]  ( .G(clk), .D(N10199), .Q(
        cacheDataOut_WEST[14]) );
  TLATXLTS \dataOut_Concatenated_reg[3][13]  ( .G(clk), .D(N10198), .Q(
        cacheDataOut_WEST[13]) );
  TLATXLTS \dataOut_Concatenated_reg[3][12]  ( .G(clk), .D(N10197), .Q(
        cacheDataOut_WEST[12]) );
  TLATXLTS \dataOut_Concatenated_reg[3][11]  ( .G(clk), .D(N10196), .Q(
        cacheDataOut_WEST[11]) );
  TLATXLTS \dataOut_Concatenated_reg[3][10]  ( .G(clk), .D(N10195), .Q(
        cacheDataOut_WEST[10]) );
  TLATXLTS \dataOut_Concatenated_reg[3][9]  ( .G(clk), .D(N10194), .Q(
        cacheDataOut_WEST[9]) );
  TLATXLTS \dataOut_Concatenated_reg[3][8]  ( .G(clk), .D(N10193), .Q(
        cacheDataOut_WEST[8]) );
  TLATXLTS \dataOut_Concatenated_reg[3][7]  ( .G(clk), .D(N10192), .Q(
        cacheDataOut_WEST[7]) );
  TLATXLTS \dataOut_Concatenated_reg[3][6]  ( .G(clk), .D(N10191), .Q(
        cacheDataOut_WEST[6]) );
  TLATXLTS \dataOut_Concatenated_reg[3][5]  ( .G(clk), .D(N10190), .Q(
        cacheDataOut_WEST[5]) );
  TLATXLTS \dataOut_Concatenated_reg[3][4]  ( .G(clk), .D(N10189), .Q(
        cacheDataOut_WEST[4]) );
  TLATXLTS \dataOut_Concatenated_reg[3][3]  ( .G(clk), .D(N10188), .Q(
        cacheDataOut_WEST[3]) );
  TLATXLTS \dataOut_Concatenated_reg[3][2]  ( .G(clk), .D(N10187), .Q(
        cacheDataOut_WEST[2]) );
  TLATXLTS \dataOut_Concatenated_reg[3][1]  ( .G(clk), .D(N10186), .Q(
        cacheDataOut_WEST[1]) );
  TLATXLTS \dataOut_Concatenated_reg[3][0]  ( .G(clk), .D(N10185), .Q(
        cacheDataOut_WEST[0]) );
  TLATXLTS \dataOut_Concatenated_reg[0][31]  ( .G(clk), .D(N10114), .Q(
        cacheDataOut_NORTH[31]) );
  TLATXLTS \dataOut_Concatenated_reg[0][30]  ( .G(clk), .D(N10113), .Q(
        cacheDataOut_NORTH[30]) );
  TLATXLTS \dataOut_Concatenated_reg[0][29]  ( .G(clk), .D(N10112), .Q(
        cacheDataOut_NORTH[29]) );
  TLATXLTS \dataOut_Concatenated_reg[0][28]  ( .G(clk), .D(N10111), .Q(
        cacheDataOut_NORTH[28]) );
  TLATXLTS \dataOut_Concatenated_reg[0][27]  ( .G(clk), .D(N10110), .Q(
        cacheDataOut_NORTH[27]) );
  TLATXLTS \dataOut_Concatenated_reg[0][26]  ( .G(clk), .D(N10109), .Q(
        cacheDataOut_NORTH[26]) );
  TLATXLTS \dataOut_Concatenated_reg[0][25]  ( .G(clk), .D(N10108), .Q(
        cacheDataOut_NORTH[25]) );
  TLATXLTS \dataOut_Concatenated_reg[0][24]  ( .G(clk), .D(N10107), .Q(
        cacheDataOut_NORTH[24]) );
  TLATXLTS \dataOut_Concatenated_reg[0][23]  ( .G(clk), .D(N10106), .Q(
        cacheDataOut_NORTH[23]) );
  TLATXLTS \dataOut_Concatenated_reg[0][22]  ( .G(clk), .D(N10105), .Q(
        cacheDataOut_NORTH[22]) );
  TLATXLTS \dataOut_Concatenated_reg[0][21]  ( .G(clk), .D(N10104), .Q(
        cacheDataOut_NORTH[21]) );
  TLATXLTS \dataOut_Concatenated_reg[0][20]  ( .G(clk), .D(N10103), .Q(
        cacheDataOut_NORTH[20]) );
  TLATXLTS \dataOut_Concatenated_reg[0][19]  ( .G(clk), .D(N10102), .Q(
        cacheDataOut_NORTH[19]) );
  TLATXLTS \dataOut_Concatenated_reg[0][18]  ( .G(clk), .D(N10101), .Q(
        cacheDataOut_NORTH[18]) );
  TLATXLTS \dataOut_Concatenated_reg[0][17]  ( .G(clk), .D(N10100), .Q(
        cacheDataOut_NORTH[17]) );
  TLATXLTS \dataOut_Concatenated_reg[0][16]  ( .G(clk), .D(N10099), .Q(
        cacheDataOut_NORTH[16]) );
  TLATXLTS \dataOut_Concatenated_reg[0][15]  ( .G(clk), .D(N10098), .Q(
        cacheDataOut_NORTH[15]) );
  TLATXLTS \dataOut_Concatenated_reg[0][14]  ( .G(clk), .D(N10097), .Q(
        cacheDataOut_NORTH[14]) );
  TLATXLTS \dataOut_Concatenated_reg[0][13]  ( .G(clk), .D(N10096), .Q(
        cacheDataOut_NORTH[13]) );
  TLATXLTS \dataOut_Concatenated_reg[0][12]  ( .G(clk), .D(N10095), .Q(
        cacheDataOut_NORTH[12]) );
  TLATXLTS \dataOut_Concatenated_reg[0][11]  ( .G(clk), .D(N10094), .Q(
        cacheDataOut_NORTH[11]) );
  TLATXLTS \dataOut_Concatenated_reg[0][10]  ( .G(clk), .D(N10093), .Q(
        cacheDataOut_NORTH[10]) );
  TLATXLTS \dataOut_Concatenated_reg[0][9]  ( .G(clk), .D(N10092), .Q(
        cacheDataOut_NORTH[9]) );
  TLATXLTS \dataOut_Concatenated_reg[0][8]  ( .G(clk), .D(N10091), .Q(
        cacheDataOut_NORTH[8]) );
  TLATXLTS \dataOut_Concatenated_reg[0][7]  ( .G(clk), .D(N10090), .Q(
        cacheDataOut_NORTH[7]) );
  TLATXLTS \dataOut_Concatenated_reg[0][6]  ( .G(clk), .D(N10089), .Q(
        cacheDataOut_NORTH[6]) );
  TLATXLTS \dataOut_Concatenated_reg[0][5]  ( .G(clk), .D(N10088), .Q(
        cacheDataOut_NORTH[5]) );
  TLATXLTS \dataOut_Concatenated_reg[0][4]  ( .G(clk), .D(N10087), .Q(
        cacheDataOut_NORTH[4]) );
  TLATXLTS \dataOut_Concatenated_reg[0][3]  ( .G(clk), .D(N10086), .Q(
        cacheDataOut_NORTH[3]) );
  TLATXLTS \dataOut_Concatenated_reg[0][2]  ( .G(clk), .D(N10085), .Q(
        cacheDataOut_NORTH[2]) );
  TLATXLTS \dataOut_Concatenated_reg[0][1]  ( .G(clk), .D(N10084), .Q(
        cacheDataOut_NORTH[1]) );
  TLATXLTS \dataOut_Concatenated_reg[0][0]  ( .G(clk), .D(N10083), .Q(
        cacheDataOut_NORTH[0]) );
  EDFFX2TS \readReady_Concatenated_reg[1]  ( .D(N10020), .E(n2496), .CK(clk), 
        .Q(readReady_SOUTH) );
  EDFFX2TS \readReady_Concatenated_reg[3]  ( .D(N10040), .E(n2494), .CK(clk), 
        .Q(readReady_WEST) );
  DFFNSRX2TS \nextEmptyBuffer_reg[2]  ( .D(n3642), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n4), .QN(n880) );
  DFFNSRXLTS \requesterPortBuffer_reg[2][1]  ( .D(n2098), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n2096) );
  DFFNSRXLTS \requesterPortBuffer_reg[3][1]  ( .D(n2101), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n2081) );
  DFFNSRXLTS \requesterPortBuffer_reg[3][0]  ( .D(n2103), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n2083) );
  DFFNSRXLTS \addressToWriteBuffer_reg[7][7]  ( .D(n3278), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n2079) );
  DFFNSRXLTS \dataToWriteBuffer_reg[7][8]  ( .D(n3409), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n2017) );
  DFFNSRXLTS \dataToWriteBuffer_reg[7][7]  ( .D(n3410), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n2015) );
  DFFNSRXLTS \dataToWriteBuffer_reg[7][6]  ( .D(n3411), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n2013) );
  DFFNSRXLTS \dataToWriteBuffer_reg[7][5]  ( .D(n3412), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n2012) );
  DFFNSRXLTS \dataToWriteBuffer_reg[7][4]  ( .D(n3413), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n2011) );
  DFFNSRXLTS \dataToWriteBuffer_reg[7][3]  ( .D(n3414), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n2010) );
  DFFNSRXLTS \dataToWriteBuffer_reg[7][2]  ( .D(n3415), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n2009) );
  DFFNSRXLTS \dataToWriteBuffer_reg[7][1]  ( .D(n3416), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n2008) );
  DFFNSRXLTS \dataToWriteBuffer_reg[7][0]  ( .D(n3417), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n2007) );
  DFFNSRXLTS \dataToWriteBuffer_reg[7][28]  ( .D(n3389), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n2057) );
  DFFNSRXLTS \dataToWriteBuffer_reg[7][27]  ( .D(n3390), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n2055) );
  DFFNSRXLTS \dataToWriteBuffer_reg[7][26]  ( .D(n3391), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n2053) );
  DFFNSRXLTS \dataToWriteBuffer_reg[7][25]  ( .D(n3392), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n2051) );
  DFFNSRXLTS \dataToWriteBuffer_reg[7][24]  ( .D(n3393), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n2049) );
  DFFNSRXLTS \dataToWriteBuffer_reg[7][23]  ( .D(n3394), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n2047) );
  DFFNSRXLTS \dataToWriteBuffer_reg[7][22]  ( .D(n3395), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n2045) );
  DFFNSRXLTS \dataToWriteBuffer_reg[7][11]  ( .D(n3406), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n2023) );
  DFFNSRXLTS \dataToWriteBuffer_reg[7][21]  ( .D(n3396), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n2043) );
  DFFNSRXLTS \dataToWriteBuffer_reg[7][20]  ( .D(n3397), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n2041) );
  DFFNSRXLTS \dataToWriteBuffer_reg[7][19]  ( .D(n3398), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n2039) );
  DFFNSRXLTS \dataToWriteBuffer_reg[7][18]  ( .D(n3399), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n2037) );
  DFFNSRXLTS \dataToWriteBuffer_reg[7][17]  ( .D(n3400), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n2035) );
  DFFNSRXLTS \dataToWriteBuffer_reg[7][16]  ( .D(n3401), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n2033) );
  DFFNSRXLTS \dataToWriteBuffer_reg[7][15]  ( .D(n3402), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n2031) );
  DFFNSRXLTS \dataToWriteBuffer_reg[7][14]  ( .D(n3403), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n2029) );
  DFFNSRXLTS \dataToWriteBuffer_reg[7][13]  ( .D(n3404), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n2027) );
  DFFNSRXLTS \dataToWriteBuffer_reg[7][12]  ( .D(n3405), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n2025) );
  DFFNSRXLTS \dataToWriteBuffer_reg[7][10]  ( .D(n3407), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n2021) );
  DFFNSRXLTS \dataToWriteBuffer_reg[7][9]  ( .D(n3408), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n2019) );
  DFFNSRXLTS \dataToWriteBuffer_reg[7][31]  ( .D(n3386), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n2063) );
  DFFNSRXLTS \dataToWriteBuffer_reg[7][30]  ( .D(n3387), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n2061) );
  DFFNSRXLTS \dataToWriteBuffer_reg[7][29]  ( .D(n3388), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n2059) );
  DFFNSRXLTS \addressToWriteBuffer_reg[7][6]  ( .D(n3279), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n2077) );
  DFFNSRXLTS \addressToWriteBuffer_reg[7][5]  ( .D(n3280), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n2075) );
  DFFNSRXLTS \addressToWriteBuffer_reg[7][4]  ( .D(n3281), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n2073) );
  DFFNSRXLTS \addressToWriteBuffer_reg[7][3]  ( .D(n3282), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n2071) );
  DFFNSRXLTS \addressToWriteBuffer_reg[7][2]  ( .D(n3283), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n2069) );
  DFFNSRXLTS \addressToWriteBuffer_reg[7][1]  ( .D(n3284), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n2067) );
  DFFNSRXLTS \addressToWriteBuffer_reg[7][0]  ( .D(n3285), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n2065) );
  DFFNSRXLTS \requesterPortBuffer_reg[1][0]  ( .D(n3267), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n46) );
  DFFNSRXLTS \requesterPortBuffer_reg[1][1]  ( .D(n3266), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n47) );
  DFFNSRXLTS \isRead_reg[0]  ( .D(n3343), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .QN(n45) );
  DFFNSRXLTS \dataToWriteBuffer_reg[6][15]  ( .D(n3434), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1828) );
  DFFNSRXLTS \dataToWriteBuffer_reg[6][14]  ( .D(n3435), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1827) );
  DFFNSRXLTS \dataToWriteBuffer_reg[6][13]  ( .D(n3436), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1826) );
  DFFNSRXLTS \dataToWriteBuffer_reg[6][12]  ( .D(n3437), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1825) );
  DFFNSRXLTS \dataToWriteBuffer_reg[6][11]  ( .D(n3438), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1823) );
  DFFNSRXLTS \dataToWriteBuffer_reg[6][10]  ( .D(n3439), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1822) );
  DFFNSRXLTS \dataToWriteBuffer_reg[6][9]  ( .D(n3440), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1821) );
  DFFNSRXLTS \dataToWriteBuffer_reg[6][8]  ( .D(n3441), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1820) );
  DFFNSRXLTS \dataToWriteBuffer_reg[6][7]  ( .D(n3442), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1818) );
  DFFNSRXLTS \dataToWriteBuffer_reg[6][6]  ( .D(n3443), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1817) );
  DFFNSRXLTS \dataToWriteBuffer_reg[6][5]  ( .D(n3444), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1816) );
  DFFNSRXLTS \dataToWriteBuffer_reg[6][4]  ( .D(n3445), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n1815) );
  DFFNSRXLTS \isWrite_reg[2]  ( .D(n3383), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .QN(n932) );
  DFFNSRXLTS \isWrite_reg[6]  ( .D(n3379), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .QN(n930) );
  DFFNSRXLTS \requesterPortBuffer_reg[5][1]  ( .D(n2100), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n653) );
  DFFNSRXLTS \requesterPortBuffer_reg[5][0]  ( .D(n2102), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n654) );
  DFFNSRXLTS \isWrite_reg[4]  ( .D(n3381), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .QN(n931) );
  DFFNSRXLTS \requesterPortBuffer_reg[6][1]  ( .D(n2104), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n655) );
  DFFNSRXLTS \requesterPortBuffer_reg[4][1]  ( .D(n2099), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n650) );
  DFFNSRXLTS \requesterPortBuffer_reg[2][0]  ( .D(n652), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[2][0] ) );
  DFFNSRXLTS \isWrite_reg[5]  ( .D(n758), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        n2093) );
  DFFNSRXLTS \requesterPortBuffer_reg[4][0]  ( .D(n651), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[4][0] ) );
  DFFNSRXLTS \requesterPortBuffer_reg[6][0]  ( .D(n656), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[6][0] ) );
  DFFNSRXLTS \isWrite_reg[3]  ( .D(n814), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        n2091) );
  DFFNSRXLTS \requesterPortBuffer_reg[7][1]  ( .D(n3252), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n658) );
  DFFNSRXLTS \requesterPortBuffer_reg[7][0]  ( .D(n3253), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n657) );
  DFFNSRXLTS \isWrite_reg[7]  ( .D(n3378), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n2094) );
  DFFNSRXLTS prevMemRead_A_reg ( .D(n2106), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .QN(n818) );
  DFFNSRXLTS prevMemRead_B_reg ( .D(n3344), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .QN(n817) );
  DFFNSRXLTS \requesterPortBuffer_reg[0][0]  ( .D(n2105), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[0][0] ) );
  DFFNSRXLTS \requesterPortBuffer_reg[0][1]  ( .D(n3268), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(\requesterPortBuffer[0][1] ), .QN(n674) );
  DFFNSRXLTS \isRead_reg[1]  ( .D(n3345), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .QN(n659) );
  DFFNSRXLTS \prevRequesterPort_B_reg[1]  ( .D(n3264), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2), .QN(n14) );
  DFFNSRXLTS \prevRequesterPort_A_reg[1]  ( .D(n3251), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3), .QN(n13) );
  DFFNSRXLTS \prevRequesterPort_A_reg[0]  ( .D(n3250), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n740), .QN(n938) );
  DFFNSRXLTS \addressToWriteBuffer_reg[0][3]  ( .D(n3338), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n779), .QN(n945) );
  DFFNSRXLTS \isWrite_reg[0]  ( .D(n3385), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n2089), .QN(n933) );
  DFFNSRXLTS \addressToWriteBuffer_reg[0][7]  ( .D(n3334), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n775), .QN(n943) );
  DFFNSRXLTS \addressToWriteBuffer_reg[0][6]  ( .D(n3335), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n776), .QN(n939) );
  DFFNSRXLTS \addressToWriteBuffer_reg[0][5]  ( .D(n3336), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n777), .QN(n944) );
  DFFNSRXLTS \addressToWriteBuffer_reg[0][4]  ( .D(n3337), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n778), .QN(n940) );
  DFFNSRXLTS \addressToWriteBuffer_reg[0][2]  ( .D(n3339), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n780), .QN(n941) );
  DFFNSRXLTS \addressToWriteBuffer_reg[0][1]  ( .D(n3340), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n781), .QN(n942) );
  DFFNSRXLTS \addressToWriteBuffer_reg[0][0]  ( .D(n3341), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n782), .QN(n934) );
  DFFNSRXLTS \requesterAddressBuffer_reg[1][1]  ( .D(n3204), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n672) );
  DFFNSRXLTS \requesterAddressBuffer_reg[1][0]  ( .D(n3203), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n673) );
  DFFNSRXLTS \isWrite_reg[1]  ( .D(n3384), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .QN(n946) );
  DFFNSRXLTS \prevRequesterAddress_B_reg[2]  ( .D(n3200), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_B[2]), .QN(n822) );
  DFFNSRXLTS \prevRequesterAddress_B_reg[1]  ( .D(n3201), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_B[1]), .QN(n823) );
  DFFNSRXLTS \prevRequesterAddress_B_reg[0]  ( .D(n3202), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_B[0]), .QN(n824) );
  DFFNSRXLTS \requesterAddressBuffer_reg[1][5]  ( .D(n3208), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n668) );
  DFFNSRXLTS \requesterAddressBuffer_reg[1][4]  ( .D(n3207), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n669) );
  DFFNSRXLTS \requesterAddressBuffer_reg[1][3]  ( .D(n3206), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n670) );
  DFFNSRXLTS \requesterAddressBuffer_reg[1][2]  ( .D(n3205), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n671) );
  DFFNSRXLTS \prevRequesterAddress_A_reg[2]  ( .D(n3188), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_A[2]), .QN(n828) );
  DFFNSRXLTS \prevRequesterAddress_A_reg[1]  ( .D(n3189), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_A[1]), .QN(n829) );
  DFFNSRXLTS \prevRequesterAddress_A_reg[0]  ( .D(n3190), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_A[0]), .QN(n830) );
  DFFNSRXLTS \prevRequesterAddress_B_reg[5]  ( .D(n3197), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_B[5]), .QN(n819) );
  DFFNSRXLTS \prevRequesterAddress_B_reg[4]  ( .D(n3198), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_B[4]), .QN(n820) );
  DFFNSRXLTS \prevRequesterAddress_B_reg[3]  ( .D(n3199), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_B[3]), .QN(n821) );
  DFFNSRXLTS \prevRequesterAddress_A_reg[5]  ( .D(n3185), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_A[5]), .QN(n825) );
  DFFNSRXLTS \prevRequesterAddress_A_reg[4]  ( .D(n3186), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_A[4]), .QN(n826) );
  DFFNSRXLTS \prevRequesterAddress_A_reg[3]  ( .D(n3187), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(prevRequesterAddress_A[3]), .QN(n827) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][31]  ( .D(n3610), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n783), .QN(n897) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][30]  ( .D(n3611), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n784), .QN(n905) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][29]  ( .D(n3612), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n785), .QN(n906) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][28]  ( .D(n3613), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n786), .QN(n907) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][27]  ( .D(n3614), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n787), .QN(n908) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][26]  ( .D(n3615), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n788), .QN(n909) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][25]  ( .D(n3616), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n789), .QN(n911) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][24]  ( .D(n3617), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n790), .QN(n898) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][23]  ( .D(n3618), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n791), .QN(n912) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][22]  ( .D(n3619), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n792), .QN(n913) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][21]  ( .D(n3620), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n793), .QN(n899) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][20]  ( .D(n3621), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n716), .QN(n914) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][19]  ( .D(n3622), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n717), .QN(n915) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][18]  ( .D(n3623), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n718), .QN(n916) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][17]  ( .D(n3624), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n719), .QN(n917) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][16]  ( .D(n3625), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n720), .QN(n900) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][15]  ( .D(n3626), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n721), .QN(n918) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][14]  ( .D(n3627), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n722), .QN(n919) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][13]  ( .D(n3628), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n723), .QN(n920) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][12]  ( .D(n3629), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n724), .QN(n901) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][11]  ( .D(n3630), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n725), .QN(n921) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][10]  ( .D(n3631), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n726), .QN(n922) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][9]  ( .D(n3632), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n727), .QN(n923) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][8]  ( .D(n3633), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n728), .QN(n902) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][7]  ( .D(n3634), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n729), .QN(n924) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][6]  ( .D(n3635), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n730), .QN(n925) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][5]  ( .D(n3636), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n731), .QN(n926) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][4]  ( .D(n3637), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n732), .QN(n903) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][3]  ( .D(n3638), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n733), .QN(n927) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][2]  ( .D(n3639), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n734), .QN(n928) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][1]  ( .D(n3640), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n735), .QN(n929) );
  DFFNSRXLTS \dataToWriteBuffer_reg[0][0]  ( .D(n3641), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n736), .QN(n904) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][15]  ( .D(n3562), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1907), .QN(n848) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][14]  ( .D(n3563), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1906), .QN(n849) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][13]  ( .D(n3564), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1905), .QN(n850) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][12]  ( .D(n3565), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1904), .QN(n851) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][11]  ( .D(n3566), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1903), .QN(n852) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][10]  ( .D(n3567), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1902), .QN(n853) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][9]  ( .D(n3568), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1901), .QN(n854) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][8]  ( .D(n3569), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1900), .QN(n855) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][7]  ( .D(n3570), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1899), .QN(n856) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][6]  ( .D(n3571), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1898), .QN(n857) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][5]  ( .D(n3572), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1897), .QN(n858) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][4]  ( .D(n3573), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1896), .QN(n859) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][3]  ( .D(n3574), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1895), .QN(n860) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][2]  ( .D(n3575), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1894), .QN(n861) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][0]  ( .D(n3577), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1892), .QN(n863) );
  DFFNSRXLTS \requesterAddressBuffer_reg[0][1]  ( .D(n774), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressBuffer[0][1] ) );
  DFFNSRXLTS \requesterAddressBuffer_reg[0][0]  ( .D(n773), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressBuffer[0][0] ) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][30]  ( .D(n3547), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1890), .QN(n833) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][29]  ( .D(n3548), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1889), .QN(n834) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][28]  ( .D(n3549), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1888), .QN(n835) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][27]  ( .D(n3550), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1887), .QN(n836) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][26]  ( .D(n3551), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1886), .QN(n837) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][25]  ( .D(n3552), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1885), .QN(n838) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][24]  ( .D(n3553), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1884), .QN(n839) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][23]  ( .D(n3554), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1883), .QN(n840) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][22]  ( .D(n3555), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1882), .QN(n841) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][21]  ( .D(n3556), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1881), .QN(n842) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][20]  ( .D(n3557), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1924), .QN(n843) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][19]  ( .D(n3558), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1923), .QN(n844) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][18]  ( .D(n3559), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1910), .QN(n845) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][17]  ( .D(n3560), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1909), .QN(n846) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][16]  ( .D(n3561), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1908), .QN(n847) );
  DFFNSRXLTS \requesterAddressBuffer_reg[0][5]  ( .D(n797), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressBuffer[0][5] ) );
  DFFNSRXLTS \requesterAddressBuffer_reg[0][4]  ( .D(n796), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressBuffer[0][4] ) );
  DFFNSRXLTS \requesterAddressBuffer_reg[0][3]  ( .D(n795), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressBuffer[0][3] ) );
  DFFNSRXLTS \requesterAddressBuffer_reg[0][2]  ( .D(n794), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressBuffer[0][2] ) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][31]  ( .D(n3546), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1891), .QN(n832) );
  DFFNSRXLTS \dataToWriteBuffer_reg[2][1]  ( .D(n3576), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1893), .QN(n862) );
  DFFNSRXLTS \addressToWriteBuffer_reg[2][7]  ( .D(n3318), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n947) );
  DFFNSRXLTS \addressToWriteBuffer_reg[2][6]  ( .D(n3319), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n948) );
  DFFNSRXLTS \addressToWriteBuffer_reg[2][5]  ( .D(n3320), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n949) );
  DFFNSRXLTS \addressToWriteBuffer_reg[2][4]  ( .D(n3321), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n950) );
  DFFNSRXLTS \addressToWriteBuffer_reg[2][3]  ( .D(n3322), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n951) );
  DFFNSRXLTS \addressToWriteBuffer_reg[2][2]  ( .D(n3323), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n952) );
  DFFNSRXLTS \addressToWriteBuffer_reg[2][1]  ( .D(n3324), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n953) );
  DFFNSRXLTS \addressToWriteBuffer_reg[2][0]  ( .D(n3325), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(n954) );
  DFFNSRXLTS \addressToWriteBuffer_reg[1][5]  ( .D(n3328), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1930), .QN(n662) );
  DFFNSRXLTS \addressToWriteBuffer_reg[1][4]  ( .D(n3329), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1929), .QN(n663) );
  DFFNSRXLTS \addressToWriteBuffer_reg[1][2]  ( .D(n3331), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1927), .QN(n665) );
  DFFNSRXLTS \addressToWriteBuffer_reg[1][1]  ( .D(n3332), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1926), .QN(n666) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][31]  ( .D(n3578), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1964), .QN(n864) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][30]  ( .D(n3579), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1963), .QN(n865) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][29]  ( .D(n3580), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1962), .QN(n866) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][28]  ( .D(n3581), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1961), .QN(n867) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][27]  ( .D(n3582), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1960), .QN(n868) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][26]  ( .D(n3583), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1959), .QN(n869) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][25]  ( .D(n3584), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1958), .QN(n870) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][24]  ( .D(n3585), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1957), .QN(n871) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][23]  ( .D(n3586), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1956), .QN(n872) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][22]  ( .D(n3587), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1955), .QN(n873) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][21]  ( .D(n3588), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1954), .QN(n874) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][20]  ( .D(n3589), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1953), .QN(n875) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][0]  ( .D(n3609), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1933), .QN(n896) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][19]  ( .D(n3590), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1952), .QN(n876) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][18]  ( .D(n3591), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1951), .QN(n877) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][17]  ( .D(n3592), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1950), .QN(n878) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][16]  ( .D(n3593), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1949), .QN(n879) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][15]  ( .D(n3594), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1948), .QN(n881) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][14]  ( .D(n3595), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1947), .QN(n882) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][13]  ( .D(n3596), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1946), .QN(n883) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][12]  ( .D(n3597), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1945), .QN(n884) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][11]  ( .D(n3598), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1944), .QN(n885) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][10]  ( .D(n3599), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1943), .QN(n886) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][9]  ( .D(n3600), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1942), .QN(n887) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][8]  ( .D(n3601), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1941), .QN(n888) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][7]  ( .D(n3602), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1940), .QN(n889) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][6]  ( .D(n3603), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1939), .QN(n890) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][5]  ( .D(n3604), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1938), .QN(n891) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][4]  ( .D(n3605), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1937), .QN(n892) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][3]  ( .D(n3606), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1936), .QN(n893) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][2]  ( .D(n3607), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1935), .QN(n894) );
  DFFNSRXLTS \dataToWriteBuffer_reg[1][1]  ( .D(n3608), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1934), .QN(n895) );
  DFFNSRXLTS \addressToWriteBuffer_reg[1][7]  ( .D(n3326), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1932), .QN(n660) );
  DFFNSRXLTS \addressToWriteBuffer_reg[1][6]  ( .D(n3327), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1931), .QN(n661) );
  DFFNSRXLTS \addressToWriteBuffer_reg[1][3]  ( .D(n3330), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1928), .QN(n664) );
  DFFNSRXLTS \addressToWriteBuffer_reg[1][0]  ( .D(n3333), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(n1925), .QN(n667) );
  DFFNSRXLTS \dataToWriteBuffer_reg[3][31]  ( .D(n3514), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1922) );
  DFFNSRXLTS \dataToWriteBuffer_reg[3][30]  ( .D(n3515), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1921) );
  DFFNSRXLTS \dataToWriteBuffer_reg[3][29]  ( .D(n3516), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1920) );
  DFFNSRXLTS \dataToWriteBuffer_reg[3][28]  ( .D(n3517), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1919) );
  DFFNSRXLTS \dataToWriteBuffer_reg[3][27]  ( .D(n3518), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1918) );
  DFFNSRXLTS \dataToWriteBuffer_reg[3][26]  ( .D(n3519), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1917) );
  DFFNSRXLTS \dataToWriteBuffer_reg[3][25]  ( .D(n3520), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1916) );
  DFFNSRXLTS \dataToWriteBuffer_reg[3][24]  ( .D(n3521), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1915) );
  DFFNSRXLTS \dataToWriteBuffer_reg[3][23]  ( .D(n3522), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1914) );
  DFFNSRXLTS \dataToWriteBuffer_reg[3][22]  ( .D(n3523), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1913) );
  DFFNSRXLTS \dataToWriteBuffer_reg[3][21]  ( .D(n3524), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1912) );
  DFFNSRXLTS \dataToWriteBuffer_reg[3][20]  ( .D(n3525), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n1911) );
  AOI22X1TS U2 ( .A0(n1515), .A1(n378), .B0(n964), .B1(n1729), .Y(n1465) );
  NOR2BX1TS U3 ( .AN(n1499), .B(n102), .Y(n1195) );
  NOR2X1TS U4 ( .A(n1568), .B(n1478), .Y(n1530) );
  NAND2X1TS U5 ( .A(n976), .B(n977), .Y(n1515) );
  NOR2X1TS U6 ( .A(memRead_NORTH), .B(memWrite_NORTH), .Y(n1476) );
  AND3X2TS U7 ( .A(n961), .B(n1025), .C(n1465), .Y(n6) );
  AND2X2TS U8 ( .A(n35), .B(n31), .Y(n7) );
  NAND3X1TS U9 ( .A(n963), .B(n1490), .C(n1531), .Y(n8) );
  AND2X2TS U10 ( .A(n93), .B(n1709), .Y(n9) );
  AND2X2TS U11 ( .A(n810), .B(n92), .Y(n10) );
  OR2X2TS U12 ( .A(n1490), .B(n1465), .Y(n11) );
  AND3X2TS U13 ( .A(n1516), .B(n353), .C(n89), .Y(n12) );
  OR3X1TS U14 ( .A(n1762), .B(n2485), .C(n1763), .Y(n15) );
  OR3X1TS U15 ( .A(n1773), .B(n2485), .C(n1774), .Y(n16) );
  CLKBUFX2TS U16 ( .A(memWrite_WEST), .Y(n25) );
  INVXLTS U17 ( .A(n13), .Y(n26) );
  INVXLTS U18 ( .A(n53), .Y(n27) );
  INVXLTS U19 ( .A(n1606), .Y(n28) );
  INVXLTS U20 ( .A(n28), .Y(n29) );
  INVXLTS U21 ( .A(n1466), .Y(n30) );
  INVXLTS U22 ( .A(n30), .Y(n31) );
  INVXLTS U23 ( .A(n8), .Y(n32) );
  INVXLTS U24 ( .A(n8), .Y(n33) );
  INVXLTS U25 ( .A(n1602), .Y(n34) );
  INVXLTS U26 ( .A(n34), .Y(n35) );
  INVXLTS U27 ( .A(n12), .Y(n36) );
  INVXLTS U28 ( .A(n12), .Y(n37) );
  INVXLTS U29 ( .A(n7), .Y(n38) );
  INVXLTS U30 ( .A(n7), .Y(n39) );
  INVXLTS U31 ( .A(n1610), .Y(n40) );
  INVXLTS U32 ( .A(n40), .Y(n41) );
  INVXLTS U33 ( .A(n1131), .Y(n42) );
  INVXLTS U34 ( .A(n42), .Y(n43) );
  INVXLTS U35 ( .A(n10), .Y(n44) );
  INVXLTS U36 ( .A(n10), .Y(n49) );
  INVXLTS U37 ( .A(n14), .Y(n51) );
  INVXLTS U38 ( .A(n5), .Y(n53) );
  INVXLTS U39 ( .A(n910), .Y(n55) );
  INVXLTS U40 ( .A(n55), .Y(n57) );
  INVX2TS U41 ( .A(n1517), .Y(n59) );
  INVXLTS U42 ( .A(n59), .Y(n61) );
  CLKBUFX2TS U43 ( .A(n1490), .Y(n63) );
  INVXLTS U44 ( .A(n6), .Y(n64) );
  INVXLTS U45 ( .A(n6), .Y(n65) );
  INVXLTS U46 ( .A(n16), .Y(n66) );
  INVXLTS U47 ( .A(n16), .Y(n67) );
  INVXLTS U48 ( .A(n1740), .Y(n68) );
  INVXLTS U49 ( .A(n68), .Y(n69) );
  INVXLTS U50 ( .A(n15), .Y(n70) );
  INVXLTS U51 ( .A(n15), .Y(n71) );
  INVXLTS U52 ( .A(n1134), .Y(n80) );
  INVXLTS U53 ( .A(n80), .Y(n81) );
  INVXLTS U54 ( .A(n9), .Y(n82) );
  INVXLTS U55 ( .A(n9), .Y(n83) );
  INVX1TS U56 ( .A(n11), .Y(n84) );
  INVXLTS U57 ( .A(n11), .Y(n85) );
  INVXLTS U58 ( .A(n1130), .Y(n86) );
  INVXLTS U59 ( .A(n86), .Y(n87) );
  INVXLTS U60 ( .A(n1569), .Y(n88) );
  INVXLTS U61 ( .A(n1569), .Y(n89) );
  INVXLTS U62 ( .A(n1730), .Y(n90) );
  INVXLTS U63 ( .A(n90), .Y(n91) );
  INVXLTS U64 ( .A(n95), .Y(n92) );
  INVXLTS U65 ( .A(n1680), .Y(n93) );
  INVXLTS U66 ( .A(n1680), .Y(n94) );
  INVXLTS U67 ( .A(n94), .Y(n95) );
  INVXLTS U68 ( .A(n94), .Y(n96) );
  INVXLTS U69 ( .A(n880), .Y(n97) );
  INVXLTS U70 ( .A(n97), .Y(n98) );
  INVXLTS U71 ( .A(n97), .Y(n99) );
  INVXLTS U72 ( .A(n813), .Y(n100) );
  INVXLTS U73 ( .A(n100), .Y(n101) );
  INVXLTS U74 ( .A(n100), .Y(n102) );
  CLKBUFX2TS U314 ( .A(n1714), .Y(n342) );
  CLKBUFX2TS U315 ( .A(n1712), .Y(n343) );
  CLKBUFX2TS U316 ( .A(n1693), .Y(n344) );
  CLKBUFX2TS U317 ( .A(n1694), .Y(n345) );
  CLKBUFX2TS U318 ( .A(n1713), .Y(n346) );
  CLKBUFX2TS U319 ( .A(n964), .Y(n349) );
  CLKBUFX2TS U320 ( .A(n1742), .Y(n350) );
  INVX2TS U321 ( .A(n801), .Y(n351) );
  INVX2TS U322 ( .A(n802), .Y(n352) );
  CLKBUFX2TS U323 ( .A(n1515), .Y(n353) );
  CLKBUFX2TS U324 ( .A(n1533), .Y(n354) );
  CLKBUFX2TS U325 ( .A(n1533), .Y(n355) );
  CLKBUFX2TS U326 ( .A(n1411), .Y(n356) );
  CLKBUFX2TS U327 ( .A(n1764), .Y(n357) );
  CLKBUFX2TS U328 ( .A(n1743), .Y(n358) );
  CLKBUFX2TS U329 ( .A(n1754), .Y(n359) );
  CLKBUFX2TS U330 ( .A(n1732), .Y(n360) );
  CLKBUFX2TS U331 ( .A(n1702), .Y(n361) );
  CLKBUFX2TS U332 ( .A(n1415), .Y(n362) );
  OR2X2TS U333 ( .A(n92), .B(n805), .Y(n1609) );
  INVX2TS U334 ( .A(n1609), .Y(n363) );
  INVX2TS U335 ( .A(n1609), .Y(n364) );
  AND2X2TS U336 ( .A(n383), .B(n96), .Y(n1601) );
  INVX2TS U337 ( .A(n1601), .Y(n365) );
  INVX2TS U338 ( .A(n1601), .Y(n366) );
  CLKBUFX2TS U339 ( .A(n1505), .Y(n367) );
  CLKBUFX2TS U340 ( .A(n1505), .Y(n368) );
  NAND2X1TS U341 ( .A(n1528), .B(n1527), .Y(n1519) );
  INVX2TS U342 ( .A(n1519), .Y(n369) );
  INVX2TS U343 ( .A(n1519), .Y(n370) );
  INVX2TS U344 ( .A(n755), .Y(n371) );
  INVX2TS U345 ( .A(n963), .Y(n372) );
  NAND2X1TS U346 ( .A(n1487), .B(n1488), .Y(n373) );
  NAND2X1TS U347 ( .A(n1487), .B(n1488), .Y(n374) );
  CLKBUFX2TS U348 ( .A(n1755), .Y(n375) );
  CLKBUFX2TS U349 ( .A(n1765), .Y(n376) );
  CLKBUFX2TS U350 ( .A(n1733), .Y(n377) );
  AO21X1TS U351 ( .A0(n53), .A1(n961), .B0(n1572), .Y(n1490) );
  INVX2TS U352 ( .A(n1460), .Y(n378) );
  CLKBUFX2TS U353 ( .A(n1456), .Y(n379) );
  NOR3BX1TS U354 ( .AN(n64), .B(n1456), .C(n96), .Y(n1568) );
  AND3X2TS U355 ( .A(n1566), .B(n1131), .C(n1565), .Y(n1556) );
  INVX2TS U356 ( .A(n1556), .Y(n380) );
  INVX2TS U357 ( .A(n1556), .Y(n381) );
  INVX2TS U358 ( .A(n805), .Y(n382) );
  INVX2TS U359 ( .A(n1604), .Y(n383) );
  INVX2TS U360 ( .A(n1604), .Y(n384) );
  AND2X2TS U361 ( .A(n1514), .B(n811), .Y(n1503) );
  INVX2TS U362 ( .A(n1503), .Y(n385) );
  INVX2TS U363 ( .A(n1503), .Y(n386) );
  CLKBUFX2TS U364 ( .A(n1517), .Y(n387) );
  OAI211X1TS U365 ( .A0(n910), .A1(n1501), .B0(n2502), .C0(n1529), .Y(n1517)
         );
  NAND3X1TS U366 ( .A(n1190), .B(n37), .C(n2206), .Y(n1412) );
  INVX2TS U367 ( .A(n1412), .Y(n388) );
  INVX2TS U368 ( .A(n1412), .Y(n389) );
  INVX2TS U369 ( .A(n1412), .Y(n390) );
  AND2X2TS U370 ( .A(n770), .B(n101), .Y(n1413) );
  INVX2TS U371 ( .A(n1413), .Y(n391) );
  INVX2TS U372 ( .A(n1413), .Y(n392) );
  INVX2TS U373 ( .A(n1413), .Y(n393) );
  NOR2X1TS U374 ( .A(n961), .B(n1), .Y(n1572) );
  CLKAND2X2TS U375 ( .A(n1531), .B(n84), .Y(n1299) );
  AO21XLTS U376 ( .A0(n98), .A1(n1530), .B0(n1528), .Y(n1529) );
  NOR2X1TS U377 ( .A(n59), .B(n2487), .Y(n1527) );
  CLKBUFX2TS U378 ( .A(n2209), .Y(n2207) );
  CLKBUFX2TS U379 ( .A(n522), .Y(n520) );
  CLKBUFX2TS U380 ( .A(n520), .Y(n519) );
  CLKBUFX2TS U381 ( .A(n2209), .Y(n2206) );
  INVXLTS U382 ( .A(n568), .Y(n560) );
  INVXLTS U383 ( .A(n568), .Y(n559) );
  CLKBUFX2TS U384 ( .A(n2210), .Y(n2205) );
  OAI21X1TS U385 ( .A0(n2489), .A1(n1725), .B0(n1139), .Y(n1709) );
  NOR3XLTS U386 ( .A(n2265), .B(n32), .C(n1122), .Y(n1231) );
  NAND3XLTS U387 ( .A(n33), .B(n812), .C(n1513), .Y(n1229) );
  CLKINVX2TS U388 ( .A(n1008), .Y(n1007) );
  CLKBUFX2TS U389 ( .A(n570), .Y(n567) );
  NOR2X1TS U390 ( .A(n44), .B(n1466), .Y(n1605) );
  NAND2XLTS U391 ( .A(n1568), .B(n1490), .Y(n1134) );
  NAND3X1TS U392 ( .A(n1463), .B(n1025), .C(n372), .Y(n1466) );
  NOR3X1TS U393 ( .A(n1336), .B(n761), .C(n1123), .Y(n1303) );
  NOR3XLTS U394 ( .A(n748), .B(n568), .C(n1132), .Y(n1376) );
  XOR2X1TS U395 ( .A(n964), .B(n1729), .Y(n1463) );
  NAND2XLTS U396 ( .A(n85), .B(n1568), .Y(n1598) );
  NAND3XLTS U397 ( .A(n65), .B(n1025), .C(n63), .Y(n1190) );
  NAND3XLTS U398 ( .A(n85), .B(n813), .C(n1499), .Y(n1192) );
  NAND3X1TS U399 ( .A(n36), .B(n1134), .C(n2208), .Y(n1191) );
  NAND3BXLTS U400 ( .AN(n85), .B(n102), .C(n1499), .Y(n1193) );
  NAND2XLTS U401 ( .A(n1565), .B(n42), .Y(n1373) );
  CLKBUFX2TS U402 ( .A(n617), .Y(n614) );
  OAI21X1TS U403 ( .A0(n965), .A1(n1700), .B0(n1515), .Y(n1602) );
  NAND2XLTS U404 ( .A(n378), .B(n964), .Y(n1569) );
  OR4XLTS U405 ( .A(n1700), .B(n88), .C(n975), .D(n965), .Y(n1606) );
  NOR2XLTS U406 ( .A(n63), .B(n95), .Y(n1488) );
  NAND3XLTS U407 ( .A(n963), .B(n1025), .C(n1463), .Y(n1153) );
  NOR2XLTS U408 ( .A(n743), .B(n975), .Y(n1472) );
  XOR2XLTS U409 ( .A(n1572), .B(n55), .Y(n1531) );
  OAI31XLTS U410 ( .A0(n349), .A1(n1478), .A2(n378), .B0(n1691), .Y(n1690) );
  NOR3XLTS U411 ( .A(n1299), .B(n59), .C(n1130), .Y(n1267) );
  NAND2XLTS U412 ( .A(n84), .B(n1544), .Y(n1553) );
  NAND2XLTS U413 ( .A(n1527), .B(n97), .Y(n1264) );
  AND2XLTS U414 ( .A(n1544), .B(n63), .Y(n1336) );
  NAND2XLTS U415 ( .A(n1336), .B(n803), .Y(n1543) );
  AOI21XLTS U416 ( .A0(n85), .A1(n803), .B0(n1416), .Y(n1502) );
  OAI211XLTS U417 ( .A0(n1530), .A1(n1553), .B0(n1555), .C0(n1128), .Y(n1341)
         );
  AND3X2TS U418 ( .A(n43), .B(n2506), .C(n1567), .Y(n394) );
  XNOR2XLTS U419 ( .A(n1463), .B(n379), .Y(n1154) );
  NOR2XLTS U420 ( .A(n966), .B(n1476), .Y(n1700) );
  OAI21X1TS U421 ( .A0(n1464), .A1(n372), .B0(n1466), .Y(n1155) );
  NOR2XLTS U422 ( .A(n379), .B(n961), .Y(n1464) );
  NAND2XLTS U423 ( .A(n1476), .B(n966), .Y(n1610) );
  NAND2XLTS U424 ( .A(n1691), .B(n353), .Y(n1459) );
  NAND2XLTS U425 ( .A(n1477), .B(n966), .Y(n1474) );
  NAND2X1TS U426 ( .A(n101), .B(n53), .Y(n1680) );
  NOR2X1TS U427 ( .A(n1516), .B(n102), .Y(n1127) );
  NAND2X1TS U428 ( .A(n55), .B(n4), .Y(n1128) );
  AOI22XLTS U429 ( .A0(n985), .A1(n2475), .B0(n2273), .B1(n1918), .Y(n1294) );
  AOI22XLTS U430 ( .A0(n984), .A1(n2477), .B0(n2273), .B1(n1919), .Y(n1295) );
  AOI22XLTS U431 ( .A0(n984), .A1(n2479), .B0(n2274), .B1(n1920), .Y(n1296) );
  AOI22XLTS U432 ( .A0(n984), .A1(n2481), .B0(n2274), .B1(n1921), .Y(n1297) );
  AOI22XLTS U433 ( .A0(n984), .A1(n2483), .B0(n2274), .B1(n1922), .Y(n1298) );
  AOI22XLTS U434 ( .A0(n993), .A1(n2461), .B0(n2271), .B1(n1911), .Y(n1287) );
  AOI22XLTS U435 ( .A0(n993), .A1(n2463), .B0(n2272), .B1(n1912), .Y(n1288) );
  AOI22XLTS U436 ( .A0(n992), .A1(n2465), .B0(n2272), .B1(n1913), .Y(n1289) );
  AOI22XLTS U437 ( .A0(n991), .A1(n2467), .B0(n2272), .B1(n1914), .Y(n1290) );
  AOI22XLTS U438 ( .A0(n985), .A1(n2469), .B0(n2272), .B1(n1915), .Y(n1291) );
  AOI22XLTS U439 ( .A0(n985), .A1(n2471), .B0(n2273), .B1(n1916), .Y(n1292) );
  AOI22XLTS U440 ( .A0(n990), .A1(n2423), .B0(n2275), .B1(n738), .Y(n1268) );
  AOI22XLTS U441 ( .A0(n369), .A1(n2281), .B0(n1007), .B1(n681), .Y(n1520) );
  AOI22XLTS U442 ( .A0(n369), .A1(n2283), .B0(n1007), .B1(n680), .Y(n1521) );
  AOI22XLTS U443 ( .A0(n369), .A1(n2285), .B0(n1007), .B1(n679), .Y(n1522) );
  AOI22XLTS U444 ( .A0(n369), .A1(n2287), .B0(n1006), .B1(n678), .Y(n1523) );
  AOI22XLTS U445 ( .A0(n370), .A1(n2289), .B0(n1006), .B1(n677), .Y(n1524) );
  AOI22XLTS U446 ( .A0(n370), .A1(n2291), .B0(n1006), .B1(n676), .Y(n1525) );
  AOI22XLTS U447 ( .A0(n370), .A1(n2293), .B0(n1006), .B1(n675), .Y(n1526) );
  AOI22XLTS U448 ( .A0(n1023), .A1(n2423), .B0(n2265), .B1(n1893), .Y(n1232)
         );
  AOI22XLTS U449 ( .A0(n1018), .A1(n2483), .B0(n2265), .B1(n1891), .Y(n1262)
         );
  XNOR2X1TS U450 ( .A(n1570), .B(n1571), .Y(n1544) );
  OAI2BB1XLTS U451 ( .A0N(n372), .A1N(n1572), .B0(n1573), .Y(n1570) );
  OAI21XLTS U452 ( .A0(n1572), .A1(n1465), .B0(n347), .Y(n1573) );
  NOR2X1TS U453 ( .A(memRead_WEST), .B(memWrite_WEST), .Y(n1456) );
  OAI222XLTS U454 ( .A0(memWrite_SOUTH), .A1(n38), .B0(memWrite_EAST), .B1(
        n1602), .C0(memWrite_WEST), .C1(n31), .Y(n1462) );
  OAI222XLTS U455 ( .A0(memWrite_EAST), .A1(n29), .B0(n1727), .B1(n1728), .C0(
        memWrite_WEST), .C1(n65), .Y(n1140) );
  OA22XLTS U456 ( .A0(n965), .A1(memWrite_NORTH), .B0(n41), .B1(memWrite_SOUTH), .Y(n1727) );
  NOR3XLTS U457 ( .A(n975), .B(n99), .C(n1569), .Y(n1542) );
  OAI21XLTS U458 ( .A0(n1458), .A1(n771), .B0(n976), .Y(n1457) );
  AOI21XLTS U459 ( .A0(memRead_NORTH), .A1(n1460), .B0(memRead_SOUTH), .Y(
        n1458) );
  OAI22XLTS U460 ( .A0(n809), .A1(n976), .B0(n1471), .B1(n1024), .Y(n1470) );
  NAND3XLTS U461 ( .A(n5), .B(n353), .C(n89), .Y(n1501) );
  NOR2X1TS U462 ( .A(n26), .B(n740), .Y(n1773) );
  NOR2X1TS U463 ( .A(n938), .B(n3), .Y(n1762) );
  NOR2X1TS U464 ( .A(n348), .B(n2), .Y(n1763) );
  AOI211X1TS U465 ( .A0(\prevRequesterPort_B[0] ), .A1(n51), .B0(n460), .C0(
        n2493), .Y(n1730) );
  OAI21XLTS U466 ( .A0(n1472), .A1(n1473), .B0(n976), .Y(n1469) );
  AOI21XLTS U467 ( .A0(memRead_NORTH), .A1(n1474), .B0(memRead_SOUTH), .Y(
        n1473) );
  NOR2X1TS U468 ( .A(n51), .B(\prevRequesterPort_B[0] ), .Y(n1774) );
  OAI21X1TS U469 ( .A0(n880), .A1(n1), .B0(n1128), .Y(n1125) );
  XOR2X1TS U470 ( .A(n57), .B(n4), .Y(n1148) );
  NAND2X1TS U471 ( .A(n755), .B(n27), .Y(n1131) );
  NOR2X1TS U472 ( .A(n4), .B(n27), .Y(n1516) );
  NOR3X1TS U473 ( .A(n27), .B(n57), .C(n1148), .Y(n1477) );
  INVX2TS U474 ( .A(n2502), .Y(n2489) );
  INVX2TS U475 ( .A(n2506), .Y(n2485) );
  INVX2TS U476 ( .A(n2498), .Y(n2487) );
  INVX2TS U477 ( .A(n2504), .Y(n2486) );
  INVX2TS U478 ( .A(n2498), .Y(n2488) );
  INVX2TS U479 ( .A(n2494), .Y(n2493) );
  INVX2TS U480 ( .A(n2497), .Y(n2490) );
  INVX2TS U481 ( .A(n2496), .Y(n2491) );
  INVX2TS U482 ( .A(n2495), .Y(n2492) );
  CLKBUFX2TS U483 ( .A(n2504), .Y(n2494) );
  CLKBUFX2TS U484 ( .A(n2499), .Y(n2498) );
  CLKBUFX2TS U485 ( .A(n2504), .Y(n2495) );
  CLKBUFX2TS U486 ( .A(n2494), .Y(n2496) );
  CLKBUFX2TS U487 ( .A(n2506), .Y(n2497) );
  CLKBUFX2TS U488 ( .A(n2240), .Y(n2236) );
  CLKBUFX2TS U489 ( .A(n2240), .Y(n2235) );
  CLKBUFX2TS U490 ( .A(n2241), .Y(n2233) );
  CLKBUFX2TS U491 ( .A(n2241), .Y(n2234) );
  CLKBUFX2TS U492 ( .A(n2503), .Y(n2499) );
  CLKBUFX2TS U493 ( .A(n2503), .Y(n2500) );
  CLKBUFX2TS U494 ( .A(n2503), .Y(n2501) );
  CLKBUFX2TS U495 ( .A(n2503), .Y(n2502) );
  CLKBUFX2TS U496 ( .A(n2499), .Y(n2504) );
  CLKBUFX2TS U497 ( .A(n2244), .Y(n2237) );
  CLKBUFX2TS U498 ( .A(n2244), .Y(n2238) );
  CLKBUFX2TS U499 ( .A(n2243), .Y(n2240) );
  CLKBUFX2TS U500 ( .A(n2243), .Y(n2241) );
  CLKBUFX2TS U501 ( .A(n2244), .Y(n2239) );
  CLKBUFX2TS U502 ( .A(n472), .Y(n461) );
  CLKBUFX2TS U503 ( .A(n472), .Y(n462) );
  CLKBUFX2TS U504 ( .A(n471), .Y(n463) );
  CLKBUFX2TS U505 ( .A(n471), .Y(n464) );
  CLKBUFX2TS U506 ( .A(n470), .Y(n465) );
  CLKBUFX2TS U507 ( .A(n470), .Y(n466) );
  CLKBUFX2TS U508 ( .A(n469), .Y(n467) );
  CLKBUFX2TS U509 ( .A(n469), .Y(n468) );
  CLKBUFX2TS U510 ( .A(n2242), .Y(n2232) );
  CLKBUFX2TS U511 ( .A(n2243), .Y(n2242) );
  CLKBUFX2TS U512 ( .A(n544), .Y(n535) );
  CLKBUFX2TS U513 ( .A(n541), .Y(n536) );
  CLKBUFX2TS U514 ( .A(n541), .Y(n537) );
  CLKBUFX2TS U515 ( .A(n540), .Y(n538) );
  CLKBUFX2TS U516 ( .A(n540), .Y(n539) );
  CLKBUFX2TS U517 ( .A(n2505), .Y(n2503) );
  CLKBUFX2TS U518 ( .A(n2506), .Y(n2505) );
  INVX2TS U519 ( .A(n585), .Y(n582) );
  CLKBUFX2TS U520 ( .A(n1229), .Y(n1030) );
  CLKBUFX2TS U521 ( .A(n684), .Y(n683) );
  CLKBUFX2TS U522 ( .A(n684), .Y(n649) );
  CLKBUFX2TS U523 ( .A(n685), .Y(n648) );
  CLKBUFX2TS U524 ( .A(n685), .Y(n647) );
  CLKBUFX2TS U525 ( .A(n685), .Y(n646) );
  CLKBUFX2TS U526 ( .A(n686), .Y(n645) );
  CLKBUFX2TS U527 ( .A(n686), .Y(n644) );
  CLKBUFX2TS U528 ( .A(n1041), .Y(n1037) );
  CLKBUFX2TS U529 ( .A(n1038), .Y(n1036) );
  CLKBUFX2TS U530 ( .A(n1038), .Y(n1035) );
  CLKBUFX2TS U531 ( .A(n1039), .Y(n1034) );
  CLKBUFX2TS U532 ( .A(n1039), .Y(n1033) );
  CLKBUFX2TS U533 ( .A(n1040), .Y(n1032) );
  CLKBUFX2TS U534 ( .A(n1040), .Y(n1031) );
  CLKBUFX2TS U535 ( .A(n545), .Y(n544) );
  CLKBUFX2TS U536 ( .A(n545), .Y(n543) );
  CLKBUFX2TS U537 ( .A(n545), .Y(n542) );
  CLKBUFX2TS U538 ( .A(n1580), .Y(n472) );
  CLKBUFX2TS U539 ( .A(n1580), .Y(n471) );
  CLKBUFX2TS U540 ( .A(n546), .Y(n541) );
  CLKBUFX2TS U541 ( .A(n546), .Y(n540) );
  CLKBUFX2TS U542 ( .A(n1580), .Y(n470) );
  CLKBUFX2TS U543 ( .A(n472), .Y(n469) );
  CLKBUFX2TS U544 ( .A(n800), .Y(n2244) );
  CLKBUFX2TS U545 ( .A(n800), .Y(n2243) );
  CLKBUFX2TS U546 ( .A(n2138), .Y(n2128) );
  CLKBUFX2TS U547 ( .A(n2137), .Y(n2129) );
  CLKBUFX2TS U548 ( .A(n2137), .Y(n2130) );
  CLKBUFX2TS U549 ( .A(n2136), .Y(n2131) );
  CLKBUFX2TS U550 ( .A(n2136), .Y(n2132) );
  CLKBUFX2TS U551 ( .A(n2255), .Y(n2245) );
  CLKBUFX2TS U552 ( .A(n2254), .Y(n2246) );
  CLKBUFX2TS U553 ( .A(n2254), .Y(n2247) );
  CLKBUFX2TS U554 ( .A(n2253), .Y(n2248) );
  CLKBUFX2TS U555 ( .A(n2253), .Y(n2249) );
  CLKBUFX2TS U556 ( .A(n2135), .Y(n2133) );
  CLKBUFX2TS U557 ( .A(n2252), .Y(n2250) );
  CLKBUFX2TS U558 ( .A(n481), .Y(n473) );
  CLKBUFX2TS U559 ( .A(n483), .Y(n474) );
  CLKBUFX2TS U560 ( .A(n483), .Y(n475) );
  CLKBUFX2TS U561 ( .A(n482), .Y(n476) );
  CLKBUFX2TS U562 ( .A(n481), .Y(n477) );
  CLKBUFX2TS U563 ( .A(n480), .Y(n478) );
  CLKBUFX2TS U564 ( .A(n480), .Y(n479) );
  CLKBUFX2TS U565 ( .A(n2135), .Y(n2134) );
  CLKBUFX2TS U566 ( .A(n2252), .Y(n2251) );
  INVX2TS U567 ( .A(n2210), .Y(n2202) );
  INVX2TS U568 ( .A(n2208), .Y(n2203) );
  INVX2TS U569 ( .A(n2207), .Y(n2204) );
  INVX2TS U570 ( .A(reset), .Y(n2506) );
  CLKBUFX2TS U571 ( .A(n555), .Y(n551) );
  CLKBUFX2TS U572 ( .A(n555), .Y(n550) );
  CLKBUFX2TS U573 ( .A(n557), .Y(n549) );
  CLKBUFX2TS U574 ( .A(n556), .Y(n548) );
  CLKBUFX2TS U575 ( .A(n556), .Y(n547) );
  CLKBUFX2TS U576 ( .A(n507), .Y(n497) );
  CLKBUFX2TS U577 ( .A(n1577), .Y(n498) );
  CLKBUFX2TS U578 ( .A(n506), .Y(n499) );
  CLKBUFX2TS U579 ( .A(n505), .Y(n500) );
  CLKBUFX2TS U580 ( .A(n505), .Y(n501) );
  CLKBUFX2TS U581 ( .A(n504), .Y(n502) );
  CLKBUFX2TS U582 ( .A(n504), .Y(n503) );
  CLKBUFX2TS U583 ( .A(n554), .Y(n553) );
  CLKBUFX2TS U584 ( .A(n554), .Y(n552) );
  CLKBUFX2TS U585 ( .A(n532), .Y(n528) );
  CLKBUFX2TS U586 ( .A(n532), .Y(n527) );
  CLKBUFX2TS U587 ( .A(n531), .Y(n526) );
  CLKBUFX2TS U588 ( .A(n533), .Y(n525) );
  CLKBUFX2TS U589 ( .A(n533), .Y(n524) );
  CLKBUFX2TS U590 ( .A(n533), .Y(n523) );
  CLKBUFX2TS U591 ( .A(n531), .Y(n530) );
  CLKBUFX2TS U592 ( .A(n531), .Y(n529) );
  INVX2TS U593 ( .A(n521), .Y(n509) );
  INVX2TS U594 ( .A(n520), .Y(n511) );
  INVX2TS U595 ( .A(n520), .Y(n512) );
  INVX2TS U596 ( .A(n520), .Y(n513) );
  INVX2TS U597 ( .A(n519), .Y(n514) );
  INVX2TS U598 ( .A(n519), .Y(n515) );
  INVX2TS U599 ( .A(n519), .Y(n516) );
  INVX2TS U600 ( .A(n519), .Y(n517) );
  INVX2TS U601 ( .A(n522), .Y(n518) );
  INVX2TS U602 ( .A(n521), .Y(n510) );
  INVX2TS U603 ( .A(n2206), .Y(n2195) );
  INVX2TS U604 ( .A(n2206), .Y(n2196) );
  INVX2TS U605 ( .A(n2206), .Y(n2197) );
  INVX2TS U606 ( .A(n2207), .Y(n2198) );
  INVX2TS U607 ( .A(n2207), .Y(n2199) );
  INVX2TS U608 ( .A(n2210), .Y(n2200) );
  INVX2TS U609 ( .A(n395), .Y(n2201) );
  INVX2TS U610 ( .A(n2190), .Y(n2152) );
  INVX2TS U611 ( .A(n2166), .Y(n2151) );
  INVX2TS U612 ( .A(n2162), .Y(n2154) );
  INVX2TS U613 ( .A(n2166), .Y(n2153) );
  INVX2TS U614 ( .A(n2187), .Y(n2155) );
  INVX2TS U615 ( .A(n2165), .Y(n2156) );
  INVX2TS U616 ( .A(n2164), .Y(n2157) );
  INVX2TS U617 ( .A(n2163), .Y(n2158) );
  INVX2TS U618 ( .A(n2162), .Y(n2159) );
  INVX2TS U619 ( .A(n2164), .Y(n2150) );
  INVX2TS U620 ( .A(n2161), .Y(n2160) );
  NOR2X1TS U621 ( .A(n2266), .B(n2486), .Y(n1513) );
  CLKBUFX2TS U622 ( .A(n592), .Y(n585) );
  CLKBUFX2TS U623 ( .A(n1229), .Y(n1039) );
  CLKBUFX2TS U624 ( .A(n1229), .Y(n1040) );
  CLKBUFX2TS U625 ( .A(n687), .Y(n686) );
  CLKBUFX2TS U626 ( .A(n1041), .Y(n1038) );
  CLKBUFX2TS U627 ( .A(n688), .Y(n684) );
  CLKBUFX2TS U628 ( .A(n688), .Y(n685) );
  CLKBUFX2TS U629 ( .A(n1784), .Y(n1739) );
  CLKBUFX2TS U630 ( .A(n1781), .Y(n1752) );
  CLKBUFX2TS U631 ( .A(n1783), .Y(n1767) );
  CLKBUFX2TS U632 ( .A(n1026), .Y(n1023) );
  CLKBUFX2TS U633 ( .A(n1026), .Y(n1022) );
  CLKBUFX2TS U634 ( .A(n1028), .Y(n1021) );
  CLKBUFX2TS U635 ( .A(n1028), .Y(n1020) );
  CLKBUFX2TS U636 ( .A(n1029), .Y(n1019) );
  CLKBUFX2TS U637 ( .A(n1029), .Y(n1018) );
  CLKBUFX2TS U638 ( .A(n1782), .Y(n1778) );
  CLKBUFX2TS U639 ( .A(n1783), .Y(n1777) );
  CLKBUFX2TS U640 ( .A(n630), .Y(n620) );
  CLKBUFX2TS U641 ( .A(n631), .Y(n621) );
  CLKBUFX2TS U642 ( .A(n627), .Y(n622) );
  CLKBUFX2TS U643 ( .A(n627), .Y(n623) );
  CLKBUFX2TS U644 ( .A(n1782), .Y(n1779) );
  CLKBUFX2TS U645 ( .A(n1781), .Y(n1780) );
  CLKBUFX2TS U646 ( .A(n626), .Y(n624) );
  CLKBUFX2TS U647 ( .A(n626), .Y(n625) );
  INVX2TS U648 ( .A(n584), .Y(n583) );
  CLKBUFX2TS U649 ( .A(n591), .Y(n589) );
  CLKBUFX2TS U650 ( .A(n592), .Y(n588) );
  CLKBUFX2TS U651 ( .A(n592), .Y(n587) );
  CLKBUFX2TS U652 ( .A(n592), .Y(n586) );
  CLKBUFX2TS U653 ( .A(n591), .Y(n590) );
  CLKBUFX2TS U654 ( .A(n1228), .Y(n1042) );
  CLKBUFX2TS U655 ( .A(n2121), .Y(n2120) );
  CLKBUFX2TS U656 ( .A(n2121), .Y(n2119) );
  CLKBUFX2TS U657 ( .A(n2122), .Y(n2118) );
  CLKBUFX2TS U658 ( .A(n2122), .Y(n2117) );
  CLKBUFX2TS U659 ( .A(n2123), .Y(n2116) );
  CLKBUFX2TS U660 ( .A(n1053), .Y(n1049) );
  CLKBUFX2TS U661 ( .A(n1050), .Y(n1048) );
  CLKBUFX2TS U662 ( .A(n1050), .Y(n1047) );
  CLKBUFX2TS U663 ( .A(n1051), .Y(n1046) );
  CLKBUFX2TS U664 ( .A(n1051), .Y(n1045) );
  CLKBUFX2TS U665 ( .A(n1052), .Y(n1044) );
  CLKBUFX2TS U666 ( .A(n1052), .Y(n1043) );
  CLKBUFX2TS U667 ( .A(n601), .Y(n600) );
  CLKBUFX2TS U668 ( .A(n601), .Y(n599) );
  CLKBUFX2TS U669 ( .A(n602), .Y(n598) );
  CLKBUFX2TS U670 ( .A(n602), .Y(n597) );
  CLKBUFX2TS U671 ( .A(n602), .Y(n596) );
  CLKBUFX2TS U672 ( .A(n603), .Y(n595) );
  CLKBUFX2TS U673 ( .A(n603), .Y(n594) );
  CLKBUFX2TS U674 ( .A(n831), .Y(n816) );
  CLKBUFX2TS U675 ( .A(n831), .Y(n815) );
  CLKBUFX2TS U676 ( .A(n935), .Y(n807) );
  CLKBUFX2TS U677 ( .A(n935), .Y(n806) );
  CLKBUFX2TS U678 ( .A(n955), .Y(n804) );
  CLKBUFX2TS U679 ( .A(n2109), .Y(n2108) );
  CLKBUFX2TS U680 ( .A(n2109), .Y(n2107) );
  CLKBUFX2TS U681 ( .A(n2110), .Y(n2087) );
  CLKBUFX2TS U682 ( .A(n2110), .Y(n2085) );
  CLKBUFX2TS U683 ( .A(n2111), .Y(n1966) );
  CLKBUFX2TS U684 ( .A(n639), .Y(n638) );
  CLKBUFX2TS U685 ( .A(n639), .Y(n637) );
  CLKBUFX2TS U686 ( .A(n640), .Y(n636) );
  CLKBUFX2TS U687 ( .A(n640), .Y(n635) );
  CLKBUFX2TS U688 ( .A(n642), .Y(n634) );
  CLKBUFX2TS U689 ( .A(n641), .Y(n633) );
  CLKBUFX2TS U690 ( .A(n641), .Y(n632) );
  CLKBUFX2TS U691 ( .A(n522), .Y(n521) );
  INVX2TS U692 ( .A(n1678), .Y(n800) );
  CLKBUFX2TS U693 ( .A(n2138), .Y(n2137) );
  CLKBUFX2TS U694 ( .A(n2255), .Y(n2254) );
  CLKBUFX2TS U695 ( .A(n1579), .Y(n483) );
  CLKBUFX2TS U696 ( .A(n1579), .Y(n482) );
  CLKBUFX2TS U697 ( .A(n2139), .Y(n2136) );
  CLKBUFX2TS U698 ( .A(n2256), .Y(n2253) );
  CLKBUFX2TS U699 ( .A(n2256), .Y(n2252) );
  CLKBUFX2TS U700 ( .A(n2139), .Y(n2135) );
  CLKBUFX2TS U701 ( .A(n484), .Y(n481) );
  CLKBUFX2TS U702 ( .A(n484), .Y(n480) );
  CLKBUFX2TS U703 ( .A(n1421), .Y(n545) );
  CLKBUFX2TS U704 ( .A(n2262), .Y(n2257) );
  CLKBUFX2TS U705 ( .A(n2262), .Y(n2258) );
  CLKBUFX2TS U706 ( .A(n2261), .Y(n2259) );
  CLKBUFX2TS U707 ( .A(n1421), .Y(n546) );
  CLKBUFX2TS U708 ( .A(n2261), .Y(n2260) );
  CLKBUFX2TS U709 ( .A(n2146), .Y(n2145) );
  CLKBUFX2TS U710 ( .A(n2146), .Y(n2144) );
  CLKBUFX2TS U711 ( .A(n2147), .Y(n2143) );
  CLKBUFX2TS U712 ( .A(n2147), .Y(n2142) );
  CLKBUFX2TS U713 ( .A(n2149), .Y(n2141) );
  CLKBUFX2TS U714 ( .A(n2149), .Y(n2140) );
  CLKBUFX2TS U715 ( .A(n2209), .Y(n2208) );
  NAND2BX1TS U716 ( .AN(n413), .B(n2501), .Y(n1765) );
  INVX2TS U717 ( .A(n2205), .Y(n2192) );
  CLKBUFX2TS U718 ( .A(n557), .Y(n556) );
  CLKBUFX2TS U719 ( .A(n1422), .Y(n533) );
  CLKBUFX2TS U720 ( .A(n507), .Y(n506) );
  CLKBUFX2TS U721 ( .A(n558), .Y(n554) );
  CLKBUFX2TS U722 ( .A(n534), .Y(n531) );
  CLKBUFX2TS U723 ( .A(n558), .Y(n555) );
  CLKBUFX2TS U724 ( .A(n534), .Y(n532) );
  CLKBUFX2TS U725 ( .A(n508), .Y(n505) );
  CLKBUFX2TS U726 ( .A(n508), .Y(n504) );
  CLKBUFX2TS U727 ( .A(n495), .Y(n486) );
  CLKBUFX2TS U728 ( .A(n495), .Y(n485) );
  CLKBUFX2TS U729 ( .A(n493), .Y(n492) );
  CLKBUFX2TS U730 ( .A(n493), .Y(n491) );
  CLKBUFX2TS U731 ( .A(n494), .Y(n490) );
  CLKBUFX2TS U732 ( .A(n494), .Y(n489) );
  CLKBUFX2TS U733 ( .A(n495), .Y(n488) );
  CLKBUFX2TS U734 ( .A(n494), .Y(n487) );
  CLKBUFX2TS U735 ( .A(n2188), .Y(n2166) );
  CLKBUFX2TS U736 ( .A(n2187), .Y(n2165) );
  CLKBUFX2TS U737 ( .A(n2187), .Y(n2164) );
  CLKBUFX2TS U738 ( .A(n2187), .Y(n2163) );
  CLKBUFX2TS U739 ( .A(n2188), .Y(n2162) );
  CLKBUFX2TS U740 ( .A(n2188), .Y(n2161) );
  INVX2TS U741 ( .A(n2205), .Y(n2193) );
  INVX2TS U742 ( .A(n2205), .Y(n2194) );
  CLKBUFX2TS U743 ( .A(n2186), .Y(n2168) );
  CLKBUFX2TS U744 ( .A(n2186), .Y(n2167) );
  CLKBUFX2TS U745 ( .A(n2186), .Y(n2169) );
  CLKBUFX2TS U746 ( .A(n2183), .Y(n2179) );
  CLKBUFX2TS U747 ( .A(n2183), .Y(n2181) );
  CLKBUFX2TS U748 ( .A(n2183), .Y(n2180) );
  CLKBUFX2TS U749 ( .A(n2184), .Y(n2178) );
  CLKBUFX2TS U750 ( .A(n2184), .Y(n2177) );
  CLKBUFX2TS U751 ( .A(n2184), .Y(n2176) );
  CLKBUFX2TS U752 ( .A(n2184), .Y(n2175) );
  CLKBUFX2TS U753 ( .A(n2186), .Y(n2170) );
  CLKBUFX2TS U754 ( .A(n2185), .Y(n2171) );
  CLKBUFX2TS U755 ( .A(n2185), .Y(n2172) );
  CLKBUFX2TS U756 ( .A(n2185), .Y(n2173) );
  CLKBUFX2TS U757 ( .A(n2185), .Y(n2174) );
  CLKBUFX2TS U758 ( .A(n2183), .Y(n2182) );
  NOR2X1TS U759 ( .A(n2485), .B(n568), .Y(n1565) );
  NOR2X1TS U760 ( .A(n761), .B(n2487), .Y(n1541) );
  NOR2X1TS U761 ( .A(n619), .B(n2487), .Y(n1554) );
  NOR2X1TS U762 ( .A(n1196), .B(n2486), .Y(n1499) );
  CLKBUFX2TS U763 ( .A(n593), .Y(n584) );
  CLKBUFX2TS U764 ( .A(n1374), .Y(n593) );
  CLKBUFX2TS U765 ( .A(n2266), .Y(n2265) );
  CLKBUFX2TS U766 ( .A(n1231), .Y(n1026) );
  CLKBUFX2TS U767 ( .A(n1231), .Y(n1027) );
  CLKBUFX2TS U768 ( .A(n1231), .Y(n1028) );
  CLKBUFX2TS U769 ( .A(n1231), .Y(n1029) );
  CLKBUFX2TS U770 ( .A(n1195), .Y(n1783) );
  CLKBUFX2TS U771 ( .A(n1195), .Y(n1784) );
  CLKBUFX2TS U772 ( .A(n630), .Y(n629) );
  CLKBUFX2TS U773 ( .A(n630), .Y(n628) );
  CLKBUFX2TS U774 ( .A(n967), .Y(n955) );
  CLKBUFX2TS U775 ( .A(n967), .Y(n956) );
  CLKBUFX2TS U776 ( .A(n2114), .Y(n2111) );
  CLKBUFX2TS U777 ( .A(n2126), .Y(n2123) );
  CLKBUFX2TS U778 ( .A(n2114), .Y(n2112) );
  CLKBUFX2TS U779 ( .A(n2126), .Y(n2124) );
  CLKBUFX2TS U780 ( .A(n1228), .Y(n1051) );
  CLKBUFX2TS U781 ( .A(n1228), .Y(n1052) );
  CLKBUFX2TS U782 ( .A(n967), .Y(n959) );
  CLKBUFX2TS U783 ( .A(n2114), .Y(n2113) );
  CLKBUFX2TS U784 ( .A(n2126), .Y(n2125) );
  CLKBUFX2TS U785 ( .A(n604), .Y(n603) );
  CLKBUFX2TS U786 ( .A(n642), .Y(n641) );
  CLKBUFX2TS U787 ( .A(n1965), .Y(n1781) );
  CLKBUFX2TS U788 ( .A(n631), .Y(n626) );
  CLKBUFX2TS U789 ( .A(n1965), .Y(n1782) );
  CLKBUFX2TS U790 ( .A(n631), .Y(n627) );
  CLKBUFX2TS U791 ( .A(n968), .Y(n831) );
  CLKBUFX2TS U792 ( .A(n968), .Y(n935) );
  CLKBUFX2TS U793 ( .A(n2115), .Y(n2109) );
  CLKBUFX2TS U794 ( .A(n2127), .Y(n2121) );
  CLKBUFX2TS U795 ( .A(n2115), .Y(n2110) );
  CLKBUFX2TS U796 ( .A(n2127), .Y(n2122) );
  CLKBUFX2TS U797 ( .A(n1053), .Y(n1050) );
  CLKBUFX2TS U798 ( .A(n605), .Y(n601) );
  CLKBUFX2TS U799 ( .A(n605), .Y(n602) );
  CLKBUFX2TS U800 ( .A(n643), .Y(n639) );
  CLKBUFX2TS U801 ( .A(n643), .Y(n640) );
  CLKBUFX2TS U802 ( .A(n1337), .Y(n687) );
  CLKBUFX2TS U803 ( .A(n1303), .Y(n768) );
  CLKBUFX2TS U804 ( .A(n769), .Y(n767) );
  CLKBUFX2TS U805 ( .A(n769), .Y(n766) );
  CLKBUFX2TS U806 ( .A(n769), .Y(n765) );
  CLKBUFX2TS U807 ( .A(n772), .Y(n764) );
  CLKBUFX2TS U808 ( .A(n772), .Y(n763) );
  CLKBUFX2TS U809 ( .A(n799), .Y(n762) );
  CLKBUFX2TS U810 ( .A(n579), .Y(n578) );
  CLKBUFX2TS U811 ( .A(n579), .Y(n577) );
  CLKBUFX2TS U812 ( .A(n580), .Y(n576) );
  CLKBUFX2TS U813 ( .A(n580), .Y(n575) );
  CLKBUFX2TS U814 ( .A(n580), .Y(n574) );
  CLKBUFX2TS U815 ( .A(n581), .Y(n573) );
  CLKBUFX2TS U816 ( .A(n581), .Y(n572) );
  CLKBUFX2TS U817 ( .A(n2277), .Y(n2268) );
  CLKBUFX2TS U818 ( .A(n2277), .Y(n2269) );
  CLKBUFX2TS U819 ( .A(n2277), .Y(n2270) );
  CLKBUFX2TS U820 ( .A(n2276), .Y(n2271) );
  CLKBUFX2TS U821 ( .A(n2276), .Y(n2272) );
  CLKBUFX2TS U822 ( .A(n2275), .Y(n2273) );
  CLKBUFX2TS U823 ( .A(n1229), .Y(n1041) );
  CLKBUFX2TS U824 ( .A(n1337), .Y(n688) );
  INVX2TS U825 ( .A(n972), .Y(n969) );
  INVX2TS U826 ( .A(n1017), .Y(n1006) );
  CLKBUFX2TS U827 ( .A(n1374), .Y(n591) );
  CLKBUFX2TS U828 ( .A(n1374), .Y(n592) );
  CLKBUFX2TS U829 ( .A(n2275), .Y(n2274) );
  INVX2TS U830 ( .A(n618), .Y(n610) );
  INVX2TS U831 ( .A(n618), .Y(n609) );
  INVX2TS U832 ( .A(n614), .Y(n608) );
  INVX2TS U833 ( .A(n618), .Y(n607) );
  INVX2TS U834 ( .A(n616), .Y(n606) );
  NOR2BX1TS U835 ( .AN(n1677), .B(n83), .Y(n1713) );
  NOR3X1TS U836 ( .A(n2192), .B(n89), .C(n39), .Y(n1678) );
  NOR3BX1TS U837 ( .AN(n1677), .B(n2204), .C(n521), .Y(n1580) );
  NOR3X1TS U838 ( .A(n2192), .B(n1678), .C(n38), .Y(n1421) );
  OAI21X1TS U839 ( .A0(n1708), .A1(n809), .B0(n2189), .Y(n1702) );
  INVX2TS U840 ( .A(n1709), .Y(n805) );
  NOR2X1TS U841 ( .A(n49), .B(n39), .Y(n1693) );
  CLKBUFX2TS U842 ( .A(n1156), .Y(n2146) );
  CLKBUFX2TS U843 ( .A(n1156), .Y(n2147) );
  CLKBUFX2TS U844 ( .A(n1156), .Y(n2148) );
  CLKBUFX2TS U845 ( .A(n1156), .Y(n2149) );
  CLKBUFX2TS U846 ( .A(n2266), .Y(n2264) );
  CLKBUFX2TS U847 ( .A(n2266), .Y(n2263) );
  CLKBUFX2TS U848 ( .A(n2267), .Y(n2262) );
  CLKBUFX2TS U849 ( .A(n2267), .Y(n2261) );
  CLKBUFX2TS U850 ( .A(n1158), .Y(n2138) );
  CLKBUFX2TS U851 ( .A(n798), .Y(n2255) );
  INVX2TS U852 ( .A(n1574), .Y(n522) );
  CLKBUFX2TS U853 ( .A(n1579), .Y(n484) );
  CLKBUFX2TS U854 ( .A(n1158), .Y(n2139) );
  CLKBUFX2TS U855 ( .A(n798), .Y(n2256) );
  CLKBUFX2TS U856 ( .A(n1377), .Y(n1263) );
  CLKBUFX2TS U857 ( .A(n1489), .Y(n1137) );
  CLKBUFX2TS U858 ( .A(n1489), .Y(n1136) );
  CLKBUFX2TS U859 ( .A(n1500), .Y(n1057) );
  CLKBUFX2TS U860 ( .A(n1500), .Y(n1056) );
  CLKBUFX2TS U861 ( .A(n1607), .Y(n1055) );
  CLKBUFX2TS U862 ( .A(n1681), .Y(n1054) );
  INVX2TS U863 ( .A(n752), .Y(n689) );
  INVX2TS U864 ( .A(n752), .Y(n690) );
  INVX2TS U865 ( .A(n753), .Y(n741) );
  INVX2TS U866 ( .A(n753), .Y(n744) );
  INVX2TS U867 ( .A(n752), .Y(n745) );
  INVX2TS U868 ( .A(n753), .Y(n746) );
  INVX2TS U869 ( .A(n753), .Y(n747) );
  INVX2TS U870 ( .A(n760), .Y(n749) );
  INVX2TS U871 ( .A(n567), .Y(n563) );
  INVX2TS U872 ( .A(n567), .Y(n562) );
  INVX2TS U873 ( .A(n567), .Y(n561) );
  INVX2TS U874 ( .A(n752), .Y(n750) );
  INVX2TS U875 ( .A(n760), .Y(n751) );
  NOR2X1TS U876 ( .A(n418), .B(n2488), .Y(n1755) );
  CLKBUFX2TS U877 ( .A(n395), .Y(n2210) );
  CLKBUFX2TS U878 ( .A(n1578), .Y(n495) );
  CLKBUFX2TS U879 ( .A(n496), .Y(n493) );
  CLKBUFX2TS U880 ( .A(n496), .Y(n494) );
  CLKBUFX2TS U881 ( .A(n395), .Y(n2209) );
  CLKBUFX2TS U882 ( .A(n1420), .Y(n557) );
  CLKBUFX2TS U883 ( .A(n1577), .Y(n507) );
  CLKBUFX2TS U884 ( .A(n416), .Y(n408) );
  CLKBUFX2TS U885 ( .A(n416), .Y(n409) );
  CLKBUFX2TS U886 ( .A(n415), .Y(n410) );
  CLKBUFX2TS U887 ( .A(n415), .Y(n411) );
  CLKBUFX2TS U888 ( .A(n414), .Y(n412) );
  CLKBUFX2TS U889 ( .A(n425), .Y(n422) );
  CLKBUFX2TS U890 ( .A(n425), .Y(n421) );
  CLKBUFX2TS U891 ( .A(n427), .Y(n420) );
  CLKBUFX2TS U892 ( .A(n427), .Y(n419) );
  CLKBUFX2TS U893 ( .A(n443), .Y(n441) );
  CLKBUFX2TS U894 ( .A(n444), .Y(n440) );
  CLKBUFX2TS U895 ( .A(n444), .Y(n439) );
  CLKBUFX2TS U896 ( .A(n1422), .Y(n534) );
  CLKBUFX2TS U897 ( .A(n1420), .Y(n558) );
  CLKBUFX2TS U898 ( .A(n1577), .Y(n508) );
  INVX2TS U899 ( .A(n1122), .Y(n811) );
  CLKBUFX2TS U900 ( .A(n424), .Y(n423) );
  CLKBUFX2TS U901 ( .A(n443), .Y(n442) );
  CLKBUFX2TS U902 ( .A(n414), .Y(n413) );
  INVX2TS U903 ( .A(n1605), .Y(n802) );
  INVX2TS U904 ( .A(n1612), .Y(n801) );
  NOR2X1TS U905 ( .A(n2231), .B(n2486), .Y(n1754) );
  NOR2X1TS U906 ( .A(n449), .B(n2487), .Y(n1732) );
  NOR2X1TS U907 ( .A(n447), .B(n2488), .Y(n1743) );
  CLKBUFX2TS U908 ( .A(n2218), .Y(n2212) );
  CLKBUFX2TS U909 ( .A(n2218), .Y(n2213) );
  CLKBUFX2TS U910 ( .A(n2217), .Y(n2214) );
  CLKBUFX2TS U911 ( .A(n2217), .Y(n2215) );
  CLKBUFX2TS U912 ( .A(n2228), .Y(n2226) );
  CLKBUFX2TS U913 ( .A(n2228), .Y(n2225) );
  CLKBUFX2TS U914 ( .A(n2229), .Y(n2223) );
  CLKBUFX2TS U915 ( .A(n2229), .Y(n2224) );
  CLKBUFX2TS U916 ( .A(n2230), .Y(n2222) );
  CLKBUFX2TS U917 ( .A(n2230), .Y(n2221) );
  CLKBUFX2TS U918 ( .A(n2217), .Y(n2216) );
  CLKBUFX2TS U919 ( .A(n2189), .Y(n2187) );
  CLKBUFX2TS U920 ( .A(n2191), .Y(n2184) );
  CLKBUFX2TS U921 ( .A(n2190), .Y(n2186) );
  CLKBUFX2TS U922 ( .A(n2190), .Y(n2185) );
  CLKBUFX2TS U923 ( .A(n2191), .Y(n2183) );
  CLKBUFX2TS U924 ( .A(n2189), .Y(n2188) );
  INVX2TS U925 ( .A(n1465), .Y(n963) );
  NAND2X1TS U926 ( .A(n1565), .B(n748), .Y(n1374) );
  CLKBUFX2TS U927 ( .A(n570), .Y(n568) );
  INVX2TS U928 ( .A(n1463), .Y(n961) );
  CLKBUFX2TS U929 ( .A(n1300), .Y(n972) );
  NAND2X1TS U930 ( .A(n1554), .B(n755), .Y(n1337) );
  INVX2TS U931 ( .A(n1530), .Y(n803) );
  CLKBUFX2TS U932 ( .A(n1303), .Y(n769) );
  CLKBUFX2TS U933 ( .A(n1303), .Y(n772) );
  CLKBUFX2TS U934 ( .A(n1303), .Y(n799) );
  CLKBUFX2TS U935 ( .A(n1376), .Y(n579) );
  CLKBUFX2TS U936 ( .A(n1376), .Y(n580) );
  CLKBUFX2TS U937 ( .A(n1376), .Y(n581) );
  CLKBUFX2TS U938 ( .A(n2278), .Y(n2277) );
  CLKBUFX2TS U939 ( .A(n2278), .Y(n2276) );
  CLKBUFX2TS U940 ( .A(n2278), .Y(n2275) );
  CLKBUFX2TS U941 ( .A(n1193), .Y(n2114) );
  CLKBUFX2TS U942 ( .A(n1338), .Y(n642) );
  CLKBUFX2TS U943 ( .A(n1192), .Y(n2126) );
  CLKBUFX2TS U944 ( .A(n1301), .Y(n967) );
  CLKBUFX2TS U945 ( .A(n1373), .Y(n604) );
  CLKBUFX2TS U946 ( .A(n1340), .Y(n630) );
  CLKBUFX2TS U947 ( .A(n1503), .Y(n2266) );
  CLKBUFX2TS U948 ( .A(n991), .Y(n990) );
  CLKBUFX2TS U949 ( .A(n991), .Y(n989) );
  CLKBUFX2TS U950 ( .A(n992), .Y(n988) );
  CLKBUFX2TS U951 ( .A(n992), .Y(n987) );
  CLKBUFX2TS U952 ( .A(n993), .Y(n986) );
  CLKBUFX2TS U953 ( .A(n992), .Y(n985) );
  CLKBUFX2TS U954 ( .A(n993), .Y(n984) );
  CLKBUFX2TS U955 ( .A(n1193), .Y(n2115) );
  CLKBUFX2TS U956 ( .A(n1338), .Y(n643) );
  CLKBUFX2TS U957 ( .A(n1192), .Y(n2127) );
  CLKBUFX2TS U958 ( .A(n1301), .Y(n968) );
  CLKBUFX2TS U959 ( .A(n1195), .Y(n1965) );
  CLKBUFX2TS U960 ( .A(n1373), .Y(n605) );
  CLKBUFX2TS U961 ( .A(n1228), .Y(n1053) );
  CLKBUFX2TS U962 ( .A(n1340), .Y(n631) );
  INVX2TS U963 ( .A(n971), .Y(n970) );
  CLKBUFX2TS U964 ( .A(n982), .Y(n981) );
  CLKBUFX2TS U965 ( .A(n982), .Y(n980) );
  CLKBUFX2TS U966 ( .A(n982), .Y(n979) );
  CLKBUFX2TS U967 ( .A(n982), .Y(n978) );
  CLKBUFX2TS U968 ( .A(n983), .Y(n974) );
  CLKBUFX2TS U969 ( .A(n1300), .Y(n973) );
  CLKBUFX2TS U970 ( .A(n1016), .Y(n1014) );
  CLKBUFX2TS U971 ( .A(n1016), .Y(n1013) );
  CLKBUFX2TS U972 ( .A(n1016), .Y(n1012) );
  CLKBUFX2TS U973 ( .A(n1017), .Y(n1011) );
  CLKBUFX2TS U974 ( .A(n1264), .Y(n1010) );
  CLKBUFX2TS U975 ( .A(n1264), .Y(n1009) );
  CLKBUFX2TS U976 ( .A(n1016), .Y(n1015) );
  CLKBUFX2TS U977 ( .A(n1003), .Y(n994) );
  CLKBUFX2TS U978 ( .A(n999), .Y(n998) );
  CLKBUFX2TS U979 ( .A(n999), .Y(n997) );
  CLKBUFX2TS U980 ( .A(n1000), .Y(n996) );
  CLKBUFX2TS U981 ( .A(n1000), .Y(n995) );
  INVX2TS U982 ( .A(n614), .Y(n613) );
  INVX2TS U983 ( .A(n614), .Y(n612) );
  INVX2TS U984 ( .A(n614), .Y(n611) );
  NOR2X1TS U985 ( .A(n82), .B(n1606), .Y(n1714) );
  NOR2X1TS U986 ( .A(n82), .B(n64), .Y(n1612) );
  NAND3X1TS U987 ( .A(n1190), .B(n1191), .C(n2208), .Y(n1156) );
  NAND2X1TS U988 ( .A(n1725), .B(n2208), .Y(n1574) );
  NOR2X1TS U989 ( .A(n64), .B(n2202), .Y(n1579) );
  NOR2X1TS U990 ( .A(n388), .B(n2486), .Y(n1487) );
  NOR2X1TS U991 ( .A(n1708), .B(n81), .Y(n1158) );
  CLKBUFX2TS U992 ( .A(n760), .Y(n752) );
  CLKBUFX2TS U993 ( .A(n760), .Y(n753) );
  NAND2X1TS U994 ( .A(n2495), .B(n1191), .Y(n1708) );
  CLKBUFX2TS U995 ( .A(n1411), .Y(n397) );
  NOR2BX1TS U996 ( .AN(n1487), .B(n81), .Y(n1411) );
  NOR2X1TS U997 ( .A(n44), .B(n35), .Y(n1694) );
  NAND2X1TS U998 ( .A(n29), .B(n65), .Y(n1728) );
  NOR2X1TS U999 ( .A(n1728), .B(n965), .Y(n1677) );
  INVX2TS U1000 ( .A(n1604), .Y(n810) );
  NAND2X1TS U1001 ( .A(n1487), .B(n1488), .Y(n1409) );
  CLKBUFX2TS U1002 ( .A(n1681), .Y(n1377) );
  CLKBUFX2TS U1003 ( .A(n1681), .Y(n1489) );
  CLKBUFX2TS U1004 ( .A(n1681), .Y(n1500) );
  CLKBUFX2TS U1005 ( .A(n1607), .Y(n1599) );
  CLKBUFX2TS U1006 ( .A(n571), .Y(n569) );
  CLKBUFX2TS U1007 ( .A(n617), .Y(n615) );
  CLKBUFX2TS U1008 ( .A(n1503), .Y(n2267) );
  INVX2TS U1009 ( .A(n1191), .Y(n798) );
  CLKBUFX2TS U1010 ( .A(n617), .Y(n616) );
  INVX2TS U1011 ( .A(n571), .Y(n566) );
  INVX2TS U1012 ( .A(n394), .Y(n565) );
  INVX2TS U1013 ( .A(n394), .Y(n564) );
  NAND2X1TS U1014 ( .A(n2496), .B(n391), .Y(n1415) );
  NAND2X1TS U1015 ( .A(n812), .B(n2499), .Y(n1122) );
  NOR2X1TS U1016 ( .A(n1602), .B(n2203), .Y(n1422) );
  NOR2X1TS U1017 ( .A(n31), .B(n2192), .Y(n1420) );
  NOR2X1TS U1018 ( .A(n1606), .B(n2203), .Y(n1577) );
  INVX2TS U1019 ( .A(n396), .Y(n449) );
  CLKBUFX2TS U1020 ( .A(n415), .Y(n416) );
  CLKBUFX2TS U1021 ( .A(n447), .Y(n445) );
  CLKBUFX2TS U1022 ( .A(n447), .Y(n446) );
  CLKBUFX2TS U1023 ( .A(n417), .Y(n414) );
  CLKBUFX2TS U1024 ( .A(n417), .Y(n415) );
  CLKBUFX2TS U1025 ( .A(n427), .Y(n425) );
  CLKBUFX2TS U1026 ( .A(n448), .Y(n444) );
  CLKBUFX2TS U1027 ( .A(n427), .Y(n424) );
  CLKBUFX2TS U1028 ( .A(n448), .Y(n443) );
  CLKBUFX2TS U1029 ( .A(n426), .Y(n418) );
  CLKBUFX2TS U1030 ( .A(n1761), .Y(n426) );
  CLKBUFX2TS U1031 ( .A(n937), .Y(n2211) );
  CLKBUFX2TS U1032 ( .A(n404), .Y(n399) );
  CLKBUFX2TS U1033 ( .A(n407), .Y(n400) );
  CLKBUFX2TS U1034 ( .A(n404), .Y(n401) );
  CLKBUFX2TS U1035 ( .A(n403), .Y(n402) );
  INVX2TS U1036 ( .A(n1598), .Y(n808) );
  CLKBUFX2TS U1037 ( .A(n1578), .Y(n496) );
  INVX2TS U1038 ( .A(n1488), .Y(n809) );
  AND2X2TS U1039 ( .A(n93), .B(n2499), .Y(n395) );
  NOR2X1TS U1040 ( .A(n436), .B(n2488), .Y(n1742) );
  CLKBUFX2TS U1041 ( .A(n1139), .Y(n2189) );
  CLKBUFX2TS U1042 ( .A(n1139), .Y(n2190) );
  CLKBUFX2TS U1043 ( .A(n1139), .Y(n2191) );
  CLKBUFX2TS U1044 ( .A(n2220), .Y(n2219) );
  CLKBUFX2TS U1045 ( .A(n2220), .Y(n2218) );
  CLKBUFX2TS U1046 ( .A(n2231), .Y(n2229) );
  CLKBUFX2TS U1047 ( .A(n2227), .Y(n2230) );
  CLKBUFX2TS U1048 ( .A(n2220), .Y(n2217) );
  CLKBUFX2TS U1049 ( .A(n2231), .Y(n2227) );
  CLKBUFX2TS U1050 ( .A(n2231), .Y(n2228) );
  CLKBUFX2TS U1051 ( .A(n432), .Y(n430) );
  CLKBUFX2TS U1052 ( .A(n433), .Y(n429) );
  CLKBUFX2TS U1053 ( .A(n433), .Y(n428) );
  INVX2TS U1054 ( .A(n460), .Y(n450) );
  INVX2TS U1055 ( .A(n460), .Y(n455) );
  INVX2TS U1056 ( .A(n458), .Y(n454) );
  INVX2TS U1057 ( .A(n396), .Y(n452) );
  INVX2TS U1058 ( .A(n458), .Y(n453) );
  INVX2TS U1059 ( .A(n396), .Y(n451) );
  INVX2TS U1060 ( .A(n459), .Y(n456) );
  CLKBUFX2TS U1061 ( .A(n432), .Y(n431) );
  INVX2TS U1062 ( .A(n458), .Y(n457) );
  INVX2TS U1063 ( .A(n2314), .Y(n2313) );
  INVX2TS U1064 ( .A(n2317), .Y(n2316) );
  INVX2TS U1065 ( .A(n1123), .Y(n756) );
  NOR3BX1TS U1066 ( .AN(n1513), .B(n32), .C(n1127), .Y(n1505) );
  XNOR2X1TS U1067 ( .A(n966), .B(n975), .Y(n1729) );
  NAND3BX1TS U1068 ( .AN(n1553), .B(n371), .C(n1554), .Y(n1338) );
  NAND3X1TS U1069 ( .A(n1336), .B(n757), .C(n1541), .Y(n1301) );
  INVX2TS U1070 ( .A(n1515), .Y(n975) );
  CLKBUFX2TS U1071 ( .A(n983), .Y(n971) );
  CLKBUFX2TS U1072 ( .A(n1300), .Y(n983) );
  CLKBUFX2TS U1073 ( .A(n1017), .Y(n1008) );
  CLKBUFX2TS U1074 ( .A(n1264), .Y(n1017) );
  AND3X2TS U1075 ( .A(n1553), .B(n1128), .C(n1554), .Y(n1340) );
  INVX2TS U1076 ( .A(n1566), .Y(n748) );
  NAND2X1TS U1077 ( .A(n1513), .B(n1127), .Y(n1228) );
  CLKBUFX2TS U1078 ( .A(n1267), .Y(n991) );
  CLKBUFX2TS U1079 ( .A(n1267), .Y(n992) );
  CLKBUFX2TS U1080 ( .A(n1267), .Y(n993) );
  CLKBUFX2TS U1081 ( .A(n1004), .Y(n1001) );
  CLKBUFX2TS U1082 ( .A(n1004), .Y(n1002) );
  CLKBUFX2TS U1083 ( .A(n1004), .Y(n1003) );
  CLKBUFX2TS U1084 ( .A(n1005), .Y(n999) );
  CLKBUFX2TS U1085 ( .A(n1005), .Y(n1000) );
  CLKBUFX2TS U1086 ( .A(n394), .Y(n570) );
  CLKBUFX2TS U1087 ( .A(n619), .Y(n618) );
  CLKBUFX2TS U1088 ( .A(n1196), .Y(n1607) );
  CLKBUFX2TS U1089 ( .A(n59), .Y(n2278) );
  CLKBUFX2TS U1090 ( .A(n1300), .Y(n982) );
  CLKBUFX2TS U1091 ( .A(n1264), .Y(n1016) );
  NOR2BX1TS U1092 ( .AN(n1677), .B(n349), .Y(n1725) );
  OAI31X1TS U1093 ( .A0(n38), .A1(n88), .A2(n96), .B0(n2502), .Y(n1604) );
  CLKBUFX2TS U1094 ( .A(n394), .Y(n571) );
  NOR2X1TS U1095 ( .A(n83), .B(n1610), .Y(n1712) );
  INVX2TS U1096 ( .A(n41), .Y(n965) );
  NOR2BX1TS U1097 ( .AN(n1141), .B(n1142), .Y(n3644) );
  NOR2BX1TS U1098 ( .AN(n1144), .B(n1142), .Y(n3642) );
  INVX2TS U1099 ( .A(n1155), .Y(n960) );
  CLKBUFX2TS U1100 ( .A(n619), .Y(n617) );
  CLKBUFX2TS U1101 ( .A(n1196), .Y(n1681) );
  CLKBUFX2TS U1102 ( .A(n761), .Y(n760) );
  NOR2X1TS U1103 ( .A(n1143), .B(n1142), .Y(n3643) );
  NOR3BX1TS U1104 ( .AN(n1153), .B(n1154), .C(n1155), .Y(n1138) );
  NAND2X1TS U1105 ( .A(n95), .B(n2500), .Y(n1139) );
  NOR2X1TS U1106 ( .A(n1610), .B(n2204), .Y(n1578) );
  INVX2TS U1107 ( .A(n1154), .Y(n962) );
  CLKBUFX2TS U1108 ( .A(n437), .Y(n436) );
  CLKBUFX2TS U1109 ( .A(n407), .Y(n404) );
  CLKBUFX2TS U1110 ( .A(n407), .Y(n403) );
  CLKBUFX2TS U1111 ( .A(n1749), .Y(n447) );
  CLKBUFX2TS U1112 ( .A(n405), .Y(n398) );
  CLKBUFX2TS U1113 ( .A(n406), .Y(n405) );
  CLKBUFX2TS U1114 ( .A(n1749), .Y(n448) );
  CLKBUFX2TS U1115 ( .A(n1775), .Y(n417) );
  CLKBUFX2TS U1116 ( .A(n1761), .Y(n427) );
  INVX2TS U1117 ( .A(n1455), .Y(n770) );
  NAND2X1TS U1118 ( .A(n757), .B(n2500), .Y(n1123) );
  CLKBUFX2TS U1119 ( .A(n460), .Y(n458) );
  NAND2X1TS U1120 ( .A(n371), .B(n2494), .Y(n1129) );
  CLKBUFX2TS U1121 ( .A(n458), .Y(n459) );
  CLKBUFX2TS U1122 ( .A(n437), .Y(n434) );
  CLKBUFX2TS U1123 ( .A(n437), .Y(n435) );
  CLKBUFX2TS U1124 ( .A(n438), .Y(n432) );
  CLKBUFX2TS U1125 ( .A(n438), .Y(n433) );
  CLKBUFX2TS U1126 ( .A(n2315), .Y(n2314) );
  CLKBUFX2TS U1127 ( .A(n2318), .Y(n2317) );
  CLKBUFX2TS U1128 ( .A(n937), .Y(n2220) );
  CLKBUFX2TS U1129 ( .A(n936), .Y(n2231) );
  INVX2TS U1130 ( .A(n2280), .Y(n2279) );
  INVX2TS U1131 ( .A(n2282), .Y(n2281) );
  INVX2TS U1132 ( .A(n2284), .Y(n2283) );
  INVX2TS U1133 ( .A(n2286), .Y(n2285) );
  INVX2TS U1134 ( .A(n2288), .Y(n2287) );
  INVX2TS U1135 ( .A(n2290), .Y(n2289) );
  INVX2TS U1136 ( .A(n2292), .Y(n2291) );
  INVX2TS U1137 ( .A(n2294), .Y(n2293) );
  INVX2TS U1138 ( .A(n2296), .Y(n2295) );
  INVX2TS U1139 ( .A(n2299), .Y(n2298) );
  INVX2TS U1140 ( .A(n2302), .Y(n2301) );
  INVX2TS U1141 ( .A(n2306), .Y(n2304) );
  INVX2TS U1142 ( .A(n2308), .Y(n2307) );
  INVX2TS U1143 ( .A(n2312), .Y(n2310) );
  INVX2TS U1144 ( .A(n1459), .Y(n771) );
  INVX2TS U1145 ( .A(n2326), .Y(n2325) );
  INVX2TS U1146 ( .A(n2330), .Y(n2328) );
  INVX2TS U1147 ( .A(n2332), .Y(n2331) );
  INVX2TS U1148 ( .A(n2336), .Y(n2334) );
  INVX2TS U1149 ( .A(n2338), .Y(n2337) );
  INVX2TS U1150 ( .A(n2341), .Y(n2340) );
  INVX2TS U1151 ( .A(n2344), .Y(n2343) );
  INVX2TS U1152 ( .A(n2348), .Y(n2346) );
  INVX2TS U1153 ( .A(n2350), .Y(n2349) );
  INVX2TS U1154 ( .A(n2353), .Y(n2352) );
  INVX2TS U1155 ( .A(n2357), .Y(n2355) );
  INVX2TS U1156 ( .A(n2359), .Y(n2358) );
  INVX2TS U1157 ( .A(n2362), .Y(n2361) );
  INVX2TS U1158 ( .A(n2366), .Y(n2364) );
  INVX2TS U1159 ( .A(n2368), .Y(n2367) );
  INVX2TS U1160 ( .A(n2372), .Y(n2370) );
  INVX2TS U1161 ( .A(n2374), .Y(n2373) );
  INVX2TS U1162 ( .A(n2377), .Y(n2376) );
  INVX2TS U1163 ( .A(n2380), .Y(n2379) );
  INVX2TS U1164 ( .A(n2384), .Y(n2382) );
  INVX2TS U1165 ( .A(n2387), .Y(n2385) );
  INVX2TS U1166 ( .A(n2390), .Y(n2388) );
  INVX2TS U1167 ( .A(n2392), .Y(n2391) );
  INVX2TS U1168 ( .A(n2395), .Y(n2394) );
  INVX2TS U1169 ( .A(n2399), .Y(n2397) );
  INVX2TS U1170 ( .A(n2401), .Y(n2400) );
  INVX2TS U1171 ( .A(n2404), .Y(n2403) );
  INVX2TS U1172 ( .A(n2407), .Y(n2406) );
  INVX2TS U1173 ( .A(n2410), .Y(n2409) );
  INVX2TS U1174 ( .A(n2413), .Y(n2412) );
  INVX2TS U1175 ( .A(n2416), .Y(n2415) );
  INVX2TS U1176 ( .A(n2419), .Y(n2418) );
  INVX2TS U1177 ( .A(n1132), .Y(n754) );
  INVX2TS U1178 ( .A(n1127), .Y(n812) );
  INVX2TS U1179 ( .A(n1128), .Y(n755) );
  NOR3BX1TS U1180 ( .AN(n1541), .B(n1125), .C(n1336), .Y(n1533) );
  NAND2X1TS U1181 ( .A(n1541), .B(n1125), .Y(n1300) );
  INVX2TS U1182 ( .A(n1460), .Y(n966) );
  NAND2X1TS U1183 ( .A(n33), .B(n1544), .Y(n1566) );
  AOI32X1TS U1184 ( .A0(n353), .A1(n347), .A2(n88), .B0(n32), .B1(n803), .Y(
        n1514) );
  AND3X2TS U1185 ( .A(n1501), .B(n2501), .C(n1502), .Y(n1196) );
  NOR2X1TS U1186 ( .A(n4), .B(n1299), .Y(n1528) );
  INVX2TS U1187 ( .A(n1476), .Y(n964) );
  CLKBUFX2TS U1188 ( .A(n1265), .Y(n1004) );
  INVX2TS U1189 ( .A(n1304), .Y(n761) );
  NAND4BX1TS U1190 ( .AN(n1542), .B(n1543), .C(n757), .D(n2504), .Y(n1304) );
  CLKBUFX2TS U1191 ( .A(n1265), .Y(n1005) );
  AOI22X1TS U1192 ( .A0(n1542), .A1(n55), .B0(n748), .B1(n803), .Y(n1567) );
  INVX2TS U1193 ( .A(n1341), .Y(n619) );
  OAI2BB1X1TS U1194 ( .A0N(n2502), .A1N(n1501), .B0(n87), .Y(n1555) );
  NAND3X1TS U1195 ( .A(n1145), .B(n2505), .C(n1146), .Y(n1142) );
  XOR2X1TS U1196 ( .A(n1147), .B(n101), .Y(n1146) );
  NAND3BX1TS U1197 ( .AN(n1143), .B(n1141), .C(n1144), .Y(n1145) );
  NAND2X1TS U1198 ( .A(n1148), .B(n1149), .Y(n1147) );
  AOI21X1TS U1199 ( .A0(n1477), .A1(n1478), .B0(n80), .Y(n1471) );
  NOR2X1TS U1200 ( .A(n1456), .B(n92), .Y(n1478) );
  INVX2TS U1201 ( .A(n1456), .Y(n1025) );
  XOR2X1TS U1202 ( .A(n1150), .B(n1151), .Y(n1143) );
  XOR2X1TS U1203 ( .A(n347), .B(n960), .Y(n1150) );
  XOR2X1TS U1204 ( .A(n1149), .B(n1148), .Y(n1144) );
  OAI211X1TS U1205 ( .A0(n743), .A1(n1476), .B0(n1471), .C0(n36), .Y(n1475) );
  OAI221XLTS U1206 ( .A0(n365), .A1(n673), .B0(n810), .B1(n824), .C0(n1692), 
        .Y(n3202) );
  AOI222XLTS U1207 ( .A0(n1605), .A1(requesterAddressIn_WEST[0]), .B0(
        requesterAddressIn_SOUTH[0]), .B1(n1693), .C0(
        requesterAddressIn_EAST[0]), .C1(n1694), .Y(n1692) );
  OAI221XLTS U1208 ( .A0(n365), .A1(n672), .B0(n383), .B1(n823), .C0(n1695), 
        .Y(n3201) );
  AOI222XLTS U1209 ( .A0(n1605), .A1(requesterAddressIn_WEST[1]), .B0(
        requesterAddressIn_SOUTH[1]), .B1(n1693), .C0(
        requesterAddressIn_EAST[1]), .C1(n1694), .Y(n1695) );
  OAI221XLTS U1210 ( .A0(n366), .A1(n671), .B0(n384), .B1(n822), .C0(n1696), 
        .Y(n3200) );
  AOI222XLTS U1211 ( .A0(n1605), .A1(requesterAddressIn_WEST[2]), .B0(
        requesterAddressIn_SOUTH[2]), .B1(n1693), .C0(
        requesterAddressIn_EAST[2]), .C1(n1694), .Y(n1696) );
  OAI221XLTS U1212 ( .A0(n366), .A1(n670), .B0(n810), .B1(n821), .C0(n1697), 
        .Y(n3199) );
  AOI222XLTS U1213 ( .A0(n352), .A1(requesterAddressIn_WEST[3]), .B0(
        requesterAddressIn_SOUTH[3]), .B1(n344), .C0(
        requesterAddressIn_EAST[3]), .C1(n345), .Y(n1697) );
  OAI221XLTS U1214 ( .A0(n366), .A1(n669), .B0(n383), .B1(n820), .C0(n1698), 
        .Y(n3198) );
  AOI222XLTS U1215 ( .A0(n352), .A1(requesterAddressIn_WEST[4]), .B0(
        requesterAddressIn_SOUTH[4]), .B1(n344), .C0(
        requesterAddressIn_EAST[4]), .C1(n345), .Y(n1698) );
  OAI221XLTS U1216 ( .A0(n366), .A1(n668), .B0(n384), .B1(n819), .C0(n1699), 
        .Y(n3197) );
  AOI222XLTS U1217 ( .A0(n352), .A1(requesterAddressIn_WEST[5]), .B0(
        requesterAddressIn_SOUTH[5]), .B1(n344), .C0(
        requesterAddressIn_EAST[5]), .C1(n345), .Y(n1699) );
  OAI22X1TS U1218 ( .A0(n2211), .A1(n1089), .B0(n417), .B1(n1121), .Y(N10083)
         );
  OAI22X1TS U1219 ( .A0(n2211), .A1(n1088), .B0(n1775), .B1(n1120), .Y(N10084)
         );
  OAI22X1TS U1220 ( .A0(n2219), .A1(n1087), .B0(n1775), .B1(n1119), .Y(N10085)
         );
  OAI22X1TS U1221 ( .A0(n2219), .A1(n1086), .B0(n408), .B1(n1118), .Y(N10086)
         );
  OAI22X1TS U1222 ( .A0(n937), .A1(n1085), .B0(n408), .B1(n1117), .Y(N10087)
         );
  OAI22X1TS U1223 ( .A0(n937), .A1(n1084), .B0(n408), .B1(n1116), .Y(N10088)
         );
  OAI22X1TS U1224 ( .A0(n2219), .A1(n1083), .B0(n408), .B1(n1115), .Y(N10089)
         );
  OAI22X1TS U1225 ( .A0(n2217), .A1(n1082), .B0(n409), .B1(n1114), .Y(N10090)
         );
  OAI22X1TS U1226 ( .A0(n2220), .A1(n1081), .B0(n409), .B1(n1113), .Y(N10091)
         );
  OAI22X1TS U1227 ( .A0(n2218), .A1(n1080), .B0(n409), .B1(n1112), .Y(N10092)
         );
  OAI22X1TS U1228 ( .A0(n2212), .A1(n1079), .B0(n409), .B1(n1111), .Y(N10093)
         );
  OAI22X1TS U1229 ( .A0(n2212), .A1(n1078), .B0(n415), .B1(n1110), .Y(N10094)
         );
  OAI22X1TS U1230 ( .A0(n2212), .A1(n1077), .B0(n414), .B1(n1109), .Y(N10095)
         );
  OAI22X1TS U1231 ( .A0(n2212), .A1(n1076), .B0(n1775), .B1(n1108), .Y(N10096)
         );
  OAI22X1TS U1232 ( .A0(n2213), .A1(n1075), .B0(n414), .B1(n1107), .Y(N10097)
         );
  OAI22X1TS U1233 ( .A0(n2213), .A1(n1074), .B0(n413), .B1(n1106), .Y(N10098)
         );
  OAI22X1TS U1234 ( .A0(n2213), .A1(n1073), .B0(n416), .B1(n1105), .Y(N10099)
         );
  OAI22X1TS U1235 ( .A0(n2213), .A1(n1072), .B0(n417), .B1(n1104), .Y(N10100)
         );
  OAI22X1TS U1236 ( .A0(n2216), .A1(n1071), .B0(n416), .B1(n1103), .Y(N10101)
         );
  OAI22X1TS U1237 ( .A0(n2216), .A1(n1070), .B0(n410), .B1(n1102), .Y(N10102)
         );
  OAI22X1TS U1238 ( .A0(n2219), .A1(n1069), .B0(n410), .B1(n1101), .Y(N10103)
         );
  OAI22X1TS U1239 ( .A0(n2218), .A1(n1068), .B0(n410), .B1(n1100), .Y(N10104)
         );
  OAI22X1TS U1240 ( .A0(n2214), .A1(n1067), .B0(n410), .B1(n1099), .Y(N10105)
         );
  OAI22X1TS U1241 ( .A0(n2214), .A1(n1066), .B0(n411), .B1(n1098), .Y(N10106)
         );
  OAI22X1TS U1242 ( .A0(n2214), .A1(n1065), .B0(n411), .B1(n1097), .Y(N10107)
         );
  OAI22X1TS U1243 ( .A0(n2214), .A1(n1064), .B0(n411), .B1(n1096), .Y(N10108)
         );
  OAI22X1TS U1244 ( .A0(n2215), .A1(n1063), .B0(n411), .B1(n1095), .Y(N10109)
         );
  OAI22X1TS U1245 ( .A0(n2215), .A1(n1062), .B0(n412), .B1(n1094), .Y(N10110)
         );
  OAI22X1TS U1246 ( .A0(n2215), .A1(n1061), .B0(n412), .B1(n1093), .Y(N10111)
         );
  OAI22X1TS U1247 ( .A0(n2215), .A1(n1060), .B0(n412), .B1(n1092), .Y(N10112)
         );
  OAI22X1TS U1248 ( .A0(n2216), .A1(n1059), .B0(n412), .B1(n1091), .Y(N10113)
         );
  OAI22X1TS U1249 ( .A0(n2216), .A1(n1058), .B0(n413), .B1(n1090), .Y(N10114)
         );
  OAI22X1TS U1250 ( .A0(n2228), .A1(n1089), .B0(n423), .B1(n1121), .Y(N10117)
         );
  OAI22X1TS U1251 ( .A0(n2228), .A1(n1088), .B0(n426), .B1(n1120), .Y(N10118)
         );
  OAI22X1TS U1252 ( .A0(n2229), .A1(n1087), .B0(n426), .B1(n1119), .Y(N10119)
         );
  OAI22X1TS U1253 ( .A0(n2230), .A1(n1086), .B0(n426), .B1(n1118), .Y(N10120)
         );
  OAI22X1TS U1254 ( .A0(n2227), .A1(n1085), .B0(n424), .B1(n1117), .Y(N10121)
         );
  OAI22X1TS U1255 ( .A0(n2227), .A1(n1084), .B0(n422), .B1(n1116), .Y(N10122)
         );
  OAI22X1TS U1256 ( .A0(n2227), .A1(n1083), .B0(n422), .B1(n1115), .Y(N10123)
         );
  OAI22X1TS U1257 ( .A0(n2226), .A1(n1082), .B0(n422), .B1(n1114), .Y(N10124)
         );
  OAI22X1TS U1258 ( .A0(n2226), .A1(n1081), .B0(n422), .B1(n1113), .Y(N10125)
         );
  OAI22X1TS U1259 ( .A0(n2226), .A1(n1080), .B0(n421), .B1(n1112), .Y(N10126)
         );
  OAI22X1TS U1260 ( .A0(n2226), .A1(n1079), .B0(n421), .B1(n1111), .Y(N10127)
         );
  OAI22X1TS U1261 ( .A0(n2225), .A1(n1078), .B0(n421), .B1(n1110), .Y(N10128)
         );
  OAI22X1TS U1262 ( .A0(n2225), .A1(n1077), .B0(n421), .B1(n1109), .Y(N10129)
         );
  OAI22X1TS U1263 ( .A0(n2225), .A1(n1076), .B0(n423), .B1(n1108), .Y(N10130)
         );
  OAI22X1TS U1264 ( .A0(n2225), .A1(n1075), .B0(n424), .B1(n1107), .Y(N10131)
         );
  OAI22X1TS U1265 ( .A0(n2224), .A1(n1074), .B0(n1761), .B1(n1106), .Y(N10132)
         );
  OAI22X1TS U1266 ( .A0(n2224), .A1(n1073), .B0(n423), .B1(n1105), .Y(N10133)
         );
  OAI22X1TS U1267 ( .A0(n2224), .A1(n1072), .B0(n425), .B1(n1104), .Y(N10134)
         );
  OAI22X1TS U1268 ( .A0(n2223), .A1(n1071), .B0(n1761), .B1(n1103), .Y(N10135)
         );
  OAI22X1TS U1269 ( .A0(n2223), .A1(n1070), .B0(n424), .B1(n1102), .Y(N10136)
         );
  OAI22X1TS U1270 ( .A0(n2223), .A1(n1069), .B0(n425), .B1(n1101), .Y(N10137)
         );
  OAI22X1TS U1271 ( .A0(n2223), .A1(n1068), .B0(n420), .B1(n1100), .Y(N10138)
         );
  OAI22X1TS U1272 ( .A0(n2222), .A1(n1067), .B0(n420), .B1(n1099), .Y(N10139)
         );
  OAI22X1TS U1273 ( .A0(n2222), .A1(n1066), .B0(n420), .B1(n1098), .Y(N10140)
         );
  OAI22X1TS U1274 ( .A0(n2224), .A1(n1065), .B0(n420), .B1(n1097), .Y(N10141)
         );
  OAI22X1TS U1275 ( .A0(n2222), .A1(n1064), .B0(n419), .B1(n1096), .Y(N10142)
         );
  OAI22X1TS U1276 ( .A0(n2222), .A1(n1063), .B0(n419), .B1(n1095), .Y(N10143)
         );
  OAI22X1TS U1277 ( .A0(n2221), .A1(n1062), .B0(n419), .B1(n1094), .Y(N10144)
         );
  OAI22X1TS U1278 ( .A0(n2221), .A1(n1061), .B0(n419), .B1(n1093), .Y(N10145)
         );
  OAI22X1TS U1279 ( .A0(n2221), .A1(n1060), .B0(n418), .B1(n1092), .Y(N10146)
         );
  OAI22X1TS U1280 ( .A0(n2221), .A1(n1059), .B0(n418), .B1(n1091), .Y(N10147)
         );
  OAI22X1TS U1281 ( .A0(n2230), .A1(n1058), .B0(n418), .B1(n1090), .Y(N10148)
         );
  OAI22X1TS U1282 ( .A0(n431), .A1(n1089), .B0(n442), .B1(n1121), .Y(N10151)
         );
  OAI22X1TS U1283 ( .A0(n431), .A1(n1088), .B0(n441), .B1(n1120), .Y(N10152)
         );
  OAI22X1TS U1284 ( .A0(n431), .A1(n1087), .B0(n441), .B1(n1119), .Y(N10153)
         );
  OAI22X1TS U1285 ( .A0(n430), .A1(n1086), .B0(n441), .B1(n1118), .Y(N10154)
         );
  OAI22X1TS U1286 ( .A0(n430), .A1(n1085), .B0(n441), .B1(n1117), .Y(N10155)
         );
  OAI22X1TS U1287 ( .A0(n430), .A1(n1084), .B0(n440), .B1(n1116), .Y(N10156)
         );
  OAI22X1TS U1288 ( .A0(n430), .A1(n1083), .B0(n440), .B1(n1115), .Y(N10157)
         );
  OAI22X1TS U1289 ( .A0(n429), .A1(n1082), .B0(n440), .B1(n1114), .Y(N10158)
         );
  OAI22X1TS U1290 ( .A0(n429), .A1(n1081), .B0(n440), .B1(n1113), .Y(N10159)
         );
  OAI22X1TS U1291 ( .A0(n429), .A1(n1080), .B0(n439), .B1(n1112), .Y(N10160)
         );
  OAI22X1TS U1292 ( .A0(n429), .A1(n1079), .B0(n439), .B1(n1111), .Y(N10161)
         );
  OAI22X1TS U1293 ( .A0(n428), .A1(n1078), .B0(n439), .B1(n1110), .Y(N10162)
         );
  OAI22X1TS U1294 ( .A0(n428), .A1(n1077), .B0(n439), .B1(n1109), .Y(N10163)
         );
  OAI22X1TS U1295 ( .A0(n428), .A1(n1076), .B0(n445), .B1(n1108), .Y(N10164)
         );
  OAI22X1TS U1296 ( .A0(n428), .A1(n1075), .B0(n443), .B1(n1107), .Y(N10165)
         );
  OAI22X1TS U1297 ( .A0(n434), .A1(n1074), .B0(n443), .B1(n1106), .Y(N10166)
         );
  OAI22X1TS U1298 ( .A0(n438), .A1(n1073), .B0(n1749), .B1(n1105), .Y(N10167)
         );
  OAI22X1TS U1299 ( .A0(n438), .A1(n1072), .B0(n445), .B1(n1104), .Y(N10168)
         );
  OAI22X1TS U1300 ( .A0(n434), .A1(n1071), .B0(n442), .B1(n1103), .Y(N10169)
         );
  OAI22X1TS U1301 ( .A0(n432), .A1(n1070), .B0(n448), .B1(n1102), .Y(N10170)
         );
  OAI22X1TS U1302 ( .A0(n437), .A1(n1069), .B0(n1749), .B1(n1101), .Y(N10171)
         );
  OAI22X1TS U1303 ( .A0(n1750), .A1(n1068), .B0(n446), .B1(n1100), .Y(N10172)
         );
  OAI22X1TS U1304 ( .A0(n435), .A1(n1067), .B0(n446), .B1(n1099), .Y(N10173)
         );
  OAI22X1TS U1305 ( .A0(n435), .A1(n1066), .B0(n442), .B1(n1098), .Y(N10174)
         );
  OAI22X1TS U1306 ( .A0(n435), .A1(n1065), .B0(n448), .B1(n1097), .Y(N10175)
         );
  OAI22X1TS U1307 ( .A0(n432), .A1(n1064), .B0(n446), .B1(n1096), .Y(N10176)
         );
  OAI22X1TS U1308 ( .A0(n433), .A1(n1063), .B0(n445), .B1(n1095), .Y(N10177)
         );
  OAI22X1TS U1309 ( .A0(n435), .A1(n1062), .B0(n446), .B1(n1094), .Y(N10178)
         );
  OAI22X1TS U1310 ( .A0(n434), .A1(n1061), .B0(n445), .B1(n1093), .Y(N10179)
         );
  OAI22X1TS U1311 ( .A0(n433), .A1(n1060), .B0(n444), .B1(n1092), .Y(N10180)
         );
  OAI22X1TS U1312 ( .A0(n436), .A1(n1059), .B0(n447), .B1(n1091), .Y(N10181)
         );
  OAI22X1TS U1313 ( .A0(n434), .A1(n1058), .B0(n444), .B1(n1090), .Y(N10182)
         );
  OAI22X1TS U1314 ( .A0(n457), .A1(n1089), .B0(n398), .B1(n1121), .Y(N10185)
         );
  OAI22X1TS U1315 ( .A0(n457), .A1(n1088), .B0(n398), .B1(n1120), .Y(N10186)
         );
  OAI22X1TS U1316 ( .A0(n457), .A1(n1087), .B0(n398), .B1(n1119), .Y(N10187)
         );
  OAI22X1TS U1317 ( .A0(n456), .A1(n1086), .B0(n406), .B1(n1118), .Y(N10188)
         );
  OAI22X1TS U1318 ( .A0(n456), .A1(n1085), .B0(n406), .B1(n1117), .Y(N10189)
         );
  OAI22X1TS U1319 ( .A0(n456), .A1(n1084), .B0(n406), .B1(n1116), .Y(N10190)
         );
  OAI22X1TS U1320 ( .A0(n456), .A1(n1083), .B0(n403), .B1(n1115), .Y(N10191)
         );
  OAI22X1TS U1321 ( .A0(n455), .A1(n1082), .B0(n404), .B1(n1114), .Y(N10192)
         );
  OAI22X1TS U1322 ( .A0(n455), .A1(n1081), .B0(n1776), .B1(n1113), .Y(N10193)
         );
  OAI22X1TS U1323 ( .A0(n455), .A1(n1080), .B0(n403), .B1(n1112), .Y(N10194)
         );
  OAI22X1TS U1324 ( .A0(n455), .A1(n1079), .B0(n407), .B1(n1111), .Y(N10195)
         );
  OAI22X1TS U1325 ( .A0(n454), .A1(n1078), .B0(n399), .B1(n1110), .Y(N10196)
         );
  OAI22X1TS U1326 ( .A0(n454), .A1(n1077), .B0(n399), .B1(n1109), .Y(N10197)
         );
  OAI22X1TS U1327 ( .A0(n454), .A1(n1076), .B0(n399), .B1(n1108), .Y(N10198)
         );
  OAI22X1TS U1328 ( .A0(n454), .A1(n1075), .B0(n399), .B1(n1107), .Y(N10199)
         );
  OAI22X1TS U1329 ( .A0(n453), .A1(n1074), .B0(n400), .B1(n1106), .Y(N10200)
         );
  OAI22X1TS U1330 ( .A0(n453), .A1(n1073), .B0(n400), .B1(n1105), .Y(N10201)
         );
  OAI22X1TS U1331 ( .A0(n453), .A1(n1072), .B0(n400), .B1(n1104), .Y(N10202)
         );
  OAI22X1TS U1332 ( .A0(n452), .A1(n1071), .B0(n400), .B1(n1103), .Y(N10203)
         );
  OAI22X1TS U1333 ( .A0(n452), .A1(n1070), .B0(n401), .B1(n1102), .Y(N10204)
         );
  OAI22X1TS U1334 ( .A0(n452), .A1(n1069), .B0(n401), .B1(n1101), .Y(N10205)
         );
  OAI22X1TS U1335 ( .A0(n452), .A1(n1068), .B0(n401), .B1(n1100), .Y(N10206)
         );
  OAI22X1TS U1336 ( .A0(n451), .A1(n1067), .B0(n401), .B1(n1099), .Y(N10207)
         );
  OAI22X1TS U1337 ( .A0(n451), .A1(n1066), .B0(n404), .B1(n1098), .Y(N10208)
         );
  OAI22X1TS U1338 ( .A0(n453), .A1(n1065), .B0(n405), .B1(n1097), .Y(N10209)
         );
  OAI22X1TS U1339 ( .A0(n451), .A1(n1064), .B0(n405), .B1(n1096), .Y(N10210)
         );
  OAI22X1TS U1340 ( .A0(n451), .A1(n1063), .B0(n1776), .B1(n1095), .Y(N10211)
         );
  OAI22X1TS U1341 ( .A0(n450), .A1(n1062), .B0(n402), .B1(n1094), .Y(N10212)
         );
  OAI22X1TS U1342 ( .A0(n450), .A1(n1061), .B0(n402), .B1(n1093), .Y(N10213)
         );
  OAI22X1TS U1343 ( .A0(n450), .A1(n1060), .B0(n402), .B1(n1092), .Y(N10214)
         );
  OAI22X1TS U1344 ( .A0(n450), .A1(n1059), .B0(n402), .B1(n1091), .Y(N10215)
         );
  OAI22X1TS U1345 ( .A0(n449), .A1(n1058), .B0(n403), .B1(n1090), .Y(N10216)
         );
  NAND4X1TS U1346 ( .A(n1690), .B(n1598), .C(n1459), .D(n2498), .Y(n1455) );
  OAI22X1TS U1347 ( .A0(n2229), .A1(n818), .B0(n423), .B1(n817), .Y(N10020) );
  OAI22X1TS U1348 ( .A0(n436), .A1(n818), .B0(n442), .B1(n817), .Y(N10030) );
  OAI22X1TS U1349 ( .A0(n449), .A1(n818), .B0(n398), .B1(n817), .Y(N10040) );
  OAI22X1TS U1350 ( .A0(n392), .A1(n673), .B0(n1415), .B1(n2319), .Y(n3203) );
  INVX2TS U1351 ( .A(requesterAddressIn_WEST[0]), .Y(n2319) );
  OAI22X1TS U1352 ( .A0(n393), .A1(n672), .B0(n1415), .B1(n2320), .Y(n3204) );
  INVX2TS U1353 ( .A(requesterAddressIn_WEST[1]), .Y(n2320) );
  OAI22X1TS U1354 ( .A0(n392), .A1(n671), .B0(n362), .B1(n2321), .Y(n3205) );
  INVX2TS U1355 ( .A(requesterAddressIn_WEST[2]), .Y(n2321) );
  OAI22X1TS U1356 ( .A0(n393), .A1(n670), .B0(n362), .B1(n2322), .Y(n3206) );
  INVX2TS U1357 ( .A(requesterAddressIn_WEST[3]), .Y(n2322) );
  OAI22X1TS U1358 ( .A0(n392), .A1(n669), .B0(n362), .B1(n2323), .Y(n3207) );
  INVX2TS U1359 ( .A(requesterAddressIn_WEST[4]), .Y(n2323) );
  OAI22X1TS U1360 ( .A0(n393), .A1(n668), .B0(n362), .B1(n2324), .Y(n3208) );
  INVX2TS U1361 ( .A(requesterAddressIn_WEST[5]), .Y(n2324) );
  NAND2X1TS U1362 ( .A(n1751), .B(n1750), .Y(n1749) );
  XOR2X1TS U1363 ( .A(n962), .B(n1), .Y(n1141) );
  NAND2X1TS U1364 ( .A(n1774), .B(n2211), .Y(n1775) );
  NAND2X1TS U1365 ( .A(n1763), .B(n936), .Y(n1761) );
  CLKBUFX2TS U1366 ( .A(n1776), .Y(n406) );
  CLKBUFX2TS U1367 ( .A(n1750), .Y(n437) );
  OAI32X1TS U1368 ( .A0(n1461), .A1(n1138), .A2(n958), .B0(n2182), .B1(n659), 
        .Y(n3344) );
  OAI21X1TS U1369 ( .A0(n962), .A1(n1155), .B0(n2205), .Y(n1461) );
  INVX2TS U1370 ( .A(n1462), .Y(n958) );
  INVX2TS U1371 ( .A(n1773), .Y(n937) );
  CLKBUFX2TS U1372 ( .A(n1776), .Y(n407) );
  CLKBUFX2TS U1373 ( .A(n396), .Y(n460) );
  INVX2TS U1374 ( .A(n1762), .Y(n936) );
  NOR3X1TS U1375 ( .A(n459), .B(n2485), .C(n91), .Y(n1733) );
  NOR3BX1TS U1376 ( .AN(n431), .B(n2489), .C(n1751), .Y(n1740) );
  NAND2X1TS U1377 ( .A(n1131), .B(n2497), .Y(n1132) );
  OAI22X1TS U1378 ( .A0(n2211), .A1(n818), .B0(n413), .B1(n817), .Y(N10010) );
  NAND2X1TS U1379 ( .A(n1773), .B(n2495), .Y(n1764) );
  CLKBUFX2TS U1380 ( .A(n2327), .Y(n2326) );
  CLKBUFX2TS U1381 ( .A(n2333), .Y(n2332) );
  CLKBUFX2TS U1382 ( .A(n2339), .Y(n2338) );
  CLKBUFX2TS U1383 ( .A(n2342), .Y(n2341) );
  CLKBUFX2TS U1384 ( .A(n2345), .Y(n2344) );
  CLKBUFX2TS U1385 ( .A(n2351), .Y(n2350) );
  CLKBUFX2TS U1386 ( .A(n2354), .Y(n2353) );
  CLKBUFX2TS U1387 ( .A(n2360), .Y(n2359) );
  CLKBUFX2TS U1388 ( .A(n2363), .Y(n2362) );
  CLKBUFX2TS U1389 ( .A(n2369), .Y(n2368) );
  CLKBUFX2TS U1390 ( .A(n2375), .Y(n2374) );
  CLKBUFX2TS U1391 ( .A(n2378), .Y(n2377) );
  CLKBUFX2TS U1392 ( .A(n2381), .Y(n2380) );
  CLKBUFX2TS U1393 ( .A(n2393), .Y(n2392) );
  CLKBUFX2TS U1394 ( .A(n2396), .Y(n2395) );
  CLKBUFX2TS U1395 ( .A(n2402), .Y(n2401) );
  CLKBUFX2TS U1396 ( .A(n2405), .Y(n2404) );
  CLKBUFX2TS U1397 ( .A(n2408), .Y(n2407) );
  CLKBUFX2TS U1398 ( .A(n2411), .Y(n2410) );
  CLKBUFX2TS U1399 ( .A(n2414), .Y(n2413) );
  CLKBUFX2TS U1400 ( .A(n2417), .Y(n2416) );
  CLKBUFX2TS U1401 ( .A(n2420), .Y(n2419) );
  CLKBUFX2TS U1402 ( .A(n2297), .Y(n2296) );
  CLKBUFX2TS U1403 ( .A(n2300), .Y(n2299) );
  CLKBUFX2TS U1404 ( .A(n2303), .Y(n2302) );
  CLKBUFX2TS U1405 ( .A(n2309), .Y(n2308) );
  CLKBUFX2TS U1406 ( .A(n1750), .Y(n438) );
  NOR2X1TS U1407 ( .A(n658), .B(n2203), .Y(n3252) );
  NOR2X1TS U1408 ( .A(n657), .B(n2202), .Y(n3253) );
  INVX2TS U1409 ( .A(n2422), .Y(n2421) );
  INVX2TS U1410 ( .A(n2424), .Y(n2423) );
  INVX2TS U1411 ( .A(n2426), .Y(n2425) );
  INVX2TS U1412 ( .A(n2428), .Y(n2427) );
  INVX2TS U1413 ( .A(n2430), .Y(n2429) );
  INVX2TS U1414 ( .A(n2432), .Y(n2431) );
  INVX2TS U1415 ( .A(n2434), .Y(n2433) );
  INVX2TS U1416 ( .A(n2436), .Y(n2435) );
  INVX2TS U1417 ( .A(n2438), .Y(n2437) );
  INVX2TS U1418 ( .A(n2440), .Y(n2439) );
  INVX2TS U1419 ( .A(n2442), .Y(n2441) );
  INVX2TS U1420 ( .A(n2444), .Y(n2443) );
  INVX2TS U1421 ( .A(n2446), .Y(n2445) );
  INVX2TS U1422 ( .A(n2448), .Y(n2447) );
  INVX2TS U1423 ( .A(n2450), .Y(n2449) );
  INVX2TS U1424 ( .A(n2452), .Y(n2451) );
  INVX2TS U1425 ( .A(n2454), .Y(n2453) );
  INVX2TS U1426 ( .A(n2456), .Y(n2455) );
  INVX2TS U1427 ( .A(n2458), .Y(n2457) );
  INVX2TS U1428 ( .A(n2460), .Y(n2459) );
  INVX2TS U1429 ( .A(n2462), .Y(n2461) );
  INVX2TS U1430 ( .A(n2464), .Y(n2463) );
  INVX2TS U1431 ( .A(n2466), .Y(n2465) );
  INVX2TS U1432 ( .A(n2468), .Y(n2467) );
  INVX2TS U1433 ( .A(n2470), .Y(n2469) );
  INVX2TS U1434 ( .A(n2472), .Y(n2471) );
  INVX2TS U1435 ( .A(n2474), .Y(n2473) );
  INVX2TS U1436 ( .A(n2476), .Y(n2475) );
  INVX2TS U1437 ( .A(n2478), .Y(n2477) );
  INVX2TS U1438 ( .A(n2480), .Y(n2479) );
  INVX2TS U1439 ( .A(n2482), .Y(n2481) );
  INVX2TS U1440 ( .A(n2484), .Y(n2483) );
  INVX2TS U1441 ( .A(cacheAddressIn_WEST[6]), .Y(n2315) );
  INVX2TS U1442 ( .A(cacheAddressIn_WEST[7]), .Y(n2318) );
  CLKBUFX2TS U1443 ( .A(n2330), .Y(n2329) );
  CLKBUFX2TS U1444 ( .A(n2336), .Y(n2335) );
  CLKBUFX2TS U1445 ( .A(n2348), .Y(n2347) );
  CLKBUFX2TS U1446 ( .A(n2357), .Y(n2356) );
  CLKBUFX2TS U1447 ( .A(n2366), .Y(n2365) );
  CLKBUFX2TS U1448 ( .A(n2372), .Y(n2371) );
  CLKBUFX2TS U1449 ( .A(n2384), .Y(n2383) );
  CLKBUFX2TS U1450 ( .A(n2387), .Y(n2386) );
  CLKBUFX2TS U1451 ( .A(n2390), .Y(n2389) );
  CLKBUFX2TS U1452 ( .A(n2399), .Y(n2398) );
  CLKBUFX2TS U1453 ( .A(n2306), .Y(n2305) );
  CLKBUFX2TS U1454 ( .A(n2312), .Y(n2311) );
  OAI32X1TS U1455 ( .A0(n674), .A1(n2491), .A2(n43), .B0(n655), .B1(n1132), 
        .Y(n2104) );
  OAI32X1TS U1456 ( .A0(n655), .A1(n2493), .A2(n757), .B0(n650), .B1(n1123), 
        .Y(n2099) );
  OAI32X1TS U1457 ( .A0(n931), .A1(n2490), .A2(n811), .B0(n1122), .B1(n932), 
        .Y(n3383) );
  OAI32X1TS U1458 ( .A0(n930), .A1(n2491), .A2(n756), .B0(n1123), .B1(n931), 
        .Y(n3381) );
  OAI32X1TS U1459 ( .A0(n933), .A1(n2492), .A2(n754), .B0(n1132), .B1(n930), 
        .Y(n3379) );
  OAI32X1TS U1460 ( .A0(n657), .A1(n2491), .A2(n371), .B0(n1129), .B1(n654), 
        .Y(n2102) );
  OAI32X1TS U1461 ( .A0(n658), .A1(n2492), .A2(n371), .B0(n1129), .B1(n653), 
        .Y(n2100) );
  INVX2TS U1462 ( .A(n1416), .Y(n813) );
  INVX2TS U1463 ( .A(n1125), .Y(n757) );
  INVX2TS U1464 ( .A(n1477), .Y(n743) );
  XOR2X1TS U1465 ( .A(n880), .B(n372), .Y(n1571) );
  NOR2X1TS U1466 ( .A(memWrite_SOUTH), .B(memRead_SOUTH), .Y(n1460) );
  NAND3X1TS U1467 ( .A(n1527), .B(n98), .C(n1299), .Y(n1265) );
  INVX2TS U1468 ( .A(memRead_EAST), .Y(n976) );
  OAI221XLTS U1469 ( .A0(n1005), .A1(n2296), .B0(n72), .B1(n61), .C0(n1518), 
        .Y(n3317) );
  AOI22X1TS U1470 ( .A0(n370), .A1(n2279), .B0(n1007), .B1(n682), .Y(n1518) );
  OAI221XLTS U1471 ( .A0(n1003), .A1(n2299), .B0(n73), .B1(n61), .C0(n1520), 
        .Y(n3316) );
  OAI221XLTS U1472 ( .A0(n1003), .A1(n2302), .B0(n74), .B1(n61), .C0(n1521), 
        .Y(n3315) );
  OAI221XLTS U1473 ( .A0(n1003), .A1(n2305), .B0(n75), .B1(n61), .C0(n1522), 
        .Y(n3314) );
  OAI221XLTS U1474 ( .A0(n994), .A1(n2308), .B0(n76), .B1(n387), .C0(n1523), 
        .Y(n3313) );
  OAI221XLTS U1475 ( .A0(n994), .A1(n2311), .B0(n77), .B1(n387), .C0(n1524), 
        .Y(n3312) );
  OAI221XLTS U1476 ( .A0(n994), .A1(n2314), .B0(n78), .B1(n387), .C0(n1525), 
        .Y(n3311) );
  OAI221XLTS U1477 ( .A0(n994), .A1(n2317), .B0(n79), .B1(n387), .C0(n1526), 
        .Y(n3310) );
  OAI221XLTS U1478 ( .A0(n1041), .A1(n2296), .B0(n386), .B1(n954), .C0(n1504), 
        .Y(n3325) );
  AOI2BB2X1TS U1479 ( .B0(n367), .B1(n2279), .A0N(n1053), .A1N(n48), .Y(n1504)
         );
  OAI221XLTS U1480 ( .A0(n1038), .A1(n2299), .B0(n385), .B1(n953), .C0(n1506), 
        .Y(n3324) );
  AOI2BB2X1TS U1481 ( .B0(n367), .B1(n2281), .A0N(n1053), .A1N(n50), .Y(n1506)
         );
  OAI221XLTS U1482 ( .A0(n1039), .A1(n2302), .B0(n386), .B1(n952), .C0(n1507), 
        .Y(n3323) );
  AOI2BB2X1TS U1483 ( .B0(n367), .B1(n2283), .A0N(n1051), .A1N(n52), .Y(n1507)
         );
  OAI221XLTS U1484 ( .A0(n1041), .A1(n2305), .B0(n385), .B1(n951), .C0(n1508), 
        .Y(n3322) );
  AOI2BB2X1TS U1485 ( .B0(n367), .B1(n2285), .A0N(n1052), .A1N(n54), .Y(n1508)
         );
  OAI221XLTS U1486 ( .A0(n1030), .A1(n2308), .B0(n386), .B1(n950), .C0(n1509), 
        .Y(n3321) );
  AOI2BB2X1TS U1487 ( .B0(n368), .B1(n2287), .A0N(n1042), .A1N(n56), .Y(n1509)
         );
  OAI221XLTS U1488 ( .A0(n1030), .A1(n2311), .B0(n385), .B1(n949), .C0(n1510), 
        .Y(n3320) );
  AOI2BB2X1TS U1489 ( .B0(n368), .B1(n2289), .A0N(n1042), .A1N(n58), .Y(n1510)
         );
  OAI221XLTS U1490 ( .A0(n1030), .A1(n2314), .B0(n386), .B1(n948), .C0(n1511), 
        .Y(n3319) );
  AOI2BB2X1TS U1491 ( .B0(n368), .B1(n2291), .A0N(n1042), .A1N(n60), .Y(n1511)
         );
  OAI221XLTS U1492 ( .A0(n1030), .A1(n2317), .B0(n385), .B1(n947), .C0(n1512), 
        .Y(n3318) );
  AOI2BB2X1TS U1493 ( .B0(n368), .B1(n2293), .A0N(n1042), .A1N(n62), .Y(n1512)
         );
  OAI221XLTS U1494 ( .A0(n959), .A1(n2297), .B0(n48), .B1(n750), .C0(n1532), 
        .Y(n3309) );
  AOI22X1TS U1495 ( .A0(n354), .A1(n2279), .B0(n970), .B1(n698), .Y(n1532) );
  OAI221XLTS U1496 ( .A0(n967), .A1(n2300), .B0(n50), .B1(n750), .C0(n1534), 
        .Y(n3308) );
  AOI22X1TS U1497 ( .A0(n354), .A1(n2281), .B0(n970), .B1(n697), .Y(n1534) );
  OAI221XLTS U1498 ( .A0(n968), .A1(n2303), .B0(n52), .B1(n750), .C0(n1535), 
        .Y(n3307) );
  AOI22X1TS U1499 ( .A0(n354), .A1(n2283), .B0(n970), .B1(n696), .Y(n1535) );
  OAI221XLTS U1500 ( .A0(n1301), .A1(n2305), .B0(n54), .B1(n750), .C0(n1536), 
        .Y(n3306) );
  AOI22X1TS U1501 ( .A0(n354), .A1(n2285), .B0(n970), .B1(n695), .Y(n1536) );
  OAI221XLTS U1502 ( .A0(n959), .A1(n2309), .B0(n56), .B1(n751), .C0(n1537), 
        .Y(n3305) );
  AOI22X1TS U1503 ( .A0(n355), .A1(n2287), .B0(n969), .B1(n694), .Y(n1537) );
  OAI221XLTS U1504 ( .A0(n959), .A1(n2311), .B0(n58), .B1(n751), .C0(n1538), 
        .Y(n3304) );
  AOI22X1TS U1505 ( .A0(n355), .A1(n2289), .B0(n969), .B1(n693), .Y(n1538) );
  OAI221XLTS U1506 ( .A0(n959), .A1(n2315), .B0(n60), .B1(n751), .C0(n1539), 
        .Y(n3303) );
  AOI22X1TS U1507 ( .A0(n355), .A1(n2291), .B0(n969), .B1(n692), .Y(n1539) );
  OAI221XLTS U1508 ( .A0(n968), .A1(n2318), .B0(n62), .B1(n751), .C0(n1540), 
        .Y(n3302) );
  AOI22X1TS U1509 ( .A0(n355), .A1(n2293), .B0(n969), .B1(n691), .Y(n1540) );
  OAI221XLTS U1510 ( .A0(n1810), .A1(n983), .B0(n2326), .B1(n816), .C0(n1302), 
        .Y(n3513) );
  AOI2BB2X1TS U1511 ( .B0(n768), .B1(n2421), .A0N(n689), .A1N(n1809), .Y(n1302) );
  OAI221XLTS U1512 ( .A0(n1811), .A1(n983), .B0(n2329), .B1(n816), .C0(n1305), 
        .Y(n3512) );
  AOI2BB2X1TS U1513 ( .B0(n768), .B1(n2423), .A0N(n689), .A1N(n1785), .Y(n1305) );
  OAI221XLTS U1514 ( .A0(n1812), .A1(n981), .B0(n2332), .B1(n816), .C0(n1306), 
        .Y(n3511) );
  AOI2BB2X1TS U1515 ( .B0(n768), .B1(n2425), .A0N(n689), .A1N(n1786), .Y(n1306) );
  OAI221XLTS U1516 ( .A0(n1813), .A1(n981), .B0(n2335), .B1(n816), .C0(n1307), 
        .Y(n3510) );
  AOI2BB2X1TS U1517 ( .B0(n768), .B1(n2427), .A0N(n689), .A1N(n1787), .Y(n1307) );
  OAI221XLTS U1518 ( .A0(n1815), .A1(n981), .B0(n2338), .B1(n815), .C0(n1308), 
        .Y(n3509) );
  AOI2BB2X1TS U1519 ( .B0(n767), .B1(n2429), .A0N(n690), .A1N(n1814), .Y(n1308) );
  OAI221XLTS U1520 ( .A0(n1816), .A1(n981), .B0(n2341), .B1(n815), .C0(n1309), 
        .Y(n3508) );
  AOI2BB2X1TS U1521 ( .B0(n767), .B1(n2431), .A0N(n690), .A1N(n1788), .Y(n1309) );
  OAI221XLTS U1522 ( .A0(n1817), .A1(n980), .B0(n2344), .B1(n815), .C0(n1310), 
        .Y(n3507) );
  AOI2BB2X1TS U1523 ( .B0(n767), .B1(n2433), .A0N(n690), .A1N(n1789), .Y(n1310) );
  OAI221XLTS U1524 ( .A0(n1818), .A1(n980), .B0(n2347), .B1(n815), .C0(n1311), 
        .Y(n3506) );
  AOI2BB2X1TS U1525 ( .B0(n767), .B1(n2435), .A0N(n690), .A1N(n1790), .Y(n1311) );
  OAI221XLTS U1526 ( .A0(n1820), .A1(n980), .B0(n2350), .B1(n807), .C0(n1312), 
        .Y(n3505) );
  AOI2BB2X1TS U1527 ( .B0(n766), .B1(n2437), .A0N(n741), .A1N(n1819), .Y(n1312) );
  OAI221XLTS U1528 ( .A0(n1821), .A1(n980), .B0(n2353), .B1(n807), .C0(n1313), 
        .Y(n3504) );
  AOI2BB2X1TS U1529 ( .B0(n766), .B1(n2439), .A0N(n741), .A1N(n1791), .Y(n1313) );
  OAI221XLTS U1530 ( .A0(n1822), .A1(n979), .B0(n2356), .B1(n807), .C0(n1314), 
        .Y(n3503) );
  AOI2BB2X1TS U1531 ( .B0(n766), .B1(n2441), .A0N(n741), .A1N(n1792), .Y(n1314) );
  OAI221XLTS U1532 ( .A0(n1823), .A1(n979), .B0(n2359), .B1(n807), .C0(n1315), 
        .Y(n3502) );
  AOI2BB2X1TS U1533 ( .B0(n766), .B1(n2443), .A0N(n741), .A1N(n1793), .Y(n1315) );
  OAI221XLTS U1534 ( .A0(n1825), .A1(n979), .B0(n2362), .B1(n806), .C0(n1316), 
        .Y(n3501) );
  AOI2BB2X1TS U1535 ( .B0(n765), .B1(n2445), .A0N(n744), .A1N(n1824), .Y(n1316) );
  OAI221XLTS U1536 ( .A0(n1826), .A1(n979), .B0(n2365), .B1(n806), .C0(n1317), 
        .Y(n3500) );
  AOI2BB2X1TS U1537 ( .B0(n765), .B1(n2447), .A0N(n744), .A1N(n1794), .Y(n1317) );
  OAI221XLTS U1538 ( .A0(n1827), .A1(n978), .B0(n2368), .B1(n806), .C0(n1318), 
        .Y(n3499) );
  AOI2BB2X1TS U1539 ( .B0(n765), .B1(n2449), .A0N(n744), .A1N(n1795), .Y(n1318) );
  OAI221XLTS U1540 ( .A0(n1828), .A1(n978), .B0(n2371), .B1(n806), .C0(n1319), 
        .Y(n3498) );
  AOI2BB2X1TS U1541 ( .B0(n765), .B1(n2451), .A0N(n744), .A1N(n1796), .Y(n1319) );
  OAI221XLTS U1542 ( .A0(n1830), .A1(n978), .B0(n2374), .B1(n804), .C0(n1320), 
        .Y(n3497) );
  AOI2BB2X1TS U1543 ( .B0(n764), .B1(n2453), .A0N(n745), .A1N(n1829), .Y(n1320) );
  OAI221XLTS U1544 ( .A0(n1831), .A1(n978), .B0(n2377), .B1(n804), .C0(n1321), 
        .Y(n3496) );
  AOI2BB2X1TS U1545 ( .B0(n764), .B1(n2455), .A0N(n745), .A1N(n1797), .Y(n1321) );
  OAI221XLTS U1546 ( .A0(n1832), .A1(n974), .B0(n2380), .B1(n804), .C0(n1322), 
        .Y(n3495) );
  AOI2BB2X1TS U1547 ( .B0(n764), .B1(n2457), .A0N(n745), .A1N(n1798), .Y(n1322) );
  OAI221XLTS U1548 ( .A0(n1833), .A1(n974), .B0(n2383), .B1(n804), .C0(n1323), 
        .Y(n3494) );
  AOI2BB2X1TS U1549 ( .B0(n764), .B1(n2459), .A0N(n745), .A1N(n1799), .Y(n1323) );
  OAI221XLTS U1550 ( .A0(n1835), .A1(n974), .B0(n2386), .B1(n955), .C0(n1324), 
        .Y(n3493) );
  AOI2BB2X1TS U1551 ( .B0(n763), .B1(n2461), .A0N(n746), .A1N(n1834), .Y(n1324) );
  OAI221XLTS U1552 ( .A0(n1836), .A1(n974), .B0(n2389), .B1(n955), .C0(n1325), 
        .Y(n3492) );
  AOI2BB2X1TS U1553 ( .B0(n763), .B1(n2463), .A0N(n746), .A1N(n1800), .Y(n1325) );
  OAI221XLTS U1554 ( .A0(n1837), .A1(n973), .B0(n2392), .B1(n831), .C0(n1326), 
        .Y(n3491) );
  AOI2BB2X1TS U1555 ( .B0(n763), .B1(n2465), .A0N(n746), .A1N(n1801), .Y(n1326) );
  OAI221XLTS U1556 ( .A0(n1838), .A1(n973), .B0(n2395), .B1(n1301), .C0(n1327), 
        .Y(n3490) );
  AOI2BB2X1TS U1557 ( .B0(n763), .B1(n2467), .A0N(n746), .A1N(n1802), .Y(n1327) );
  OAI221XLTS U1558 ( .A0(n1840), .A1(n973), .B0(n2398), .B1(n956), .C0(n1328), 
        .Y(n3489) );
  AOI2BB2X1TS U1559 ( .B0(n799), .B1(n2469), .A0N(n747), .A1N(n1839), .Y(n1328) );
  OAI221XLTS U1560 ( .A0(n1841), .A1(n973), .B0(n2401), .B1(n956), .C0(n1329), 
        .Y(n3488) );
  AOI2BB2X1TS U1561 ( .B0(n799), .B1(n2471), .A0N(n747), .A1N(n1803), .Y(n1329) );
  OAI221XLTS U1562 ( .A0(n1842), .A1(n972), .B0(n2404), .B1(n935), .C0(n1330), 
        .Y(n3487) );
  AOI2BB2X1TS U1563 ( .B0(n772), .B1(n2473), .A0N(n747), .A1N(n1804), .Y(n1330) );
  OAI221XLTS U1564 ( .A0(n1843), .A1(n972), .B0(n2407), .B1(n935), .C0(n1331), 
        .Y(n3486) );
  AOI2BB2X1TS U1565 ( .B0(n799), .B1(n2475), .A0N(n747), .A1N(n1805), .Y(n1331) );
  OAI221XLTS U1566 ( .A0(n1845), .A1(n972), .B0(n2410), .B1(n956), .C0(n1332), 
        .Y(n3485) );
  AOI2BB2X1TS U1567 ( .B0(n762), .B1(n2477), .A0N(n749), .A1N(n1844), .Y(n1332) );
  OAI221XLTS U1568 ( .A0(n1846), .A1(n971), .B0(n2413), .B1(n956), .C0(n1333), 
        .Y(n3484) );
  AOI2BB2X1TS U1569 ( .B0(n762), .B1(n2479), .A0N(n749), .A1N(n1806), .Y(n1333) );
  OAI221XLTS U1570 ( .A0(n1847), .A1(n971), .B0(n2416), .B1(n955), .C0(n1334), 
        .Y(n3483) );
  AOI2BB2X1TS U1571 ( .B0(n762), .B1(n2481), .A0N(n749), .A1N(n1807), .Y(n1334) );
  OAI221XLTS U1572 ( .A0(n1848), .A1(n971), .B0(n2419), .B1(n831), .C0(n1335), 
        .Y(n3482) );
  AOI2BB2X1TS U1573 ( .B0(n762), .B1(n2483), .A0N(n749), .A1N(n1808), .Y(n1335) );
  OAI221XLTS U1574 ( .A0(n1809), .A1(n1051), .B0(n2327), .B1(n1040), .C0(n1230), .Y(n3577) );
  AOI22X1TS U1575 ( .A0(n1023), .A1(n2421), .B0(n2260), .B1(n1892), .Y(n1230)
         );
  OAI221XLTS U1576 ( .A0(n1785), .A1(n1052), .B0(n2329), .B1(n1040), .C0(n1232), .Y(n3576) );
  OAI221XLTS U1577 ( .A0(n1786), .A1(n1050), .B0(n2333), .B1(n1039), .C0(n1233), .Y(n3575) );
  AOI22X1TS U1578 ( .A0(n1023), .A1(n2425), .B0(n2264), .B1(n1894), .Y(n1233)
         );
  OAI221XLTS U1579 ( .A0(n1787), .A1(n1050), .B0(n2335), .B1(n1038), .C0(n1234), .Y(n3574) );
  AOI22X1TS U1580 ( .A0(n1023), .A1(n2427), .B0(n2262), .B1(n1895), .Y(n1234)
         );
  OAI221XLTS U1581 ( .A0(n1814), .A1(n1049), .B0(n2339), .B1(n1037), .C0(n1235), .Y(n3573) );
  AOI22X1TS U1582 ( .A0(n1022), .A1(n2429), .B0(n2262), .B1(n1896), .Y(n1235)
         );
  OAI221XLTS U1583 ( .A0(n1788), .A1(n1049), .B0(n2342), .B1(n1037), .C0(n1236), .Y(n3572) );
  AOI22X1TS U1584 ( .A0(n1022), .A1(n2431), .B0(n2261), .B1(n1897), .Y(n1236)
         );
  OAI221XLTS U1585 ( .A0(n1789), .A1(n1049), .B0(n2345), .B1(n1037), .C0(n1237), .Y(n3571) );
  AOI22X1TS U1586 ( .A0(n1022), .A1(n2433), .B0(n2267), .B1(n1898), .Y(n1237)
         );
  OAI221XLTS U1587 ( .A0(n1790), .A1(n1049), .B0(n2347), .B1(n1037), .C0(n1238), .Y(n3570) );
  AOI22X1TS U1588 ( .A0(n1022), .A1(n2435), .B0(n2264), .B1(n1899), .Y(n1238)
         );
  OAI221XLTS U1589 ( .A0(n1819), .A1(n1048), .B0(n2351), .B1(n1036), .C0(n1239), .Y(n3569) );
  AOI22X1TS U1590 ( .A0(n1027), .A1(n2437), .B0(n2264), .B1(n1900), .Y(n1239)
         );
  OAI221XLTS U1591 ( .A0(n1791), .A1(n1048), .B0(n2354), .B1(n1036), .C0(n1240), .Y(n3568) );
  AOI22X1TS U1592 ( .A0(n1027), .A1(n2439), .B0(n2261), .B1(n1901), .Y(n1240)
         );
  OAI221XLTS U1593 ( .A0(n1792), .A1(n1048), .B0(n2356), .B1(n1036), .C0(n1241), .Y(n3567) );
  AOI22X1TS U1594 ( .A0(n1026), .A1(n2441), .B0(n2263), .B1(n1902), .Y(n1241)
         );
  OAI221XLTS U1595 ( .A0(n1793), .A1(n1048), .B0(n2360), .B1(n1036), .C0(n1242), .Y(n3566) );
  AOI22X1TS U1596 ( .A0(n1029), .A1(n2443), .B0(n2263), .B1(n1903), .Y(n1242)
         );
  OAI221XLTS U1597 ( .A0(n1824), .A1(n1047), .B0(n2363), .B1(n1035), .C0(n1243), .Y(n3565) );
  AOI22X1TS U1598 ( .A0(n1027), .A1(n2445), .B0(n2263), .B1(n1904), .Y(n1243)
         );
  OAI221XLTS U1599 ( .A0(n1794), .A1(n1047), .B0(n2365), .B1(n1035), .C0(n1244), .Y(n3564) );
  AOI22X1TS U1600 ( .A0(n1028), .A1(n2447), .B0(n2264), .B1(n1905), .Y(n1244)
         );
  OAI221XLTS U1601 ( .A0(n1795), .A1(n1047), .B0(n2369), .B1(n1035), .C0(n1245), .Y(n3563) );
  AOI22X1TS U1602 ( .A0(n1027), .A1(n2449), .B0(n2260), .B1(n1906), .Y(n1245)
         );
  OAI221XLTS U1603 ( .A0(n1796), .A1(n1047), .B0(n2371), .B1(n1035), .C0(n1246), .Y(n3562) );
  AOI22X1TS U1604 ( .A0(n1028), .A1(n2451), .B0(n2267), .B1(n1907), .Y(n1246)
         );
  OAI221XLTS U1605 ( .A0(n1829), .A1(n1046), .B0(n2375), .B1(n1034), .C0(n1247), .Y(n3561) );
  AOI22X1TS U1606 ( .A0(n1021), .A1(n2453), .B0(n2263), .B1(n1908), .Y(n1247)
         );
  OAI221XLTS U1607 ( .A0(n1797), .A1(n1046), .B0(n2378), .B1(n1034), .C0(n1248), .Y(n3560) );
  AOI22X1TS U1608 ( .A0(n1021), .A1(n2455), .B0(n2257), .B1(n1909), .Y(n1248)
         );
  OAI221XLTS U1609 ( .A0(n1798), .A1(n1046), .B0(n2381), .B1(n1034), .C0(n1249), .Y(n3559) );
  AOI22X1TS U1610 ( .A0(n1021), .A1(n2457), .B0(n2257), .B1(n1910), .Y(n1249)
         );
  OAI221XLTS U1611 ( .A0(n1799), .A1(n1046), .B0(n2383), .B1(n1034), .C0(n1250), .Y(n3558) );
  AOI22X1TS U1612 ( .A0(n1021), .A1(n2459), .B0(n2257), .B1(n1923), .Y(n1250)
         );
  OAI221XLTS U1613 ( .A0(n1834), .A1(n1045), .B0(n2386), .B1(n1033), .C0(n1251), .Y(n3557) );
  AOI22X1TS U1614 ( .A0(n1020), .A1(n2461), .B0(n2257), .B1(n1924), .Y(n1251)
         );
  OAI221XLTS U1615 ( .A0(n1800), .A1(n1045), .B0(n2389), .B1(n1033), .C0(n1252), .Y(n3556) );
  AOI22X1TS U1616 ( .A0(n1020), .A1(n2463), .B0(n2258), .B1(n1881), .Y(n1252)
         );
  OAI221XLTS U1617 ( .A0(n1801), .A1(n1045), .B0(n2393), .B1(n1033), .C0(n1253), .Y(n3555) );
  AOI22X1TS U1618 ( .A0(n1020), .A1(n2465), .B0(n2258), .B1(n1882), .Y(n1253)
         );
  OAI221XLTS U1619 ( .A0(n1802), .A1(n1045), .B0(n2396), .B1(n1033), .C0(n1254), .Y(n3554) );
  AOI22X1TS U1620 ( .A0(n1020), .A1(n2467), .B0(n2258), .B1(n1883), .Y(n1254)
         );
  OAI221XLTS U1621 ( .A0(n1839), .A1(n1044), .B0(n2398), .B1(n1032), .C0(n1255), .Y(n3553) );
  AOI22X1TS U1622 ( .A0(n1019), .A1(n2469), .B0(n2258), .B1(n1884), .Y(n1255)
         );
  OAI221XLTS U1623 ( .A0(n1803), .A1(n1044), .B0(n2402), .B1(n1032), .C0(n1256), .Y(n3552) );
  AOI22X1TS U1624 ( .A0(n1019), .A1(n2471), .B0(n2259), .B1(n1885), .Y(n1256)
         );
  OAI221XLTS U1625 ( .A0(n1804), .A1(n1044), .B0(n2405), .B1(n1032), .C0(n1257), .Y(n3551) );
  AOI22X1TS U1626 ( .A0(n1019), .A1(n2473), .B0(n2259), .B1(n1886), .Y(n1257)
         );
  OAI221XLTS U1627 ( .A0(n1805), .A1(n1044), .B0(n2408), .B1(n1032), .C0(n1258), .Y(n3550) );
  AOI22X1TS U1628 ( .A0(n1019), .A1(n2475), .B0(n2259), .B1(n1887), .Y(n1258)
         );
  OAI221XLTS U1629 ( .A0(n1844), .A1(n1043), .B0(n2411), .B1(n1031), .C0(n1259), .Y(n3549) );
  AOI22X1TS U1630 ( .A0(n1018), .A1(n2477), .B0(n2259), .B1(n1888), .Y(n1259)
         );
  OAI221XLTS U1631 ( .A0(n1806), .A1(n1043), .B0(n2414), .B1(n1031), .C0(n1260), .Y(n3548) );
  AOI22X1TS U1632 ( .A0(n1018), .A1(n2479), .B0(n2260), .B1(n1889), .Y(n1260)
         );
  OAI221XLTS U1633 ( .A0(n1807), .A1(n1043), .B0(n2417), .B1(n1031), .C0(n1261), .Y(n3547) );
  AOI22X1TS U1634 ( .A0(n1018), .A1(n2481), .B0(n2260), .B1(n1890), .Y(n1261)
         );
  OAI221XLTS U1635 ( .A0(n1808), .A1(n1043), .B0(n2420), .B1(n1031), .C0(n1262), .Y(n3546) );
  OAI221XLTS U1636 ( .A0(n1849), .A1(n1015), .B0(n2327), .B1(n998), .C0(n1266), 
        .Y(n3545) );
  AOI22X1TS U1637 ( .A0(n990), .A1(n2421), .B0(n2277), .B1(n739), .Y(n1266) );
  OAI221XLTS U1638 ( .A0(n1850), .A1(n1015), .B0(n2329), .B1(n998), .C0(n1268), 
        .Y(n3544) );
  OAI221XLTS U1639 ( .A0(n1851), .A1(n1014), .B0(n2333), .B1(n998), .C0(n1269), 
        .Y(n3543) );
  AOI22X1TS U1640 ( .A0(n990), .A1(n2425), .B0(n2268), .B1(n737), .Y(n1269) );
  OAI221XLTS U1641 ( .A0(n1852), .A1(n1014), .B0(n2335), .B1(n998), .C0(n1270), 
        .Y(n3542) );
  AOI22X1TS U1642 ( .A0(n990), .A1(n2427), .B0(n2268), .B1(n715), .Y(n1270) );
  OAI221XLTS U1643 ( .A0(n1853), .A1(n1014), .B0(n2339), .B1(n997), .C0(n1271), 
        .Y(n3541) );
  AOI22X1TS U1644 ( .A0(n989), .A1(n2429), .B0(n2268), .B1(n714), .Y(n1271) );
  OAI221XLTS U1645 ( .A0(n1854), .A1(n1014), .B0(n2342), .B1(n997), .C0(n1272), 
        .Y(n3540) );
  AOI22X1TS U1646 ( .A0(n989), .A1(n2431), .B0(n2268), .B1(n713), .Y(n1272) );
  OAI221XLTS U1647 ( .A0(n1855), .A1(n1013), .B0(n2345), .B1(n997), .C0(n1273), 
        .Y(n3539) );
  AOI22X1TS U1648 ( .A0(n989), .A1(n2433), .B0(n2269), .B1(n712), .Y(n1273) );
  OAI221XLTS U1649 ( .A0(n1856), .A1(n1013), .B0(n2347), .B1(n997), .C0(n1274), 
        .Y(n3538) );
  AOI22X1TS U1650 ( .A0(n989), .A1(n2435), .B0(n2269), .B1(n711), .Y(n1274) );
  OAI221XLTS U1651 ( .A0(n1857), .A1(n1013), .B0(n2351), .B1(n996), .C0(n1275), 
        .Y(n3537) );
  AOI22X1TS U1652 ( .A0(n988), .A1(n2437), .B0(n2269), .B1(n710), .Y(n1275) );
  OAI221XLTS U1653 ( .A0(n1858), .A1(n1013), .B0(n2354), .B1(n996), .C0(n1276), 
        .Y(n3536) );
  AOI22X1TS U1654 ( .A0(n988), .A1(n2439), .B0(n2269), .B1(n709), .Y(n1276) );
  OAI221XLTS U1655 ( .A0(n1859), .A1(n1012), .B0(n2356), .B1(n996), .C0(n1277), 
        .Y(n3535) );
  AOI22X1TS U1656 ( .A0(n988), .A1(n2441), .B0(n2270), .B1(n708), .Y(n1277) );
  OAI221XLTS U1657 ( .A0(n1860), .A1(n1012), .B0(n2360), .B1(n996), .C0(n1278), 
        .Y(n3534) );
  AOI22X1TS U1658 ( .A0(n988), .A1(n2443), .B0(n2270), .B1(n707), .Y(n1278) );
  OAI221XLTS U1659 ( .A0(n1861), .A1(n1012), .B0(n2363), .B1(n995), .C0(n1279), 
        .Y(n3533) );
  AOI22X1TS U1660 ( .A0(n987), .A1(n2445), .B0(n2270), .B1(n706), .Y(n1279) );
  OAI221XLTS U1661 ( .A0(n1862), .A1(n1012), .B0(n2365), .B1(n995), .C0(n1280), 
        .Y(n3532) );
  AOI22X1TS U1662 ( .A0(n987), .A1(n2447), .B0(n2270), .B1(n705), .Y(n1280) );
  OAI221XLTS U1663 ( .A0(n1863), .A1(n1011), .B0(n2369), .B1(n995), .C0(n1281), 
        .Y(n3531) );
  AOI22X1TS U1664 ( .A0(n987), .A1(n2449), .B0(n2274), .B1(n704), .Y(n1281) );
  OAI221XLTS U1665 ( .A0(n1864), .A1(n1011), .B0(n2371), .B1(n995), .C0(n1282), 
        .Y(n3530) );
  AOI22X1TS U1666 ( .A0(n987), .A1(n2451), .B0(n2276), .B1(n703), .Y(n1282) );
  OAI221XLTS U1667 ( .A0(n1865), .A1(n1011), .B0(n2375), .B1(n1001), .C0(n1283), .Y(n3529) );
  AOI22X1TS U1668 ( .A0(n986), .A1(n2453), .B0(n2275), .B1(n702), .Y(n1283) );
  OAI221XLTS U1669 ( .A0(n1866), .A1(n1011), .B0(n2378), .B1(n1000), .C0(n1284), .Y(n3528) );
  AOI22X1TS U1670 ( .A0(n986), .A1(n2455), .B0(n2271), .B1(n701), .Y(n1284) );
  OAI221XLTS U1671 ( .A0(n1867), .A1(n1010), .B0(n2381), .B1(n1265), .C0(n1285), .Y(n3527) );
  AOI22X1TS U1672 ( .A0(n986), .A1(n2457), .B0(n2271), .B1(n700), .Y(n1285) );
  OAI221XLTS U1673 ( .A0(n1868), .A1(n1010), .B0(n2383), .B1(n1265), .C0(n1286), .Y(n3526) );
  AOI22X1TS U1674 ( .A0(n986), .A1(n2459), .B0(n2271), .B1(n699), .Y(n1286) );
  OAI221XLTS U1675 ( .A0(n1869), .A1(n1010), .B0(n2386), .B1(n1001), .C0(n1287), .Y(n3525) );
  OAI221XLTS U1676 ( .A0(n1870), .A1(n1010), .B0(n2389), .B1(n1001), .C0(n1288), .Y(n3524) );
  OAI221XLTS U1677 ( .A0(n1871), .A1(n1009), .B0(n2393), .B1(n1001), .C0(n1289), .Y(n3523) );
  OAI221XLTS U1678 ( .A0(n1872), .A1(n1009), .B0(n2396), .B1(n999), .C0(n1290), 
        .Y(n3522) );
  OAI221XLTS U1679 ( .A0(n1873), .A1(n1009), .B0(n2398), .B1(n1002), .C0(n1291), .Y(n3521) );
  OAI221XLTS U1680 ( .A0(n1874), .A1(n1009), .B0(n2402), .B1(n1002), .C0(n1292), .Y(n3520) );
  OAI221XLTS U1681 ( .A0(n1875), .A1(n1017), .B0(n2405), .B1(n1000), .C0(n1293), .Y(n3519) );
  AOI22X1TS U1682 ( .A0(n985), .A1(n2473), .B0(n2273), .B1(n1917), .Y(n1293)
         );
  OAI221XLTS U1683 ( .A0(n1876), .A1(n1015), .B0(n2408), .B1(n999), .C0(n1294), 
        .Y(n3518) );
  OAI221XLTS U1684 ( .A0(n1877), .A1(n1015), .B0(n2411), .B1(n1002), .C0(n1295), .Y(n3517) );
  OAI221XLTS U1685 ( .A0(n1878), .A1(n1008), .B0(n2414), .B1(n1002), .C0(n1296), .Y(n3516) );
  OAI221XLTS U1686 ( .A0(n1879), .A1(n1008), .B0(n2417), .B1(n1005), .C0(n1297), .Y(n3515) );
  OAI221XLTS U1687 ( .A0(n1880), .A1(n1008), .B0(n2420), .B1(n1004), .C0(n1298), .Y(n3514) );
  OAI221XLTS U1688 ( .A0(n2329), .A1(n2120), .B0(n2424), .B1(n2108), .C0(n1197), .Y(n3608) );
  AOI22X1TS U1689 ( .A0(n1784), .A1(n738), .B0(n1934), .B1(n1263), .Y(n1197)
         );
  OAI221XLTS U1690 ( .A0(n2333), .A1(n2120), .B0(n2426), .B1(n2108), .C0(n1198), .Y(n3607) );
  AOI22X1TS U1691 ( .A0(n1781), .A1(n737), .B0(n1935), .B1(n1263), .Y(n1198)
         );
  OAI221XLTS U1692 ( .A0(n2335), .A1(n2120), .B0(n2428), .B1(n2108), .C0(n1199), .Y(n3606) );
  AOI22X1TS U1693 ( .A0(n1781), .A1(n715), .B0(n1936), .B1(n1263), .Y(n1199)
         );
  OAI221XLTS U1694 ( .A0(n2339), .A1(n2119), .B0(n2430), .B1(n2107), .C0(n1200), .Y(n3605) );
  AOI22X1TS U1695 ( .A0(n1739), .A1(n714), .B0(n1937), .B1(n1263), .Y(n1200)
         );
  OAI221XLTS U1696 ( .A0(n2342), .A1(n2119), .B0(n2432), .B1(n2107), .C0(n1201), .Y(n3604) );
  AOI22X1TS U1697 ( .A0(n1739), .A1(n713), .B0(n1938), .B1(n1137), .Y(n1201)
         );
  OAI221XLTS U1698 ( .A0(n2345), .A1(n2119), .B0(n2434), .B1(n2107), .C0(n1202), .Y(n3603) );
  AOI22X1TS U1699 ( .A0(n1739), .A1(n712), .B0(n1939), .B1(n1137), .Y(n1202)
         );
  OAI221XLTS U1700 ( .A0(n2347), .A1(n2119), .B0(n2436), .B1(n2107), .C0(n1203), .Y(n3602) );
  AOI22X1TS U1701 ( .A0(n1739), .A1(n711), .B0(n1940), .B1(n1137), .Y(n1203)
         );
  OAI221XLTS U1702 ( .A0(n2351), .A1(n2118), .B0(n2438), .B1(n2087), .C0(n1204), .Y(n3601) );
  AOI22X1TS U1703 ( .A0(n1965), .A1(n710), .B0(n1941), .B1(n1137), .Y(n1204)
         );
  OAI221XLTS U1704 ( .A0(n2354), .A1(n2118), .B0(n2440), .B1(n2087), .C0(n1205), .Y(n3600) );
  AOI22X1TS U1705 ( .A0(n1965), .A1(n709), .B0(n1942), .B1(n1136), .Y(n1205)
         );
  OAI221XLTS U1706 ( .A0(n2356), .A1(n2118), .B0(n2442), .B1(n2087), .C0(n1206), .Y(n3599) );
  AOI22X1TS U1707 ( .A0(n1782), .A1(n708), .B0(n1943), .B1(n1136), .Y(n1206)
         );
  OAI221XLTS U1708 ( .A0(n2360), .A1(n2118), .B0(n2444), .B1(n2087), .C0(n1207), .Y(n3598) );
  AOI22X1TS U1709 ( .A0(n1195), .A1(n707), .B0(n1944), .B1(n1136), .Y(n1207)
         );
  OAI221XLTS U1710 ( .A0(n2363), .A1(n2117), .B0(n2446), .B1(n2085), .C0(n1208), .Y(n3597) );
  AOI22X1TS U1711 ( .A0(n1752), .A1(n706), .B0(n1945), .B1(n1136), .Y(n1208)
         );
  OAI221XLTS U1712 ( .A0(n2365), .A1(n2117), .B0(n2448), .B1(n2085), .C0(n1209), .Y(n3596) );
  AOI22X1TS U1713 ( .A0(n1752), .A1(n705), .B0(n1946), .B1(n1057), .Y(n1209)
         );
  OAI221XLTS U1714 ( .A0(n2369), .A1(n2117), .B0(n2450), .B1(n2085), .C0(n1210), .Y(n3595) );
  AOI22X1TS U1715 ( .A0(n1752), .A1(n704), .B0(n1947), .B1(n1057), .Y(n1210)
         );
  OAI221XLTS U1716 ( .A0(n2371), .A1(n2117), .B0(n2452), .B1(n2085), .C0(n1211), .Y(n3594) );
  AOI22X1TS U1717 ( .A0(n1752), .A1(n703), .B0(n1948), .B1(n1057), .Y(n1211)
         );
  OAI221XLTS U1718 ( .A0(n2375), .A1(n2116), .B0(n2454), .B1(n1966), .C0(n1212), .Y(n3593) );
  AOI22X1TS U1719 ( .A0(n1767), .A1(n702), .B0(n1949), .B1(n1057), .Y(n1212)
         );
  OAI221XLTS U1720 ( .A0(n2378), .A1(n2116), .B0(n2456), .B1(n1966), .C0(n1213), .Y(n3592) );
  AOI22X1TS U1721 ( .A0(n1767), .A1(n701), .B0(n1950), .B1(n1056), .Y(n1213)
         );
  OAI221XLTS U1722 ( .A0(n2381), .A1(n2116), .B0(n2458), .B1(n1966), .C0(n1214), .Y(n3591) );
  AOI22X1TS U1723 ( .A0(n1767), .A1(n700), .B0(n1951), .B1(n1056), .Y(n1214)
         );
  OAI221XLTS U1724 ( .A0(n2383), .A1(n2116), .B0(n2460), .B1(n1966), .C0(n1215), .Y(n3590) );
  AOI22X1TS U1725 ( .A0(n1767), .A1(n699), .B0(n1952), .B1(n1056), .Y(n1215)
         );
  OAI221XLTS U1726 ( .A0(n2386), .A1(n2122), .B0(n2462), .B1(n2110), .C0(n1216), .Y(n3589) );
  AOI22X1TS U1727 ( .A0(n1911), .A1(n1779), .B0(n1953), .B1(n1056), .Y(n1216)
         );
  OAI221XLTS U1728 ( .A0(n2389), .A1(n2123), .B0(n2464), .B1(n2111), .C0(n1217), .Y(n3588) );
  AOI22X1TS U1729 ( .A0(n1912), .A1(n1779), .B0(n1954), .B1(n1599), .Y(n1217)
         );
  OAI221XLTS U1730 ( .A0(n2393), .A1(n1192), .B0(n2466), .B1(n1193), .C0(n1218), .Y(n3587) );
  AOI22X1TS U1731 ( .A0(n1913), .A1(n1783), .B0(n1955), .B1(n1599), .Y(n1218)
         );
  OAI221XLTS U1732 ( .A0(n2396), .A1(n1192), .B0(n2468), .B1(n1193), .C0(n1219), .Y(n3586) );
  AOI22X1TS U1733 ( .A0(n1914), .A1(n1784), .B0(n1956), .B1(n1500), .Y(n1219)
         );
  OAI221XLTS U1734 ( .A0(n2398), .A1(n2124), .B0(n2470), .B1(n2112), .C0(n1220), .Y(n3585) );
  AOI22X1TS U1735 ( .A0(n1915), .A1(n1779), .B0(n1957), .B1(n1377), .Y(n1220)
         );
  OAI221XLTS U1736 ( .A0(n2402), .A1(n2124), .B0(n2472), .B1(n2112), .C0(n1221), .Y(n3584) );
  AOI22X1TS U1737 ( .A0(n1916), .A1(n1779), .B0(n1958), .B1(n1599), .Y(n1221)
         );
  OAI221XLTS U1738 ( .A0(n2405), .A1(n2123), .B0(n2474), .B1(n2111), .C0(n1222), .Y(n3583) );
  AOI22X1TS U1739 ( .A0(n1917), .A1(n1780), .B0(n1959), .B1(n1599), .Y(n1222)
         );
  OAI221XLTS U1740 ( .A0(n2408), .A1(n2121), .B0(n2476), .B1(n2109), .C0(n1223), .Y(n3582) );
  AOI22X1TS U1741 ( .A0(n1918), .A1(n1783), .B0(n1960), .B1(n1489), .Y(n1223)
         );
  OAI221XLTS U1742 ( .A0(n2411), .A1(n2124), .B0(n2478), .B1(n2112), .C0(n1224), .Y(n3581) );
  AOI22X1TS U1743 ( .A0(n1919), .A1(n1784), .B0(n1961), .B1(n1489), .Y(n1224)
         );
  OAI221XLTS U1744 ( .A0(n2414), .A1(n2124), .B0(n2480), .B1(n2112), .C0(n1225), .Y(n3580) );
  AOI22X1TS U1745 ( .A0(n1920), .A1(n1780), .B0(n1962), .B1(n1055), .Y(n1225)
         );
  OAI221XLTS U1746 ( .A0(n2417), .A1(n2121), .B0(n2482), .B1(n2109), .C0(n1226), .Y(n3579) );
  AOI22X1TS U1747 ( .A0(n1921), .A1(n1780), .B0(n1963), .B1(n1055), .Y(n1226)
         );
  OAI221XLTS U1748 ( .A0(n2420), .A1(n2122), .B0(n2484), .B1(n2110), .C0(n1227), .Y(n3578) );
  AOI22X1TS U1749 ( .A0(n1922), .A1(n1780), .B0(n1964), .B1(n1055), .Y(n1227)
         );
  OAI221XLTS U1750 ( .A0(n2280), .A1(n380), .B0(n604), .B1(n934), .C0(n1557), 
        .Y(n3293) );
  AOI22X1TS U1751 ( .A0(n2295), .A1(n583), .B0(n569), .B1(n698), .Y(n1557) );
  OAI221XLTS U1752 ( .A0(n2282), .A1(n380), .B0(n601), .B1(n942), .C0(n1558), 
        .Y(n3292) );
  AOI22X1TS U1753 ( .A0(n2298), .A1(n583), .B0(n569), .B1(n697), .Y(n1558) );
  OAI221XLTS U1754 ( .A0(n2284), .A1(n380), .B0(n1373), .B1(n941), .C0(n1559), 
        .Y(n3291) );
  AOI22X1TS U1755 ( .A0(n2301), .A1(n583), .B0(n569), .B1(n696), .Y(n1559) );
  OAI221XLTS U1756 ( .A0(n2286), .A1(n380), .B0(n601), .B1(n945), .C0(n1560), 
        .Y(n3290) );
  AOI22X1TS U1757 ( .A0(n2304), .A1(n583), .B0(n567), .B1(n695), .Y(n1560) );
  OAI221XLTS U1758 ( .A0(n2288), .A1(n381), .B0(n603), .B1(n940), .C0(n1561), 
        .Y(n3289) );
  AOI22X1TS U1759 ( .A0(n2307), .A1(n582), .B0(n571), .B1(n694), .Y(n1561) );
  OAI221XLTS U1760 ( .A0(n2290), .A1(n381), .B0(n603), .B1(n944), .C0(n1562), 
        .Y(n3288) );
  AOI22X1TS U1761 ( .A0(n2310), .A1(n582), .B0(n571), .B1(n693), .Y(n1562) );
  OAI221XLTS U1762 ( .A0(n2292), .A1(n381), .B0(n1373), .B1(n939), .C0(n1563), 
        .Y(n3287) );
  AOI22X1TS U1763 ( .A0(n2313), .A1(n582), .B0(n570), .B1(n692), .Y(n1563) );
  OAI221XLTS U1764 ( .A0(n2294), .A1(n381), .B0(n604), .B1(n943), .C0(n1564), 
        .Y(n3286) );
  AOI22X1TS U1765 ( .A0(n2316), .A1(n582), .B0(n569), .B1(n691), .Y(n1564) );
  OAI221XLTS U1766 ( .A0(n2065), .A1(n687), .B0(n642), .B1(n2297), .C0(n1545), 
        .Y(n3301) );
  AOI22X1TS U1767 ( .A0(n2279), .A1(n624), .B0(n616), .B1(n682), .Y(n1545) );
  OAI221XLTS U1768 ( .A0(n2067), .A1(n686), .B0(n642), .B1(n2300), .C0(n1546), 
        .Y(n3300) );
  AOI22X1TS U1769 ( .A0(n2281), .A1(n624), .B0(n616), .B1(n681), .Y(n1546) );
  OAI221XLTS U1770 ( .A0(n2069), .A1(n687), .B0(n643), .B1(n2303), .C0(n1547), 
        .Y(n3299) );
  AOI22X1TS U1771 ( .A0(n2283), .A1(n624), .B0(n616), .B1(n680), .Y(n1547) );
  OAI221XLTS U1772 ( .A0(n2071), .A1(n684), .B0(n1338), .B1(n2305), .C0(n1548), 
        .Y(n3298) );
  AOI22X1TS U1773 ( .A0(n2285), .A1(n624), .B0(n615), .B1(n679), .Y(n1548) );
  OAI221XLTS U1774 ( .A0(n2073), .A1(n687), .B0(n639), .B1(n2309), .C0(n1549), 
        .Y(n3297) );
  AOI22X1TS U1775 ( .A0(n2287), .A1(n625), .B0(n615), .B1(n678), .Y(n1549) );
  OAI221XLTS U1776 ( .A0(n2075), .A1(n1337), .B0(n640), .B1(n2311), .C0(n1550), 
        .Y(n3296) );
  AOI22X1TS U1777 ( .A0(n2289), .A1(n625), .B0(n615), .B1(n677), .Y(n1550) );
  OAI221XLTS U1778 ( .A0(n2077), .A1(n686), .B0(n643), .B1(n2315), .C0(n1551), 
        .Y(n3295) );
  AOI22X1TS U1779 ( .A0(n2291), .A1(n625), .B0(n615), .B1(n676), .Y(n1551) );
  OAI221XLTS U1780 ( .A0(n2079), .A1(n1337), .B0(n1338), .B1(n2318), .C0(n1552), .Y(n3294) );
  AOI22X1TS U1781 ( .A0(n2293), .A1(n625), .B0(n618), .B1(n675), .Y(n1552) );
  OAI221XLTS U1782 ( .A0(n2125), .A1(n2296), .B0(n2113), .B1(n2280), .C0(n1491), .Y(n3333) );
  AOI22X1TS U1783 ( .A0(n1777), .A1(n17), .B0(n1925), .B1(n1055), .Y(n1491) );
  OAI221XLTS U1784 ( .A0(n2125), .A1(n2299), .B0(n2113), .B1(n2282), .C0(n1492), .Y(n3332) );
  AOI22X1TS U1785 ( .A0(n1778), .A1(n18), .B0(n1926), .B1(n1054), .Y(n1492) );
  OAI221XLTS U1786 ( .A0(n2126), .A1(n2302), .B0(n2114), .B1(n2284), .C0(n1493), .Y(n3331) );
  AOI22X1TS U1787 ( .A0(n1778), .A1(n19), .B0(n1927), .B1(n1054), .Y(n1493) );
  OAI221XLTS U1788 ( .A0(n2123), .A1(n2306), .B0(n2111), .B1(n2286), .C0(n1494), .Y(n3330) );
  AOI22X1TS U1789 ( .A0(n1777), .A1(n20), .B0(n1928), .B1(n1054), .Y(n1494) );
  OAI221XLTS U1790 ( .A0(n2125), .A1(n2308), .B0(n2113), .B1(n2288), .C0(n1495), .Y(n3329) );
  AOI22X1TS U1791 ( .A0(n1778), .A1(n21), .B0(n1929), .B1(n1054), .Y(n1495) );
  OAI221XLTS U1792 ( .A0(n2127), .A1(n2312), .B0(n2115), .B1(n2290), .C0(n1496), .Y(n3328) );
  AOI22X1TS U1793 ( .A0(n1778), .A1(n22), .B0(n1930), .B1(n1500), .Y(n1496) );
  OAI221XLTS U1794 ( .A0(n2125), .A1(n2314), .B0(n2113), .B1(n2292), .C0(n1497), .Y(n3327) );
  AOI22X1TS U1795 ( .A0(n1777), .A1(n23), .B0(n1931), .B1(n1607), .Y(n1497) );
  OAI221XLTS U1796 ( .A0(n2127), .A1(n2317), .B0(n2115), .B1(n2294), .C0(n1498), .Y(n3326) );
  AOI22X1TS U1797 ( .A0(n1782), .A1(n24), .B0(n1932), .B1(n1607), .Y(n1498) );
  OAI221XLTS U1798 ( .A0(n904), .A1(n600), .B0(n2326), .B1(n590), .C0(n1375), 
        .Y(n3449) );
  AOI2BB2X1TS U1799 ( .B0(n578), .B1(dataIn_EAST[0]), .A0N(n566), .A1N(n1810), 
        .Y(n1375) );
  OAI221XLTS U1800 ( .A0(n929), .A1(n600), .B0(n2330), .B1(n590), .C0(n1378), 
        .Y(n3448) );
  AOI2BB2X1TS U1801 ( .B0(n578), .B1(dataIn_EAST[1]), .A0N(n566), .A1N(n1811), 
        .Y(n1378) );
  OAI221XLTS U1802 ( .A0(n928), .A1(n600), .B0(n2332), .B1(n591), .C0(n1379), 
        .Y(n3447) );
  AOI2BB2X1TS U1803 ( .B0(n578), .B1(dataIn_EAST[2]), .A0N(n566), .A1N(n1812), 
        .Y(n1379) );
  OAI221XLTS U1804 ( .A0(n927), .A1(n600), .B0(n2336), .B1(n593), .C0(n1380), 
        .Y(n3446) );
  AOI2BB2X1TS U1805 ( .B0(n578), .B1(dataIn_EAST[3]), .A0N(n566), .A1N(n1813), 
        .Y(n1380) );
  OAI221XLTS U1806 ( .A0(n903), .A1(n599), .B0(n2338), .B1(n593), .C0(n1381), 
        .Y(n3445) );
  AOI2BB2X1TS U1807 ( .B0(n577), .B1(dataIn_EAST[4]), .A0N(n565), .A1N(n1815), 
        .Y(n1381) );
  OAI221XLTS U1808 ( .A0(n926), .A1(n599), .B0(n2341), .B1(n1374), .C0(n1382), 
        .Y(n3444) );
  AOI2BB2X1TS U1809 ( .B0(n577), .B1(dataIn_EAST[5]), .A0N(n565), .A1N(n1816), 
        .Y(n1382) );
  OAI221XLTS U1810 ( .A0(n925), .A1(n599), .B0(n2344), .B1(n590), .C0(n1383), 
        .Y(n3443) );
  AOI2BB2X1TS U1811 ( .B0(n577), .B1(dataIn_EAST[6]), .A0N(n565), .A1N(n1817), 
        .Y(n1383) );
  OAI221XLTS U1812 ( .A0(n924), .A1(n599), .B0(n2348), .B1(n590), .C0(n1384), 
        .Y(n3442) );
  AOI2BB2X1TS U1813 ( .B0(n577), .B1(dataIn_EAST[7]), .A0N(n565), .A1N(n1818), 
        .Y(n1384) );
  OAI221XLTS U1814 ( .A0(n902), .A1(n598), .B0(n2350), .B1(n591), .C0(n1385), 
        .Y(n3441) );
  AOI2BB2X1TS U1815 ( .B0(n576), .B1(dataIn_EAST[8]), .A0N(n564), .A1N(n1820), 
        .Y(n1385) );
  OAI221XLTS U1816 ( .A0(n923), .A1(n598), .B0(n2353), .B1(n593), .C0(n1386), 
        .Y(n3440) );
  AOI2BB2X1TS U1817 ( .B0(n576), .B1(dataIn_EAST[9]), .A0N(n564), .A1N(n1821), 
        .Y(n1386) );
  OAI221XLTS U1818 ( .A0(n922), .A1(n598), .B0(n2357), .B1(n589), .C0(n1387), 
        .Y(n3439) );
  AOI2BB2X1TS U1819 ( .B0(n576), .B1(dataIn_EAST[10]), .A0N(n564), .A1N(n1822), 
        .Y(n1387) );
  OAI221XLTS U1820 ( .A0(n921), .A1(n598), .B0(n2359), .B1(n589), .C0(n1388), 
        .Y(n3438) );
  AOI2BB2X1TS U1821 ( .B0(n576), .B1(dataIn_EAST[11]), .A0N(n564), .A1N(n1823), 
        .Y(n1388) );
  OAI221XLTS U1822 ( .A0(n901), .A1(n597), .B0(n2362), .B1(n589), .C0(n1389), 
        .Y(n3437) );
  AOI2BB2X1TS U1823 ( .B0(n575), .B1(dataIn_EAST[12]), .A0N(n563), .A1N(n1825), 
        .Y(n1389) );
  OAI221XLTS U1824 ( .A0(n920), .A1(n597), .B0(n2366), .B1(n589), .C0(n1390), 
        .Y(n3436) );
  AOI2BB2X1TS U1825 ( .B0(n575), .B1(dataIn_EAST[13]), .A0N(n563), .A1N(n1826), 
        .Y(n1390) );
  OAI221XLTS U1826 ( .A0(n919), .A1(n597), .B0(n2368), .B1(n588), .C0(n1391), 
        .Y(n3435) );
  AOI2BB2X1TS U1827 ( .B0(n575), .B1(dataIn_EAST[14]), .A0N(n563), .A1N(n1827), 
        .Y(n1391) );
  OAI221XLTS U1828 ( .A0(n918), .A1(n597), .B0(n2372), .B1(n588), .C0(n1392), 
        .Y(n3434) );
  AOI2BB2X1TS U1829 ( .B0(n575), .B1(dataIn_EAST[15]), .A0N(n563), .A1N(n1828), 
        .Y(n1392) );
  OAI221XLTS U1830 ( .A0(n900), .A1(n602), .B0(n2374), .B1(n588), .C0(n1393), 
        .Y(n3433) );
  AOI2BB2X1TS U1831 ( .B0(n580), .B1(dataIn_EAST[16]), .A0N(n562), .A1N(n1830), 
        .Y(n1393) );
  OAI221XLTS U1832 ( .A0(n917), .A1(n605), .B0(n2377), .B1(n588), .C0(n1394), 
        .Y(n3432) );
  AOI2BB2X1TS U1833 ( .B0(n581), .B1(dataIn_EAST[17]), .A0N(n562), .A1N(n1831), 
        .Y(n1394) );
  OAI221XLTS U1834 ( .A0(n916), .A1(n604), .B0(n2380), .B1(n587), .C0(n1395), 
        .Y(n3431) );
  AOI2BB2X1TS U1835 ( .B0(n579), .B1(dataIn_EAST[18]), .A0N(n562), .A1N(n1832), 
        .Y(n1395) );
  OAI221XLTS U1836 ( .A0(n915), .A1(n605), .B0(n2384), .B1(n587), .C0(n1396), 
        .Y(n3430) );
  AOI2BB2X1TS U1837 ( .B0(n579), .B1(dataIn_EAST[19]), .A0N(n562), .A1N(n1833), 
        .Y(n1396) );
  OAI221XLTS U1838 ( .A0(n914), .A1(n596), .B0(n2387), .B1(n587), .C0(n1397), 
        .Y(n3429) );
  AOI2BB2X1TS U1839 ( .B0(n574), .B1(dataIn_EAST[20]), .A0N(n561), .A1N(n1835), 
        .Y(n1397) );
  OAI221XLTS U1840 ( .A0(n899), .A1(n596), .B0(n2390), .B1(n587), .C0(n1398), 
        .Y(n3428) );
  AOI2BB2X1TS U1841 ( .B0(n574), .B1(dataIn_EAST[21]), .A0N(n561), .A1N(n1836), 
        .Y(n1398) );
  OAI221XLTS U1842 ( .A0(n913), .A1(n596), .B0(n2392), .B1(n586), .C0(n1399), 
        .Y(n3427) );
  AOI2BB2X1TS U1843 ( .B0(n574), .B1(dataIn_EAST[22]), .A0N(n561), .A1N(n1837), 
        .Y(n1399) );
  OAI221XLTS U1844 ( .A0(n912), .A1(n596), .B0(n2395), .B1(n586), .C0(n1400), 
        .Y(n3426) );
  AOI2BB2X1TS U1845 ( .B0(n574), .B1(dataIn_EAST[23]), .A0N(n561), .A1N(n1838), 
        .Y(n1400) );
  OAI221XLTS U1846 ( .A0(n898), .A1(n595), .B0(n2399), .B1(n586), .C0(n1401), 
        .Y(n3425) );
  AOI2BB2X1TS U1847 ( .B0(n573), .B1(dataIn_EAST[24]), .A0N(n560), .A1N(n1840), 
        .Y(n1401) );
  OAI221XLTS U1848 ( .A0(n911), .A1(n595), .B0(n2401), .B1(n586), .C0(n1402), 
        .Y(n3424) );
  AOI2BB2X1TS U1849 ( .B0(n573), .B1(dataIn_EAST[25]), .A0N(n560), .A1N(n1841), 
        .Y(n1402) );
  OAI221XLTS U1850 ( .A0(n909), .A1(n595), .B0(n2404), .B1(n585), .C0(n1403), 
        .Y(n3423) );
  AOI2BB2X1TS U1851 ( .B0(n573), .B1(dataIn_EAST[26]), .A0N(n560), .A1N(n1842), 
        .Y(n1403) );
  OAI221XLTS U1852 ( .A0(n908), .A1(n595), .B0(n2407), .B1(n585), .C0(n1404), 
        .Y(n3422) );
  AOI2BB2X1TS U1853 ( .B0(n573), .B1(dataIn_EAST[27]), .A0N(n560), .A1N(n1843), 
        .Y(n1404) );
  OAI221XLTS U1854 ( .A0(n907), .A1(n594), .B0(n2410), .B1(n585), .C0(n1405), 
        .Y(n3421) );
  AOI2BB2X1TS U1855 ( .B0(n572), .B1(dataIn_EAST[28]), .A0N(n559), .A1N(n1845), 
        .Y(n1405) );
  OAI221XLTS U1856 ( .A0(n906), .A1(n594), .B0(n2413), .B1(n584), .C0(n1406), 
        .Y(n3420) );
  AOI2BB2X1TS U1857 ( .B0(n572), .B1(dataIn_EAST[29]), .A0N(n559), .A1N(n1846), 
        .Y(n1406) );
  OAI221XLTS U1858 ( .A0(n905), .A1(n594), .B0(n2416), .B1(n584), .C0(n1407), 
        .Y(n3419) );
  AOI2BB2X1TS U1859 ( .B0(n572), .B1(dataIn_EAST[30]), .A0N(n559), .A1N(n1847), 
        .Y(n1407) );
  OAI221XLTS U1860 ( .A0(n897), .A1(n594), .B0(n2419), .B1(n584), .C0(n1408), 
        .Y(n3418) );
  AOI2BB2X1TS U1861 ( .B0(n572), .B1(dataIn_EAST[31]), .A0N(n559), .A1N(n1848), 
        .Y(n1408) );
  OAI221XLTS U1862 ( .A0(n2007), .A1(n683), .B0(n2326), .B1(n638), .C0(n1339), 
        .Y(n3481) );
  AOI2BB2X1TS U1863 ( .B0(n629), .B1(n2421), .A0N(n613), .A1N(n1849), .Y(n1339) );
  OAI221XLTS U1864 ( .A0(n2008), .A1(n683), .B0(n2330), .B1(n638), .C0(n1342), 
        .Y(n3480) );
  AOI2BB2X1TS U1865 ( .B0(n629), .B1(n2423), .A0N(n613), .A1N(n1850), .Y(n1342) );
  OAI221XLTS U1866 ( .A0(n2009), .A1(n683), .B0(n2332), .B1(n638), .C0(n1343), 
        .Y(n3479) );
  AOI2BB2X1TS U1867 ( .B0(n626), .B1(n2425), .A0N(n613), .A1N(n1851), .Y(n1343) );
  OAI221XLTS U1868 ( .A0(n2010), .A1(n683), .B0(n2336), .B1(n638), .C0(n1344), 
        .Y(n3478) );
  AOI2BB2X1TS U1869 ( .B0(n631), .B1(n2427), .A0N(n613), .A1N(n1852), .Y(n1344) );
  OAI221XLTS U1870 ( .A0(n2011), .A1(n649), .B0(n2338), .B1(n637), .C0(n1345), 
        .Y(n3477) );
  AOI2BB2X1TS U1871 ( .B0(n629), .B1(n2429), .A0N(n612), .A1N(n1853), .Y(n1345) );
  OAI221XLTS U1872 ( .A0(n2012), .A1(n649), .B0(n2341), .B1(n637), .C0(n1346), 
        .Y(n3476) );
  AOI2BB2X1TS U1873 ( .B0(n629), .B1(n2431), .A0N(n612), .A1N(n1854), .Y(n1346) );
  OAI221XLTS U1874 ( .A0(n2013), .A1(n649), .B0(n2344), .B1(n637), .C0(n1347), 
        .Y(n3475) );
  AOI2BB2X1TS U1875 ( .B0(n630), .B1(n2433), .A0N(n612), .A1N(n1855), .Y(n1347) );
  OAI221XLTS U1876 ( .A0(n2015), .A1(n649), .B0(n2348), .B1(n637), .C0(n1348), 
        .Y(n3474) );
  AOI2BB2X1TS U1877 ( .B0(n627), .B1(n2435), .A0N(n612), .A1N(n1856), .Y(n1348) );
  OAI221XLTS U1878 ( .A0(n2017), .A1(n648), .B0(n2350), .B1(n636), .C0(n1349), 
        .Y(n3473) );
  AOI2BB2X1TS U1879 ( .B0(n628), .B1(n2437), .A0N(n611), .A1N(n1857), .Y(n1349) );
  OAI221XLTS U1880 ( .A0(n2019), .A1(n648), .B0(n2353), .B1(n636), .C0(n1350), 
        .Y(n3472) );
  AOI2BB2X1TS U1881 ( .B0(n628), .B1(n2439), .A0N(n611), .A1N(n1858), .Y(n1350) );
  OAI221XLTS U1882 ( .A0(n2021), .A1(n648), .B0(n2357), .B1(n636), .C0(n1351), 
        .Y(n3471) );
  AOI2BB2X1TS U1883 ( .B0(n628), .B1(n2441), .A0N(n611), .A1N(n1859), .Y(n1351) );
  OAI221XLTS U1884 ( .A0(n2023), .A1(n648), .B0(n2359), .B1(n636), .C0(n1352), 
        .Y(n3470) );
  AOI2BB2X1TS U1885 ( .B0(n626), .B1(n2443), .A0N(n611), .A1N(n1860), .Y(n1352) );
  OAI221XLTS U1886 ( .A0(n2025), .A1(n647), .B0(n2362), .B1(n635), .C0(n1353), 
        .Y(n3469) );
  AOI2BB2X1TS U1887 ( .B0(n627), .B1(n2445), .A0N(n610), .A1N(n1861), .Y(n1353) );
  OAI221XLTS U1888 ( .A0(n2029), .A1(n647), .B0(n2368), .B1(n635), .C0(n1355), 
        .Y(n3467) );
  AOI2BB2X1TS U1889 ( .B0(n628), .B1(n2449), .A0N(n610), .A1N(n1863), .Y(n1355) );
  OAI221XLTS U1890 ( .A0(n2031), .A1(n647), .B0(n2372), .B1(n635), .C0(n1356), 
        .Y(n3466) );
  AOI2BB2X1TS U1891 ( .B0(n1340), .B1(n2451), .A0N(n610), .A1N(n1864), .Y(
        n1356) );
  OAI221XLTS U1892 ( .A0(n2033), .A1(n688), .B0(n2374), .B1(n634), .C0(n1357), 
        .Y(n3465) );
  AOI2BB2X1TS U1893 ( .B0(n620), .B1(n2453), .A0N(n609), .A1N(n1865), .Y(n1357) );
  OAI221XLTS U1894 ( .A0(n2035), .A1(n685), .B0(n2377), .B1(n634), .C0(n1358), 
        .Y(n3464) );
  AOI2BB2X1TS U1895 ( .B0(n620), .B1(n2455), .A0N(n609), .A1N(n1866), .Y(n1358) );
  OAI221XLTS U1896 ( .A0(n2039), .A1(n688), .B0(n2384), .B1(n634), .C0(n1360), 
        .Y(n3462) );
  AOI2BB2X1TS U1897 ( .B0(n620), .B1(n2459), .A0N(n609), .A1N(n1868), .Y(n1360) );
  OAI221XLTS U1898 ( .A0(n2041), .A1(n646), .B0(n2387), .B1(n633), .C0(n1361), 
        .Y(n3461) );
  AOI2BB2X1TS U1899 ( .B0(n621), .B1(n2461), .A0N(n608), .A1N(n1869), .Y(n1361) );
  OAI221XLTS U1900 ( .A0(n2043), .A1(n646), .B0(n2390), .B1(n633), .C0(n1362), 
        .Y(n3460) );
  AOI2BB2X1TS U1901 ( .B0(n621), .B1(n2463), .A0N(n608), .A1N(n1870), .Y(n1362) );
  OAI221XLTS U1902 ( .A0(n2045), .A1(n646), .B0(n2392), .B1(n633), .C0(n1363), 
        .Y(n3459) );
  AOI2BB2X1TS U1903 ( .B0(n621), .B1(n2465), .A0N(n608), .A1N(n1871), .Y(n1363) );
  OAI221XLTS U1904 ( .A0(n2047), .A1(n646), .B0(n2395), .B1(n633), .C0(n1364), 
        .Y(n3458) );
  AOI2BB2X1TS U1905 ( .B0(n621), .B1(n2467), .A0N(n608), .A1N(n1872), .Y(n1364) );
  OAI221XLTS U1906 ( .A0(n2049), .A1(n645), .B0(n2399), .B1(n632), .C0(n1365), 
        .Y(n3457) );
  AOI2BB2X1TS U1907 ( .B0(n622), .B1(n2469), .A0N(n607), .A1N(n1873), .Y(n1365) );
  OAI221XLTS U1908 ( .A0(n2051), .A1(n645), .B0(n2401), .B1(n632), .C0(n1366), 
        .Y(n3456) );
  AOI2BB2X1TS U1909 ( .B0(n622), .B1(n2471), .A0N(n607), .A1N(n1874), .Y(n1366) );
  OAI221XLTS U1910 ( .A0(n2053), .A1(n645), .B0(n2404), .B1(n632), .C0(n1367), 
        .Y(n3455) );
  AOI2BB2X1TS U1911 ( .B0(n622), .B1(n2473), .A0N(n607), .A1N(n1875), .Y(n1367) );
  OAI221XLTS U1912 ( .A0(n2055), .A1(n645), .B0(n2407), .B1(n632), .C0(n1368), 
        .Y(n3454) );
  AOI2BB2X1TS U1913 ( .B0(n622), .B1(n2475), .A0N(n607), .A1N(n1876), .Y(n1368) );
  OAI221XLTS U1914 ( .A0(n2057), .A1(n644), .B0(n2410), .B1(n641), .C0(n1369), 
        .Y(n3453) );
  AOI2BB2X1TS U1915 ( .B0(n623), .B1(n2477), .A0N(n606), .A1N(n1877), .Y(n1369) );
  OAI221XLTS U1916 ( .A0(n2059), .A1(n644), .B0(n2413), .B1(n641), .C0(n1370), 
        .Y(n3452) );
  AOI2BB2X1TS U1917 ( .B0(n623), .B1(n2479), .A0N(n606), .A1N(n1878), .Y(n1370) );
  OAI221XLTS U1918 ( .A0(n2061), .A1(n644), .B0(n2416), .B1(n640), .C0(n1371), 
        .Y(n3451) );
  AOI2BB2X1TS U1919 ( .B0(n623), .B1(n2481), .A0N(n606), .A1N(n1879), .Y(n1371) );
  OAI221XLTS U1920 ( .A0(n2063), .A1(n644), .B0(n2419), .B1(n639), .C0(n1372), 
        .Y(n3450) );
  AOI2BB2X1TS U1921 ( .B0(n623), .B1(n2483), .A0N(n606), .A1N(n1880), .Y(n1372) );
  OAI221XLTS U1922 ( .A0(n2327), .A1(n2120), .B0(n2422), .B1(n2108), .C0(n1194), .Y(n3609) );
  AOI22X1TS U1923 ( .A0(n1777), .A1(n739), .B0(n1933), .B1(n1377), .Y(n1194)
         );
  OAI221XLTS U1924 ( .A0(n2027), .A1(n647), .B0(n2366), .B1(n635), .C0(n1354), 
        .Y(n3468) );
  AOI2BB2X1TS U1925 ( .B0(n1340), .B1(n2447), .A0N(n610), .A1N(n1862), .Y(
        n1354) );
  OAI221XLTS U1926 ( .A0(n2037), .A1(n684), .B0(n2380), .B1(n634), .C0(n1359), 
        .Y(n3463) );
  AOI2BB2X1TS U1927 ( .B0(n620), .B1(n2457), .A0N(n609), .A1N(n1867), .Y(n1359) );
  INVX2TS U1928 ( .A(memWrite_EAST), .Y(n977) );
  OAI211X1TS U1929 ( .A0(n960), .A1(n1151), .B0(n1152), .C0(n1153), .Y(n1149)
         );
  OAI2BB1X1TS U1930 ( .A0N(n1151), .A1N(n960), .B0(n910), .Y(n1152) );
  INVX2TS U1931 ( .A(memRead_WEST), .Y(n1024) );
  OAI22X1TS U1932 ( .A0(n2095), .A1(n509), .B0(n521), .B1(n1726), .Y(n3184) );
  AOI221X1TS U1933 ( .A0(n96), .A1(n933), .B0(n92), .B1(n1140), .C0(n2493), 
        .Y(n1726) );
  OAI22X1TS U1934 ( .A0(n2097), .A1(n2232), .B0(n1678), .B1(n1679), .Y(n3217)
         );
  AOI221X1TS U1935 ( .A0(n95), .A1(n946), .B0(n93), .B1(n1462), .C0(n2493), 
        .Y(n1679) );
  OAI22X1TS U1936 ( .A0(n45), .A1(n742), .B0(n1467), .B1(n1468), .Y(n3343) );
  INVX2TS U1937 ( .A(n1467), .Y(n742) );
  AOI32X1TS U1938 ( .A0(n2160), .A1(n1469), .A2(n379), .B0(n1470), .B1(n2501), 
        .Y(n1468) );
  NOR4BX1TS U1939 ( .AN(n1474), .B(n1472), .C(n2488), .D(n1475), .Y(n1467) );
  OAI211X1TS U1940 ( .A0(n1999), .A1(n515), .B0(n1627), .C0(n1628), .Y(n3242)
         );
  AOI222XLTS U1941 ( .A0(n500), .A1(dataIn_EAST[24]), .B0(n488), .B1(
        dataIn_SOUTH[24]), .C0(n483), .C1(n2397), .Y(n1628) );
  AOI22X1TS U1942 ( .A0(dataIn_NORTH[24]), .A1(n465), .B0(n790), .B1(n2155), 
        .Y(n1627) );
  OAI211X1TS U1943 ( .A0(n2000), .A1(n515), .B0(n1625), .C0(n1626), .Y(n3243)
         );
  AOI222XLTS U1944 ( .A0(n500), .A1(dataIn_EAST[25]), .B0(n488), .B1(
        dataIn_SOUTH[25]), .C0(n482), .C1(n2400), .Y(n1626) );
  AOI22X1TS U1945 ( .A0(dataIn_NORTH[25]), .A1(n465), .B0(n789), .B1(n2155), 
        .Y(n1625) );
  OAI211X1TS U1946 ( .A0(n2001), .A1(n515), .B0(n1623), .C0(n1624), .Y(n3244)
         );
  AOI222XLTS U1947 ( .A0(n500), .A1(dataIn_EAST[26]), .B0(n488), .B1(
        dataIn_SOUTH[26]), .C0(n483), .C1(n2403), .Y(n1624) );
  AOI22X1TS U1948 ( .A0(dataIn_NORTH[26]), .A1(n465), .B0(n788), .B1(n2155), 
        .Y(n1623) );
  OAI211X1TS U1949 ( .A0(n2002), .A1(n516), .B0(n1621), .C0(n1622), .Y(n3245)
         );
  AOI222XLTS U1950 ( .A0(n500), .A1(dataIn_EAST[27]), .B0(n488), .B1(
        dataIn_SOUTH[27]), .C0(n482), .C1(n2406), .Y(n1622) );
  AOI22X1TS U1951 ( .A0(dataIn_NORTH[27]), .A1(n465), .B0(n787), .B1(n2156), 
        .Y(n1621) );
  OAI211X1TS U1952 ( .A0(n2003), .A1(n516), .B0(n1619), .C0(n1620), .Y(n3246)
         );
  AOI222XLTS U1953 ( .A0(n501), .A1(dataIn_EAST[28]), .B0(n487), .B1(
        dataIn_SOUTH[28]), .C0(n477), .C1(n2409), .Y(n1620) );
  AOI22X1TS U1954 ( .A0(dataIn_NORTH[28]), .A1(n466), .B0(n786), .B1(n2158), 
        .Y(n1619) );
  OAI211X1TS U1955 ( .A0(n2004), .A1(n516), .B0(n1617), .C0(n1618), .Y(n3247)
         );
  AOI222XLTS U1956 ( .A0(n501), .A1(dataIn_EAST[29]), .B0(n487), .B1(
        dataIn_SOUTH[29]), .C0(n477), .C1(n2412), .Y(n1618) );
  AOI22X1TS U1957 ( .A0(dataIn_NORTH[29]), .A1(n466), .B0(n785), .B1(n2158), 
        .Y(n1617) );
  OAI211X1TS U1958 ( .A0(n2005), .A1(n516), .B0(n1615), .C0(n1616), .Y(n3248)
         );
  AOI222XLTS U1959 ( .A0(n501), .A1(dataIn_EAST[30]), .B0(n487), .B1(
        dataIn_SOUTH[30]), .C0(n477), .C1(n2415), .Y(n1616) );
  AOI22X1TS U1960 ( .A0(dataIn_NORTH[30]), .A1(n466), .B0(n784), .B1(n2158), 
        .Y(n1615) );
  OAI211X1TS U1961 ( .A0(n2006), .A1(n517), .B0(n1613), .C0(n1614), .Y(n3249)
         );
  AOI222XLTS U1962 ( .A0(n501), .A1(dataIn_EAST[31]), .B0(n487), .B1(
        dataIn_SOUTH[31]), .C0(n477), .C1(n2418), .Y(n1614) );
  AOI22X1TS U1963 ( .A0(dataIn_NORTH[31]), .A1(n466), .B0(n783), .B1(n2159), 
        .Y(n1613) );
  OAI211X1TS U1964 ( .A0(n1967), .A1(n517), .B0(n1593), .C0(n1594), .Y(n3270)
         );
  AOI222XLTS U1965 ( .A0(n502), .A1(cacheAddressIn_EAST[0]), .B0(
        cacheAddressIn_SOUTH[0]), .B1(n486), .C0(n478), .C1(n2295), .Y(n1594)
         );
  AOI22X1TS U1966 ( .A0(cacheAddressIn_NORTH[0]), .A1(n467), .B0(n782), .B1(
        n2157), .Y(n1593) );
  OAI211X1TS U1967 ( .A0(n1968), .A1(n517), .B0(n1591), .C0(n1592), .Y(n3271)
         );
  AOI222XLTS U1968 ( .A0(n502), .A1(cacheAddressIn_EAST[1]), .B0(
        cacheAddressIn_SOUTH[1]), .B1(n486), .C0(n478), .C1(n2298), .Y(n1592)
         );
  AOI22X1TS U1969 ( .A0(cacheAddressIn_NORTH[1]), .A1(n467), .B0(n781), .B1(
        n2157), .Y(n1591) );
  OAI211X1TS U1970 ( .A0(n1969), .A1(n517), .B0(n1589), .C0(n1590), .Y(n3272)
         );
  AOI222XLTS U1971 ( .A0(n502), .A1(cacheAddressIn_EAST[2]), .B0(
        cacheAddressIn_SOUTH[2]), .B1(n486), .C0(n478), .C1(n2301), .Y(n1590)
         );
  AOI22X1TS U1972 ( .A0(cacheAddressIn_NORTH[2]), .A1(n467), .B0(n780), .B1(
        n2157), .Y(n1589) );
  OAI211X1TS U1973 ( .A0(n1970), .A1(n518), .B0(n1587), .C0(n1588), .Y(n3273)
         );
  AOI222XLTS U1974 ( .A0(n502), .A1(cacheAddressIn_EAST[3]), .B0(
        cacheAddressIn_SOUTH[3]), .B1(n486), .C0(n478), .C1(n2304), .Y(n1588)
         );
  AOI22X1TS U1975 ( .A0(cacheAddressIn_NORTH[3]), .A1(n467), .B0(n779), .B1(
        n2158), .Y(n1587) );
  OAI211X1TS U1976 ( .A0(n1971), .A1(n518), .B0(n1585), .C0(n1586), .Y(n3274)
         );
  AOI222XLTS U1977 ( .A0(n503), .A1(cacheAddressIn_EAST[4]), .B0(
        cacheAddressIn_SOUTH[4]), .B1(n485), .C0(n479), .C1(n2307), .Y(n1586)
         );
  AOI22X1TS U1978 ( .A0(cacheAddressIn_NORTH[4]), .A1(n468), .B0(n778), .B1(
        n2159), .Y(n1585) );
  OAI211X1TS U1979 ( .A0(n1972), .A1(n518), .B0(n1583), .C0(n1584), .Y(n3275)
         );
  AOI222XLTS U1980 ( .A0(n503), .A1(cacheAddressIn_EAST[5]), .B0(
        cacheAddressIn_SOUTH[5]), .B1(n485), .C0(n479), .C1(n2310), .Y(n1584)
         );
  AOI22X1TS U1981 ( .A0(cacheAddressIn_NORTH[5]), .A1(n468), .B0(n777), .B1(
        n2159), .Y(n1583) );
  OAI211X1TS U1982 ( .A0(n1973), .A1(n518), .B0(n1581), .C0(n1582), .Y(n3276)
         );
  AOI222XLTS U1983 ( .A0(n503), .A1(cacheAddressIn_EAST[6]), .B0(
        cacheAddressIn_SOUTH[6]), .B1(n485), .C0(n479), .C1(n2313), .Y(n1582)
         );
  AOI22X1TS U1984 ( .A0(cacheAddressIn_NORTH[6]), .A1(n468), .B0(n776), .B1(
        n2159), .Y(n1581) );
  OAI211X1TS U1985 ( .A0(n1974), .A1(n1574), .B0(n1575), .C0(n1576), .Y(n3277)
         );
  AOI222XLTS U1986 ( .A0(n503), .A1(cacheAddressIn_EAST[7]), .B0(
        cacheAddressIn_SOUTH[7]), .B1(n485), .C0(n479), .C1(n2316), .Y(n1576)
         );
  AOI22X1TS U1987 ( .A0(cacheAddressIn_NORTH[7]), .A1(n468), .B0(n775), .B1(
        n2150), .Y(n1575) );
  OAI211X1TS U1988 ( .A0(n41), .A1(n82), .B0(n801), .C0(n1611), .Y(n3250) );
  AOI22X1TS U1989 ( .A0(n364), .A1(\requesterPortBuffer[0][0] ), .B0(n740), 
        .B1(n805), .Y(n1611) );
  OAI221XLTS U1990 ( .A0(n2180), .A1(n667), .B0(n2014), .B1(n2233), .C0(n1689), 
        .Y(n3209) );
  AOI222XLTS U1991 ( .A0(n2295), .A1(n553), .B0(cacheAddressIn_SOUTH[0]), .B1(
        n535), .C0(cacheAddressIn_EAST[0]), .C1(n530), .Y(n1689) );
  OAI221XLTS U1992 ( .A0(n2181), .A1(n666), .B0(n2016), .B1(n2237), .C0(n1688), 
        .Y(n3210) );
  AOI222XLTS U1993 ( .A0(n2298), .A1(n553), .B0(cacheAddressIn_SOUTH[1]), .B1(
        n535), .C0(cacheAddressIn_EAST[1]), .C1(n530), .Y(n1688) );
  OAI221XLTS U1994 ( .A0(n2181), .A1(n665), .B0(n2018), .B1(n2237), .C0(n1687), 
        .Y(n3211) );
  AOI222XLTS U1995 ( .A0(n2301), .A1(n553), .B0(cacheAddressIn_SOUTH[2]), .B1(
        n535), .C0(cacheAddressIn_EAST[2]), .C1(n530), .Y(n1687) );
  OAI221XLTS U1996 ( .A0(n2181), .A1(n664), .B0(n2020), .B1(n2237), .C0(n1686), 
        .Y(n3212) );
  AOI222XLTS U1997 ( .A0(n2304), .A1(n553), .B0(cacheAddressIn_SOUTH[3]), .B1(
        n535), .C0(cacheAddressIn_EAST[3]), .C1(n530), .Y(n1686) );
  OAI221XLTS U1998 ( .A0(n2179), .A1(n663), .B0(n2022), .B1(n2241), .C0(n1685), 
        .Y(n3213) );
  AOI222XLTS U1999 ( .A0(n2307), .A1(n552), .B0(cacheAddressIn_SOUTH[4]), .B1(
        n540), .C0(cacheAddressIn_EAST[4]), .C1(n529), .Y(n1685) );
  OAI221XLTS U2000 ( .A0(n2181), .A1(n662), .B0(n2024), .B1(n2242), .C0(n1684), 
        .Y(n3214) );
  AOI222XLTS U2001 ( .A0(n2310), .A1(n552), .B0(cacheAddressIn_SOUTH[5]), .B1(
        n544), .C0(cacheAddressIn_EAST[5]), .C1(n529), .Y(n1684) );
  OAI221XLTS U2002 ( .A0(n2180), .A1(n661), .B0(n2026), .B1(n2238), .C0(n1683), 
        .Y(n3215) );
  AOI222XLTS U2003 ( .A0(n2313), .A1(n552), .B0(cacheAddressIn_SOUTH[6]), .B1(
        n1421), .C0(cacheAddressIn_EAST[6]), .C1(n529), .Y(n1683) );
  OAI221XLTS U2004 ( .A0(n2180), .A1(n660), .B0(n2028), .B1(n2238), .C0(n1682), 
        .Y(n3216) );
  AOI222XLTS U2005 ( .A0(n2316), .A1(n552), .B0(cacheAddressIn_SOUTH[7]), .B1(
        n1421), .C0(cacheAddressIn_EAST[7]), .C1(n529), .Y(n1682) );
  OAI221XLTS U2006 ( .A0(n2178), .A1(n896), .B0(n2030), .B1(n2242), .C0(n1453), 
        .Y(n3346) );
  AOI222XLTS U2007 ( .A0(n551), .A1(n2325), .B0(dataIn_SOUTH[0]), .B1(n543), 
        .C0(n528), .C1(dataIn_EAST[0]), .Y(n1453) );
  OAI221XLTS U2008 ( .A0(n2177), .A1(n895), .B0(n2032), .B1(n2240), .C0(n1452), 
        .Y(n3347) );
  AOI222XLTS U2009 ( .A0(n551), .A1(n2328), .B0(dataIn_SOUTH[1]), .B1(n543), 
        .C0(n528), .C1(dataIn_EAST[1]), .Y(n1452) );
  OAI221XLTS U2010 ( .A0(n2176), .A1(n894), .B0(n2034), .B1(n2240), .C0(n1451), 
        .Y(n3348) );
  AOI222XLTS U2011 ( .A0(n551), .A1(n2331), .B0(dataIn_SOUTH[2]), .B1(n544), 
        .C0(n528), .C1(dataIn_EAST[2]), .Y(n1451) );
  OAI221XLTS U2012 ( .A0(n2177), .A1(n893), .B0(n2036), .B1(n2241), .C0(n1450), 
        .Y(n3349) );
  AOI222XLTS U2013 ( .A0(n551), .A1(n2334), .B0(dataIn_SOUTH[3]), .B1(n541), 
        .C0(n528), .C1(dataIn_EAST[3]), .Y(n1450) );
  OAI221XLTS U2014 ( .A0(n2177), .A1(n892), .B0(n2038), .B1(n2238), .C0(n1449), 
        .Y(n3350) );
  AOI222XLTS U2015 ( .A0(n550), .A1(n2337), .B0(dataIn_SOUTH[4]), .B1(n544), 
        .C0(n527), .C1(dataIn_EAST[4]), .Y(n1449) );
  OAI221XLTS U2016 ( .A0(n2176), .A1(n891), .B0(n2040), .B1(n2237), .C0(n1448), 
        .Y(n3351) );
  AOI222XLTS U2017 ( .A0(n550), .A1(n2340), .B0(dataIn_SOUTH[5]), .B1(n541), 
        .C0(n527), .C1(dataIn_EAST[5]), .Y(n1448) );
  OAI221XLTS U2018 ( .A0(n2176), .A1(n890), .B0(n2042), .B1(n2239), .C0(n1447), 
        .Y(n3352) );
  AOI222XLTS U2019 ( .A0(n550), .A1(n2343), .B0(dataIn_SOUTH[6]), .B1(n540), 
        .C0(n527), .C1(dataIn_EAST[6]), .Y(n1447) );
  OAI221XLTS U2020 ( .A0(n2176), .A1(n889), .B0(n2044), .B1(n2239), .C0(n1446), 
        .Y(n3353) );
  AOI222XLTS U2021 ( .A0(n550), .A1(n2346), .B0(dataIn_SOUTH[7]), .B1(n543), 
        .C0(n527), .C1(dataIn_EAST[7]), .Y(n1446) );
  OAI221XLTS U2022 ( .A0(n2175), .A1(n888), .B0(n2046), .B1(n2238), .C0(n1445), 
        .Y(n3354) );
  AOI222XLTS U2023 ( .A0(n557), .A1(n2349), .B0(dataIn_SOUTH[8]), .B1(n542), 
        .C0(n533), .C1(dataIn_EAST[8]), .Y(n1445) );
  OAI221XLTS U2024 ( .A0(n2175), .A1(n887), .B0(n2048), .B1(n2244), .C0(n1444), 
        .Y(n3355) );
  AOI222XLTS U2025 ( .A0(n1420), .A1(n2352), .B0(dataIn_SOUTH[9]), .B1(n542), 
        .C0(n534), .C1(dataIn_EAST[9]), .Y(n1444) );
  OAI221XLTS U2026 ( .A0(n2175), .A1(n886), .B0(n2050), .B1(n2239), .C0(n1443), 
        .Y(n3356) );
  AOI222XLTS U2027 ( .A0(n556), .A1(n2355), .B0(dataIn_SOUTH[10]), .B1(n545), 
        .C0(n534), .C1(dataIn_EAST[10]), .Y(n1443) );
  OAI221XLTS U2028 ( .A0(n2175), .A1(n885), .B0(n2052), .B1(n2242), .C0(n1442), 
        .Y(n3357) );
  AOI222XLTS U2029 ( .A0(n555), .A1(n2358), .B0(dataIn_SOUTH[11]), .B1(n543), 
        .C0(n531), .C1(dataIn_EAST[11]), .Y(n1442) );
  OAI221XLTS U2030 ( .A0(n2174), .A1(n884), .B0(n2054), .B1(n2239), .C0(n1441), 
        .Y(n3358) );
  AOI222XLTS U2031 ( .A0(n1420), .A1(n2361), .B0(dataIn_SOUTH[12]), .B1(n546), 
        .C0(n532), .C1(dataIn_EAST[12]), .Y(n1441) );
  OAI221XLTS U2032 ( .A0(n2174), .A1(n883), .B0(n2056), .B1(n2236), .C0(n1440), 
        .Y(n3359) );
  AOI222XLTS U2033 ( .A0(n558), .A1(n2364), .B0(dataIn_SOUTH[13]), .B1(n542), 
        .C0(n1422), .C1(dataIn_EAST[13]), .Y(n1440) );
  OAI221XLTS U2034 ( .A0(n2169), .A1(n882), .B0(n2058), .B1(n2236), .C0(n1439), 
        .Y(n3360) );
  AOI222XLTS U2035 ( .A0(n556), .A1(n2367), .B0(dataIn_SOUTH[14]), .B1(n546), 
        .C0(n532), .C1(dataIn_EAST[14]), .Y(n1439) );
  OAI221XLTS U2036 ( .A0(n2170), .A1(n881), .B0(n2060), .B1(n2236), .C0(n1438), 
        .Y(n3361) );
  AOI222XLTS U2037 ( .A0(n554), .A1(n2370), .B0(dataIn_SOUTH[15]), .B1(n542), 
        .C0(n1422), .C1(dataIn_EAST[15]), .Y(n1438) );
  OAI221XLTS U2038 ( .A0(n2170), .A1(n879), .B0(n2062), .B1(n2236), .C0(n1437), 
        .Y(n3362) );
  AOI222XLTS U2039 ( .A0(n555), .A1(n2373), .B0(dataIn_SOUTH[16]), .B1(n536), 
        .C0(n526), .C1(dataIn_EAST[16]), .Y(n1437) );
  OAI221XLTS U2040 ( .A0(n2170), .A1(n878), .B0(n2064), .B1(n2235), .C0(n1436), 
        .Y(n3363) );
  AOI222XLTS U2041 ( .A0(n554), .A1(n2376), .B0(dataIn_SOUTH[17]), .B1(n536), 
        .C0(n526), .C1(dataIn_EAST[17]), .Y(n1436) );
  OAI221XLTS U2042 ( .A0(n2170), .A1(n877), .B0(n2066), .B1(n2235), .C0(n1435), 
        .Y(n3364) );
  AOI222XLTS U2043 ( .A0(n558), .A1(n2379), .B0(dataIn_SOUTH[18]), .B1(n536), 
        .C0(n526), .C1(dataIn_EAST[18]), .Y(n1435) );
  OAI221XLTS U2044 ( .A0(n2171), .A1(n876), .B0(n2068), .B1(n2235), .C0(n1434), 
        .Y(n3365) );
  AOI222XLTS U2045 ( .A0(n557), .A1(n2382), .B0(dataIn_SOUTH[19]), .B1(n536), 
        .C0(n526), .C1(dataIn_EAST[19]), .Y(n1434) );
  OAI221XLTS U2046 ( .A0(n2171), .A1(n875), .B0(n2070), .B1(n2235), .C0(n1433), 
        .Y(n3366) );
  AOI222XLTS U2047 ( .A0(n549), .A1(n2385), .B0(dataIn_SOUTH[20]), .B1(n537), 
        .C0(n525), .C1(dataIn_EAST[20]), .Y(n1433) );
  OAI221XLTS U2048 ( .A0(n2171), .A1(n874), .B0(n2072), .B1(n2234), .C0(n1432), 
        .Y(n3367) );
  AOI222XLTS U2049 ( .A0(n549), .A1(n2388), .B0(dataIn_SOUTH[21]), .B1(n537), 
        .C0(n525), .C1(dataIn_EAST[21]), .Y(n1432) );
  OAI221XLTS U2050 ( .A0(n2171), .A1(n873), .B0(n2074), .B1(n2234), .C0(n1431), 
        .Y(n3368) );
  AOI222XLTS U2051 ( .A0(n549), .A1(n2391), .B0(dataIn_SOUTH[22]), .B1(n537), 
        .C0(n525), .C1(dataIn_EAST[22]), .Y(n1431) );
  OAI221XLTS U2052 ( .A0(n2172), .A1(n872), .B0(n2076), .B1(n2234), .C0(n1430), 
        .Y(n3369) );
  AOI222XLTS U2053 ( .A0(n549), .A1(n2394), .B0(dataIn_SOUTH[23]), .B1(n537), 
        .C0(n525), .C1(dataIn_EAST[23]), .Y(n1430) );
  OAI221XLTS U2054 ( .A0(n2172), .A1(n871), .B0(n2078), .B1(n2233), .C0(n1429), 
        .Y(n3370) );
  AOI222XLTS U2055 ( .A0(n548), .A1(n2397), .B0(dataIn_SOUTH[24]), .B1(n538), 
        .C0(n524), .C1(dataIn_EAST[24]), .Y(n1429) );
  OAI221XLTS U2056 ( .A0(n2172), .A1(n870), .B0(n2080), .B1(n2233), .C0(n1428), 
        .Y(n3371) );
  AOI222XLTS U2057 ( .A0(n548), .A1(n2400), .B0(dataIn_SOUTH[25]), .B1(n538), 
        .C0(n524), .C1(dataIn_EAST[25]), .Y(n1428) );
  OAI221XLTS U2058 ( .A0(n2172), .A1(n869), .B0(n2082), .B1(n2233), .C0(n1427), 
        .Y(n3372) );
  AOI222XLTS U2059 ( .A0(n548), .A1(n2403), .B0(dataIn_SOUTH[26]), .B1(n538), 
        .C0(n524), .C1(dataIn_EAST[26]), .Y(n1427) );
  OAI221XLTS U2060 ( .A0(n2173), .A1(n868), .B0(n2084), .B1(n2234), .C0(n1426), 
        .Y(n3373) );
  AOI222XLTS U2061 ( .A0(n548), .A1(n2406), .B0(dataIn_SOUTH[27]), .B1(n538), 
        .C0(n524), .C1(dataIn_EAST[27]), .Y(n1426) );
  OAI221XLTS U2062 ( .A0(n2173), .A1(n867), .B0(n2086), .B1(n2232), .C0(n1425), 
        .Y(n3374) );
  AOI222XLTS U2063 ( .A0(n547), .A1(n2409), .B0(dataIn_SOUTH[28]), .B1(n539), 
        .C0(n523), .C1(dataIn_EAST[28]), .Y(n1425) );
  OAI221XLTS U2064 ( .A0(n2173), .A1(n866), .B0(n2088), .B1(n2232), .C0(n1424), 
        .Y(n3375) );
  AOI222XLTS U2065 ( .A0(n547), .A1(n2412), .B0(dataIn_SOUTH[29]), .B1(n539), 
        .C0(n523), .C1(dataIn_EAST[29]), .Y(n1424) );
  OAI221XLTS U2066 ( .A0(n2173), .A1(n865), .B0(n2090), .B1(n2232), .C0(n1423), 
        .Y(n3376) );
  AOI222XLTS U2067 ( .A0(n547), .A1(n2415), .B0(dataIn_SOUTH[30]), .B1(n539), 
        .C0(n523), .C1(dataIn_EAST[30]), .Y(n1423) );
  OAI221XLTS U2068 ( .A0(n2174), .A1(n864), .B0(n2092), .B1(n2243), .C0(n1419), 
        .Y(n3377) );
  AOI222XLTS U2069 ( .A0(n547), .A1(n2418), .B0(dataIn_SOUTH[31]), .B1(n539), 
        .C0(n523), .C1(dataIn_EAST[31]), .Y(n1419) );
  OAI221XLTS U2070 ( .A0(n2145), .A1(n2424), .B0(n2162), .B1(n862), .C0(n1159), 
        .Y(n3640) );
  AOI22X1TS U2071 ( .A0(n2328), .A1(n2138), .B0(n735), .B1(n2255), .Y(n1159)
         );
  OAI221XLTS U2072 ( .A0(n2145), .A1(n2426), .B0(n2163), .B1(n861), .C0(n1160), 
        .Y(n3639) );
  AOI22X1TS U2073 ( .A0(n2331), .A1(n2139), .B0(n734), .B1(n2251), .Y(n1160)
         );
  OAI221XLTS U2074 ( .A0(n2145), .A1(n2428), .B0(n2164), .B1(n860), .C0(n1161), 
        .Y(n3638) );
  AOI22X1TS U2075 ( .A0(n2334), .A1(n2137), .B0(n733), .B1(n2251), .Y(n1161)
         );
  OAI221XLTS U2076 ( .A0(n2144), .A1(n2432), .B0(n2189), .B1(n858), .C0(n1163), 
        .Y(n3636) );
  AOI22X1TS U2077 ( .A0(n2340), .A1(n1158), .B0(n731), .B1(n798), .Y(n1163) );
  OAI221XLTS U2078 ( .A0(n2144), .A1(n2434), .B0(n2163), .B1(n857), .C0(n1164), 
        .Y(n3635) );
  AOI22X1TS U2079 ( .A0(n2343), .A1(n2137), .B0(n730), .B1(n2256), .Y(n1164)
         );
  OAI221XLTS U2080 ( .A0(n2144), .A1(n2436), .B0(n2165), .B1(n856), .C0(n1165), 
        .Y(n3634) );
  AOI22X1TS U2081 ( .A0(n2346), .A1(n1158), .B0(n729), .B1(n2256), .Y(n1165)
         );
  OAI221XLTS U2082 ( .A0(n2143), .A1(n2440), .B0(n2166), .B1(n854), .C0(n1167), 
        .Y(n3632) );
  AOI22X1TS U2083 ( .A0(n2352), .A1(n2136), .B0(n727), .B1(n2253), .Y(n1167)
         );
  OAI221XLTS U2084 ( .A0(n2143), .A1(n2442), .B0(n2166), .B1(n853), .C0(n1168), 
        .Y(n3631) );
  AOI22X1TS U2085 ( .A0(n2355), .A1(n2139), .B0(n726), .B1(n2255), .Y(n1168)
         );
  OAI221XLTS U2086 ( .A0(n2145), .A1(n2422), .B0(n2161), .B1(n863), .C0(n1157), 
        .Y(n3641) );
  AOI22X1TS U2087 ( .A0(n2325), .A1(n2134), .B0(n736), .B1(n798), .Y(n1157) );
  OAI221XLTS U2088 ( .A0(n2144), .A1(n2430), .B0(n2165), .B1(n859), .C0(n1162), 
        .Y(n3637) );
  AOI22X1TS U2089 ( .A0(n2337), .A1(n2134), .B0(n732), .B1(n2254), .Y(n1162)
         );
  OAI221XLTS U2090 ( .A0(n2143), .A1(n2438), .B0(n2182), .B1(n855), .C0(n1166), 
        .Y(n3633) );
  AOI22X1TS U2091 ( .A0(n2349), .A1(n2138), .B0(n728), .B1(n2253), .Y(n1166)
         );
  OAI221XLTS U2092 ( .A0(n2143), .A1(n2444), .B0(n2164), .B1(n852), .C0(n1169), 
        .Y(n3630) );
  AOI22X1TS U2093 ( .A0(n2358), .A1(n2136), .B0(n725), .B1(n2254), .Y(n1169)
         );
  OAI221XLTS U2094 ( .A0(n2142), .A1(n2446), .B0(n2163), .B1(n851), .C0(n1170), 
        .Y(n3629) );
  AOI22X1TS U2095 ( .A0(n2361), .A1(n2128), .B0(n724), .B1(n2245), .Y(n1170)
         );
  OAI221XLTS U2096 ( .A0(n2179), .A1(n951), .B0(n1409), .B1(n2286), .C0(n1482), 
        .Y(n3338) );
  AOI22X1TS U2097 ( .A0(n2304), .A1(n397), .B0(n779), .B1(n388), .Y(n1482) );
  OAI221XLTS U2098 ( .A0(n2179), .A1(n949), .B0(n373), .B1(n2290), .C0(n1484), 
        .Y(n3336) );
  AOI22X1TS U2099 ( .A0(n2310), .A1(n356), .B0(n777), .B1(n390), .Y(n1484) );
  OAI221XLTS U2100 ( .A0(n2180), .A1(n947), .B0(n374), .B1(n2294), .C0(n1486), 
        .Y(n3334) );
  AOI22X1TS U2101 ( .A0(n2316), .A1(n356), .B0(n775), .B1(n389), .Y(n1486) );
  OAI221XLTS U2102 ( .A0(n2178), .A1(n953), .B0(n1409), .B1(n2282), .C0(n1480), 
        .Y(n3340) );
  AOI22X1TS U2103 ( .A0(n2298), .A1(n397), .B0(n781), .B1(n390), .Y(n1480) );
  OAI221XLTS U2104 ( .A0(n2178), .A1(n952), .B0(n373), .B1(n2284), .C0(n1481), 
        .Y(n3339) );
  AOI22X1TS U2105 ( .A0(n2301), .A1(n1411), .B0(n780), .B1(n389), .Y(n1481) );
  OAI221XLTS U2106 ( .A0(n2178), .A1(n950), .B0(n374), .B1(n2288), .C0(n1483), 
        .Y(n3337) );
  AOI22X1TS U2107 ( .A0(n2307), .A1(n356), .B0(n778), .B1(n390), .Y(n1483) );
  OAI221XLTS U2108 ( .A0(n2179), .A1(n948), .B0(n1409), .B1(n2292), .C0(n1485), 
        .Y(n3335) );
  AOI22X1TS U2109 ( .A0(n2313), .A1(n397), .B0(n776), .B1(n389), .Y(n1485) );
  OAI221XLTS U2110 ( .A0(n2177), .A1(n954), .B0(n373), .B1(n2280), .C0(n1479), 
        .Y(n3341) );
  AOI22X1TS U2111 ( .A0(n2295), .A1(n397), .B0(n782), .B1(n390), .Y(n1479) );
  OAI221XLTS U2112 ( .A0(n2174), .A1(n932), .B0(n374), .B1(n977), .C0(n1410), 
        .Y(n3385) );
  AOI22X1TS U2113 ( .A0(n25), .A1(n356), .B0(n2089), .B1(n389), .Y(n1410) );
  OAI221XLTS U2114 ( .A0(n2142), .A1(n2448), .B0(n2191), .B1(n850), .C0(n1171), 
        .Y(n3628) );
  AOI22X1TS U2115 ( .A0(n2364), .A1(n2128), .B0(n723), .B1(n2245), .Y(n1171)
         );
  OAI221XLTS U2116 ( .A0(n2142), .A1(n2450), .B0(n2191), .B1(n849), .C0(n1172), 
        .Y(n3627) );
  AOI22X1TS U2117 ( .A0(n2367), .A1(n2128), .B0(n722), .B1(n2245), .Y(n1172)
         );
  OAI221XLTS U2118 ( .A0(n2142), .A1(n2452), .B0(n2190), .B1(n848), .C0(n1173), 
        .Y(n3626) );
  AOI22X1TS U2119 ( .A0(n2370), .A1(n2128), .B0(n721), .B1(n2245), .Y(n1173)
         );
  OAI221XLTS U2120 ( .A0(n2148), .A1(n2456), .B0(n2161), .B1(n846), .C0(n1175), 
        .Y(n3624) );
  AOI22X1TS U2121 ( .A0(n2376), .A1(n2129), .B0(n719), .B1(n2246), .Y(n1175)
         );
  OAI221XLTS U2122 ( .A0(n2148), .A1(n2458), .B0(n2165), .B1(n845), .C0(n1176), 
        .Y(n3623) );
  AOI22X1TS U2123 ( .A0(n2379), .A1(n2129), .B0(n718), .B1(n2246), .Y(n1176)
         );
  OAI221XLTS U2124 ( .A0(n2146), .A1(n2460), .B0(n2162), .B1(n844), .C0(n1177), 
        .Y(n3622) );
  AOI22X1TS U2125 ( .A0(n2382), .A1(n2129), .B0(n717), .B1(n2246), .Y(n1177)
         );
  OAI221XLTS U2126 ( .A0(n2148), .A1(n2462), .B0(n2188), .B1(n843), .C0(n1178), 
        .Y(n3621) );
  AOI22X1TS U2127 ( .A0(n2385), .A1(n2130), .B0(n716), .B1(n2247), .Y(n1178)
         );
  OAI221XLTS U2128 ( .A0(n2148), .A1(n2466), .B0(n2167), .B1(n841), .C0(n1180), 
        .Y(n3619) );
  AOI22X1TS U2129 ( .A0(n2391), .A1(n2130), .B0(n792), .B1(n2247), .Y(n1180)
         );
  OAI221XLTS U2130 ( .A0(n2147), .A1(n2468), .B0(n2169), .B1(n840), .C0(n1181), 
        .Y(n3618) );
  AOI22X1TS U2131 ( .A0(n2394), .A1(n2130), .B0(n791), .B1(n2247), .Y(n1181)
         );
  OAI221XLTS U2132 ( .A0(n2141), .A1(n2472), .B0(n2167), .B1(n838), .C0(n1183), 
        .Y(n3616) );
  AOI22X1TS U2133 ( .A0(n2400), .A1(n2131), .B0(n789), .B1(n2248), .Y(n1183)
         );
  OAI221XLTS U2134 ( .A0(n2141), .A1(n2474), .B0(n2168), .B1(n837), .C0(n1184), 
        .Y(n3615) );
  AOI22X1TS U2135 ( .A0(n2403), .A1(n2131), .B0(n788), .B1(n2248), .Y(n1184)
         );
  OAI221XLTS U2136 ( .A0(n2141), .A1(n2476), .B0(n2168), .B1(n836), .C0(n1185), 
        .Y(n3614) );
  AOI22X1TS U2137 ( .A0(n2406), .A1(n2131), .B0(n787), .B1(n2248), .Y(n1185)
         );
  OAI221XLTS U2138 ( .A0(n2140), .A1(n2478), .B0(n2168), .B1(n835), .C0(n1186), 
        .Y(n3613) );
  AOI22X1TS U2139 ( .A0(n2409), .A1(n2132), .B0(n786), .B1(n2249), .Y(n1186)
         );
  OAI221XLTS U2140 ( .A0(n2140), .A1(n2480), .B0(n2168), .B1(n834), .C0(n1187), 
        .Y(n3612) );
  AOI22X1TS U2141 ( .A0(n2412), .A1(n2132), .B0(n785), .B1(n2249), .Y(n1187)
         );
  OAI221XLTS U2142 ( .A0(n2140), .A1(n2482), .B0(n2169), .B1(n833), .C0(n1188), 
        .Y(n3611) );
  AOI22X1TS U2143 ( .A0(n2415), .A1(n2132), .B0(n784), .B1(n2249), .Y(n1188)
         );
  OAI221XLTS U2144 ( .A0(n2146), .A1(n2454), .B0(n2161), .B1(n847), .C0(n1174), 
        .Y(n3625) );
  AOI22X1TS U2145 ( .A0(n2373), .A1(n2129), .B0(n720), .B1(n2246), .Y(n1174)
         );
  OAI221XLTS U2146 ( .A0(n2149), .A1(n2464), .B0(n2167), .B1(n842), .C0(n1179), 
        .Y(n3620) );
  AOI22X1TS U2147 ( .A0(n2388), .A1(n2130), .B0(n793), .B1(n2247), .Y(n1179)
         );
  OAI221XLTS U2148 ( .A0(n2141), .A1(n2470), .B0(n2167), .B1(n839), .C0(n1182), 
        .Y(n3617) );
  AOI22X1TS U2149 ( .A0(n2397), .A1(n2131), .B0(n790), .B1(n2248), .Y(n1182)
         );
  OAI221XLTS U2150 ( .A0(n2140), .A1(n2484), .B0(n2169), .B1(n832), .C0(n1189), 
        .Y(n3610) );
  AOI22X1TS U2151 ( .A0(n2418), .A1(n2132), .B0(n783), .B1(n2249), .Y(n1189)
         );
  OAI211X1TS U2152 ( .A0(n1709), .A1(n830), .B0(n1710), .C0(n1711), .Y(n3190)
         );
  AOI22X1TS U2153 ( .A0(requesterAddressIn_NORTH[0]), .A1(n1713), .B0(n1714), 
        .B1(requesterAddressIn_EAST[0]), .Y(n1710) );
  AOI222XLTS U2154 ( .A0(n1712), .A1(requesterAddressIn_SOUTH[0]), .B0(n1612), 
        .B1(requesterAddressIn_WEST[0]), .C0(\requesterAddressBuffer[0][0] ), 
        .C1(n363), .Y(n1711) );
  OAI211X1TS U2155 ( .A0(n1709), .A1(n829), .B0(n1715), .C0(n1716), .Y(n3189)
         );
  AOI22X1TS U2156 ( .A0(requesterAddressIn_NORTH[1]), .A1(n1713), .B0(n1714), 
        .B1(requesterAddressIn_EAST[1]), .Y(n1715) );
  AOI222XLTS U2157 ( .A0(n1712), .A1(requesterAddressIn_SOUTH[1]), .B0(n1612), 
        .B1(requesterAddressIn_WEST[1]), .C0(\requesterAddressBuffer[0][1] ), 
        .C1(n363), .Y(n1716) );
  OAI211X1TS U2158 ( .A0(n382), .A1(n828), .B0(n1717), .C0(n1718), .Y(n3188)
         );
  AOI22X1TS U2159 ( .A0(requesterAddressIn_NORTH[2]), .A1(n1713), .B0(n1714), 
        .B1(requesterAddressIn_EAST[2]), .Y(n1717) );
  AOI222XLTS U2160 ( .A0(n1712), .A1(requesterAddressIn_SOUTH[2]), .B0(n1612), 
        .B1(requesterAddressIn_WEST[2]), .C0(\requesterAddressBuffer[0][2] ), 
        .C1(n363), .Y(n1718) );
  OAI211X1TS U2161 ( .A0(n382), .A1(n827), .B0(n1719), .C0(n1720), .Y(n3187)
         );
  AOI22X1TS U2162 ( .A0(requesterAddressIn_NORTH[3]), .A1(n346), .B0(n342), 
        .B1(requesterAddressIn_EAST[3]), .Y(n1719) );
  AOI222XLTS U2163 ( .A0(n343), .A1(requesterAddressIn_SOUTH[3]), .B0(n351), 
        .B1(requesterAddressIn_WEST[3]), .C0(\requesterAddressBuffer[0][3] ), 
        .C1(n363), .Y(n1720) );
  OAI211X1TS U2164 ( .A0(n382), .A1(n826), .B0(n1721), .C0(n1722), .Y(n3186)
         );
  AOI22X1TS U2165 ( .A0(requesterAddressIn_NORTH[4]), .A1(n346), .B0(n342), 
        .B1(requesterAddressIn_EAST[4]), .Y(n1721) );
  AOI222XLTS U2166 ( .A0(n343), .A1(requesterAddressIn_SOUTH[4]), .B0(n351), 
        .B1(requesterAddressIn_WEST[4]), .C0(\requesterAddressBuffer[0][4] ), 
        .C1(n364), .Y(n1722) );
  OAI211X1TS U2167 ( .A0(n382), .A1(n825), .B0(n1723), .C0(n1724), .Y(n3185)
         );
  AOI22X1TS U2168 ( .A0(requesterAddressIn_NORTH[5]), .A1(n346), .B0(n342), 
        .B1(requesterAddressIn_EAST[5]), .Y(n1723) );
  AOI222XLTS U2169 ( .A0(n343), .A1(requesterAddressIn_SOUTH[5]), .B0(n351), 
        .B1(requesterAddressIn_WEST[5]), .C0(\requesterAddressBuffer[0][5] ), 
        .C1(n364), .Y(n1724) );
  OAI211X1TS U2170 ( .A0(n1975), .A1(n509), .B0(n1675), .C0(n1676), .Y(n3218)
         );
  AOI222XLTS U2171 ( .A0(n1577), .A1(dataIn_EAST[0]), .B0(n492), .B1(
        dataIn_SOUTH[0]), .C0(n484), .C1(n2325), .Y(n1676) );
  AOI22X1TS U2172 ( .A0(dataIn_NORTH[0]), .A1(n461), .B0(n736), .B1(n2155), 
        .Y(n1675) );
  OAI211X1TS U2173 ( .A0(n1976), .A1(n509), .B0(n1673), .C0(n1674), .Y(n3219)
         );
  AOI222XLTS U2174 ( .A0(n507), .A1(dataIn_EAST[1]), .B0(n492), .B1(
        dataIn_SOUTH[1]), .C0(n480), .C1(n2328), .Y(n1674) );
  AOI22X1TS U2175 ( .A0(dataIn_NORTH[1]), .A1(n461), .B0(n735), .B1(n2150), 
        .Y(n1673) );
  OAI211X1TS U2176 ( .A0(n1977), .A1(n509), .B0(n1671), .C0(n1672), .Y(n3220)
         );
  AOI222XLTS U2177 ( .A0(n507), .A1(dataIn_EAST[2]), .B0(n492), .B1(
        dataIn_SOUTH[2]), .C0(n484), .C1(n2331), .Y(n1672) );
  AOI22X1TS U2178 ( .A0(dataIn_NORTH[2]), .A1(n461), .B0(n734), .B1(n2150), 
        .Y(n1671) );
  OAI211X1TS U2179 ( .A0(n1978), .A1(n510), .B0(n1669), .C0(n1670), .Y(n3221)
         );
  AOI222XLTS U2180 ( .A0(n506), .A1(dataIn_EAST[3]), .B0(n492), .B1(
        dataIn_SOUTH[3]), .C0(n1579), .C1(n2334), .Y(n1670) );
  AOI22X1TS U2181 ( .A0(dataIn_NORTH[3]), .A1(n461), .B0(n733), .B1(n2150), 
        .Y(n1669) );
  OAI211X1TS U2182 ( .A0(n1979), .A1(n510), .B0(n1667), .C0(n1668), .Y(n3222)
         );
  AOI222XLTS U2183 ( .A0(n508), .A1(dataIn_EAST[4]), .B0(n491), .B1(
        dataIn_SOUTH[4]), .C0(n473), .C1(n2337), .Y(n1668) );
  AOI22X1TS U2184 ( .A0(dataIn_NORTH[4]), .A1(n462), .B0(n732), .B1(n2152), 
        .Y(n1667) );
  OAI211X1TS U2185 ( .A0(n1980), .A1(n510), .B0(n1665), .C0(n1666), .Y(n3223)
         );
  AOI222XLTS U2186 ( .A0(n505), .A1(dataIn_EAST[5]), .B0(n491), .B1(
        dataIn_SOUTH[5]), .C0(n473), .C1(n2340), .Y(n1666) );
  AOI22X1TS U2187 ( .A0(dataIn_NORTH[5]), .A1(n462), .B0(n731), .B1(n2152), 
        .Y(n1665) );
  OAI211X1TS U2188 ( .A0(n1981), .A1(n510), .B0(n1663), .C0(n1664), .Y(n3224)
         );
  AOI222XLTS U2189 ( .A0(n508), .A1(dataIn_EAST[6]), .B0(n491), .B1(
        dataIn_SOUTH[6]), .C0(n473), .C1(n2343), .Y(n1664) );
  AOI22X1TS U2190 ( .A0(dataIn_NORTH[6]), .A1(n462), .B0(n730), .B1(n2152), 
        .Y(n1663) );
  OAI211X1TS U2191 ( .A0(n1982), .A1(n511), .B0(n1661), .C0(n1662), .Y(n3225)
         );
  AOI222XLTS U2192 ( .A0(n504), .A1(dataIn_EAST[7]), .B0(n491), .B1(
        dataIn_SOUTH[7]), .C0(n473), .C1(n2346), .Y(n1662) );
  AOI22X1TS U2193 ( .A0(dataIn_NORTH[7]), .A1(n462), .B0(n729), .B1(n2152), 
        .Y(n1661) );
  OAI211X1TS U2194 ( .A0(n1983), .A1(n511), .B0(n1659), .C0(n1660), .Y(n3226)
         );
  AOI222XLTS U2195 ( .A0(n497), .A1(dataIn_EAST[8]), .B0(n490), .B1(
        dataIn_SOUTH[8]), .C0(n474), .C1(n2349), .Y(n1660) );
  AOI22X1TS U2196 ( .A0(dataIn_NORTH[8]), .A1(n463), .B0(n728), .B1(n2151), 
        .Y(n1659) );
  OAI211X1TS U2197 ( .A0(n1984), .A1(n511), .B0(n1657), .C0(n1658), .Y(n3227)
         );
  AOI222XLTS U2198 ( .A0(n497), .A1(dataIn_EAST[9]), .B0(n490), .B1(
        dataIn_SOUTH[9]), .C0(n474), .C1(n2352), .Y(n1658) );
  AOI22X1TS U2199 ( .A0(dataIn_NORTH[9]), .A1(n463), .B0(n727), .B1(n2151), 
        .Y(n1657) );
  OAI211X1TS U2200 ( .A0(n1985), .A1(n511), .B0(n1655), .C0(n1656), .Y(n3228)
         );
  AOI222XLTS U2201 ( .A0(n497), .A1(dataIn_EAST[10]), .B0(n490), .B1(
        dataIn_SOUTH[10]), .C0(n474), .C1(n2355), .Y(n1656) );
  AOI22X1TS U2202 ( .A0(dataIn_NORTH[10]), .A1(n463), .B0(n726), .B1(n2151), 
        .Y(n1655) );
  OAI211X1TS U2203 ( .A0(n1986), .A1(n512), .B0(n1653), .C0(n1654), .Y(n3229)
         );
  AOI222XLTS U2204 ( .A0(n497), .A1(dataIn_EAST[11]), .B0(n490), .B1(
        dataIn_SOUTH[11]), .C0(n474), .C1(n2358), .Y(n1654) );
  AOI22X1TS U2205 ( .A0(dataIn_NORTH[11]), .A1(n463), .B0(n725), .B1(n2151), 
        .Y(n1653) );
  OAI211X1TS U2206 ( .A0(n1987), .A1(n512), .B0(n1651), .C0(n1652), .Y(n3230)
         );
  AOI222XLTS U2207 ( .A0(n498), .A1(dataIn_EAST[12]), .B0(n489), .B1(
        dataIn_SOUTH[12]), .C0(n475), .C1(n2361), .Y(n1652) );
  AOI22X1TS U2208 ( .A0(dataIn_NORTH[12]), .A1(n464), .B0(n724), .B1(n2154), 
        .Y(n1651) );
  OAI211X1TS U2209 ( .A0(n1988), .A1(n512), .B0(n1649), .C0(n1650), .Y(n3231)
         );
  AOI222XLTS U2210 ( .A0(n498), .A1(dataIn_EAST[13]), .B0(n489), .B1(
        dataIn_SOUTH[13]), .C0(n475), .C1(n2364), .Y(n1650) );
  AOI22X1TS U2211 ( .A0(dataIn_NORTH[13]), .A1(n464), .B0(n723), .B1(n2154), 
        .Y(n1649) );
  OAI211X1TS U2212 ( .A0(n1989), .A1(n512), .B0(n1647), .C0(n1648), .Y(n3232)
         );
  AOI222XLTS U2213 ( .A0(n498), .A1(dataIn_EAST[14]), .B0(n489), .B1(
        dataIn_SOUTH[14]), .C0(n475), .C1(n2367), .Y(n1648) );
  AOI22X1TS U2214 ( .A0(dataIn_NORTH[14]), .A1(n464), .B0(n722), .B1(n2154), 
        .Y(n1647) );
  OAI211X1TS U2215 ( .A0(n1990), .A1(n513), .B0(n1645), .C0(n1646), .Y(n3233)
         );
  AOI222XLTS U2216 ( .A0(n498), .A1(dataIn_EAST[15]), .B0(n489), .B1(
        dataIn_SOUTH[15]), .C0(n475), .C1(n2370), .Y(n1646) );
  AOI22X1TS U2217 ( .A0(dataIn_NORTH[15]), .A1(n464), .B0(n721), .B1(n2154), 
        .Y(n1645) );
  OAI211X1TS U2218 ( .A0(n1991), .A1(n513), .B0(n1643), .C0(n1644), .Y(n3234)
         );
  AOI222XLTS U2219 ( .A0(n499), .A1(dataIn_EAST[16]), .B0(n493), .B1(
        dataIn_SOUTH[16]), .C0(n476), .C1(n2373), .Y(n1644) );
  AOI22X1TS U2220 ( .A0(dataIn_NORTH[16]), .A1(n1580), .B0(n720), .B1(n2153), 
        .Y(n1643) );
  OAI211X1TS U2221 ( .A0(n1992), .A1(n513), .B0(n1641), .C0(n1642), .Y(n3235)
         );
  AOI222XLTS U2222 ( .A0(n499), .A1(dataIn_EAST[17]), .B0(n494), .B1(
        dataIn_SOUTH[17]), .C0(n476), .C1(n2376), .Y(n1642) );
  AOI22X1TS U2223 ( .A0(dataIn_NORTH[17]), .A1(n472), .B0(n719), .B1(n2153), 
        .Y(n1641) );
  OAI211X1TS U2224 ( .A0(n1993), .A1(n513), .B0(n1639), .C0(n1640), .Y(n3236)
         );
  AOI222XLTS U2225 ( .A0(n499), .A1(dataIn_EAST[18]), .B0(n1578), .B1(
        dataIn_SOUTH[18]), .C0(n476), .C1(n2379), .Y(n1640) );
  AOI22X1TS U2226 ( .A0(dataIn_NORTH[18]), .A1(n471), .B0(n718), .B1(n2153), 
        .Y(n1639) );
  OAI211X1TS U2227 ( .A0(n1994), .A1(n514), .B0(n1637), .C0(n1638), .Y(n3237)
         );
  AOI222XLTS U2228 ( .A0(n499), .A1(dataIn_EAST[19]), .B0(n1578), .B1(
        dataIn_SOUTH[19]), .C0(n476), .C1(n2382), .Y(n1638) );
  AOI22X1TS U2229 ( .A0(dataIn_NORTH[19]), .A1(n470), .B0(n717), .B1(n2153), 
        .Y(n1637) );
  OAI211X1TS U2230 ( .A0(n1995), .A1(n514), .B0(n1635), .C0(n1636), .Y(n3238)
         );
  AOI222XLTS U2231 ( .A0(n506), .A1(dataIn_EAST[20]), .B0(n496), .B1(
        dataIn_SOUTH[20]), .C0(n482), .C1(n2385), .Y(n1636) );
  AOI22X1TS U2232 ( .A0(dataIn_NORTH[20]), .A1(n469), .B0(n716), .B1(n2156), 
        .Y(n1635) );
  OAI211X1TS U2233 ( .A0(n1996), .A1(n514), .B0(n1633), .C0(n1634), .Y(n3239)
         );
  AOI222XLTS U2234 ( .A0(n506), .A1(dataIn_EAST[21]), .B0(n495), .B1(
        dataIn_SOUTH[21]), .C0(n481), .C1(n2388), .Y(n1634) );
  AOI22X1TS U2235 ( .A0(dataIn_NORTH[21]), .A1(n471), .B0(n793), .B1(n2156), 
        .Y(n1633) );
  OAI211X1TS U2236 ( .A0(n1997), .A1(n514), .B0(n1631), .C0(n1632), .Y(n3240)
         );
  AOI222XLTS U2237 ( .A0(n505), .A1(dataIn_EAST[22]), .B0(n496), .B1(
        dataIn_SOUTH[22]), .C0(n481), .C1(n2391), .Y(n1632) );
  AOI22X1TS U2238 ( .A0(dataIn_NORTH[22]), .A1(n470), .B0(n792), .B1(n2156), 
        .Y(n1631) );
  OAI211X1TS U2239 ( .A0(n1998), .A1(n515), .B0(n1629), .C0(n1630), .Y(n3241)
         );
  AOI222XLTS U2240 ( .A0(n504), .A1(dataIn_EAST[23]), .B0(n493), .B1(
        dataIn_SOUTH[23]), .C0(n480), .C1(n2394), .Y(n1630) );
  AOI22X1TS U2241 ( .A0(dataIn_NORTH[23]), .A1(n469), .B0(n791), .B1(n2157), 
        .Y(n1629) );
  OAI211X1TS U2242 ( .A0(n29), .A1(n83), .B0(n801), .C0(n1608), .Y(n3251) );
  AOI22X1TS U2243 ( .A0(n364), .A1(\requesterPortBuffer[0][1] ), .B0(n26), 
        .B1(n805), .Y(n1608) );
  INVX2TS U2244 ( .A(n1707), .Y(n773) );
  AOI222XLTS U2245 ( .A0(n2134), .A1(requesterAddressIn_WEST[0]), .B0(n1702), 
        .B1(requesterAddressIn_EAST[0]), .C0(n2251), .C1(
        \requesterAddressBuffer[0][0] ), .Y(n1707) );
  INVX2TS U2246 ( .A(n1706), .Y(n774) );
  AOI222XLTS U2247 ( .A0(n2134), .A1(requesterAddressIn_WEST[1]), .B0(n1702), 
        .B1(requesterAddressIn_EAST[1]), .C0(n2251), .C1(
        \requesterAddressBuffer[0][1] ), .Y(n1706) );
  INVX2TS U2248 ( .A(n1704), .Y(n795) );
  AOI222XLTS U2249 ( .A0(n2133), .A1(requesterAddressIn_WEST[3]), .B0(n1702), 
        .B1(requesterAddressIn_EAST[3]), .C0(n2250), .C1(
        \requesterAddressBuffer[0][3] ), .Y(n1704) );
  INVX2TS U2250 ( .A(n1705), .Y(n794) );
  AOI222XLTS U2251 ( .A0(n2133), .A1(requesterAddressIn_WEST[2]), .B0(n361), 
        .B1(requesterAddressIn_EAST[2]), .C0(n2250), .C1(
        \requesterAddressBuffer[0][2] ), .Y(n1705) );
  INVX2TS U2252 ( .A(n1703), .Y(n796) );
  AOI222XLTS U2253 ( .A0(n2133), .A1(requesterAddressIn_WEST[4]), .B0(n361), 
        .B1(requesterAddressIn_EAST[4]), .C0(n2250), .C1(
        \requesterAddressBuffer[0][4] ), .Y(n1703) );
  INVX2TS U2254 ( .A(n1701), .Y(n797) );
  AOI222XLTS U2255 ( .A0(n2133), .A1(requesterAddressIn_WEST[5]), .B0(n361), 
        .B1(requesterAddressIn_EAST[5]), .C0(n2250), .C1(
        \requesterAddressBuffer[0][5] ), .Y(n1701) );
  NAND2X1TS U2256 ( .A(n99), .B(n2500), .Y(n1130) );
  OAI22X1TS U2257 ( .A0(n46), .A1(n391), .B0(n2489), .B1(n1596), .Y(n3267) );
  AOI2BB1X1TS U2258 ( .A0N(n102), .A1N(n2083), .B0(n808), .Y(n1596) );
  OAI22X1TS U2259 ( .A0(n47), .A1(n393), .B0(n2489), .B1(n1597), .Y(n3266) );
  AOI2BB1X1TS U2260 ( .A0N(n813), .A1N(n2081), .B0(n808), .Y(n1597) );
  OAI22X1TS U2261 ( .A0(n392), .A1(n946), .B0(n1414), .B1(n1415), .Y(n3384) );
  AOI22X1TS U2262 ( .A0(n808), .A1(n25), .B0(n2091), .B1(n1416), .Y(n1414) );
  NAND2X1TS U2263 ( .A(n5), .B(n1154), .Y(n1151) );
  NAND3X1TS U2264 ( .A(\prevRequesterPort_B[0] ), .B(n449), .C(n51), .Y(n1776)
         );
  NAND2X1TS U2265 ( .A(n26), .B(n938), .Y(n1750) );
  OAI21X1TS U2266 ( .A0(n2490), .A1(n81), .B0(n1135), .Y(n2105) );
  AOI32X1TS U2267 ( .A0(\requesterPortBuffer[0][0] ), .A1(n36), .A2(n2210), 
        .B0(n2160), .B1(\requesterPortBuffer[2][0] ), .Y(n1135) );
  OAI2BB1X1TS U2268 ( .A0N(requesterAddressOut_SOUTH[0]), .A1N(n70), .B0(n1760), .Y(n3166) );
  AOI22X1TS U2269 ( .A0(n1754), .A1(prevRequesterAddress_A[0]), .B0(n1755), 
        .B1(prevRequesterAddress_B[0]), .Y(n1760) );
  OAI2BB1X1TS U2270 ( .A0N(requesterAddressOut_SOUTH[1]), .A1N(n71), .B0(n1759), .Y(n3167) );
  AOI22X1TS U2271 ( .A0(n1754), .A1(prevRequesterAddress_A[1]), .B0(n1755), 
        .B1(prevRequesterAddress_B[1]), .Y(n1759) );
  OAI2BB1X1TS U2272 ( .A0N(requesterAddressOut_SOUTH[2]), .A1N(n70), .B0(n1758), .Y(n3168) );
  AOI22X1TS U2273 ( .A0(n359), .A1(prevRequesterAddress_A[2]), .B0(n375), .B1(
        prevRequesterAddress_B[2]), .Y(n1758) );
  OAI2BB1X1TS U2274 ( .A0N(requesterAddressOut_SOUTH[3]), .A1N(n71), .B0(n1757), .Y(n3169) );
  AOI22X1TS U2275 ( .A0(n359), .A1(prevRequesterAddress_A[3]), .B0(n375), .B1(
        prevRequesterAddress_B[3]), .Y(n1757) );
  OAI2BB1X1TS U2276 ( .A0N(requesterAddressOut_SOUTH[4]), .A1N(n70), .B0(n1756), .Y(n3170) );
  AOI22X1TS U2277 ( .A0(n1754), .A1(prevRequesterAddress_A[4]), .B0(n1755), 
        .B1(prevRequesterAddress_B[4]), .Y(n1756) );
  OAI2BB1X1TS U2278 ( .A0N(requesterAddressOut_SOUTH[5]), .A1N(n71), .B0(n1753), .Y(n3171) );
  AOI22X1TS U2279 ( .A0(n359), .A1(prevRequesterAddress_A[5]), .B0(n375), .B1(
        prevRequesterAddress_B[5]), .Y(n1753) );
  OAI32X1TS U2280 ( .A0(n770), .A1(n2491), .A2(n1454), .B0(n1455), .B1(n659), 
        .Y(n3345) );
  AOI21X1TS U2281 ( .A0(n379), .A1(n1457), .B0(memRead_WEST), .Y(n1454) );
  OAI32X1TS U2282 ( .A0(n2204), .A1(n957), .A2(n1138), .B0(n45), .B1(n2182), 
        .Y(n2106) );
  INVX2TS U2283 ( .A(n1140), .Y(n957) );
  OAI221XLTS U2284 ( .A0(n830), .A1(n1764), .B0(n824), .B1(n1765), .C0(n1772), 
        .Y(n3160) );
  NAND2X1TS U2285 ( .A(requesterAddressOut_NORTH[0]), .B(n66), .Y(n1772) );
  OAI221XLTS U2286 ( .A0(n829), .A1(n1764), .B0(n823), .B1(n1765), .C0(n1771), 
        .Y(n3161) );
  NAND2X1TS U2287 ( .A(requesterAddressOut_NORTH[1]), .B(n67), .Y(n1771) );
  OAI221XLTS U2288 ( .A0(n828), .A1(n1764), .B0(n822), .B1(n1765), .C0(n1770), 
        .Y(n3162) );
  NAND2X1TS U2289 ( .A(requesterAddressOut_NORTH[2]), .B(n66), .Y(n1770) );
  OAI221XLTS U2290 ( .A0(n827), .A1(n357), .B0(n821), .B1(n376), .C0(n1769), 
        .Y(n3163) );
  NAND2X1TS U2291 ( .A(requesterAddressOut_NORTH[3]), .B(n67), .Y(n1769) );
  OAI221XLTS U2292 ( .A0(n826), .A1(n357), .B0(n820), .B1(n376), .C0(n1768), 
        .Y(n3164) );
  NAND2X1TS U2293 ( .A(requesterAddressOut_NORTH[4]), .B(n66), .Y(n1768) );
  OAI221XLTS U2294 ( .A0(n825), .A1(n357), .B0(n819), .B1(n376), .C0(n1766), 
        .Y(n3165) );
  NAND2X1TS U2295 ( .A(requesterAddressOut_NORTH[5]), .B(n67), .Y(n1766) );
  OAI221XLTS U2296 ( .A0(n2096), .A1(n2182), .B0(n2490), .B1(n1134), .C0(n1595), .Y(n3268) );
  OAI2BB1X1TS U2297 ( .A0N(n37), .A1N(n674), .B0(n2207), .Y(n1595) );
  OAI211X1TS U2298 ( .A0(n1569), .A1(n49), .B0(n802), .C0(n1600), .Y(n3265) );
  OA22X1TS U2299 ( .A0(n348), .A1(n384), .B0(n365), .B1(n46), .Y(n1600) );
  OAI211X1TS U2300 ( .A0(n35), .A1(n44), .B0(n802), .C0(n1603), .Y(n3264) );
  AOI2BB2X1TS U2301 ( .B0(n51), .B1(n1604), .A0N(n365), .A1N(n47), .Y(n1603)
         );
  AND2X2TS U2302 ( .A(n740), .B(n3), .Y(n396) );
  NOR2BX1TS U2303 ( .AN(n2), .B(\prevRequesterPort_B[0] ), .Y(n1751) );
  OAI2BB1X1TS U2304 ( .A0N(requesterAddressOut_WEST[0]), .A1N(n1730), .B0(
        n1738), .Y(n3178) );
  AOI22X1TS U2305 ( .A0(n1732), .A1(prevRequesterAddress_A[0]), .B0(n1733), 
        .B1(prevRequesterAddress_B[0]), .Y(n1738) );
  OAI2BB1X1TS U2306 ( .A0N(requesterAddressOut_WEST[1]), .A1N(n91), .B0(n1737), 
        .Y(n3179) );
  AOI22X1TS U2307 ( .A0(n1732), .A1(prevRequesterAddress_A[1]), .B0(n1733), 
        .B1(prevRequesterAddress_B[1]), .Y(n1737) );
  OAI2BB1X1TS U2308 ( .A0N(requesterAddressOut_WEST[2]), .A1N(n1730), .B0(
        n1736), .Y(n3180) );
  AOI22X1TS U2309 ( .A0(n1732), .A1(prevRequesterAddress_A[2]), .B0(n1733), 
        .B1(prevRequesterAddress_B[2]), .Y(n1736) );
  OAI2BB1X1TS U2310 ( .A0N(requesterAddressOut_WEST[3]), .A1N(n91), .B0(n1735), 
        .Y(n3181) );
  AOI22X1TS U2311 ( .A0(n360), .A1(prevRequesterAddress_A[3]), .B0(n377), .B1(
        prevRequesterAddress_B[3]), .Y(n1735) );
  OAI2BB1X1TS U2312 ( .A0N(requesterAddressOut_WEST[4]), .A1N(n1730), .B0(
        n1734), .Y(n3182) );
  AOI22X1TS U2313 ( .A0(n360), .A1(prevRequesterAddress_A[4]), .B0(n377), .B1(
        prevRequesterAddress_B[4]), .Y(n1734) );
  OAI2BB1X1TS U2314 ( .A0N(requesterAddressOut_WEST[5]), .A1N(n91), .B0(n1731), 
        .Y(n3183) );
  AOI22X1TS U2315 ( .A0(n360), .A1(prevRequesterAddress_A[5]), .B0(n377), .B1(
        prevRequesterAddress_B[5]), .Y(n1731) );
  INVX2TS U2316 ( .A(dataIn_EAST[0]), .Y(n2422) );
  INVX2TS U2317 ( .A(dataIn_EAST[1]), .Y(n2424) );
  INVX2TS U2318 ( .A(dataIn_EAST[2]), .Y(n2426) );
  INVX2TS U2319 ( .A(dataIn_EAST[3]), .Y(n2428) );
  INVX2TS U2320 ( .A(dataIn_EAST[4]), .Y(n2430) );
  INVX2TS U2321 ( .A(dataIn_EAST[5]), .Y(n2432) );
  INVX2TS U2322 ( .A(dataIn_EAST[6]), .Y(n2434) );
  INVX2TS U2323 ( .A(dataIn_EAST[7]), .Y(n2436) );
  INVX2TS U2324 ( .A(dataIn_EAST[8]), .Y(n2438) );
  INVX2TS U2325 ( .A(dataIn_EAST[9]), .Y(n2440) );
  INVX2TS U2326 ( .A(dataIn_EAST[10]), .Y(n2442) );
  INVX2TS U2327 ( .A(dataIn_EAST[11]), .Y(n2444) );
  INVX2TS U2328 ( .A(dataIn_EAST[12]), .Y(n2446) );
  INVX2TS U2329 ( .A(dataIn_EAST[13]), .Y(n2448) );
  INVX2TS U2330 ( .A(dataIn_EAST[14]), .Y(n2450) );
  INVX2TS U2331 ( .A(dataIn_EAST[15]), .Y(n2452) );
  INVX2TS U2332 ( .A(dataIn_EAST[16]), .Y(n2454) );
  INVX2TS U2333 ( .A(dataIn_EAST[17]), .Y(n2456) );
  INVX2TS U2334 ( .A(dataIn_EAST[18]), .Y(n2458) );
  INVX2TS U2335 ( .A(dataIn_EAST[19]), .Y(n2460) );
  INVX2TS U2336 ( .A(dataIn_EAST[20]), .Y(n2462) );
  INVX2TS U2337 ( .A(dataIn_EAST[21]), .Y(n2464) );
  INVX2TS U2338 ( .A(dataIn_EAST[22]), .Y(n2466) );
  INVX2TS U2339 ( .A(dataIn_EAST[23]), .Y(n2468) );
  INVX2TS U2340 ( .A(dataIn_EAST[24]), .Y(n2470) );
  INVX2TS U2341 ( .A(dataIn_EAST[25]), .Y(n2472) );
  INVX2TS U2342 ( .A(dataIn_EAST[26]), .Y(n2474) );
  INVX2TS U2343 ( .A(dataIn_EAST[27]), .Y(n2476) );
  INVX2TS U2344 ( .A(dataIn_EAST[28]), .Y(n2478) );
  INVX2TS U2345 ( .A(dataIn_EAST[29]), .Y(n2480) );
  INVX2TS U2346 ( .A(dataIn_EAST[30]), .Y(n2482) );
  INVX2TS U2347 ( .A(dataIn_EAST[31]), .Y(n2484) );
  NOR2BX1TS U2348 ( .AN(n2094), .B(n2204), .Y(n3378) );
  OAI2BB1X1TS U2349 ( .A0N(requesterAddressOut_EAST[0]), .A1N(n69), .B0(n1748), 
        .Y(n3172) );
  AOI22X1TS U2350 ( .A0(n1742), .A1(prevRequesterAddress_A[0]), .B0(n1743), 
        .B1(prevRequesterAddress_B[0]), .Y(n1748) );
  OAI2BB1X1TS U2351 ( .A0N(requesterAddressOut_EAST[1]), .A1N(n1740), .B0(
        n1747), .Y(n3173) );
  AOI22X1TS U2352 ( .A0(n1742), .A1(prevRequesterAddress_A[1]), .B0(n1743), 
        .B1(prevRequesterAddress_B[1]), .Y(n1747) );
  OAI2BB1X1TS U2353 ( .A0N(requesterAddressOut_EAST[2]), .A1N(n69), .B0(n1746), 
        .Y(n3174) );
  AOI22X1TS U2354 ( .A0(n1742), .A1(prevRequesterAddress_A[2]), .B0(n1743), 
        .B1(prevRequesterAddress_B[2]), .Y(n1746) );
  OAI2BB1X1TS U2355 ( .A0N(requesterAddressOut_EAST[3]), .A1N(n1740), .B0(
        n1745), .Y(n3175) );
  AOI22X1TS U2356 ( .A0(n350), .A1(prevRequesterAddress_A[3]), .B0(n358), .B1(
        prevRequesterAddress_B[3]), .Y(n1745) );
  OAI2BB1X1TS U2357 ( .A0N(requesterAddressOut_EAST[4]), .A1N(n69), .B0(n1744), 
        .Y(n3176) );
  AOI22X1TS U2358 ( .A0(n350), .A1(prevRequesterAddress_A[4]), .B0(n358), .B1(
        prevRequesterAddress_B[4]), .Y(n1744) );
  OAI2BB1X1TS U2359 ( .A0N(requesterAddressOut_EAST[5]), .A1N(n1740), .B0(
        n1741), .Y(n3177) );
  AOI22X1TS U2360 ( .A0(n350), .A1(prevRequesterAddress_A[5]), .B0(n358), .B1(
        prevRequesterAddress_B[5]), .Y(n1741) );
  NOR2X1TS U2361 ( .A(n2008), .B(n2193), .Y(n3416) );
  NOR2X1TS U2362 ( .A(n2009), .B(n2193), .Y(n3415) );
  NOR2X1TS U2363 ( .A(n2010), .B(n2193), .Y(n3414) );
  NOR2X1TS U2364 ( .A(n2011), .B(n2193), .Y(n3413) );
  NOR2X1TS U2365 ( .A(n2012), .B(n2194), .Y(n3412) );
  NOR2X1TS U2366 ( .A(n2013), .B(n2194), .Y(n3411) );
  NOR2X1TS U2367 ( .A(n2015), .B(n2194), .Y(n3410) );
  NOR2X1TS U2368 ( .A(n2017), .B(n2194), .Y(n3409) );
  NOR2X1TS U2369 ( .A(n2019), .B(n2195), .Y(n3408) );
  NOR2X1TS U2370 ( .A(n2021), .B(n2195), .Y(n3407) );
  NOR2X1TS U2371 ( .A(n2023), .B(n2198), .Y(n3406) );
  NOR2X1TS U2372 ( .A(n2025), .B(n2195), .Y(n3405) );
  NOR2X1TS U2373 ( .A(n2027), .B(n2195), .Y(n3404) );
  NOR2X1TS U2374 ( .A(n2029), .B(n2196), .Y(n3403) );
  NOR2X1TS U2375 ( .A(n2031), .B(n2196), .Y(n3402) );
  NOR2X1TS U2376 ( .A(n2033), .B(n2196), .Y(n3401) );
  NOR2X1TS U2377 ( .A(n2035), .B(n2196), .Y(n3400) );
  NOR2X1TS U2378 ( .A(n2037), .B(n2197), .Y(n3399) );
  NOR2X1TS U2379 ( .A(n2039), .B(n2197), .Y(n3398) );
  NOR2X1TS U2380 ( .A(n2041), .B(n2197), .Y(n3397) );
  NOR2X1TS U2381 ( .A(n2043), .B(n2197), .Y(n3396) );
  NOR2X1TS U2382 ( .A(n2045), .B(n2198), .Y(n3395) );
  NOR2X1TS U2383 ( .A(n2047), .B(n2198), .Y(n3394) );
  NOR2X1TS U2384 ( .A(n2049), .B(n2198), .Y(n3393) );
  NOR2X1TS U2385 ( .A(n2051), .B(n2199), .Y(n3392) );
  NOR2X1TS U2386 ( .A(n2053), .B(n2199), .Y(n3391) );
  NOR2X1TS U2387 ( .A(n2055), .B(n2199), .Y(n3390) );
  NOR2X1TS U2388 ( .A(n2057), .B(n2199), .Y(n3389) );
  NOR2X1TS U2389 ( .A(n2059), .B(n2200), .Y(n3388) );
  NOR2X1TS U2390 ( .A(n2061), .B(n2200), .Y(n3387) );
  NOR2X1TS U2391 ( .A(n2063), .B(n2200), .Y(n3386) );
  NOR2X1TS U2392 ( .A(n2065), .B(n2201), .Y(n3285) );
  NOR2X1TS U2393 ( .A(n2067), .B(n2200), .Y(n3284) );
  NOR2X1TS U2394 ( .A(n2069), .B(n2201), .Y(n3283) );
  NOR2X1TS U2395 ( .A(n2071), .B(n2202), .Y(n3282) );
  NOR2X1TS U2396 ( .A(n2073), .B(n2201), .Y(n3281) );
  NOR2X1TS U2397 ( .A(n2075), .B(n2202), .Y(n3280) );
  NOR2X1TS U2398 ( .A(n2077), .B(n2201), .Y(n3279) );
  NOR2X1TS U2399 ( .A(n2079), .B(n2203), .Y(n3278) );
  NOR2X1TS U2400 ( .A(n2007), .B(n2192), .Y(n3417) );
  INVX2TS U2401 ( .A(cacheAddressIn_EAST[0]), .Y(n2280) );
  INVX2TS U2402 ( .A(cacheAddressIn_WEST[0]), .Y(n2297) );
  INVX2TS U2403 ( .A(cacheAddressIn_EAST[1]), .Y(n2282) );
  INVX2TS U2404 ( .A(cacheAddressIn_WEST[1]), .Y(n2300) );
  INVX2TS U2405 ( .A(cacheAddressIn_EAST[2]), .Y(n2284) );
  INVX2TS U2406 ( .A(cacheAddressIn_WEST[2]), .Y(n2303) );
  INVX2TS U2407 ( .A(cacheAddressIn_EAST[3]), .Y(n2286) );
  INVX2TS U2408 ( .A(cacheAddressIn_WEST[3]), .Y(n2306) );
  INVX2TS U2409 ( .A(cacheAddressIn_EAST[4]), .Y(n2288) );
  INVX2TS U2410 ( .A(cacheAddressIn_WEST[4]), .Y(n2309) );
  INVX2TS U2411 ( .A(cacheAddressIn_EAST[5]), .Y(n2290) );
  INVX2TS U2412 ( .A(cacheAddressIn_WEST[5]), .Y(n2312) );
  INVX2TS U2413 ( .A(cacheAddressIn_EAST[6]), .Y(n2292) );
  INVX2TS U2414 ( .A(cacheAddressIn_EAST[7]), .Y(n2294) );
  INVX2TS U2415 ( .A(dataIn_WEST[0]), .Y(n2327) );
  INVX2TS U2416 ( .A(dataIn_WEST[1]), .Y(n2330) );
  INVX2TS U2417 ( .A(dataIn_WEST[2]), .Y(n2333) );
  INVX2TS U2418 ( .A(dataIn_WEST[3]), .Y(n2336) );
  INVX2TS U2419 ( .A(dataIn_WEST[4]), .Y(n2339) );
  INVX2TS U2420 ( .A(dataIn_WEST[5]), .Y(n2342) );
  INVX2TS U2421 ( .A(dataIn_WEST[6]), .Y(n2345) );
  INVX2TS U2422 ( .A(dataIn_WEST[7]), .Y(n2348) );
  INVX2TS U2423 ( .A(dataIn_WEST[8]), .Y(n2351) );
  INVX2TS U2424 ( .A(dataIn_WEST[9]), .Y(n2354) );
  INVX2TS U2425 ( .A(dataIn_WEST[10]), .Y(n2357) );
  INVX2TS U2426 ( .A(dataIn_WEST[11]), .Y(n2360) );
  INVX2TS U2427 ( .A(dataIn_WEST[12]), .Y(n2363) );
  INVX2TS U2428 ( .A(dataIn_WEST[13]), .Y(n2366) );
  INVX2TS U2429 ( .A(dataIn_WEST[14]), .Y(n2369) );
  INVX2TS U2430 ( .A(dataIn_WEST[15]), .Y(n2372) );
  INVX2TS U2431 ( .A(dataIn_WEST[16]), .Y(n2375) );
  INVX2TS U2432 ( .A(dataIn_WEST[17]), .Y(n2378) );
  INVX2TS U2433 ( .A(dataIn_WEST[18]), .Y(n2381) );
  INVX2TS U2434 ( .A(dataIn_WEST[19]), .Y(n2384) );
  INVX2TS U2435 ( .A(dataIn_WEST[20]), .Y(n2387) );
  INVX2TS U2436 ( .A(dataIn_WEST[21]), .Y(n2390) );
  INVX2TS U2437 ( .A(dataIn_WEST[22]), .Y(n2393) );
  INVX2TS U2438 ( .A(dataIn_WEST[23]), .Y(n2396) );
  INVX2TS U2439 ( .A(dataIn_WEST[24]), .Y(n2399) );
  INVX2TS U2440 ( .A(dataIn_WEST[25]), .Y(n2402) );
  INVX2TS U2441 ( .A(dataIn_WEST[26]), .Y(n2405) );
  INVX2TS U2442 ( .A(dataIn_WEST[27]), .Y(n2408) );
  INVX2TS U2443 ( .A(dataIn_WEST[28]), .Y(n2411) );
  INVX2TS U2444 ( .A(dataIn_WEST[29]), .Y(n2414) );
  INVX2TS U2445 ( .A(dataIn_WEST[30]), .Y(n2417) );
  INVX2TS U2446 ( .A(dataIn_WEST[31]), .Y(n2420) );
  INVX2TS U2447 ( .A(n1418), .Y(n758) );
  AOI32X1TS U2448 ( .A0(n2094), .A1(n2496), .A2(n1129), .B0(n759), .B1(n2093), 
        .Y(n1418) );
  INVX2TS U2449 ( .A(n1129), .Y(n759) );
  INVX2TS U2450 ( .A(n1126), .Y(n652) );
  AOI32X1TS U2451 ( .A0(\requesterPortBuffer[4][0] ), .A1(n2501), .A2(n1127), 
        .B0(n811), .B1(\requesterPortBuffer[2][0] ), .Y(n1126) );
  INVX2TS U2452 ( .A(n1124), .Y(n651) );
  AOI32X1TS U2453 ( .A0(\requesterPortBuffer[6][0] ), .A1(n2498), .A2(n1125), 
        .B0(n756), .B1(\requesterPortBuffer[4][0] ), .Y(n1124) );
  INVX2TS U2454 ( .A(n1417), .Y(n814) );
  AOI32X1TS U2455 ( .A0(n2093), .A1(n2497), .A2(n1130), .B0(n86), .B1(n2091), 
        .Y(n1417) );
  INVX2TS U2456 ( .A(n1133), .Y(n656) );
  AOI32X1TS U2457 ( .A0(\requesterPortBuffer[0][0] ), .A1(n2500), .A2(n42), 
        .B0(\requesterPortBuffer[6][0] ), .B1(n754), .Y(n1133) );
  OAI32X1TS U2458 ( .A0(n650), .A1(n2490), .A2(n812), .B0(n2096), .B1(n1122), 
        .Y(n2098) );
  OAI32X1TS U2459 ( .A0(n653), .A1(n2492), .A2(n880), .B0(n2081), .B1(n87), 
        .Y(n2101) );
  OAI32X1TS U2460 ( .A0(n654), .A1(n2492), .A2(n99), .B0(n2083), .B1(n1130), 
        .Y(n2103) );
  NAND2X1TS U2461 ( .A(n57), .B(n98), .Y(n1416) );
  NOR3X1TS U2462 ( .A(n1148), .B(n910), .C(n53), .Y(n1691) );
  INVX2TS U2463 ( .A(cacheDataOut_A[0]), .Y(n1089) );
  INVX2TS U2464 ( .A(cacheDataOut_A[1]), .Y(n1088) );
  INVX2TS U2465 ( .A(cacheDataOut_A[2]), .Y(n1087) );
  INVX2TS U2466 ( .A(cacheDataOut_A[3]), .Y(n1086) );
  INVX2TS U2467 ( .A(cacheDataOut_A[4]), .Y(n1085) );
  INVX2TS U2468 ( .A(cacheDataOut_A[5]), .Y(n1084) );
  INVX2TS U2469 ( .A(cacheDataOut_A[6]), .Y(n1083) );
  INVX2TS U2470 ( .A(cacheDataOut_A[7]), .Y(n1082) );
  INVX2TS U2471 ( .A(cacheDataOut_A[8]), .Y(n1081) );
  INVX2TS U2472 ( .A(cacheDataOut_A[9]), .Y(n1080) );
  INVX2TS U2473 ( .A(cacheDataOut_A[10]), .Y(n1079) );
  INVX2TS U2474 ( .A(cacheDataOut_A[11]), .Y(n1078) );
  INVX2TS U2475 ( .A(cacheDataOut_A[12]), .Y(n1077) );
  INVX2TS U2476 ( .A(cacheDataOut_A[13]), .Y(n1076) );
  INVX2TS U2477 ( .A(cacheDataOut_A[14]), .Y(n1075) );
  INVX2TS U2478 ( .A(cacheDataOut_A[15]), .Y(n1074) );
  INVX2TS U2479 ( .A(cacheDataOut_A[16]), .Y(n1073) );
  INVX2TS U2480 ( .A(cacheDataOut_A[17]), .Y(n1072) );
  INVX2TS U2481 ( .A(cacheDataOut_A[18]), .Y(n1071) );
  INVX2TS U2482 ( .A(cacheDataOut_A[19]), .Y(n1070) );
  INVX2TS U2483 ( .A(cacheDataOut_A[20]), .Y(n1069) );
  INVX2TS U2484 ( .A(cacheDataOut_A[21]), .Y(n1068) );
  INVX2TS U2485 ( .A(cacheDataOut_A[22]), .Y(n1067) );
  INVX2TS U2486 ( .A(cacheDataOut_A[23]), .Y(n1066) );
  INVX2TS U2487 ( .A(cacheDataOut_A[24]), .Y(n1065) );
  INVX2TS U2488 ( .A(cacheDataOut_A[25]), .Y(n1064) );
  INVX2TS U2489 ( .A(cacheDataOut_A[26]), .Y(n1063) );
  INVX2TS U2490 ( .A(cacheDataOut_A[27]), .Y(n1062) );
  INVX2TS U2491 ( .A(cacheDataOut_A[28]), .Y(n1061) );
  INVX2TS U2492 ( .A(cacheDataOut_A[29]), .Y(n1060) );
  INVX2TS U2493 ( .A(cacheDataOut_A[30]), .Y(n1059) );
  INVX2TS U2494 ( .A(cacheDataOut_A[31]), .Y(n1058) );
  INVX2TS U2495 ( .A(cacheDataOut_B[0]), .Y(n1121) );
  INVX2TS U2496 ( .A(cacheDataOut_B[1]), .Y(n1120) );
  INVX2TS U2497 ( .A(cacheDataOut_B[2]), .Y(n1119) );
  INVX2TS U2498 ( .A(cacheDataOut_B[3]), .Y(n1118) );
  INVX2TS U2499 ( .A(cacheDataOut_B[4]), .Y(n1117) );
  INVX2TS U2500 ( .A(cacheDataOut_B[5]), .Y(n1116) );
  INVX2TS U2501 ( .A(cacheDataOut_B[6]), .Y(n1115) );
  INVX2TS U2502 ( .A(cacheDataOut_B[7]), .Y(n1114) );
  INVX2TS U2503 ( .A(cacheDataOut_B[8]), .Y(n1113) );
  INVX2TS U2504 ( .A(cacheDataOut_B[9]), .Y(n1112) );
  INVX2TS U2505 ( .A(cacheDataOut_B[10]), .Y(n1111) );
  INVX2TS U2506 ( .A(cacheDataOut_B[11]), .Y(n1110) );
  INVX2TS U2507 ( .A(cacheDataOut_B[12]), .Y(n1109) );
  INVX2TS U2508 ( .A(cacheDataOut_B[13]), .Y(n1108) );
  INVX2TS U2509 ( .A(cacheDataOut_B[14]), .Y(n1107) );
  INVX2TS U2510 ( .A(cacheDataOut_B[15]), .Y(n1106) );
  INVX2TS U2511 ( .A(cacheDataOut_B[16]), .Y(n1105) );
  INVX2TS U2512 ( .A(cacheDataOut_B[17]), .Y(n1104) );
  INVX2TS U2513 ( .A(cacheDataOut_B[18]), .Y(n1103) );
  INVX2TS U2514 ( .A(cacheDataOut_B[19]), .Y(n1102) );
  INVX2TS U2515 ( .A(cacheDataOut_B[20]), .Y(n1101) );
  INVX2TS U2516 ( .A(cacheDataOut_B[21]), .Y(n1100) );
  INVX2TS U2517 ( .A(cacheDataOut_B[22]), .Y(n1099) );
  INVX2TS U2518 ( .A(cacheDataOut_B[23]), .Y(n1098) );
  INVX2TS U2519 ( .A(cacheDataOut_B[24]), .Y(n1097) );
  INVX2TS U2520 ( .A(cacheDataOut_B[25]), .Y(n1096) );
  INVX2TS U2521 ( .A(cacheDataOut_B[26]), .Y(n1095) );
  INVX2TS U2522 ( .A(cacheDataOut_B[27]), .Y(n1094) );
  INVX2TS U2523 ( .A(cacheDataOut_B[28]), .Y(n1093) );
  INVX2TS U2524 ( .A(cacheDataOut_B[29]), .Y(n1092) );
  INVX2TS U2525 ( .A(cacheDataOut_B[30]), .Y(n1091) );
  INVX2TS U2526 ( .A(cacheDataOut_B[31]), .Y(n1090) );
endmodule


module outputPortArbiter_0 ( clk, reset, selectBit_NORTH, 
        destinationAddressIn_NORTH, requesterAddressIn_NORTH, readIn_NORTH, 
        writeIn_NORTH, dataIn_NORTH, selectBit_SOUTH, 
        destinationAddressIn_SOUTH, requesterAddressIn_SOUTH, readIn_SOUTH, 
        writeIn_SOUTH, dataIn_SOUTH, selectBit_EAST, destinationAddressIn_EAST, 
        requesterAddressIn_EAST, readIn_EAST, writeIn_EAST, dataIn_EAST, 
        selectBit_WEST, destinationAddressIn_WEST, requesterAddressIn_WEST, 
        readIn_WEST, dataIn_WEST, readReady, readRequesterAddress, 
        cacheDataOut, destinationAddressOut, requesterAddressOut, readOut, 
        writeOut, dataOut, writeIn_WEST_BAR );
  input [13:0] destinationAddressIn_NORTH;
  input [5:0] requesterAddressIn_NORTH;
  input [31:0] dataIn_NORTH;
  input [13:0] destinationAddressIn_SOUTH;
  input [5:0] requesterAddressIn_SOUTH;
  input [31:0] dataIn_SOUTH;
  input [13:0] destinationAddressIn_EAST;
  input [5:0] requesterAddressIn_EAST;
  input [31:0] dataIn_EAST;
  input [13:0] destinationAddressIn_WEST;
  input [5:0] requesterAddressIn_WEST;
  input [31:0] dataIn_WEST;
  input [5:0] readRequesterAddress;
  input [31:0] cacheDataOut;
  output [13:0] destinationAddressOut;
  output [5:0] requesterAddressOut;
  output [31:0] dataOut;
  input clk, reset, selectBit_NORTH, readIn_NORTH, writeIn_NORTH,
         selectBit_SOUTH, readIn_SOUTH, writeIn_SOUTH, selectBit_EAST,
         readIn_EAST, writeIn_EAST, selectBit_WEST, readIn_WEST, readReady,
         writeIn_WEST_BAR;
  output readOut, writeOut;
  wire   writeIn_WEST, n2486, n2484, n2482, n2480, n2457, n2455, n2453, n2485,
         n2483, n2481, n2458, n2454, n2479, n2456, n2452, n2499, n2496, n2493,
         n2528, n2527, n2526, n2525, n2524, n2523, n2522, n2521, n2498, n2497,
         n2494, n2500, n2495, n2541, n2540, n2537, n2535, n2511, n2507, n2542,
         n2539, n2538, n2536, n2514, n2513, n2512, n2510, n2509, n2508, n2703,
         n2692, n2691, n2689, n2706, n2705, n2700, n2698, n2696, n2695, n2694,
         n2690, n2687, n2686, n2685, n2684, n2677, n2675, n2704, n2702, n2701,
         n2699, n2697, n2693, n2688, n2683, n2682, n2681, n2680, n2679, n2678,
         n2676, n2520, n2519, n2518, n2517, n2516, n2515, n2672, n2671, n2670,
         n2669, n2668, n2667, n2666, n2665, n2664, n2662, n2661, n2660, n2657,
         n2656, n2655, n2654, n2653, n2652, n2651, n2650, n2649, n2648, n2647,
         n2646, n2645, n2644, n2534, n2533, n2532, n2531, n2530, n2529, n2673,
         n2663, n2659, n2658, n2643, n2850, \requesterAddressbuffer[2][2] ,
         n2849, \requesterAddressbuffer[2][3] , n2847,
         \requesterAddressbuffer[2][5] , n2840, \requesterAddressbuffer[0][0] ,
         n2839, \requesterAddressbuffer[0][1] , n2838,
         \requesterAddressbuffer[0][2] , n2836, \requesterAddressbuffer[0][4] ,
         n2852, \requesterAddressbuffer[2][0] , n2851,
         \requesterAddressbuffer[2][1] , n2848, \requesterAddressbuffer[2][4] ,
         n2837, \requesterAddressbuffer[0][3] , n2835,
         \requesterAddressbuffer[0][5] , n2566, \readOutbuffer[2] ,
         readOutbuffer_7, n2569, n2568, n2564, n2870, n2869, n2868, n2867,
         n2866, n2865, n2576, n2860, n2859, n2864, n2863, n2862, n2861, n2573,
         n2731, n2968, n2770, n2768, n2764, n2754, n2748, n2746, n2739, n2834,
         n2833, n2832, n2829, n2825, n2814, n2811, n2807, n2806, n2736, n2924,
         n2734, n2944, n2733, n99, n2725, n98, n2723, n97, n2720, n96, n2718,
         n95, n2715, n94, n2713, n93, n2504, n92, n2769, n2760, n2743, n2492,
         n2491, n2489, n2488, n2487, n2464, n91, n2460, n90, n2738, n89, n2737,
         n88, n2735, n87, n2732, n86, n2730, n85, n2729, n84, n2728, n83,
         n2727, n82, n2726, n81, n2724, n80, n2722, n79, n2721, n78, n2719,
         n77, n2717, n76, n2716, n75, n2714, n74, n2712, n73, n2711, n72,
         n2710, n71, n2709, n70, n2708, n69, n2707, n68, n2506, n67, n2505,
         n66, n2503, n65, n2502, n64, n2501, n63, n2767, n2766, n2765, n2763,
         n2762, n2761, n2759, n2758, n2757, n2756, n2755, n2753, n2752, n2751,
         n2750, n2749, n2747, n2745, n2744, n2742, n2741, n2740, n2490, n2831,
         n62, n2830, n61, n2828, n60, n2827, n59, n2826, n58, n2824, n57,
         n2823, n56, n2822, n55, n2821, n54, n2820, n53, n2819, n52, n2818,
         n51, n2817, n50, n2816, n49, n2815, n48, n2813, n47, n2812, n46,
         n2810, n45, n2809, n44, n2808, n43, n2805, n42, n2804, n41, n2803,
         n40, n2463, n39, n2462, n38, n2461, n37, n2459, n36, n2571, n2574,
         n2577, n2575, n2570, n2565, n2567, n2889, N4718, n2285, n2288, n2434,
         n2284, n2431, n2283, n2450, n2286, n2440, n2361, n2439, n2370, n2438,
         n2379, n2437, n2388, n2436, n2890, n2435, n2899, n2433, n2900, n2432,
         n2901, n2430, n2902, n2429, n2903, n2428, n2912, n2427, n2921, n2426,
         n2930, n2425, n2939, n2424, n2948, n2423, n2957, n2422, n2966, n2421,
         n2975, n2420, n2984, n2419, n2993, n2418, n3002, n2417, n3011, n2416,
         n3020, n2415, n3029, n2414, n3038, n2413, n3047, n2412, n3056, n2411,
         n3065, n2410, n3074, n2409, n3083, n2408, n3092, n2407, n3101, n2406,
         n3110, n2405, n3119, n2404, n3128, n2403, n3137, n2402, n3146, n2401,
         n3155, n2400, n3164, n2399, n3173, n2398, n3182, n2397, n3191, n2448,
         n2447, n2446, n2445, n2444, n2443, n2442, n2441, n2549, n2472, n2471,
         n2470, n2469, n2468, n2467, n2466, n2558, n2802, n2610, n2609, n2608,
         n2607, n2606, n2605, n2604, n2603, n2602, n2601, n2600, n2599, n2598,
         n2597, n2596, n2595, n2594, n2593, n2592, n2591, n2590, n2589, n2588,
         n2587, n2586, n2585, n2584, n2583, n2582, n2581, n2580, n2579, n2561,
         n2560, n2559, n2557, n2801, n2799, n2798, n2796, n2795, n2793, n2791,
         n2790, n2789, n2788, n2787, n2786, n2785, n2784, n2781, n2779, n2778,
         n2777, n2776, n2774, n2773, n2772, n2771, n2478, n2477, n2476, n2475,
         n2473, n2562, n2548, n2547, n2546, n2545, n2543, n2800, n2797, n2794,
         n2792, n2783, n2782, n2780, n2775, n2544, n2552, n593, n2474, n2858,
         \requesterAddressbuffer[3][0] , n2857, \requesterAddressbuffer[3][1] ,
         n2856, \requesterAddressbuffer[3][2] , n2855,
         \requesterAddressbuffer[3][3] , n2853, \requesterAddressbuffer[3][5] ,
         n2854, \requesterAddressbuffer[3][4] , n2875,
         \requesterAddressbuffer[6][1] , n2874, \requesterAddressbuffer[6][2] ,
         n2873, \requesterAddressbuffer[6][3] , n2872,
         \requesterAddressbuffer[6][4] , n2871, \requesterAddressbuffer[6][5] ,
         n2876, \requesterAddressbuffer[6][0] , n2578, n2882, n2881, n2879,
         n2880, n2878, n2877, n2563, n2846, n2845, n2844, n2843, n2842, n2841,
         n2556, n2555, n2554, n2551, n2553, n2572, n2883, n459, n2884, n8,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2550, n2465, n2885, n2888, n5327, n2887, n6, n2886,
         n2451, n2674, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n757, n758, n759, n760, n761, n762,
         n764, n766, n767, n769, n771, n773, n774, n775, n777, n780, n784,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n936, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n960, n966, n967, n969, n970, n972, n979, n980, n981, n982,
         n996, n1029, n1084, n1130, n1131, n1132, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1798, n1799, n1800, n1801, n1802, n1804, n1805,
         n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
         n1817, n1818, n1819, n1820, n1821, n1822, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2287,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2360, n2362, n2363, n2364, n2365, n2367, n2368, n2369, n2371, n2373,
         n2374, n2375, n2376, n2377, n2378, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2449,
         n2891, n2892, n2893, n2894, n2896, n2897, n2898, n2904, n2905, n2906,
         n2908, n2910, n2911, n2915, n2916, n2917, n2918, n2919, n2920, n2922,
         n2926, n2927, n2928, n2929, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2940, n2941, n2942, n2943, n2946, n2947, n2949, n2951, n2953,
         n2954, n2955, n2956, n2958, n2960, n2962, n2963, n2964, n2965, n2967,
         n2969, n2970, n2971, n2972, n2973, n2976, n2977, n2978, n2980, n2981,
         n2982, n2983, n2987, n2988, n2989, n2990, n2991, n2994, n2995, n2997,
         n2998, n2999, n3000, n3001, n3003, n3005, n3006, n3007, n3008, n3009,
         n3010, n3012, n3013, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
         n3039, n3040, n3041, n3042, n3043, n3045, n3046, n3048, n3050, n3051,
         n3052, n3053, n3054, n3055, n3057, n3058, n3059, n3061, n3062, n3063,
         n3064, n3066, n3067, n3068, n3070, n3071, n3072, n3073, n3075, n3076,
         n3077, n3078, n3079, n3080, n3081, n3084, n3086, n3088, n3089, n3090,
         n3091, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3102, n3104,
         n3105, n3106, n3107, n3108, n3109, n3111, n3113, n3115, n3116, n3117,
         n3118, n3120, n3122, n3123, n3124, n3125, n3126, n3127, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3141, n3142, n3144, n3145, n3149,
         n3150, n3151, n3152, n3153, n3154, n3156, n3158, n3159, n3160, n3162,
         n3163, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3174, n3175,
         n3176, n3177, n3178, n3180, n3181, n3183, n3185, n3186, n3187, n3188,
         n3189, n3190, n3192, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n1, n2, n3,
         n4, n5, n7, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n710, n755,
         n756, n763, n765, n768, n770, n772, n776, n778, n779, n781, n782,
         n783, n785, n786, n787, n899, n900, n935, n937, n938, n959, n961,
         n962, n963, n964, n965, n968, n971, n973, n974, n975, n976, n977,
         n978, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1133, n1153, n1180, n1197, n1213, n1244, n1660,
         n1797, n1803, n1806, n1823, n1845, n1891, n1916, n2033, n2057, n2155,
         n2359, n2366, n2372, n2380, n2389, n2895, n2907, n2909, n2913, n2914,
         n2923, n2925, n2938, n2945, n2950, n2952, n2959, n2961, n2974, n2979,
         n2985, n2986, n2992, n2996, n3004, n3014, n3015, n3016, n3017, n3018,
         n3019, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3037,
         n3044, n3049, n3060, n3069, n3082, n3085, n3087, n3100, n3103, n3112,
         n3114, n3121, n3136, n3138, n3139, n3140, n3143, n3147, n3148, n3157,
         n3161, n3172, n3179, n3184, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504;
  assign writeIn_WEST = writeIn_WEST_BAR;

  DFFNSRX2TS \dataoutbuffer_reg[4][3]  ( .D(n2703), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3111) );
  DFFNSRX2TS \dataoutbuffer_reg[4][14]  ( .D(n2692), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3080) );
  DFFNSRX2TS \dataoutbuffer_reg[4][15]  ( .D(n2691), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3078) );
  DFFNSRX2TS \dataoutbuffer_reg[4][17]  ( .D(n2689), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3073) );
  DFFNSRX2TS \dataoutbuffer_reg[4][0]  ( .D(n2706), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3120) );
  DFFNSRX2TS \dataoutbuffer_reg[4][1]  ( .D(n2705), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3117) );
  DFFNSRX2TS \dataoutbuffer_reg[4][6]  ( .D(n2700), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3104) );
  DFFNSRX2TS \dataoutbuffer_reg[4][8]  ( .D(n2698), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3097) );
  DFFNSRX2TS \dataoutbuffer_reg[4][10]  ( .D(n2696), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3093) );
  DFFNSRX2TS \dataoutbuffer_reg[4][11]  ( .D(n2695), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3090) );
  DFFNSRX2TS \dataoutbuffer_reg[4][12]  ( .D(n2694), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3088) );
  DFFNSRX2TS \dataoutbuffer_reg[4][16]  ( .D(n2690), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3076) );
  DFFNSRX2TS \dataoutbuffer_reg[4][19]  ( .D(n2687), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3068) );
  DFFNSRX2TS \dataoutbuffer_reg[4][20]  ( .D(n2686), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3066) );
  DFFNSRX2TS \dataoutbuffer_reg[4][21]  ( .D(n2685), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3063) );
  DFFNSRX2TS \dataoutbuffer_reg[4][22]  ( .D(n2684), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3061) );
  DFFNSRX2TS \dataoutbuffer_reg[4][29]  ( .D(n2677), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3042) );
  DFFNSRX2TS \dataoutbuffer_reg[4][31]  ( .D(n2675), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3036) );
  DFFNSRX2TS \dataoutbuffer_reg[4][2]  ( .D(n2704), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3115) );
  DFFNSRX2TS \dataoutbuffer_reg[4][4]  ( .D(n2702), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3108) );
  DFFNSRX2TS \dataoutbuffer_reg[4][5]  ( .D(n2701), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3106) );
  DFFNSRX2TS \dataoutbuffer_reg[4][7]  ( .D(n2699), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3099) );
  DFFNSRX2TS \dataoutbuffer_reg[4][9]  ( .D(n2697), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3095) );
  DFFNSRX2TS \dataoutbuffer_reg[4][13]  ( .D(n2693), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3084) );
  DFFNSRX2TS \dataoutbuffer_reg[4][18]  ( .D(n2688), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3071) );
  DFFNSRX2TS \dataoutbuffer_reg[4][23]  ( .D(n2683), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3058) );
  DFFNSRX2TS \dataoutbuffer_reg[4][24]  ( .D(n2682), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3055) );
  DFFNSRX2TS \dataoutbuffer_reg[4][25]  ( .D(n2681), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3053) );
  DFFNSRX2TS \dataoutbuffer_reg[4][26]  ( .D(n2680), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3051) );
  DFFNSRX2TS \dataoutbuffer_reg[4][27]  ( .D(n2679), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3048) );
  DFFNSRX2TS \dataoutbuffer_reg[4][28]  ( .D(n2678), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3045) );
  DFFNSRX2TS \dataoutbuffer_reg[4][30]  ( .D(n2676), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3040) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][0]  ( .D(n2520), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3134) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][1]  ( .D(n2519), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3132) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][2]  ( .D(n2518), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3130) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][3]  ( .D(n2517), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3127) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][4]  ( .D(n2516), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3125) );
  DFFNSRX2TS \destinationAddressbuffer_reg[4][5]  ( .D(n2515), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3123) );
  DFFNSRX2TS \writeOutbuffer_reg[3]  ( .D(n2574), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n748) );
  DFFNSRX2TS \writeOutbuffer_reg[1]  ( .D(n2572), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n898) );
  DFFNSRX2TS \dataoutbuffer_reg[3][7]  ( .D(n2731), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n661), .QN(n2968) );
  DFFNSRX2TS \dataoutbuffer_reg[3][2]  ( .D(n2736), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n678), .QN(n2924) );
  DFFNSRX2TS \dataoutbuffer_reg[3][4]  ( .D(n2734), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n679), .QN(n2944) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][7]  ( .D(n2499), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3315), .QN(n578) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][8]  ( .D(n2498), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3313), .QN(n589) );
  DFFNSRX2TS \destinationAddressbuffer_reg[3][6]  ( .D(n2500), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3317), .QN(n592) );
  DFFNSRX2TS \destinationAddressbuffer_reg[1][6]  ( .D(n2472), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3279), .QN(n789) );
  DFFNSRX2TS \destinationAddressbuffer_reg[1][7]  ( .D(n2471), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3278), .QN(n790) );
  DFFNSRX2TS \destinationAddressbuffer_reg[1][8]  ( .D(n2470), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3277), .QN(n791) );
  DFFNSRX2TS \destinationAddressbuffer_reg[1][9]  ( .D(n2469), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3276), .QN(n792) );
  DFFNSRX2TS \destinationAddressbuffer_reg[1][10]  ( .D(n2468), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3275), .QN(n793) );
  DFFNSRX2TS \destinationAddressbuffer_reg[1][11]  ( .D(n2467), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3274), .QN(n794) );
  DFFNSRX2TS \destinationAddressbuffer_reg[1][12]  ( .D(n2466), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3273), .QN(n795) );
  DFFNSRX2TS \destinationAddressbuffer_reg[1][13]  ( .D(n2465), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3272), .QN(n934) );
  DFFNSRX2TS empty_reg_reg ( .D(n2885), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        n13), .QN(n443) );
  DFFNSRX2TS \read_reg_reg[2]  ( .D(n2884), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n8), .QN(n440) );
  DFFNSRX2TS \read_reg_reg[0]  ( .D(n2889), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n11), .QN(n430) );
  DFFNSRX2TS \read_reg_reg[1]  ( .D(n2883), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n12), .QN(n459) );
  DFFNSRX2TS \write_reg_reg[0]  ( .D(n2888), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n424), .QN(n5327) );
  DFFNSRX2TS \write_reg_reg[2]  ( .D(n2886), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n441), .QN(n10) );
  DFFNSRX2TS writeOut_reg ( .D(n659), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        writeOut), .QN(n2288) );
  DFFNSRX2TS \requesterAddressOut_reg[0]  ( .D(n2434), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[0]), .QN(n2284) );
  DFFNSRX2TS \requesterAddressOut_reg[3]  ( .D(n2431), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[3]), .QN(n2283) );
  DFFNSRX2TS readOut_reg ( .D(n2450), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        readOut), .QN(n2286) );
  DFFNSRX2TS \destinationAddressOut_reg[0]  ( .D(n2440), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[0]), .QN(n2361) );
  DFFNSRX2TS \destinationAddressOut_reg[1]  ( .D(n2439), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[1]), .QN(n2370) );
  DFFNSRX2TS \destinationAddressOut_reg[2]  ( .D(n2438), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[2]), .QN(n2379) );
  DFFNSRX2TS \destinationAddressOut_reg[3]  ( .D(n2437), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[3]), .QN(n2388) );
  DFFNSRX2TS \destinationAddressOut_reg[4]  ( .D(n2436), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[4]), .QN(n2890) );
  DFFNSRX2TS \destinationAddressOut_reg[5]  ( .D(n2435), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[5]), .QN(n2899) );
  DFFNSRX2TS \requesterAddressOut_reg[1]  ( .D(n2433), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[1]), .QN(n2900) );
  DFFNSRX2TS \requesterAddressOut_reg[2]  ( .D(n2432), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[2]), .QN(n2901) );
  DFFNSRX2TS \requesterAddressOut_reg[4]  ( .D(n2430), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[4]), .QN(n2902) );
  DFFNSRX2TS \requesterAddressOut_reg[5]  ( .D(n2429), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[5]), .QN(n2903) );
  DFFNSRX2TS \dataOut_reg[0]  ( .D(n2428), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[0]), .QN(n2912) );
  DFFNSRX2TS \dataOut_reg[1]  ( .D(n2427), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[1]), .QN(n2921) );
  DFFNSRX2TS \dataOut_reg[2]  ( .D(n2426), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[2]), .QN(n2930) );
  DFFNSRX2TS \dataOut_reg[3]  ( .D(n2425), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[3]), .QN(n2939) );
  DFFNSRX2TS \dataOut_reg[4]  ( .D(n2424), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[4]), .QN(n2948) );
  DFFNSRX2TS \dataOut_reg[5]  ( .D(n2423), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[5]), .QN(n2957) );
  DFFNSRX2TS \dataOut_reg[6]  ( .D(n2422), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[6]), .QN(n2966) );
  DFFNSRX2TS \dataOut_reg[7]  ( .D(n2421), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[7]), .QN(n2975) );
  DFFNSRX2TS \dataOut_reg[8]  ( .D(n2420), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[8]), .QN(n2984) );
  DFFNSRX2TS \dataOut_reg[9]  ( .D(n2419), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[9]), .QN(n2993) );
  DFFNSRX2TS \dataOut_reg[10]  ( .D(n2418), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[10]), .QN(n3002) );
  DFFNSRX2TS \dataOut_reg[11]  ( .D(n2417), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[11]), .QN(n3011) );
  DFFNSRX2TS \dataOut_reg[12]  ( .D(n2416), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[12]), .QN(n3020) );
  DFFNSRX2TS \dataOut_reg[13]  ( .D(n2415), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[13]), .QN(n3029) );
  DFFNSRX2TS \dataOut_reg[14]  ( .D(n2414), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[14]), .QN(n3038) );
  DFFNSRX2TS \dataOut_reg[15]  ( .D(n2413), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[15]), .QN(n3047) );
  DFFNSRX2TS \dataOut_reg[16]  ( .D(n2412), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[16]), .QN(n3056) );
  DFFNSRX2TS \dataOut_reg[17]  ( .D(n2411), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[17]), .QN(n3065) );
  DFFNSRX2TS \dataOut_reg[18]  ( .D(n2410), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[18]), .QN(n3074) );
  DFFNSRX2TS \dataOut_reg[19]  ( .D(n2409), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[19]), .QN(n3083) );
  DFFNSRX2TS \dataOut_reg[20]  ( .D(n2408), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[20]), .QN(n3092) );
  DFFNSRX2TS \dataOut_reg[21]  ( .D(n2407), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[21]), .QN(n3101) );
  DFFNSRX2TS \dataOut_reg[22]  ( .D(n2406), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[22]), .QN(n3110) );
  DFFNSRX2TS \dataOut_reg[23]  ( .D(n2405), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[23]), .QN(n3119) );
  DFFNSRX2TS \dataOut_reg[24]  ( .D(n2404), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[24]), .QN(n3128) );
  DFFNSRX2TS \dataOut_reg[25]  ( .D(n2403), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[25]), .QN(n3137) );
  DFFNSRX2TS \dataOut_reg[26]  ( .D(n2402), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[26]), .QN(n3146) );
  DFFNSRX2TS \dataOut_reg[27]  ( .D(n2401), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[27]), .QN(n3155) );
  DFFNSRX2TS \dataOut_reg[28]  ( .D(n2400), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[28]), .QN(n3164) );
  DFFNSRX2TS \dataOut_reg[29]  ( .D(n2399), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[29]), .QN(n3173) );
  DFFNSRX2TS \dataOut_reg[30]  ( .D(n2398), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[30]), .QN(n3182) );
  DFFNSRX2TS \dataOut_reg[31]  ( .D(n2397), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[31]), .QN(n3191) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][4]  ( .D(n2530), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n641) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][4]  ( .D(n2558), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n796) );
  DFFNSRXLTS \dataoutbuffer_reg[5][2]  ( .D(n2672), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n611) );
  DFFNSRXLTS \dataoutbuffer_reg[5][3]  ( .D(n2671), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n612) );
  DFFNSRXLTS \dataoutbuffer_reg[5][4]  ( .D(n2670), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n613) );
  DFFNSRXLTS \dataoutbuffer_reg[5][5]  ( .D(n2669), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n614) );
  DFFNSRXLTS \dataoutbuffer_reg[5][6]  ( .D(n2668), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n615) );
  DFFNSRXLTS \dataoutbuffer_reg[5][7]  ( .D(n2667), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n616) );
  DFFNSRXLTS \dataoutbuffer_reg[5][8]  ( .D(n2666), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n617) );
  DFFNSRXLTS \dataoutbuffer_reg[5][9]  ( .D(n2665), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n618) );
  DFFNSRXLTS \dataoutbuffer_reg[5][10]  ( .D(n2664), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n619) );
  DFFNSRXLTS \dataoutbuffer_reg[5][12]  ( .D(n2662), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n620) );
  DFFNSRXLTS \dataoutbuffer_reg[5][13]  ( .D(n2661), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n621) );
  DFFNSRXLTS \dataoutbuffer_reg[5][14]  ( .D(n2660), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n622) );
  DFFNSRXLTS \dataoutbuffer_reg[5][17]  ( .D(n2657), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n623) );
  DFFNSRXLTS \dataoutbuffer_reg[5][18]  ( .D(n2656), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n624) );
  DFFNSRXLTS \dataoutbuffer_reg[5][19]  ( .D(n2655), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n625) );
  DFFNSRXLTS \dataoutbuffer_reg[5][20]  ( .D(n2654), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n626) );
  DFFNSRXLTS \dataoutbuffer_reg[5][21]  ( .D(n2653), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n627) );
  DFFNSRXLTS \dataoutbuffer_reg[5][22]  ( .D(n2652), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n628) );
  DFFNSRXLTS \dataoutbuffer_reg[5][23]  ( .D(n2651), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n629) );
  DFFNSRXLTS \dataoutbuffer_reg[5][24]  ( .D(n2650), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n630) );
  DFFNSRXLTS \dataoutbuffer_reg[5][25]  ( .D(n2649), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n631) );
  DFFNSRXLTS \dataoutbuffer_reg[5][26]  ( .D(n2648), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n632) );
  DFFNSRXLTS \dataoutbuffer_reg[5][27]  ( .D(n2647), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n633) );
  DFFNSRXLTS \dataoutbuffer_reg[5][28]  ( .D(n2646), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n634) );
  DFFNSRXLTS \dataoutbuffer_reg[5][29]  ( .D(n2645), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n635) );
  DFFNSRXLTS \dataoutbuffer_reg[5][30]  ( .D(n2644), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n636) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][0]  ( .D(n2534), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n637) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][1]  ( .D(n2533), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n638) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][2]  ( .D(n2532), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n639) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][3]  ( .D(n2531), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n640) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][5]  ( .D(n2529), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n642) );
  DFFNSRXLTS \dataoutbuffer_reg[5][1]  ( .D(n2673), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n643) );
  DFFNSRXLTS \dataoutbuffer_reg[5][11]  ( .D(n2663), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n644) );
  DFFNSRXLTS \dataoutbuffer_reg[5][15]  ( .D(n2659), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n645) );
  DFFNSRXLTS \dataoutbuffer_reg[5][16]  ( .D(n2658), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n646) );
  DFFNSRXLTS \dataoutbuffer_reg[5][31]  ( .D(n2643), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n647) );
  DFFNSRXLTS \requesterAddressbuffer_reg[5][0]  ( .D(n2870), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n652) );
  DFFNSRXLTS \requesterAddressbuffer_reg[5][1]  ( .D(n2869), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n653) );
  DFFNSRXLTS \requesterAddressbuffer_reg[5][2]  ( .D(n2868), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n654) );
  DFFNSRXLTS \requesterAddressbuffer_reg[5][3]  ( .D(n2867), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n655) );
  DFFNSRXLTS \requesterAddressbuffer_reg[5][4]  ( .D(n2866), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n656) );
  DFFNSRXLTS \requesterAddressbuffer_reg[5][5]  ( .D(n2865), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n657) );
  DFFNSRXLTS \dataoutbuffer_reg[7][0]  ( .D(n2610), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n798) );
  DFFNSRXLTS \dataoutbuffer_reg[7][1]  ( .D(n2609), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n799) );
  DFFNSRXLTS \dataoutbuffer_reg[7][2]  ( .D(n2608), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n800) );
  DFFNSRXLTS \dataoutbuffer_reg[7][3]  ( .D(n2607), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n801) );
  DFFNSRXLTS \dataoutbuffer_reg[7][4]  ( .D(n2606), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n802) );
  DFFNSRXLTS \dataoutbuffer_reg[7][5]  ( .D(n2605), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n803) );
  DFFNSRXLTS \dataoutbuffer_reg[7][6]  ( .D(n2604), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n804) );
  DFFNSRXLTS \dataoutbuffer_reg[7][7]  ( .D(n2603), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n805) );
  DFFNSRXLTS \dataoutbuffer_reg[7][8]  ( .D(n2602), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n806) );
  DFFNSRXLTS \dataoutbuffer_reg[7][9]  ( .D(n2601), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n807) );
  DFFNSRXLTS \dataoutbuffer_reg[7][10]  ( .D(n2600), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n808) );
  DFFNSRXLTS \dataoutbuffer_reg[7][11]  ( .D(n2599), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n809) );
  DFFNSRXLTS \dataoutbuffer_reg[7][12]  ( .D(n2598), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n810) );
  DFFNSRXLTS \dataoutbuffer_reg[7][13]  ( .D(n2597), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n811) );
  DFFNSRXLTS \dataoutbuffer_reg[7][14]  ( .D(n2596), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n812) );
  DFFNSRXLTS \dataoutbuffer_reg[7][15]  ( .D(n2595), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n813) );
  DFFNSRXLTS \dataoutbuffer_reg[7][16]  ( .D(n2594), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n814) );
  DFFNSRXLTS \dataoutbuffer_reg[7][17]  ( .D(n2593), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n815) );
  DFFNSRXLTS \dataoutbuffer_reg[7][18]  ( .D(n2592), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n816) );
  DFFNSRXLTS \dataoutbuffer_reg[7][19]  ( .D(n2591), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n817) );
  DFFNSRXLTS \dataoutbuffer_reg[7][20]  ( .D(n2590), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n818) );
  DFFNSRXLTS \dataoutbuffer_reg[7][21]  ( .D(n2589), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n819) );
  DFFNSRXLTS \dataoutbuffer_reg[7][22]  ( .D(n2588), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n820) );
  DFFNSRXLTS \dataoutbuffer_reg[7][23]  ( .D(n2587), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n821) );
  DFFNSRXLTS \dataoutbuffer_reg[7][24]  ( .D(n2586), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n822) );
  DFFNSRXLTS \dataoutbuffer_reg[7][25]  ( .D(n2585), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n823) );
  DFFNSRXLTS \dataoutbuffer_reg[7][26]  ( .D(n2584), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n824) );
  DFFNSRXLTS \dataoutbuffer_reg[7][27]  ( .D(n2583), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n825) );
  DFFNSRXLTS \dataoutbuffer_reg[7][28]  ( .D(n2582), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n826) );
  DFFNSRXLTS \dataoutbuffer_reg[7][29]  ( .D(n2581), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n827) );
  DFFNSRXLTS \dataoutbuffer_reg[7][30]  ( .D(n2580), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n828) );
  DFFNSRXLTS \dataoutbuffer_reg[7][31]  ( .D(n2579), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n829) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][1]  ( .D(n2561), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n830) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][2]  ( .D(n2560), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n831) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][3]  ( .D(n2559), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n832) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][5]  ( .D(n2557), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n833) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][0]  ( .D(n2562), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n862) );
  DFFNSRXLTS \requesterAddressbuffer_reg[7][0]  ( .D(n2882), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n880) );
  DFFNSRXLTS \requesterAddressbuffer_reg[7][1]  ( .D(n2881), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n881) );
  DFFNSRXLTS \requesterAddressbuffer_reg[7][3]  ( .D(n2879), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n882) );
  DFFNSRXLTS \requesterAddressbuffer_reg[7][2]  ( .D(n2880), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n883) );
  DFFNSRXLTS \requesterAddressbuffer_reg[7][4]  ( .D(n2878), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n884) );
  DFFNSRXLTS \requesterAddressbuffer_reg[7][5]  ( .D(n2877), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n885) );
  DFFNSRXLTS \dataoutbuffer_reg[5][0]  ( .D(n2674), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n967) );
  DFFNSRXLTS \requesterAddressbuffer_reg[2][2]  ( .D(n2850), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][2] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[2][3]  ( .D(n2849), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][3] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[2][5]  ( .D(n2847), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][5] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[2][0]  ( .D(n2852), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][0] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[2][1]  ( .D(n2851), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][1] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[2][4]  ( .D(n2848), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][4] ) );
  DFFNSRXLTS \dataoutbuffer_reg[1][0]  ( .D(n2802), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3185), .QN(n797) );
  DFFNSRXLTS \dataoutbuffer_reg[1][1]  ( .D(n2801), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3183), .QN(n834) );
  DFFNSRXLTS \dataoutbuffer_reg[1][3]  ( .D(n2799), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3180), .QN(n835) );
  DFFNSRXLTS \dataoutbuffer_reg[1][4]  ( .D(n2798), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3178), .QN(n836) );
  DFFNSRXLTS \dataoutbuffer_reg[1][6]  ( .D(n2796), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3176), .QN(n837) );
  DFFNSRXLTS \dataoutbuffer_reg[1][7]  ( .D(n2795), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3175), .QN(n838) );
  DFFNSRXLTS \dataoutbuffer_reg[1][9]  ( .D(n2793), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3171), .QN(n839) );
  DFFNSRXLTS \dataoutbuffer_reg[1][11]  ( .D(n2791), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3169), .QN(n840) );
  DFFNSRXLTS \dataoutbuffer_reg[1][12]  ( .D(n2790), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3168), .QN(n841) );
  DFFNSRXLTS \dataoutbuffer_reg[1][13]  ( .D(n2789), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3167), .QN(n842) );
  DFFNSRXLTS \dataoutbuffer_reg[1][14]  ( .D(n2788), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3166), .QN(n843) );
  DFFNSRXLTS \dataoutbuffer_reg[1][15]  ( .D(n2787), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3165), .QN(n844) );
  DFFNSRXLTS \dataoutbuffer_reg[1][16]  ( .D(n2786), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3163), .QN(n845) );
  DFFNSRXLTS \dataoutbuffer_reg[1][17]  ( .D(n2785), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3162), .QN(n846) );
  DFFNSRXLTS \dataoutbuffer_reg[1][18]  ( .D(n2784), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3160), .QN(n847) );
  DFFNSRXLTS \dataoutbuffer_reg[1][21]  ( .D(n2781), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3156), .QN(n848) );
  DFFNSRXLTS \dataoutbuffer_reg[1][23]  ( .D(n2779), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3153), .QN(n849) );
  DFFNSRXLTS \dataoutbuffer_reg[1][24]  ( .D(n2778), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3152), .QN(n850) );
  DFFNSRXLTS \dataoutbuffer_reg[1][25]  ( .D(n2777), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3151), .QN(n851) );
  DFFNSRXLTS \dataoutbuffer_reg[1][26]  ( .D(n2776), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3150), .QN(n852) );
  DFFNSRXLTS \dataoutbuffer_reg[1][28]  ( .D(n2774), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3145), .QN(n853) );
  DFFNSRXLTS \dataoutbuffer_reg[1][29]  ( .D(n2773), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3144), .QN(n854) );
  DFFNSRXLTS \dataoutbuffer_reg[1][30]  ( .D(n2772), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3142), .QN(n855) );
  DFFNSRXLTS \dataoutbuffer_reg[1][31]  ( .D(n2771), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3141), .QN(n856) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][0]  ( .D(n2478), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3192), .QN(n857) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][1]  ( .D(n2477), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3190), .QN(n858) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][2]  ( .D(n2476), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3189), .QN(n859) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][3]  ( .D(n2475), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3188), .QN(n860) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][5]  ( .D(n2473), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3186), .QN(n861) );
  DFFNSRXLTS \dataoutbuffer_reg[1][2]  ( .D(n2800), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3181), .QN(n863) );
  DFFNSRXLTS \dataoutbuffer_reg[1][5]  ( .D(n2797), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3177), .QN(n864) );
  DFFNSRXLTS \dataoutbuffer_reg[1][8]  ( .D(n2794), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3174), .QN(n865) );
  DFFNSRXLTS \dataoutbuffer_reg[1][10]  ( .D(n2792), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3170), .QN(n866) );
  DFFNSRXLTS \dataoutbuffer_reg[1][19]  ( .D(n2783), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3159), .QN(n867) );
  DFFNSRXLTS \dataoutbuffer_reg[1][20]  ( .D(n2782), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3158), .QN(n868) );
  DFFNSRXLTS \dataoutbuffer_reg[1][22]  ( .D(n2780), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3154), .QN(n869) );
  DFFNSRXLTS \dataoutbuffer_reg[1][27]  ( .D(n2775), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3149), .QN(n870) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][0]  ( .D(n2846), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3013), .QN(n887) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][1]  ( .D(n2845), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3010), .QN(n888) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][2]  ( .D(n2844), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3009), .QN(n889) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][3]  ( .D(n2843), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3012), .QN(n890) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][4]  ( .D(n2842), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3008), .QN(n891) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][5]  ( .D(n2841), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3007), .QN(n892) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][4]  ( .D(n2474), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3187), .QN(n872) );
  DFFNSRX1TS \dataoutbuffer_reg[0][0]  ( .D(n2834), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n669) );
  DFFNSRX1TS \dataoutbuffer_reg[0][1]  ( .D(n2833), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n670) );
  DFFNSRX1TS \dataoutbuffer_reg[0][2]  ( .D(n2832), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n671) );
  DFFNSRX1TS \dataoutbuffer_reg[0][5]  ( .D(n2829), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n672) );
  DFFNSRX1TS \dataoutbuffer_reg[0][9]  ( .D(n2825), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n673) );
  DFFNSRX1TS \dataoutbuffer_reg[0][20]  ( .D(n2814), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n674) );
  DFFNSRX1TS \dataoutbuffer_reg[0][23]  ( .D(n2811), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n675) );
  DFFNSRX1TS \dataoutbuffer_reg[0][27]  ( .D(n2807), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n676) );
  DFFNSRX1TS \dataoutbuffer_reg[0][28]  ( .D(n2806), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n677) );
  DFFNSRXLTS \readOutbuffer_reg[0]  ( .D(n2563), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n886) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][0]  ( .D(n2548), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3135) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][1]  ( .D(n2547), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3133) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][2]  ( .D(n2546), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3131) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][3]  ( .D(n2545), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3129) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][5]  ( .D(n2543), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3124) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][4]  ( .D(n2544), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3126) );
  DFFNSRXLTS \requesterAddressbuffer_reg[6][1]  ( .D(n2875), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][1] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[6][2]  ( .D(n2874), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][2] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[6][3]  ( .D(n2873), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][3] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[6][4]  ( .D(n2872), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][4] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[6][5]  ( .D(n2871), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][5] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[6][0]  ( .D(n2876), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][0] ) );
  DFFNSRXLTS \dataoutbuffer_reg[6][31]  ( .D(n2611), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3039), .QN(n901) );
  DFFNSRXLTS \dataoutbuffer_reg[6][30]  ( .D(n2612), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3041), .QN(n902) );
  DFFNSRXLTS \dataoutbuffer_reg[6][29]  ( .D(n2613), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3043), .QN(n903) );
  DFFNSRXLTS \dataoutbuffer_reg[6][28]  ( .D(n2614), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3046), .QN(n904) );
  DFFNSRXLTS \dataoutbuffer_reg[6][27]  ( .D(n2615), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3050), .QN(n905) );
  DFFNSRXLTS \dataoutbuffer_reg[6][26]  ( .D(n2616), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3052), .QN(n906) );
  DFFNSRXLTS \dataoutbuffer_reg[6][25]  ( .D(n2617), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3054), .QN(n907) );
  DFFNSRXLTS \dataoutbuffer_reg[6][24]  ( .D(n2618), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3057), .QN(n908) );
  DFFNSRXLTS \dataoutbuffer_reg[6][23]  ( .D(n2619), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3059), .QN(n909) );
  DFFNSRXLTS \dataoutbuffer_reg[6][22]  ( .D(n2620), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3062), .QN(n910) );
  DFFNSRXLTS \dataoutbuffer_reg[6][21]  ( .D(n2621), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3064), .QN(n911) );
  DFFNSRXLTS \dataoutbuffer_reg[6][20]  ( .D(n2622), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3067), .QN(n912) );
  DFFNSRXLTS \dataoutbuffer_reg[6][19]  ( .D(n2623), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3070), .QN(n913) );
  DFFNSRXLTS \dataoutbuffer_reg[6][18]  ( .D(n2624), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3072), .QN(n914) );
  DFFNSRXLTS \dataoutbuffer_reg[6][17]  ( .D(n2625), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3075), .QN(n915) );
  DFFNSRXLTS \dataoutbuffer_reg[6][16]  ( .D(n2626), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3077), .QN(n916) );
  DFFNSRXLTS \dataoutbuffer_reg[6][15]  ( .D(n2627), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3079), .QN(n917) );
  DFFNSRXLTS \dataoutbuffer_reg[6][14]  ( .D(n2628), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3081), .QN(n918) );
  DFFNSRXLTS \dataoutbuffer_reg[6][13]  ( .D(n2629), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3086), .QN(n919) );
  DFFNSRXLTS \dataoutbuffer_reg[6][12]  ( .D(n2630), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3089), .QN(n920) );
  DFFNSRXLTS \dataoutbuffer_reg[6][11]  ( .D(n2631), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3091), .QN(n921) );
  DFFNSRXLTS \dataoutbuffer_reg[6][10]  ( .D(n2632), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3094), .QN(n922) );
  DFFNSRXLTS \dataoutbuffer_reg[6][9]  ( .D(n2633), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3096), .QN(n923) );
  DFFNSRXLTS \dataoutbuffer_reg[6][8]  ( .D(n2634), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3098), .QN(n924) );
  DFFNSRXLTS \dataoutbuffer_reg[6][7]  ( .D(n2635), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3102), .QN(n925) );
  DFFNSRXLTS \dataoutbuffer_reg[6][6]  ( .D(n2636), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3105), .QN(n926) );
  DFFNSRXLTS \dataoutbuffer_reg[6][5]  ( .D(n2637), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3107), .QN(n927) );
  DFFNSRXLTS \dataoutbuffer_reg[6][4]  ( .D(n2638), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3109), .QN(n928) );
  DFFNSRXLTS \dataoutbuffer_reg[6][3]  ( .D(n2639), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3113), .QN(n929) );
  DFFNSRXLTS \dataoutbuffer_reg[6][2]  ( .D(n2640), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3116), .QN(n930) );
  DFFNSRXLTS \dataoutbuffer_reg[6][1]  ( .D(n2641), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3118), .QN(n931) );
  DFFNSRXLTS \dataoutbuffer_reg[6][0]  ( .D(n2642), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3122), .QN(n932) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][13]  ( .D(n2507), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3280), .QN(n600) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][13]  ( .D(n2549), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3289), .QN(n788) );
  DFFNSRXLTS \writeOutbuffer_reg[4]  ( .D(n2575), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n750) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][9]  ( .D(n2511), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3284), .QN(n599) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][6]  ( .D(n2514), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3287), .QN(n605) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][7]  ( .D(n2513), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3286), .QN(n606) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][8]  ( .D(n2512), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3285), .QN(n607) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][10]  ( .D(n2510), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3283), .QN(n608) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][11]  ( .D(n2509), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3282), .QN(n609) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][12]  ( .D(n2508), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3281), .QN(n610) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][10]  ( .D(n2552), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n593), .QN(n871) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][6]  ( .D(n2556), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3302), .QN(n893) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][7]  ( .D(n2555), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3300), .QN(n894) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][8]  ( .D(n2554), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3298), .QN(n895) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][11]  ( .D(n2551), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3293), .QN(n896) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][9]  ( .D(n2553), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3296), .QN(n897) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][12]  ( .D(n2550), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3291), .QN(n933) );
  DFFNSRXLTS \writeOutbuffer_reg[7]  ( .D(n2578), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3270), .QN(n879) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][1]  ( .D(n2491), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n692) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][0]  ( .D(n2492), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n691) );
  DFFNSRXLTS \dataoutbuffer_reg[2][31]  ( .D(n2739), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n668) );
  DFFNSRXLTS \dataoutbuffer_reg[2][30]  ( .D(n2740), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n745) );
  DFFNSRXLTS \dataoutbuffer_reg[2][29]  ( .D(n2741), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n744) );
  DFFNSRXLTS \dataoutbuffer_reg[2][28]  ( .D(n2742), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n743) );
  DFFNSRXLTS \dataoutbuffer_reg[2][27]  ( .D(n2743), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n690) );
  DFFNSRXLTS \dataoutbuffer_reg[2][26]  ( .D(n2744), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n742) );
  DFFNSRXLTS \dataoutbuffer_reg[2][25]  ( .D(n2745), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n741) );
  DFFNSRXLTS \dataoutbuffer_reg[2][24]  ( .D(n2746), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n667) );
  DFFNSRXLTS \dataoutbuffer_reg[2][23]  ( .D(n2747), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n740) );
  DFFNSRXLTS \dataoutbuffer_reg[2][22]  ( .D(n2748), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n666) );
  DFFNSRXLTS \dataoutbuffer_reg[2][21]  ( .D(n2749), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n739) );
  DFFNSRXLTS \dataoutbuffer_reg[2][20]  ( .D(n2750), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n738) );
  DFFNSRXLTS \dataoutbuffer_reg[2][19]  ( .D(n2751), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n737) );
  DFFNSRXLTS \dataoutbuffer_reg[2][18]  ( .D(n2752), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n736) );
  DFFNSRXLTS \dataoutbuffer_reg[2][17]  ( .D(n2753), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n735) );
  DFFNSRXLTS \dataoutbuffer_reg[2][16]  ( .D(n2754), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n665) );
  DFFNSRXLTS \dataoutbuffer_reg[2][15]  ( .D(n2755), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n734) );
  DFFNSRXLTS \dataoutbuffer_reg[2][14]  ( .D(n2756), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n733) );
  DFFNSRXLTS \dataoutbuffer_reg[2][13]  ( .D(n2757), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n732) );
  DFFNSRXLTS \dataoutbuffer_reg[2][12]  ( .D(n2758), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n731) );
  DFFNSRXLTS \dataoutbuffer_reg[2][11]  ( .D(n2759), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n730) );
  DFFNSRXLTS \dataoutbuffer_reg[2][10]  ( .D(n2760), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n689) );
  DFFNSRXLTS \dataoutbuffer_reg[2][9]  ( .D(n2761), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n729) );
  DFFNSRXLTS \dataoutbuffer_reg[2][8]  ( .D(n2762), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n728) );
  DFFNSRXLTS \dataoutbuffer_reg[2][7]  ( .D(n2763), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n727) );
  DFFNSRXLTS \dataoutbuffer_reg[2][6]  ( .D(n2764), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n664) );
  DFFNSRXLTS \dataoutbuffer_reg[2][5]  ( .D(n2765), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n726) );
  DFFNSRXLTS \dataoutbuffer_reg[2][4]  ( .D(n2766), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n725) );
  DFFNSRXLTS \dataoutbuffer_reg[2][3]  ( .D(n2767), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n724) );
  DFFNSRXLTS \dataoutbuffer_reg[2][2]  ( .D(n2768), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n663) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][5]  ( .D(n2487), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n695) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][4]  ( .D(n2488), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n694) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][3]  ( .D(n2489), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n693) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][2]  ( .D(n2490), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n746) );
  DFFNSRXLTS \dataoutbuffer_reg[2][1]  ( .D(n2769), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n688) );
  DFFNSRXLTS \dataoutbuffer_reg[2][0]  ( .D(n2770), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n662) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][13]  ( .D(n2479), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3334), .QN(n575) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][12]  ( .D(n2480), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3333), .QN(n566) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][11]  ( .D(n2481), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3332), .QN(n572) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][10]  ( .D(n2482), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3331), .QN(n565) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][9]  ( .D(n2483), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3330), .QN(n571) );
  DFFNSRXLTS \writeOutbuffer_reg[2]  ( .D(n2573), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n660) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][8]  ( .D(n2484), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3329), .QN(n564) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][7]  ( .D(n2485), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3328), .QN(n570) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][6]  ( .D(n2486), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3327), .QN(n563) );
  DFFNSRXLTS \requesterAddressbuffer_reg[0][3]  ( .D(n2837), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][3] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[0][2]  ( .D(n2838), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][2] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[0][0]  ( .D(n2840), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][0] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[0][1]  ( .D(n2839), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][1] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[0][5]  ( .D(n2835), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][5] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[0][4]  ( .D(n2836), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][4] ) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][1]  ( .D(n2463), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n39) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][0]  ( .D(n2464), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n91) );
  DFFNSRXLTS \dataoutbuffer_reg[0][31]  ( .D(n2803), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n40) );
  DFFNSRXLTS \dataoutbuffer_reg[0][30]  ( .D(n2804), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n41) );
  DFFNSRXLTS \dataoutbuffer_reg[0][29]  ( .D(n2805), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n42) );
  DFFNSRXLTS \dataoutbuffer_reg[0][26]  ( .D(n2808), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n43) );
  DFFNSRXLTS \dataoutbuffer_reg[0][25]  ( .D(n2809), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n44) );
  DFFNSRXLTS \dataoutbuffer_reg[0][24]  ( .D(n2810), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n45) );
  DFFNSRXLTS \dataoutbuffer_reg[0][22]  ( .D(n2812), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n46) );
  DFFNSRXLTS \dataoutbuffer_reg[0][21]  ( .D(n2813), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n47) );
  DFFNSRXLTS \dataoutbuffer_reg[0][19]  ( .D(n2815), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n48) );
  DFFNSRXLTS \dataoutbuffer_reg[0][18]  ( .D(n2816), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n49) );
  DFFNSRXLTS \dataoutbuffer_reg[0][17]  ( .D(n2817), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n50) );
  DFFNSRXLTS \dataoutbuffer_reg[0][16]  ( .D(n2818), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n51) );
  DFFNSRXLTS \dataoutbuffer_reg[0][15]  ( .D(n2819), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n52) );
  DFFNSRXLTS \dataoutbuffer_reg[0][14]  ( .D(n2820), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n53) );
  DFFNSRXLTS \dataoutbuffer_reg[0][13]  ( .D(n2821), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n54) );
  DFFNSRXLTS \dataoutbuffer_reg[0][12]  ( .D(n2822), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n55) );
  DFFNSRXLTS \dataoutbuffer_reg[0][11]  ( .D(n2823), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n56) );
  DFFNSRXLTS \dataoutbuffer_reg[0][10]  ( .D(n2824), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n57) );
  DFFNSRXLTS \dataoutbuffer_reg[0][8]  ( .D(n2826), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n58) );
  DFFNSRXLTS \dataoutbuffer_reg[0][7]  ( .D(n2827), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n59) );
  DFFNSRXLTS \dataoutbuffer_reg[0][6]  ( .D(n2828), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n60) );
  DFFNSRXLTS \dataoutbuffer_reg[0][4]  ( .D(n2830), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n61) );
  DFFNSRXLTS \dataoutbuffer_reg[0][3]  ( .D(n2831), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n62) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][4]  ( .D(n2460), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n90) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][3]  ( .D(n2461), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n37) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][2]  ( .D(n2462), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n38) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][5]  ( .D(n2459), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n36) );
  DFFNSRXLTS \destinationAddressOut_reg[7]  ( .D(n2447), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[7]) );
  DFFNSRXLTS \destinationAddressOut_reg[6]  ( .D(n2448), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[6]) );
  DFFNSRXLTS \destinationAddressOut_reg[9]  ( .D(n2445), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[9]) );
  DFFNSRXLTS \destinationAddressOut_reg[8]  ( .D(n2446), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[8]) );
  DFFNSRXLTS \destinationAddressOut_reg[13]  ( .D(n2441), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[13]) );
  DFFNSRXLTS \destinationAddressOut_reg[12]  ( .D(n2442), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[12]) );
  DFFNSRXLTS \destinationAddressOut_reg[11]  ( .D(n2443), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[11]) );
  DFFNSRXLTS \destinationAddressOut_reg[10]  ( .D(n2444), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[10]) );
  DFFNSRXLTS \write_reg_reg[1]  ( .D(n2887), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n6), .QN(n9) );
  DFFNSRXLTS \readOutbuffer_reg[1]  ( .D(n2564), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n651) );
  DFFNSRXLTS \readOutbuffer_reg[5]  ( .D(n2568), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n650) );
  DFFNSRXLTS \readOutbuffer_reg[6]  ( .D(n2569), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n649) );
  DFFNSRXLTS \readOutbuffer_reg[7]  ( .D(n2570), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer_7) );
  DFFNSRXLTS full_reg_reg ( .D(N4718), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        n2285), .QN(n764) );
  DFFNSRXLTS \readOutbuffer_reg[4]  ( .D(n2567), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n752) );
  DFFNSRXLTS \readOutbuffer_reg[3]  ( .D(n2566), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n648) );
  DFFNSRXLTS \readOutbuffer_reg[2]  ( .D(n2565), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\readOutbuffer[2] ), .QN(n751) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][8]  ( .D(n2456), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3321), .QN(n576) );
  DFFNSRXLTS \writeOutbuffer_reg[0]  ( .D(n2571), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n747) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][7]  ( .D(n2457), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3320), .QN(n567) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][6]  ( .D(n2458), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3319), .QN(n573) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][9]  ( .D(n2455), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3322), .QN(n568) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][12]  ( .D(n2452), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3325), .QN(n577) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][11]  ( .D(n2453), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3324), .QN(n569) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][10]  ( .D(n2454), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3323), .QN(n574) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][13]  ( .D(n2451), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3326), .QN(n966) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][11]  ( .D(n2537), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3308), .QN(n597) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][9]  ( .D(n2539), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3312), .QN(n602) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][7]  ( .D(n2541), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3316), .QN(n595) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][6]  ( .D(n2542), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3318), .QN(n601) );
  DFFNSRXLTS \writeOutbuffer_reg[6]  ( .D(n2577), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n749) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][12]  ( .D(n2536), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3306), .QN(n604) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][10]  ( .D(n2538), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3310), .QN(n603) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][8]  ( .D(n2540), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3314), .QN(n596) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][13]  ( .D(n2535), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3304), .QN(n598) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][13]  ( .D(n2521), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3288), .QN(n588) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][12]  ( .D(n2522), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3290), .QN(n587) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][11]  ( .D(n2523), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3292), .QN(n586) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][10]  ( .D(n2524), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3294), .QN(n585) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][9]  ( .D(n2525), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3295), .QN(n584) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][5]  ( .D(n2853), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][5] ), .QN(n877) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][4]  ( .D(n2854), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][4] ), .QN(n878) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][3]  ( .D(n2855), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][3] ), .QN(n876) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][2]  ( .D(n2856), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][2] ), .QN(n875) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][1]  ( .D(n2857), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][1] ), .QN(n874) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][0]  ( .D(n2858), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][0] ), .QN(n873) );
  DFFNSRXLTS \writeOutbuffer_reg[5]  ( .D(n2576), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3271), .QN(n658) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][8]  ( .D(n2526), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3297), .QN(n583) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][7]  ( .D(n2527), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3299), .QN(n582) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][6]  ( .D(n2528), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3301), .QN(n581) );
  DFFNSRXLTS \dataoutbuffer_reg[3][1]  ( .D(n2737), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n88), .QN(n697) );
  DFFNSRXLTS \dataoutbuffer_reg[3][0]  ( .D(n2738), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n89), .QN(n696) );
  DFFNSRXLTS \requesterAddressbuffer_reg[4][2]  ( .D(n2862), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3032) );
  DFFNSRXLTS \requesterAddressbuffer_reg[4][1]  ( .D(n2863), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3033) );
  DFFNSRXLTS \requesterAddressbuffer_reg[4][3]  ( .D(n2861), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3034) );
  DFFNSRXLTS \requesterAddressbuffer_reg[4][0]  ( .D(n2864), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3035) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][5]  ( .D(n2501), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n63), .QN(n723) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][4]  ( .D(n2502), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n64), .QN(n722) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][3]  ( .D(n2503), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n65), .QN(n721) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][2]  ( .D(n2504), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n92), .QN(n687) );
  DFFNSRXLTS \requesterAddressbuffer_reg[4][5]  ( .D(n2859), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3030) );
  DFFNSRXLTS \requesterAddressbuffer_reg[4][4]  ( .D(n2860), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3031) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][1]  ( .D(n2505), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n66), .QN(n720) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][0]  ( .D(n2506), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n67), .QN(n719) );
  DFFNSRXLTS \dataoutbuffer_reg[3][31]  ( .D(n2707), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n68), .QN(n718) );
  DFFNSRXLTS \dataoutbuffer_reg[3][30]  ( .D(n2708), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n69), .QN(n717) );
  DFFNSRXLTS \dataoutbuffer_reg[3][29]  ( .D(n2709), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n70), .QN(n716) );
  DFFNSRXLTS \dataoutbuffer_reg[3][28]  ( .D(n2710), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n71), .QN(n715) );
  DFFNSRXLTS \dataoutbuffer_reg[3][27]  ( .D(n2711), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n72), .QN(n714) );
  DFFNSRXLTS \dataoutbuffer_reg[3][26]  ( .D(n2712), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n73), .QN(n713) );
  DFFNSRXLTS \dataoutbuffer_reg[3][25]  ( .D(n2713), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n93), .QN(n686) );
  DFFNSRXLTS \dataoutbuffer_reg[3][24]  ( .D(n2714), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n74), .QN(n712) );
  DFFNSRXLTS \dataoutbuffer_reg[3][23]  ( .D(n2715), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n94), .QN(n685) );
  DFFNSRXLTS \dataoutbuffer_reg[3][22]  ( .D(n2716), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n75), .QN(n711) );
  DFFNSRXLTS \dataoutbuffer_reg[3][21]  ( .D(n2717), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n76), .QN(n709) );
  DFFNSRXLTS \dataoutbuffer_reg[3][20]  ( .D(n2718), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n95), .QN(n684) );
  DFFNSRXLTS \dataoutbuffer_reg[3][19]  ( .D(n2719), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n77), .QN(n708) );
  DFFNSRXLTS \dataoutbuffer_reg[3][18]  ( .D(n2720), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n96), .QN(n683) );
  DFFNSRXLTS \dataoutbuffer_reg[3][17]  ( .D(n2721), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n78), .QN(n707) );
  DFFNSRXLTS \dataoutbuffer_reg[3][16]  ( .D(n2722), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n79), .QN(n706) );
  DFFNSRXLTS \dataoutbuffer_reg[3][15]  ( .D(n2723), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n97), .QN(n682) );
  DFFNSRXLTS \dataoutbuffer_reg[3][14]  ( .D(n2724), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n80), .QN(n705) );
  DFFNSRXLTS \dataoutbuffer_reg[3][13]  ( .D(n2725), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n98), .QN(n681) );
  DFFNSRXLTS \dataoutbuffer_reg[3][12]  ( .D(n2726), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n81), .QN(n704) );
  DFFNSRXLTS \dataoutbuffer_reg[3][11]  ( .D(n2727), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n82), .QN(n703) );
  DFFNSRXLTS \dataoutbuffer_reg[3][10]  ( .D(n2728), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n83), .QN(n702) );
  DFFNSRXLTS \dataoutbuffer_reg[3][9]  ( .D(n2729), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n84), .QN(n701) );
  DFFNSRXLTS \dataoutbuffer_reg[3][8]  ( .D(n2730), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n85), .QN(n700) );
  DFFNSRXLTS \dataoutbuffer_reg[3][6]  ( .D(n2732), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n86), .QN(n699) );
  DFFNSRXLTS \dataoutbuffer_reg[3][5]  ( .D(n2733), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n99), .QN(n680) );
  DFFNSRXLTS \dataoutbuffer_reg[3][3]  ( .D(n2735), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n87), .QN(n698) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][10]  ( .D(n2496), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3309), .QN(n579) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][9]  ( .D(n2497), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3311), .QN(n590) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][12]  ( .D(n2494), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3305), .QN(n591) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][11]  ( .D(n2495), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3307), .QN(n594) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][13]  ( .D(n2493), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3303), .QN(n580) );
  NAND2XLTS U2 ( .A(n1820), .B(n1816), .Y(n1790) );
  BUFX3TS U3 ( .A(n3746), .Y(n3745) );
  OAI22X2TS U4 ( .A0(n1833), .A1(n233), .B0(n1917), .B1(n143), .Y(n1795) );
  AOI2BB1X2TS U5 ( .A0N(n139), .A1N(n1961), .B0(n1837), .Y(n1833) );
  XOR2X2TS U6 ( .A(n972), .B(selectBit_EAST), .Y(n3006) );
  INVX1TS U7 ( .A(n421), .Y(n1) );
  CLKINVX2TS U8 ( .A(n1), .Y(n2) );
  BUFX4TS U9 ( .A(n3474), .Y(n3463) );
  BUFX4TS U10 ( .A(n3803), .Y(n3800) );
  AOI21X1TS U11 ( .A0(n446), .A1(n952), .B0(n941), .Y(n1858) );
  INVX1TS U12 ( .A(n1857), .Y(n941) );
  BUFX2TS U13 ( .A(n1247), .Y(n3228) );
  BUFX4TS U14 ( .A(n1247), .Y(n3229) );
  BUFX4TS U15 ( .A(n3087), .Y(n3085) );
  XNOR2X1TS U16 ( .A(n2058), .B(n2059), .Y(n2008) );
  OR2X2TS U17 ( .A(selectBit_NORTH), .B(selectBit_SOUTH), .Y(n2963) );
  AOI21X1TS U18 ( .A0(n958), .A1(n960), .B0(n1798), .Y(n1838) );
  XOR2X1TS U19 ( .A(n2055), .B(n123), .Y(n1940) );
  NOR2X1TS U20 ( .A(n2008), .B(n1084), .Y(n1894) );
  INVX2TS U21 ( .A(n1940), .Y(n947) );
  NOR2BX1TS U22 ( .AN(n2008), .B(n1084), .Y(n1939) );
  CLKBUFX2TS U23 ( .A(n1939), .Y(n28) );
  AOI21X1TS U24 ( .A0(n141), .A1(n142), .B0(n3793), .Y(n1830) );
  AOI21X1TS U25 ( .A0(n958), .A1(n163), .B0(n531), .Y(n1854) );
  NOR3BX1TS U26 ( .AN(n162), .B(n1865), .C(n950), .Y(n524) );
  AOI21X1TS U27 ( .A0(n1841), .A1(n952), .B0(n944), .Y(n1843) );
  NAND2X1TS U28 ( .A(n1833), .B(n1830), .Y(n1794) );
  OAI21X1TS U29 ( .A0(n1836), .A1(n2007), .B0(n2054), .Y(n1865) );
  AOI2BB1X1TS U30 ( .A0N(n955), .A1N(n1961), .B0(n1865), .Y(n1863) );
  INVX2TS U31 ( .A(writeIn_WEST), .Y(n3) );
  INVX2TS U32 ( .A(n1798), .Y(n516) );
  CLKBUFX2TS U33 ( .A(n3389), .Y(n3388) );
  OA22X2TS U34 ( .A0(n523), .A1(n428), .B0(n434), .B1(n450), .Y(n19) );
  INVX2TS U35 ( .A(n19), .Y(n127) );
  INVX2TS U36 ( .A(n1800), .Y(n224) );
  CLKBUFX2TS U37 ( .A(n1265), .Y(n2389) );
  CLKBUFX2TS U38 ( .A(n1265), .Y(n2380) );
  INVX1TS U39 ( .A(n1801), .Y(n206) );
  OA22X1TS U40 ( .A0(n1858), .A1(n16), .B0(n1889), .B1(n164), .Y(n531) );
  OA22X1TS U41 ( .A0(n1863), .A1(n232), .B0(n1917), .B1(n2024), .Y(n4) );
  OA21XLTS U42 ( .A0(n1984), .A1(n232), .B0(n1975), .Y(n1798) );
  NOR3BXLTS U43 ( .AN(n1830), .B(n1837), .C(n156), .Y(n1200) );
  NAND3XLTS U44 ( .A(n1894), .B(n445), .C(n1940), .Y(n1842) );
  AOI32X1TS U45 ( .A0(n450), .A1(n428), .A2(n423), .B0(n3006), .B1(n429), .Y(
        n3005) );
  NAND2XLTS U46 ( .A(n1863), .B(n1860), .Y(n1805) );
  NOR3BX1TS U47 ( .AN(n1860), .B(n161), .C(n940), .Y(n1265) );
  AOI21X1TS U48 ( .A0(n523), .A1(n438), .B0(n146), .Y(n2062) );
  INVX1TS U49 ( .A(n18), .Y(n146) );
  NAND3XLTS U50 ( .A(n957), .B(n1939), .C(n1940), .Y(n2054) );
  NAND3XLTS U51 ( .A(n957), .B(n1894), .C(n1940), .Y(n1852) );
  CLKBUFX2TS U52 ( .A(n2380), .Y(n2033) );
  CLKINVX2TS U53 ( .A(n516), .Y(n773) );
  INVX2TS U54 ( .A(n519), .Y(n784) );
  CLKBUFX2TS U55 ( .A(n218), .Y(n3765) );
  OAI21X1TS U56 ( .A0(n946), .A1(n949), .B0(n145), .Y(n1890) );
  CLKBUFX2TS U57 ( .A(n1186), .Y(n3510) );
  NAND2X1TS U58 ( .A(n1814), .B(n2060), .Y(n1962) );
  CLKBUFX2TS U59 ( .A(n1217), .Y(n3395) );
  CLKBUFX2TS U60 ( .A(n1200), .Y(n3477) );
  CLKBUFX2TS U61 ( .A(n1200), .Y(n3476) );
  INVX2TS U62 ( .A(n445), .Y(n957) );
  AO21X1TS U63 ( .A0(n958), .A1(n142), .B0(n530), .Y(n5) );
  NOR2X1TS U64 ( .A(n1962), .B(n450), .Y(n1892) );
  INVX2TS U65 ( .A(n947), .Y(n433) );
  CLKBUFX2TS U66 ( .A(n3822), .Y(n3821) );
  CLKBUFX2TS U67 ( .A(n1149), .Y(n3707) );
  CLKBUFX2TS U68 ( .A(n3593), .Y(n3590) );
  CLKBUFX2TS U69 ( .A(n3559), .Y(n3552) );
  OA22X1TS U70 ( .A0(n1828), .A1(n233), .B0(n1889), .B1(n1930), .Y(n530) );
  INVX2TS U71 ( .A(selectBit_EAST), .Y(n450) );
  CLKBUFX2TS U72 ( .A(n3229), .Y(n3223) );
  CLKBUFX2TS U73 ( .A(n3793), .Y(n3792) );
  CLKBUFX2TS U74 ( .A(n3475), .Y(n3469) );
  CLKBUFX2TS U75 ( .A(n3502), .Y(n3501) );
  CLKBUFX2TS U76 ( .A(n3558), .Y(n3551) );
  INVX2TS U77 ( .A(n1838), .Y(n24) );
  AO21X1TS U78 ( .A0(n1892), .A1(n948), .B0(n1835), .Y(n1837) );
  NOR3BX1TS U79 ( .AN(n1939), .B(n444), .C(n433), .Y(n1835) );
  NOR3X1TS U80 ( .A(n1819), .B(n1822), .C(n1821), .Y(n1820) );
  CLKINVX2TS U81 ( .A(n15), .Y(n215) );
  CLKBUFX2TS U82 ( .A(n3406), .Y(n3405) );
  AOI222XLTS U83 ( .A0(n3994), .A1(n2985), .B0(n3951), .B1(n2380), .C0(n4174), 
        .C1(n442), .Y(n2046) );
  AOI222XLTS U84 ( .A0(n3997), .A1(n2985), .B0(n3954), .B1(n2380), .C0(n4177), 
        .C1(n442), .Y(n2047) );
  AOI222XLTS U85 ( .A0(n4139), .A1(n2986), .B0(n4144), .B1(n1265), .C0(n4153), 
        .C1(n1808), .Y(n1807) );
  AOI222XLTS U86 ( .A0(n4000), .A1(n2985), .B0(n3957), .B1(n2033), .C0(n4180), 
        .C1(n1808), .Y(n2048) );
  AOI222XLTS U87 ( .A0(n4484), .A1(n3697), .B0(n33), .B1(n3683), .C0(n4122), 
        .C1(n3667), .Y(n1148) );
  AOI222XLTS U88 ( .A0(n4482), .A1(n3704), .B0(n458), .B1(n3678), .C0(n4386), 
        .C1(n3669), .Y(n1788) );
  AOI222XLTS U89 ( .A0(n4479), .A1(n3705), .B0(n461), .B1(n3678), .C0(n4383), 
        .C1(n3669), .Y(n1786) );
  AOI222XLTS U90 ( .A0(n4476), .A1(n3703), .B0(n463), .B1(n3679), .C0(n4380), 
        .C1(n3669), .Y(n1784) );
  AOI222XLTS U91 ( .A0(n4473), .A1(n3704), .B0(n465), .B1(n3679), .C0(n4377), 
        .C1(n3669), .Y(n1782) );
  AOI222XLTS U92 ( .A0(n4470), .A1(n3705), .B0(n467), .B1(n3679), .C0(n4374), 
        .C1(n3668), .Y(n1780) );
  AOI222XLTS U93 ( .A0(n4467), .A1(n3702), .B0(n469), .B1(n3679), .C0(n4371), 
        .C1(n3668), .Y(n1778) );
  AOI222XLTS U94 ( .A0(n4464), .A1(n3702), .B0(n471), .B1(n3680), .C0(n4368), 
        .C1(n3668), .Y(n1776) );
  AOI222XLTS U95 ( .A0(n4461), .A1(n1149), .B0(n473), .B1(n3680), .C0(n4365), 
        .C1(n3668), .Y(n1774) );
  AOI222XLTS U96 ( .A0(n4458), .A1(n3702), .B0(n475), .B1(n3680), .C0(n4362), 
        .C1(n3676), .Y(n1772) );
  AOI222XLTS U97 ( .A0(n4455), .A1(n3707), .B0(n477), .B1(n3680), .C0(n4359), 
        .C1(n3672), .Y(n1770) );
  AOI222XLTS U98 ( .A0(n4452), .A1(n3697), .B0(n479), .B1(n3681), .C0(n4356), 
        .C1(n3673), .Y(n1768) );
  AOI222XLTS U99 ( .A0(n4449), .A1(n3697), .B0(n481), .B1(n3681), .C0(n4353), 
        .C1(n3673), .Y(n1766) );
  AOI222XLTS U100 ( .A0(n4446), .A1(n3697), .B0(n483), .B1(n3681), .C0(n4350), 
        .C1(n3671), .Y(n1764) );
  AOI222XLTS U101 ( .A0(n4443), .A1(n3696), .B0(n485), .B1(n3681), .C0(n4347), 
        .C1(n3670), .Y(n1762) );
  AOI222XLTS U102 ( .A0(n4440), .A1(n3696), .B0(n487), .B1(n3685), .C0(n4344), 
        .C1(n3670), .Y(n1760) );
  AOI222XLTS U103 ( .A0(n4437), .A1(n3696), .B0(n489), .B1(n3688), .C0(n4341), 
        .C1(n3672), .Y(n1758) );
  AOI222XLTS U104 ( .A0(n4434), .A1(n3696), .B0(n491), .B1(n3689), .C0(n4338), 
        .C1(n3667), .Y(n1756) );
  AOI222XLTS U105 ( .A0(n4431), .A1(n3695), .B0(n493), .B1(n3683), .C0(n4335), 
        .C1(n3667), .Y(n1754) );
  AOI222XLTS U106 ( .A0(n4428), .A1(n3695), .B0(n495), .B1(n3685), .C0(n4332), 
        .C1(n3667), .Y(n1752) );
  AOI222XLTS U107 ( .A0(n4425), .A1(n3695), .B0(n497), .B1(n3685), .C0(n4329), 
        .C1(n3666), .Y(n1750) );
  AOI222XLTS U108 ( .A0(n4422), .A1(n3695), .B0(n499), .B1(n3687), .C0(n4326), 
        .C1(n3666), .Y(n1748) );
  AOI222XLTS U109 ( .A0(n4419), .A1(n3694), .B0(n501), .B1(n3690), .C0(n4323), 
        .C1(n3666), .Y(n1746) );
  AOI222XLTS U110 ( .A0(n4416), .A1(n3694), .B0(n503), .B1(n3684), .C0(n4320), 
        .C1(n3666), .Y(n1744) );
  AOI222XLTS U111 ( .A0(n4413), .A1(n3694), .B0(n505), .B1(n3684), .C0(n4317), 
        .C1(n3665), .Y(n1742) );
  AOI222XLTS U112 ( .A0(n4410), .A1(n3694), .B0(n452), .B1(n3686), .C0(n4314), 
        .C1(n3665), .Y(n1740) );
  AOI222XLTS U113 ( .A0(n4407), .A1(n3693), .B0(n507), .B1(n3686), .C0(n4311), 
        .C1(n3665), .Y(n1738) );
  AOI222XLTS U114 ( .A0(n4404), .A1(n3693), .B0(n509), .B1(n3684), .C0(n4308), 
        .C1(n3665), .Y(n1736) );
  AOI222XLTS U115 ( .A0(n4401), .A1(n3693), .B0(n454), .B1(n3684), .C0(n4305), 
        .C1(n3664), .Y(n1734) );
  AOI222XLTS U116 ( .A0(n4398), .A1(n3693), .B0(n511), .B1(n3687), .C0(n4302), 
        .C1(n3664), .Y(n1732) );
  AOI222XLTS U117 ( .A0(n4395), .A1(n3692), .B0(n456), .B1(n3685), .C0(n4299), 
        .C1(n3664), .Y(n1730) );
  AOI222XLTS U118 ( .A0(n4392), .A1(n3692), .B0(n515), .B1(n3682), .C0(n4296), 
        .C1(n3664), .Y(n1728) );
  AOI222XLTS U119 ( .A0(n4389), .A1(n3692), .B0(n513), .B1(n3682), .C0(n4293), 
        .C1(n3663), .Y(n1726) );
  XOR2X1TS U120 ( .A(n127), .B(n199), .Y(n2058) );
  INVX2TS U121 ( .A(n4), .Y(n128) );
  CLKBUFX2TS U122 ( .A(n784), .Y(n3751) );
  OAI22X1TS U123 ( .A0(n942), .A1(n232), .B0(n1917), .B1(n1985), .Y(n1801) );
  AND2X2TS U124 ( .A(n145), .B(n4502), .Y(n7) );
  CLKINVX2TS U125 ( .A(n224), .Y(n225) );
  CLKINVX2TS U126 ( .A(selectBit_SOUTH), .Y(n428) );
  AND3X2TS U127 ( .A(n1854), .B(n1859), .C(n1858), .Y(n14) );
  AND2X2TS U128 ( .A(n1838), .B(n955), .Y(n15) );
  OR2X2TS U129 ( .A(n2064), .B(n2285), .Y(n16) );
  INVX2TS U130 ( .A(n1893), .Y(n445) );
  CLKAND2X2TS U131 ( .A(n2063), .B(n164), .Y(n17) );
  OR2X2TS U132 ( .A(n972), .B(n438), .Y(n18) );
  AND2X2TS U133 ( .A(n6), .B(n26), .Y(n20) );
  INVX2TS U134 ( .A(n218), .Y(n219) );
  INVX1TS U135 ( .A(n1794), .Y(n229) );
  CLKINVX2TS U136 ( .A(n229), .Y(n230) );
  NOR2X1TS U137 ( .A(n126), .B(n4504), .Y(n1131) );
  OR2X2TS U138 ( .A(n1130), .B(n534), .Y(n21) );
  AND2X2TS U139 ( .A(n13), .B(n4502), .Y(n22) );
  INVX2TS U140 ( .A(selectBit_EAST), .Y(n1029) );
  INVX2TS U141 ( .A(n24), .Y(n25) );
  NOR2X1TS U142 ( .A(n956), .B(n1986), .Y(n1841) );
  CLKBUFX2TS U143 ( .A(n1846), .Y(n23) );
  AOI21X1TS U144 ( .A0(n141), .A1(n960), .B0(n3809), .Y(n1846) );
  INVX1TS U145 ( .A(n2061), .Y(n26) );
  NAND2X1TS U146 ( .A(n2062), .B(n429), .Y(n2061) );
  INVXLTS U147 ( .A(n951), .Y(n27) );
  NAND2X1TS U148 ( .A(n954), .B(n173), .Y(n1859) );
  INVXLTS U149 ( .A(readRequesterAddress[0]), .Y(n29) );
  INVXLTS U150 ( .A(n29), .Y(n30) );
  INVXLTS U151 ( .A(n29), .Y(n31) );
  INVXLTS U152 ( .A(n29), .Y(n32) );
  INVXLTS U153 ( .A(n29), .Y(n33) );
  INVXLTS U154 ( .A(readRequesterAddress[1]), .Y(n34) );
  INVXLTS U155 ( .A(n34), .Y(n35) );
  INVXLTS U156 ( .A(n34), .Y(n100) );
  INVXLTS U157 ( .A(n34), .Y(n101) );
  INVXLTS U158 ( .A(n34), .Y(n102) );
  INVXLTS U159 ( .A(readRequesterAddress[2]), .Y(n103) );
  INVXLTS U160 ( .A(n103), .Y(n104) );
  INVXLTS U161 ( .A(n103), .Y(n105) );
  INVXLTS U162 ( .A(n103), .Y(n106) );
  INVXLTS U163 ( .A(n103), .Y(n107) );
  INVXLTS U164 ( .A(readRequesterAddress[3]), .Y(n108) );
  INVXLTS U165 ( .A(n108), .Y(n109) );
  INVXLTS U166 ( .A(n108), .Y(n110) );
  INVXLTS U167 ( .A(n108), .Y(n111) );
  INVXLTS U168 ( .A(n108), .Y(n112) );
  INVXLTS U169 ( .A(readRequesterAddress[4]), .Y(n113) );
  INVXLTS U170 ( .A(n113), .Y(n114) );
  INVXLTS U171 ( .A(n113), .Y(n115) );
  INVXLTS U172 ( .A(n113), .Y(n116) );
  INVXLTS U173 ( .A(n113), .Y(n117) );
  INVXLTS U174 ( .A(readRequesterAddress[5]), .Y(n118) );
  INVXLTS U175 ( .A(n118), .Y(n119) );
  INVXLTS U176 ( .A(n118), .Y(n120) );
  INVXLTS U177 ( .A(n118), .Y(n121) );
  INVXLTS U178 ( .A(n118), .Y(n122) );
  INVXLTS U179 ( .A(n441), .Y(n123) );
  INVXLTS U180 ( .A(n123), .Y(n124) );
  INVXLTS U181 ( .A(n12), .Y(n125) );
  INVXLTS U182 ( .A(n443), .Y(n126) );
  INVX2TS U183 ( .A(n1795), .Y(n780) );
  NOR3BX1TS U184 ( .AN(n28), .B(n444), .C(n433), .Y(n129) );
  CLKBUFX2TS U185 ( .A(n1816), .Y(n130) );
  AOI21X1TS U186 ( .A0(n169), .A1(n140), .B0(n1128), .Y(n1816) );
  INVXLTS U187 ( .A(n5), .Y(n131) );
  INVXLTS U188 ( .A(n5), .Y(n132) );
  INVXLTS U189 ( .A(n1815), .Y(n133) );
  INVXLTS U190 ( .A(n133), .Y(n134) );
  OAI21X1TS U191 ( .A0(n1888), .A1(n170), .B0(n1146), .Y(n1815) );
  CLKINVX2TS U192 ( .A(n1854), .Y(n135) );
  INVX2TS U193 ( .A(n135), .Y(n136) );
  CLKBUFX2TS U194 ( .A(n1830), .Y(n137) );
  INVXLTS U195 ( .A(n17), .Y(n138) );
  INVX1TS U196 ( .A(n17), .Y(n139) );
  INVXLTS U197 ( .A(n21), .Y(n140) );
  INVXLTS U198 ( .A(n21), .Y(n141) );
  INVXLTS U199 ( .A(n1930), .Y(n142) );
  INVXLTS U200 ( .A(n142), .Y(n143) );
  INVXLTS U201 ( .A(n16), .Y(n144) );
  INVX1TS U202 ( .A(n16), .Y(n145) );
  INVX1TS U203 ( .A(n18), .Y(n147) );
  INVXLTS U204 ( .A(n7), .Y(n148) );
  INVXLTS U205 ( .A(n3897), .Y(n149) );
  INVXLTS U206 ( .A(n3787), .Y(n150) );
  INVXLTS U207 ( .A(n3787), .Y(n151) );
  INVXLTS U208 ( .A(n240), .Y(n152) );
  INVXLTS U209 ( .A(n152), .Y(n153) );
  INVXLTS U210 ( .A(n152), .Y(n154) );
  INVXLTS U211 ( .A(n950), .Y(n155) );
  INVXLTS U212 ( .A(n155), .Y(n156) );
  INVXLTS U213 ( .A(n2999), .Y(n157) );
  OAI22X1TS U214 ( .A0(n970), .A1(n2997), .B0(n2998), .B1(n2999), .Y(n2982) );
  INVXLTS U215 ( .A(n981), .Y(n158) );
  INVXLTS U216 ( .A(n158), .Y(n159) );
  INVXLTS U217 ( .A(n11), .Y(n160) );
  INVXLTS U218 ( .A(n948), .Y(n161) );
  CLKBUFX2TS U219 ( .A(n1860), .Y(n162) );
  AOI21X1TS U220 ( .A0(n140), .A1(n163), .B0(n4), .Y(n1860) );
  INVXLTS U221 ( .A(n2024), .Y(n163) );
  INVXLTS U222 ( .A(n163), .Y(n164) );
  INVXLTS U223 ( .A(n459), .Y(n165) );
  INVXLTS U224 ( .A(n160), .Y(n166) );
  INVXLTS U225 ( .A(n440), .Y(n167) );
  INVXLTS U226 ( .A(n167), .Y(n168) );
  INVXLTS U227 ( .A(n1879), .Y(n169) );
  INVXLTS U228 ( .A(n169), .Y(n170) );
  INVXLTS U229 ( .A(n22), .Y(n171) );
  INVXLTS U230 ( .A(n22), .Y(n172) );
  INVXLTS U231 ( .A(n533), .Y(n173) );
  INVXLTS U232 ( .A(n754), .Y(n174) );
  INVXLTS U233 ( .A(n174), .Y(n175) );
  INVXLTS U234 ( .A(n174), .Y(n176) );
  INVXLTS U235 ( .A(n760), .Y(n177) );
  INVXLTS U236 ( .A(n177), .Y(n178) );
  INVXLTS U237 ( .A(n177), .Y(n179) );
  INVXLTS U238 ( .A(n979), .Y(n180) );
  INVXLTS U239 ( .A(n180), .Y(n181) );
  INVXLTS U240 ( .A(n180), .Y(n182) );
  INVXLTS U241 ( .A(n980), .Y(n183) );
  INVXLTS U242 ( .A(n183), .Y(n184) );
  INVXLTS U243 ( .A(n183), .Y(n185) );
  INVXLTS U244 ( .A(destinationAddressIn_NORTH[13]), .Y(n186) );
  INVXLTS U245 ( .A(destinationAddressIn_NORTH[13]), .Y(n187) );
  INVXLTS U246 ( .A(destinationAddressIn_NORTH[11]), .Y(n188) );
  INVXLTS U247 ( .A(destinationAddressIn_NORTH[11]), .Y(n189) );
  INVXLTS U248 ( .A(destinationAddressIn_NORTH[9]), .Y(n190) );
  INVXLTS U249 ( .A(destinationAddressIn_NORTH[9]), .Y(n191) );
  INVXLTS U250 ( .A(destinationAddressIn_NORTH[12]), .Y(n192) );
  INVXLTS U251 ( .A(destinationAddressIn_NORTH[12]), .Y(n193) );
  INVXLTS U252 ( .A(destinationAddressIn_NORTH[10]), .Y(n194) );
  INVXLTS U253 ( .A(destinationAddressIn_NORTH[10]), .Y(n195) );
  INVXLTS U254 ( .A(destinationAddressIn_NORTH[8]), .Y(n196) );
  INVXLTS U255 ( .A(destinationAddressIn_NORTH[8]), .Y(n197) );
  INVXLTS U256 ( .A(n533), .Y(n198) );
  INVXLTS U257 ( .A(n198), .Y(n199) );
  INVXLTS U258 ( .A(n762), .Y(n200) );
  INVXLTS U259 ( .A(n200), .Y(n201) );
  INVXLTS U260 ( .A(n200), .Y(n202) );
  INVXLTS U261 ( .A(writeIn_NORTH), .Y(n203) );
  INVXLTS U262 ( .A(writeIn_NORTH), .Y(n204) );
  INVXLTS U263 ( .A(n3897), .Y(n205) );
  INVXLTS U264 ( .A(n206), .Y(n207) );
  INVXLTS U265 ( .A(n206), .Y(n208) );
  INVXLTS U266 ( .A(n1792), .Y(n209) );
  INVXLTS U267 ( .A(n209), .Y(n210) );
  INVXLTS U268 ( .A(n209), .Y(n211) );
  INVXLTS U269 ( .A(n14), .Y(n212) );
  INVXLTS U270 ( .A(n14), .Y(n213) );
  INVXLTS U271 ( .A(n14), .Y(n214) );
  INVXLTS U272 ( .A(n15), .Y(n216) );
  INVXLTS U273 ( .A(n15), .Y(n217) );
  INVXLTS U274 ( .A(n1790), .Y(n218) );
  INVXLTS U275 ( .A(n218), .Y(n220) );
  INVXLTS U276 ( .A(n2096), .Y(n221) );
  INVXLTS U277 ( .A(n221), .Y(n222) );
  INVXLTS U278 ( .A(n221), .Y(n223) );
  INVXLTS U279 ( .A(n224), .Y(n226) );
  INVXLTS U280 ( .A(n3930), .Y(n227) );
  INVXLTS U281 ( .A(n3930), .Y(n228) );
  INVXLTS U282 ( .A(n229), .Y(n231) );
  INVX2TS U283 ( .A(n144), .Y(n232) );
  CLKINVX1TS U284 ( .A(n145), .Y(n233) );
  INVXLTS U285 ( .A(n2079), .Y(n234) );
  INVXLTS U286 ( .A(n2079), .Y(n235) );
  INVXLTS U287 ( .A(n2084), .Y(n236) );
  INVXLTS U288 ( .A(n236), .Y(n237) );
  INVXLTS U289 ( .A(n236), .Y(n238) );
  INVXLTS U290 ( .A(n1131), .Y(n239) );
  INVXLTS U291 ( .A(n239), .Y(n240) );
  INVXLTS U292 ( .A(n239), .Y(n241) );
  INVXLTS U293 ( .A(n239), .Y(n242) );
  INVX2TS U472 ( .A(n138), .Y(n955) );
  INVXLTS U473 ( .A(selectBit_EAST), .Y(n421) );
  INVX2TS U474 ( .A(n2), .Y(n422) );
  NAND2X1TS U475 ( .A(n422), .B(n1962), .Y(n2007) );
  OAI2BB1X2TS U476 ( .A0N(n434), .A1N(n422), .B0(n3005), .Y(n2999) );
  INVX1TS U477 ( .A(n523), .Y(n423) );
  CLKINVX2TS U478 ( .A(selectBit_NORTH), .Y(n523) );
  INVX2TS U479 ( .A(selectBit_NORTH), .Y(n972) );
  INVX2TS U480 ( .A(n1084), .Y(n425) );
  INVXLTS U481 ( .A(n429), .Y(n426) );
  OAI31XLTS U482 ( .A0(n954), .A1(n147), .A2(n958), .B0(n145), .Y(n1889) );
  INVX2TS U483 ( .A(n1130), .Y(n427) );
  INVX1TS U484 ( .A(n428), .Y(n429) );
  INVX2TS U485 ( .A(readIn_SOUTH), .Y(n431) );
  CLKBUFX2TS U486 ( .A(n2962), .Y(n432) );
  OAI21XLTS U487 ( .A0(n2962), .A1(n970), .B0(n3000), .Y(n3003) );
  CLKINVX2TS U488 ( .A(n2963), .Y(n434) );
  INVXLTS U489 ( .A(n2963), .Y(n435) );
  OAI221XLTS U490 ( .A0(n124), .A1(n1853), .B0(n1850), .B1(n2007), .C0(n1852), 
        .Y(n1851) );
  CLKBUFX2TS U491 ( .A(n2082), .Y(n761) );
  INVX2TS U492 ( .A(n761), .Y(n436) );
  INVX2TS U493 ( .A(n761), .Y(n437) );
  INVX2TS U494 ( .A(n5327), .Y(n534) );
  INVX2TS U495 ( .A(n534), .Y(n438) );
  INVX2TS U496 ( .A(n534), .Y(n439) );
  NOR2X1TS U497 ( .A(n157), .B(n438), .Y(n2059) );
  OAI32X1TS U498 ( .A0(n2056), .A1(n438), .A2(n970), .B0(n19), .B1(n9), .Y(
        n2055) );
  INVXLTS U499 ( .A(n767), .Y(n442) );
  INVXLTS U500 ( .A(n524), .Y(n767) );
  XOR2X1TS U501 ( .A(n424), .B(n970), .Y(n1893) );
  CLKINVX1TS U502 ( .A(n1893), .Y(n444) );
  OR2XLTS U503 ( .A(n2011), .B(n1986), .Y(n1826) );
  INVX2TS U504 ( .A(n1826), .Y(n446) );
  INVX2TS U505 ( .A(n1826), .Y(n447) );
  AOI21X1TS U506 ( .A0(n1892), .A1(n446), .B0(n945), .Y(n1828) );
  CLKBUFX2TS U507 ( .A(n2081), .Y(n759) );
  INVX2TS U508 ( .A(n759), .Y(n448) );
  INVX2TS U509 ( .A(n759), .Y(n449) );
  CLKBUFX2TS U510 ( .A(cacheDataOut[7]), .Y(n451) );
  CLKBUFX2TS U511 ( .A(cacheDataOut[7]), .Y(n452) );
  CLKBUFX2TS U512 ( .A(cacheDataOut[4]), .Y(n453) );
  CLKBUFX2TS U513 ( .A(cacheDataOut[4]), .Y(n454) );
  CLKBUFX2TS U514 ( .A(cacheDataOut[2]), .Y(n455) );
  CLKBUFX2TS U515 ( .A(cacheDataOut[2]), .Y(n456) );
  CLKBUFX2TS U516 ( .A(cacheDataOut[31]), .Y(n457) );
  CLKBUFX2TS U517 ( .A(cacheDataOut[31]), .Y(n458) );
  CLKBUFX2TS U518 ( .A(cacheDataOut[30]), .Y(n460) );
  CLKBUFX2TS U519 ( .A(cacheDataOut[30]), .Y(n461) );
  CLKBUFX2TS U520 ( .A(cacheDataOut[29]), .Y(n462) );
  CLKBUFX2TS U521 ( .A(cacheDataOut[29]), .Y(n463) );
  CLKBUFX2TS U522 ( .A(cacheDataOut[28]), .Y(n464) );
  CLKBUFX2TS U523 ( .A(cacheDataOut[28]), .Y(n465) );
  CLKBUFX2TS U524 ( .A(cacheDataOut[27]), .Y(n466) );
  CLKBUFX2TS U525 ( .A(cacheDataOut[27]), .Y(n467) );
  CLKBUFX2TS U526 ( .A(cacheDataOut[26]), .Y(n468) );
  CLKBUFX2TS U527 ( .A(cacheDataOut[26]), .Y(n469) );
  CLKBUFX2TS U528 ( .A(cacheDataOut[25]), .Y(n470) );
  CLKBUFX2TS U529 ( .A(cacheDataOut[25]), .Y(n471) );
  CLKBUFX2TS U530 ( .A(cacheDataOut[24]), .Y(n472) );
  CLKBUFX2TS U531 ( .A(cacheDataOut[24]), .Y(n473) );
  CLKBUFX2TS U532 ( .A(cacheDataOut[23]), .Y(n474) );
  CLKBUFX2TS U533 ( .A(cacheDataOut[23]), .Y(n475) );
  CLKBUFX2TS U534 ( .A(cacheDataOut[22]), .Y(n476) );
  CLKBUFX2TS U535 ( .A(cacheDataOut[22]), .Y(n477) );
  CLKBUFX2TS U536 ( .A(cacheDataOut[21]), .Y(n478) );
  CLKBUFX2TS U537 ( .A(cacheDataOut[21]), .Y(n479) );
  CLKBUFX2TS U538 ( .A(cacheDataOut[20]), .Y(n480) );
  CLKBUFX2TS U539 ( .A(cacheDataOut[20]), .Y(n481) );
  CLKBUFX2TS U540 ( .A(cacheDataOut[19]), .Y(n482) );
  CLKBUFX2TS U541 ( .A(cacheDataOut[19]), .Y(n483) );
  CLKBUFX2TS U542 ( .A(cacheDataOut[18]), .Y(n484) );
  CLKBUFX2TS U543 ( .A(cacheDataOut[18]), .Y(n485) );
  CLKBUFX2TS U544 ( .A(cacheDataOut[17]), .Y(n486) );
  CLKBUFX2TS U545 ( .A(cacheDataOut[17]), .Y(n487) );
  CLKBUFX2TS U546 ( .A(cacheDataOut[16]), .Y(n488) );
  CLKBUFX2TS U547 ( .A(cacheDataOut[16]), .Y(n489) );
  CLKBUFX2TS U548 ( .A(cacheDataOut[15]), .Y(n490) );
  CLKBUFX2TS U549 ( .A(cacheDataOut[15]), .Y(n491) );
  CLKBUFX2TS U550 ( .A(cacheDataOut[14]), .Y(n492) );
  CLKBUFX2TS U551 ( .A(cacheDataOut[14]), .Y(n493) );
  CLKBUFX2TS U552 ( .A(cacheDataOut[13]), .Y(n494) );
  CLKBUFX2TS U553 ( .A(cacheDataOut[13]), .Y(n495) );
  CLKBUFX2TS U554 ( .A(cacheDataOut[12]), .Y(n496) );
  CLKBUFX2TS U555 ( .A(cacheDataOut[12]), .Y(n497) );
  CLKBUFX2TS U556 ( .A(cacheDataOut[11]), .Y(n498) );
  CLKBUFX2TS U557 ( .A(cacheDataOut[11]), .Y(n499) );
  CLKBUFX2TS U558 ( .A(cacheDataOut[10]), .Y(n500) );
  CLKBUFX2TS U559 ( .A(cacheDataOut[10]), .Y(n501) );
  CLKBUFX2TS U560 ( .A(cacheDataOut[9]), .Y(n502) );
  CLKBUFX2TS U561 ( .A(cacheDataOut[9]), .Y(n503) );
  CLKBUFX2TS U562 ( .A(cacheDataOut[8]), .Y(n504) );
  CLKBUFX2TS U563 ( .A(cacheDataOut[8]), .Y(n505) );
  CLKBUFX2TS U564 ( .A(cacheDataOut[6]), .Y(n506) );
  CLKBUFX2TS U565 ( .A(cacheDataOut[6]), .Y(n507) );
  CLKBUFX2TS U566 ( .A(cacheDataOut[5]), .Y(n508) );
  CLKBUFX2TS U567 ( .A(cacheDataOut[5]), .Y(n509) );
  CLKBUFX2TS U568 ( .A(cacheDataOut[3]), .Y(n510) );
  CLKBUFX2TS U569 ( .A(cacheDataOut[3]), .Y(n511) );
  CLKBUFX2TS U570 ( .A(cacheDataOut[0]), .Y(n512) );
  CLKBUFX2TS U571 ( .A(cacheDataOut[0]), .Y(n513) );
  CLKBUFX2TS U572 ( .A(cacheDataOut[1]), .Y(n514) );
  CLKBUFX2TS U573 ( .A(cacheDataOut[1]), .Y(n515) );
  INVXLTS U574 ( .A(n1798), .Y(n517) );
  INVXLTS U575 ( .A(n1798), .Y(n518) );
  OA21XLTS U576 ( .A0(n1985), .A1(n1962), .B0(n1843), .Y(n1984) );
  AND2XLTS U577 ( .A(n1819), .B(n1816), .Y(n1164) );
  CLKINVX2TS U578 ( .A(n1164), .Y(n519) );
  INVXLTS U579 ( .A(n1164), .Y(n520) );
  INVXLTS U580 ( .A(n1164), .Y(n521) );
  INVXLTS U581 ( .A(n1164), .Y(n522) );
  INVX1TS U582 ( .A(n3426), .Y(n3421) );
  INVX1TS U583 ( .A(n3424), .Y(n3423) );
  INVXLTS U584 ( .A(n3425), .Y(n3422) );
  CLKINVX2TS U585 ( .A(n3640), .Y(n3627) );
  CLKINVX2TS U586 ( .A(n3640), .Y(n3628) );
  CLKINVX2TS U587 ( .A(n3640), .Y(n3629) );
  CLKINVX2TS U588 ( .A(n3641), .Y(n3630) );
  CLKINVX2TS U589 ( .A(n3641), .Y(n3631) );
  CLKINVX2TS U590 ( .A(n3641), .Y(n3632) );
  CLKINVX2TS U591 ( .A(n3641), .Y(n3633) );
  CLKINVX2TS U592 ( .A(n3642), .Y(n3626) );
  NAND2X1TS U593 ( .A(n20), .B(n955), .Y(n1814) );
  NAND3XLTS U594 ( .A(n131), .B(n1859), .C(n1828), .Y(n1792) );
  NAND2XLTS U595 ( .A(n16), .B(n4502), .Y(n1134) );
  NAND2XLTS U596 ( .A(selectBit_WEST), .B(readReady), .Y(n3000) );
  INVX2TS U597 ( .A(n3492), .Y(n3478) );
  NOR2BX1TS U598 ( .AN(n1892), .B(n1850), .Y(n1819) );
  INVXLTS U599 ( .A(n1836), .Y(n948) );
  OAI22XLTS U600 ( .A0(n139), .A1(n981), .B0(n955), .B1(n996), .Y(n1844) );
  CLKINVX2TS U601 ( .A(n2061), .Y(n954) );
  OAI211XLTS U602 ( .A0(n3487), .A1(n4201), .B0(n1534), .C0(n1535), .Y(n2705)
         );
  OAI211XLTS U603 ( .A0(n3487), .A1(n4198), .B0(n1532), .C0(n1533), .Y(n2706)
         );
  OAI211XLTS U604 ( .A0(n3478), .A1(n3992), .B0(n1951), .C0(n1952), .Y(n2515)
         );
  OAI211XLTS U605 ( .A0(n3478), .A1(n3989), .B0(n1949), .C0(n1950), .Y(n2516)
         );
  OAI211XLTS U606 ( .A0(n3478), .A1(n3986), .B0(n1947), .C0(n1948), .Y(n2517)
         );
  OAI211XLTS U607 ( .A0(n3486), .A1(n4207), .B0(n1538), .C0(n1539), .Y(n2703)
         );
  AOI222XLTS U608 ( .A0(n3972), .A1(n3121), .B0(n4014), .B1(n3138), .C0(
        destinationAddressIn_SOUTH[13]), .C1(n3225), .Y(n2032) );
  NOR2XLTS U609 ( .A(n1853), .B(n10), .Y(n1822) );
  CLKBUFX2TS U610 ( .A(n6), .Y(n533) );
  INVXLTS U611 ( .A(n1814), .Y(n953) );
  NOR2XLTS U612 ( .A(n1814), .B(n1815), .Y(n1149) );
  INVXLTS U613 ( .A(n3491), .Y(n3486) );
  INVXLTS U614 ( .A(n3374), .Y(n3369) );
  INVXLTS U615 ( .A(n3490), .Y(n3487) );
  INVXLTS U616 ( .A(n3373), .Y(n3370) );
  INVXLTS U617 ( .A(n3489), .Y(n3488) );
  INVXLTS U618 ( .A(n3372), .Y(n3371) );
  INVX1TS U619 ( .A(n1805), .Y(n766) );
  INVX1TS U620 ( .A(n225), .Y(n775) );
  CLKBUFX2TS U621 ( .A(n3577), .Y(n3574) );
  CLKBUFX2TS U622 ( .A(n3577), .Y(n3575) );
  NOR2BXLTS U623 ( .AN(n1854), .B(n27), .Y(n1247) );
  NOR2BXLTS U624 ( .AN(n131), .B(n27), .Y(n1183) );
  CLKBUFX2TS U625 ( .A(n3247), .Y(n3244) );
  CLKBUFX2TS U626 ( .A(n3247), .Y(n3245) );
  AND2XLTS U627 ( .A(n944), .B(n25), .Y(n526) );
  INVXLTS U628 ( .A(n1859), .Y(n951) );
  CLKBUFX2TS U629 ( .A(n1116), .Y(n1111) );
  CLKBUFX2TS U630 ( .A(n1116), .Y(n1112) );
  NOR3BX1TS U631 ( .AN(n162), .B(n1865), .C(n156), .Y(n1808) );
  NAND3XLTS U632 ( .A(n947), .B(n444), .C(n1939), .Y(n1827) );
  NAND3XLTS U633 ( .A(n947), .B(n445), .C(n1894), .Y(n1812) );
  NAND2XLTS U634 ( .A(n1841), .B(n1892), .Y(n1811) );
  NOR2BXLTS U635 ( .AN(n1846), .B(n1852), .Y(n1233) );
  NOR2BXLTS U636 ( .AN(n1860), .B(n2054), .Y(n1263) );
  NOR2XLTS U637 ( .A(n1812), .B(n1815), .Y(n1152) );
  NOR2XLTS U638 ( .A(n1811), .B(n1815), .Y(n1151) );
  NOR3BX1TS U639 ( .AN(n1830), .B(n161), .C(n129), .Y(n1202) );
  NAND2XLTS U640 ( .A(n956), .B(n2010), .Y(n1961) );
  NOR2BXLTS U641 ( .AN(n1854), .B(n1857), .Y(n1249) );
  OR4XLTS U642 ( .A(n134), .B(n949), .C(n946), .D(n953), .Y(n527) );
  CLKINVX2TS U643 ( .A(n1851), .Y(n942) );
  AND3XLTS U644 ( .A(n447), .B(n1857), .C(n136), .Y(n1250) );
  AND3XLTS U645 ( .A(n1841), .B(n1842), .C(n1838), .Y(n1216) );
  CLKINVX2TS U646 ( .A(n1801), .Y(n777) );
  AND2XLTS U647 ( .A(n129), .B(n137), .Y(n528) );
  INVX1TS U648 ( .A(n1228), .Y(n3378) );
  NAND3BXLTS U649 ( .AN(n1850), .B(n23), .C(n1852), .Y(n1228) );
  NAND3XLTS U650 ( .A(n28), .B(n444), .C(n433), .Y(n1857) );
  NAND2XLTS U651 ( .A(n4141), .B(n945), .Y(n1824) );
  NAND2XLTS U652 ( .A(n4142), .B(n944), .Y(n1839) );
  NOR2X1TS U653 ( .A(n426), .B(n2062), .Y(n2010) );
  AOI21XLTS U654 ( .A0(n426), .A1(n2062), .B0(n2010), .Y(n1986) );
  AOI32XLTS U655 ( .A0(n136), .A1(n1855), .A2(n1856), .B0(n3246), .B1(n651), 
        .Y(n2564) );
  NAND2XLTS U656 ( .A(n4141), .B(n941), .Y(n1855) );
  AOI32XLTS U657 ( .A0(n447), .A1(n1857), .A2(n4147), .B0(n1858), .B1(n1829), 
        .Y(n1856) );
  XOR2XLTS U658 ( .A(n147), .B(n199), .Y(n2011) );
  AND2XLTS U659 ( .A(n1822), .B(n1816), .Y(n1167) );
  OAI2BB1X1TS U660 ( .A0N(n2995), .A1N(n525), .B0(n2987), .Y(n2972) );
  OA22X1TS U661 ( .A0(n1140), .A1(n2989), .B0(n2988), .B1(n2971), .Y(n525) );
  OAI32XLTS U662 ( .A0(n4149), .A1(n943), .A2(n1850), .B0(n1851), .B1(n159), 
        .Y(n1849) );
  OAI22XLTS U663 ( .A0(n951), .A1(n159), .B0(n27), .B1(n996), .Y(n1829) );
  AOI22XLTS U664 ( .A0(n1814), .A1(n159), .B0(n953), .B1(n996), .Y(n1813) );
  NAND2X1TS U665 ( .A(n199), .B(n124), .Y(n1879) );
  NAND2X1TS U666 ( .A(n173), .B(n441), .Y(n1930) );
  XOR2X1TS U667 ( .A(n3001), .B(n758), .Y(n1140) );
  NAND3X1TS U668 ( .A(n168), .B(n430), .C(n165), .Y(n2097) );
  OAI211XLTS U669 ( .A0(n4501), .A1(n3912), .B0(n1274), .C0(n1275), .Y(n2835)
         );
  OAI211XLTS U670 ( .A0(n4498), .A1(n3912), .B0(n1272), .C0(n1273), .Y(n2836)
         );
  OAI211XLTS U671 ( .A0(n3478), .A1(n3983), .B0(n1945), .C0(n1946), .Y(n2518)
         );
  OAI211XLTS U672 ( .A0(n3479), .A1(n3980), .B0(n1943), .C0(n1944), .Y(n2519)
         );
  OAI211XLTS U673 ( .A0(n3479), .A1(n3977), .B0(n1941), .C0(n1942), .Y(n2520)
         );
  OAI211XLTS U674 ( .A0(n3479), .A1(n4288), .B0(n1592), .C0(n1593), .Y(n2676)
         );
  OAI211XLTS U675 ( .A0(n3480), .A1(n4282), .B0(n1588), .C0(n1589), .Y(n2678)
         );
  OAI211XLTS U676 ( .A0(n3480), .A1(n4279), .B0(n1586), .C0(n1587), .Y(n2679)
         );
  OAI211XLTS U677 ( .A0(n3480), .A1(n4276), .B0(n1584), .C0(n1585), .Y(n2680)
         );
  OAI211XLTS U678 ( .A0(n3481), .A1(n4273), .B0(n1582), .C0(n1583), .Y(n2681)
         );
  OAI211XLTS U679 ( .A0(n3481), .A1(n4270), .B0(n1580), .C0(n1581), .Y(n2682)
         );
  OAI211XLTS U680 ( .A0(n3481), .A1(n4267), .B0(n1578), .C0(n1579), .Y(n2683)
         );
  OAI211XLTS U681 ( .A0(n3482), .A1(n4252), .B0(n1568), .C0(n1569), .Y(n2688)
         );
  OAI211XLTS U682 ( .A0(n3484), .A1(n4237), .B0(n1558), .C0(n1559), .Y(n2693)
         );
  OAI211XLTS U683 ( .A0(n3485), .A1(n4225), .B0(n1550), .C0(n1551), .Y(n2697)
         );
  OAI211XLTS U684 ( .A0(n3485), .A1(n4219), .B0(n1546), .C0(n1547), .Y(n2699)
         );
  OAI211XLTS U685 ( .A0(n3486), .A1(n4213), .B0(n1542), .C0(n1543), .Y(n2701)
         );
  OAI211XLTS U686 ( .A0(n3486), .A1(n4210), .B0(n1540), .C0(n1541), .Y(n2702)
         );
  OAI211XLTS U687 ( .A0(n3486), .A1(n4204), .B0(n1536), .C0(n1537), .Y(n2704)
         );
  OAI211XLTS U688 ( .A0(n3479), .A1(n4291), .B0(n1594), .C0(n1595), .Y(n2675)
         );
  OAI211XLTS U689 ( .A0(n3480), .A1(n4285), .B0(n1590), .C0(n1591), .Y(n2677)
         );
  OAI211XLTS U690 ( .A0(n3481), .A1(n4264), .B0(n1576), .C0(n1577), .Y(n2684)
         );
  OAI211XLTS U691 ( .A0(n3482), .A1(n4261), .B0(n1574), .C0(n1575), .Y(n2685)
         );
  OAI211XLTS U692 ( .A0(n3482), .A1(n4258), .B0(n1572), .C0(n1573), .Y(n2686)
         );
  OAI211XLTS U693 ( .A0(n3482), .A1(n4255), .B0(n1570), .C0(n1571), .Y(n2687)
         );
  OAI211XLTS U694 ( .A0(n3483), .A1(n4246), .B0(n1564), .C0(n1565), .Y(n2690)
         );
  OAI211XLTS U695 ( .A0(n3484), .A1(n4234), .B0(n1556), .C0(n1557), .Y(n2694)
         );
  OAI211XLTS U696 ( .A0(n3484), .A1(n4231), .B0(n1554), .C0(n1555), .Y(n2695)
         );
  OAI211XLTS U697 ( .A0(n3484), .A1(n4228), .B0(n1552), .C0(n1553), .Y(n2696)
         );
  OAI211XLTS U698 ( .A0(n3485), .A1(n4222), .B0(n1548), .C0(n1549), .Y(n2698)
         );
  OAI211XLTS U699 ( .A0(n3485), .A1(n4216), .B0(n1544), .C0(n1545), .Y(n2700)
         );
  OAI211XLTS U700 ( .A0(n3483), .A1(n4249), .B0(n1566), .C0(n1567), .Y(n2689)
         );
  OAI211XLTS U701 ( .A0(n3483), .A1(n4243), .B0(n1562), .C0(n1563), .Y(n2691)
         );
  OAI211XLTS U702 ( .A0(n3483), .A1(n4240), .B0(n1560), .C0(n1561), .Y(n2692)
         );
  OAI211XLTS U703 ( .A0(n4032), .A1(n3487), .B0(n1211), .C0(n1212), .Y(n2859)
         );
  OAI211XLTS U704 ( .A0(n4029), .A1(n3487), .B0(n1209), .C0(n1210), .Y(n2860)
         );
  OAI211XLTS U705 ( .A0(n4026), .A1(n3488), .B0(n1207), .C0(n1208), .Y(n2861)
         );
  OAI211XLTS U706 ( .A0(n4023), .A1(n3488), .B0(n1205), .C0(n1206), .Y(n2862)
         );
  OAI211XLTS U707 ( .A0(n4020), .A1(n3488), .B0(n1203), .C0(n1204), .Y(n2863)
         );
  OAI211XLTS U708 ( .A0(n4017), .A1(n3488), .B0(n1198), .C0(n1199), .Y(n2864)
         );
  OAI211XLTS U709 ( .A0(n3912), .A1(n4393), .B0(n1278), .C0(n1279), .Y(n2833)
         );
  OAI211XLTS U710 ( .A0(n3912), .A1(n4390), .B0(n1276), .C0(n1277), .Y(n2834)
         );
  OAI211XLTS U711 ( .A0(n3917), .A1(n4171), .B0(n2044), .C0(n2045), .Y(n2459)
         );
  OAI211XLTS U712 ( .A0(n3915), .A1(n4165), .B0(n2040), .C0(n2041), .Y(n2461)
         );
  OAI211XLTS U713 ( .A0(n3917), .A1(n4162), .B0(n2038), .C0(n2039), .Y(n2462)
         );
  OAI211XLTS U714 ( .A0(n3905), .A1(n4159), .B0(n2036), .C0(n2037), .Y(n2463)
         );
  OAI211XLTS U715 ( .A0(n3905), .A1(n4483), .B0(n1338), .C0(n1339), .Y(n2803)
         );
  OAI211XLTS U716 ( .A0(n3905), .A1(n4480), .B0(n1336), .C0(n1337), .Y(n2804)
         );
  OAI211XLTS U717 ( .A0(n3906), .A1(n4477), .B0(n1334), .C0(n1335), .Y(n2805)
         );
  OAI211XLTS U718 ( .A0(n3906), .A1(n4468), .B0(n1328), .C0(n1329), .Y(n2808)
         );
  OAI211XLTS U719 ( .A0(n3907), .A1(n4465), .B0(n1326), .C0(n1327), .Y(n2809)
         );
  OAI211XLTS U720 ( .A0(n3907), .A1(n4462), .B0(n1324), .C0(n1325), .Y(n2810)
         );
  OAI211XLTS U721 ( .A0(n3907), .A1(n4456), .B0(n1320), .C0(n1321), .Y(n2812)
         );
  OAI211XLTS U722 ( .A0(n3914), .A1(n4453), .B0(n1318), .C0(n1319), .Y(n2813)
         );
  OAI211XLTS U723 ( .A0(n3915), .A1(n4447), .B0(n1314), .C0(n1315), .Y(n2815)
         );
  OAI211XLTS U724 ( .A0(n3914), .A1(n4444), .B0(n1312), .C0(n1313), .Y(n2816)
         );
  OAI211XLTS U725 ( .A0(n3908), .A1(n4441), .B0(n1310), .C0(n1311), .Y(n2817)
         );
  OAI211XLTS U726 ( .A0(n3908), .A1(n4438), .B0(n1308), .C0(n1309), .Y(n2818)
         );
  OAI211XLTS U727 ( .A0(n3908), .A1(n4435), .B0(n1306), .C0(n1307), .Y(n2819)
         );
  OAI211XLTS U728 ( .A0(n3908), .A1(n4432), .B0(n1304), .C0(n1305), .Y(n2820)
         );
  OAI211XLTS U729 ( .A0(n3909), .A1(n4429), .B0(n1302), .C0(n1303), .Y(n2821)
         );
  OAI211XLTS U730 ( .A0(n3909), .A1(n4426), .B0(n1300), .C0(n1301), .Y(n2822)
         );
  OAI211XLTS U731 ( .A0(n3909), .A1(n4423), .B0(n1298), .C0(n1299), .Y(n2823)
         );
  OAI211XLTS U732 ( .A0(n3909), .A1(n4420), .B0(n1296), .C0(n1297), .Y(n2824)
         );
  OAI211XLTS U733 ( .A0(n3910), .A1(n4414), .B0(n1292), .C0(n1293), .Y(n2826)
         );
  OAI211XLTS U734 ( .A0(n3910), .A1(n4411), .B0(n1290), .C0(n1291), .Y(n2827)
         );
  OAI211XLTS U735 ( .A0(n3910), .A1(n4408), .B0(n1288), .C0(n1289), .Y(n2828)
         );
  OAI211XLTS U736 ( .A0(n3911), .A1(n4402), .B0(n1284), .C0(n1285), .Y(n2830)
         );
  OAI211XLTS U737 ( .A0(n3911), .A1(n4399), .B0(n1282), .C0(n1283), .Y(n2831)
         );
  OAI211XLTS U738 ( .A0(n3916), .A1(n4168), .B0(n2042), .C0(n2043), .Y(n2460)
         );
  OAI211XLTS U739 ( .A0(n3905), .A1(n4156), .B0(n2034), .C0(n2035), .Y(n2464)
         );
  OAI211XLTS U740 ( .A0(n3906), .A1(n4474), .B0(n1332), .C0(n1333), .Y(n2806)
         );
  OAI211XLTS U741 ( .A0(n3906), .A1(n4471), .B0(n1330), .C0(n1331), .Y(n2807)
         );
  OAI211XLTS U742 ( .A0(n3907), .A1(n4459), .B0(n1322), .C0(n1323), .Y(n2811)
         );
  OAI211XLTS U743 ( .A0(n3916), .A1(n4450), .B0(n1316), .C0(n1317), .Y(n2814)
         );
  OAI211XLTS U744 ( .A0(n3910), .A1(n4417), .B0(n1294), .C0(n1295), .Y(n2825)
         );
  OAI211XLTS U745 ( .A0(n3911), .A1(n4405), .B0(n1286), .C0(n1287), .Y(n2829)
         );
  OAI211XLTS U746 ( .A0(n3911), .A1(n4396), .B0(n1280), .C0(n1281), .Y(n2832)
         );
  AOI2BB2XLTS U747 ( .B0(n1809), .B1(n1810), .A0N(n3719), .A1N(readOutbuffer_7), .Y(n2570) );
  AOI32XLTS U748 ( .A0(n1811), .A1(n1812), .A2(n1813), .B0(n4148), .B1(n949), 
        .Y(n1810) );
  NAND2XLTS U749 ( .A(n4141), .B(n129), .Y(n1831) );
  OAI211XLTS U750 ( .A0(n522), .A1(n3938), .B0(n1897), .C0(n1898), .Y(n2547)
         );
  OAI211XLTS U751 ( .A0(n521), .A1(n3935), .B0(n1895), .C0(n1896), .Y(n2548)
         );
  OAI211XLTS U752 ( .A0(n520), .A1(n3947), .B0(n1903), .C0(n1904), .Y(n2544)
         );
  OAI211XLTS U753 ( .A0(n522), .A1(n3950), .B0(n1905), .C0(n1906), .Y(n2543)
         );
  OAI211XLTS U754 ( .A0(n521), .A1(n3944), .B0(n1901), .C0(n1902), .Y(n2545)
         );
  OAI211XLTS U755 ( .A0(n520), .A1(n3941), .B0(n1899), .C0(n1900), .Y(n2546)
         );
  OAI211XLTS U756 ( .A0(n4135), .A1(n522), .B0(n1176), .C0(n1177), .Y(n2872)
         );
  OAI211XLTS U757 ( .A0(n4132), .A1(n521), .B0(n1174), .C0(n1175), .Y(n2873)
         );
  OAI211XLTS U758 ( .A0(n4129), .A1(n520), .B0(n1172), .C0(n1173), .Y(n2874)
         );
  OAI211XLTS U759 ( .A0(n4126), .A1(n520), .B0(n1170), .C0(n1171), .Y(n2875)
         );
  OAI211XLTS U760 ( .A0(n4123), .A1(n522), .B0(n1165), .C0(n1166), .Y(n2876)
         );
  OAI211XLTS U761 ( .A0(n4138), .A1(n521), .B0(n1178), .C0(n1179), .Y(n2871)
         );
  OAI211XLTS U762 ( .A0(n4495), .A1(n3913), .B0(n1270), .C0(n1271), .Y(n2837)
         );
  OAI211XLTS U763 ( .A0(n4492), .A1(n3913), .B0(n1268), .C0(n1269), .Y(n2838)
         );
  OAI211XLTS U764 ( .A0(n1119), .A1(n903), .B0(n1719), .C0(n1720), .Y(n2613)
         );
  OAI211XLTS U765 ( .A0(n1119), .A1(n901), .B0(n1723), .C0(n1724), .Y(n2611)
         );
  OAI211XLTS U766 ( .A0(n1119), .A1(n902), .B0(n1721), .C0(n1722), .Y(n2612)
         );
  OAI211XLTS U767 ( .A0(n3232), .A1(n861), .B0(n2022), .C0(n2023), .Y(n2473)
         );
  OAI211XLTS U768 ( .A0(n3562), .A1(n655), .B0(n1191), .C0(n1192), .Y(n2867)
         );
  OAI211XLTS U769 ( .A0(n3562), .A1(n653), .B0(n1187), .C0(n1188), .Y(n2869)
         );
  OAI211XLTS U770 ( .A0(n3232), .A1(n890), .B0(n1255), .C0(n1256), .Y(n2843)
         );
  OAI211XLTS U771 ( .A0(n3232), .A1(n888), .B0(n1251), .C0(n1252), .Y(n2845)
         );
  OAI211XLTS U772 ( .A0(n3422), .A1(n4201), .B0(n1470), .C0(n1471), .Y(n2737)
         );
  OAI211XLTS U773 ( .A0(n3422), .A1(n4198), .B0(n1468), .C0(n1469), .Y(n2738)
         );
  OAI211XLTS U774 ( .A0(n4489), .A1(n3913), .B0(n1266), .C0(n1267), .Y(n2839)
         );
  OAI211XLTS U775 ( .A0(n4486), .A1(n3913), .B0(n1261), .C0(n1262), .Y(n2840)
         );
  OAI211XLTS U776 ( .A0(n3562), .A1(n642), .B0(n1928), .C0(n1929), .Y(n2529)
         );
  OAI211XLTS U777 ( .A0(n3370), .A1(n4297), .B0(n1406), .C0(n1407), .Y(n2769)
         );
  OAI211XLTS U778 ( .A0(n3370), .A1(n4294), .B0(n1404), .C0(n1405), .Y(n2770)
         );
  OAI211XLTS U779 ( .A0(n3414), .A1(n3980), .B0(n1965), .C0(n1966), .Y(n2505)
         );
  OAI211XLTS U780 ( .A0(n3414), .A1(n3977), .B0(n1963), .C0(n1964), .Y(n2506)
         );
  OAI211XLTS U781 ( .A0(n3414), .A1(n4291), .B0(n1530), .C0(n1531), .Y(n2707)
         );
  OAI211XLTS U782 ( .A0(n3414), .A1(n4288), .B0(n1528), .C0(n1529), .Y(n2708)
         );
  OAI211XLTS U783 ( .A0(n3415), .A1(n4285), .B0(n1526), .C0(n1527), .Y(n2709)
         );
  OAI211XLTS U784 ( .A0(n3415), .A1(n4282), .B0(n1524), .C0(n1525), .Y(n2710)
         );
  OAI211XLTS U785 ( .A0(n3415), .A1(n4279), .B0(n1522), .C0(n1523), .Y(n2711)
         );
  OAI211XLTS U786 ( .A0(n3415), .A1(n4276), .B0(n1520), .C0(n1521), .Y(n2712)
         );
  OAI211XLTS U787 ( .A0(n3416), .A1(n4270), .B0(n1516), .C0(n1517), .Y(n2714)
         );
  OAI211XLTS U788 ( .A0(n3416), .A1(n4264), .B0(n1512), .C0(n1513), .Y(n2716)
         );
  OAI211XLTS U789 ( .A0(n3417), .A1(n4261), .B0(n1510), .C0(n1511), .Y(n2717)
         );
  OAI211XLTS U790 ( .A0(n3417), .A1(n4255), .B0(n1506), .C0(n1507), .Y(n2719)
         );
  OAI211XLTS U791 ( .A0(n3418), .A1(n4249), .B0(n1502), .C0(n1503), .Y(n2721)
         );
  OAI211XLTS U792 ( .A0(n3418), .A1(n4246), .B0(n1500), .C0(n1501), .Y(n2722)
         );
  OAI211XLTS U793 ( .A0(n3418), .A1(n4240), .B0(n1496), .C0(n1497), .Y(n2724)
         );
  OAI211XLTS U794 ( .A0(n3419), .A1(n4234), .B0(n1492), .C0(n1493), .Y(n2726)
         );
  OAI211XLTS U795 ( .A0(n3419), .A1(n4231), .B0(n1490), .C0(n1491), .Y(n2727)
         );
  OAI211XLTS U796 ( .A0(n3419), .A1(n4228), .B0(n1488), .C0(n1489), .Y(n2728)
         );
  OAI211XLTS U797 ( .A0(n3420), .A1(n4225), .B0(n1486), .C0(n1487), .Y(n2729)
         );
  OAI211XLTS U798 ( .A0(n3420), .A1(n4222), .B0(n1484), .C0(n1485), .Y(n2730)
         );
  OAI211XLTS U799 ( .A0(n3420), .A1(n4216), .B0(n1480), .C0(n1481), .Y(n2732)
         );
  OAI211XLTS U800 ( .A0(n3421), .A1(n4207), .B0(n1474), .C0(n1475), .Y(n2735)
         );
  OAI211XLTS U801 ( .A0(n3416), .A1(n4273), .B0(n1518), .C0(n1519), .Y(n2713)
         );
  OAI211XLTS U802 ( .A0(n3416), .A1(n4267), .B0(n1514), .C0(n1515), .Y(n2715)
         );
  OAI211XLTS U803 ( .A0(n3417), .A1(n4258), .B0(n1508), .C0(n1509), .Y(n2718)
         );
  OAI211XLTS U804 ( .A0(n3417), .A1(n4252), .B0(n1504), .C0(n1505), .Y(n2720)
         );
  OAI211XLTS U805 ( .A0(n3418), .A1(n4243), .B0(n1498), .C0(n1499), .Y(n2723)
         );
  OAI211XLTS U806 ( .A0(n3419), .A1(n4237), .B0(n1494), .C0(n1495), .Y(n2725)
         );
  OAI211XLTS U807 ( .A0(n3421), .A1(n4213), .B0(n1478), .C0(n1479), .Y(n2733)
         );
  OAI211XLTS U808 ( .A0(n3421), .A1(n4210), .B0(n1476), .C0(n1477), .Y(n2734)
         );
  OAI211XLTS U809 ( .A0(n3421), .A1(n4204), .B0(n1472), .C0(n1473), .Y(n2736)
         );
  OAI211XLTS U810 ( .A0(n3420), .A1(n4219), .B0(n1482), .C0(n1483), .Y(n2731)
         );
  OAI211XLTS U811 ( .A0(n3413), .A1(n3992), .B0(n1973), .C0(n1974), .Y(n2501)
         );
  OAI211XLTS U812 ( .A0(n3413), .A1(n3989), .B0(n1971), .C0(n1972), .Y(n2502)
         );
  OAI211XLTS U813 ( .A0(n3413), .A1(n3986), .B0(n1969), .C0(n1970), .Y(n2503)
         );
  OAI211XLTS U814 ( .A0(n3413), .A1(n3983), .B0(n1967), .C0(n1968), .Y(n2504)
         );
  OAI211XLTS U815 ( .A0(n3361), .A1(n3941), .B0(n1991), .C0(n1992), .Y(n2490)
         );
  OAI211XLTS U816 ( .A0(n3362), .A1(n4384), .B0(n1464), .C0(n1465), .Y(n2740)
         );
  OAI211XLTS U817 ( .A0(n3363), .A1(n4381), .B0(n1462), .C0(n1463), .Y(n2741)
         );
  OAI211XLTS U818 ( .A0(n3363), .A1(n4378), .B0(n1460), .C0(n1461), .Y(n2742)
         );
  OAI211XLTS U819 ( .A0(n3363), .A1(n4372), .B0(n1456), .C0(n1457), .Y(n2744)
         );
  OAI211XLTS U820 ( .A0(n3364), .A1(n4369), .B0(n1454), .C0(n1455), .Y(n2745)
         );
  OAI211XLTS U821 ( .A0(n3364), .A1(n4363), .B0(n1450), .C0(n1451), .Y(n2747)
         );
  OAI211XLTS U822 ( .A0(n3365), .A1(n4357), .B0(n1446), .C0(n1447), .Y(n2749)
         );
  OAI211XLTS U823 ( .A0(n3365), .A1(n4354), .B0(n1444), .C0(n1445), .Y(n2750)
         );
  OAI211XLTS U824 ( .A0(n3365), .A1(n4351), .B0(n1442), .C0(n1443), .Y(n2751)
         );
  OAI211XLTS U825 ( .A0(n3365), .A1(n4348), .B0(n1440), .C0(n1441), .Y(n2752)
         );
  OAI211XLTS U826 ( .A0(n3366), .A1(n4345), .B0(n1438), .C0(n1439), .Y(n2753)
         );
  OAI211XLTS U827 ( .A0(n3366), .A1(n4339), .B0(n1434), .C0(n1435), .Y(n2755)
         );
  OAI211XLTS U828 ( .A0(n3366), .A1(n4336), .B0(n1432), .C0(n1433), .Y(n2756)
         );
  OAI211XLTS U829 ( .A0(n3367), .A1(n4333), .B0(n1430), .C0(n1431), .Y(n2757)
         );
  OAI211XLTS U830 ( .A0(n3367), .A1(n4330), .B0(n1428), .C0(n1429), .Y(n2758)
         );
  OAI211XLTS U831 ( .A0(n3367), .A1(n4327), .B0(n1426), .C0(n1427), .Y(n2759)
         );
  OAI211XLTS U832 ( .A0(n3368), .A1(n4321), .B0(n1422), .C0(n1423), .Y(n2761)
         );
  OAI211XLTS U833 ( .A0(n3368), .A1(n4318), .B0(n1420), .C0(n1421), .Y(n2762)
         );
  OAI211XLTS U834 ( .A0(n3368), .A1(n4315), .B0(n1418), .C0(n1419), .Y(n2763)
         );
  OAI211XLTS U835 ( .A0(n3369), .A1(n4309), .B0(n1414), .C0(n1415), .Y(n2765)
         );
  OAI211XLTS U836 ( .A0(n3369), .A1(n4306), .B0(n1412), .C0(n1413), .Y(n2766)
         );
  OAI211XLTS U837 ( .A0(n3369), .A1(n4303), .B0(n1410), .C0(n1411), .Y(n2767)
         );
  OAI211XLTS U838 ( .A0(n3361), .A1(n3950), .B0(n1997), .C0(n1998), .Y(n2487)
         );
  OAI211XLTS U839 ( .A0(n3361), .A1(n3947), .B0(n1995), .C0(n1996), .Y(n2488)
         );
  OAI211XLTS U840 ( .A0(n3361), .A1(n3944), .B0(n1993), .C0(n1994), .Y(n2489)
         );
  OAI211XLTS U841 ( .A0(n3362), .A1(n3938), .B0(n1989), .C0(n1990), .Y(n2491)
         );
  OAI211XLTS U842 ( .A0(n3362), .A1(n3935), .B0(n1987), .C0(n1988), .Y(n2492)
         );
  OAI211XLTS U843 ( .A0(n3363), .A1(n4375), .B0(n1458), .C0(n1459), .Y(n2743)
         );
  OAI211XLTS U844 ( .A0(n3367), .A1(n4324), .B0(n1424), .C0(n1425), .Y(n2760)
         );
  OAI211XLTS U845 ( .A0(n3362), .A1(n4387), .B0(n1466), .C0(n1467), .Y(n2739)
         );
  OAI211XLTS U846 ( .A0(n3364), .A1(n4366), .B0(n1452), .C0(n1453), .Y(n2746)
         );
  OAI211XLTS U847 ( .A0(n3364), .A1(n4360), .B0(n1448), .C0(n1449), .Y(n2748)
         );
  OAI211XLTS U848 ( .A0(n3366), .A1(n4342), .B0(n1436), .C0(n1437), .Y(n2754)
         );
  OAI211XLTS U849 ( .A0(n3368), .A1(n4312), .B0(n1416), .C0(n1417), .Y(n2764)
         );
  OAI211XLTS U850 ( .A0(n3369), .A1(n4300), .B0(n1408), .C0(n1409), .Y(n2768)
         );
  OAI211XLTS U851 ( .A0(n1126), .A1(n928), .B0(n1669), .C0(n1670), .Y(n2638)
         );
  OAI211XLTS U852 ( .A0(n1125), .A1(n927), .B0(n1671), .C0(n1672), .Y(n2637)
         );
  OAI211XLTS U853 ( .A0(n1125), .A1(n926), .B0(n1673), .C0(n1674), .Y(n2636)
         );
  OAI211XLTS U854 ( .A0(n1125), .A1(n925), .B0(n1675), .C0(n1676), .Y(n2635)
         );
  OAI211XLTS U855 ( .A0(n1125), .A1(n924), .B0(n1677), .C0(n1678), .Y(n2634)
         );
  OAI211XLTS U856 ( .A0(n1124), .A1(n923), .B0(n1679), .C0(n1680), .Y(n2633)
         );
  OAI211XLTS U857 ( .A0(n1124), .A1(n922), .B0(n1681), .C0(n1682), .Y(n2632)
         );
  OAI211XLTS U858 ( .A0(n1124), .A1(n921), .B0(n1683), .C0(n1684), .Y(n2631)
         );
  OAI211XLTS U859 ( .A0(n1124), .A1(n920), .B0(n1685), .C0(n1686), .Y(n2630)
         );
  OAI211XLTS U860 ( .A0(n1123), .A1(n919), .B0(n1687), .C0(n1688), .Y(n2629)
         );
  OAI211XLTS U861 ( .A0(n1123), .A1(n918), .B0(n1689), .C0(n1690), .Y(n2628)
         );
  OAI211XLTS U862 ( .A0(n1123), .A1(n917), .B0(n1691), .C0(n1692), .Y(n2627)
         );
  OAI211XLTS U863 ( .A0(n1123), .A1(n916), .B0(n1693), .C0(n1694), .Y(n2626)
         );
  OAI211XLTS U864 ( .A0(n1122), .A1(n915), .B0(n1695), .C0(n1696), .Y(n2625)
         );
  OAI211XLTS U865 ( .A0(n1122), .A1(n914), .B0(n1697), .C0(n1698), .Y(n2624)
         );
  OAI211XLTS U866 ( .A0(n1122), .A1(n913), .B0(n1699), .C0(n1700), .Y(n2623)
         );
  OAI211XLTS U867 ( .A0(n1122), .A1(n912), .B0(n1701), .C0(n1702), .Y(n2622)
         );
  OAI211XLTS U868 ( .A0(n1121), .A1(n911), .B0(n1703), .C0(n1704), .Y(n2621)
         );
  OAI211XLTS U869 ( .A0(n1121), .A1(n910), .B0(n1705), .C0(n1706), .Y(n2620)
         );
  OAI211XLTS U870 ( .A0(n1121), .A1(n909), .B0(n1707), .C0(n1708), .Y(n2619)
         );
  OAI211XLTS U871 ( .A0(n1121), .A1(n908), .B0(n1709), .C0(n1710), .Y(n2618)
         );
  OAI211XLTS U872 ( .A0(n1120), .A1(n907), .B0(n1711), .C0(n1712), .Y(n2617)
         );
  OAI211XLTS U873 ( .A0(n1120), .A1(n906), .B0(n1713), .C0(n1714), .Y(n2616)
         );
  OAI211XLTS U874 ( .A0(n1120), .A1(n905), .B0(n1715), .C0(n1716), .Y(n2615)
         );
  OAI211XLTS U875 ( .A0(n1120), .A1(n904), .B0(n1717), .C0(n1718), .Y(n2614)
         );
  OAI211XLTS U876 ( .A0(n1126), .A1(n931), .B0(n1663), .C0(n1664), .Y(n2641)
         );
  OAI211XLTS U877 ( .A0(n1126), .A1(n930), .B0(n1665), .C0(n1666), .Y(n2640)
         );
  OAI211XLTS U878 ( .A0(n1126), .A1(n929), .B0(n1667), .C0(n1668), .Y(n2639)
         );
  OAI211XLTS U879 ( .A0(n3563), .A1(n967), .B0(n1596), .C0(n1597), .Y(n2674)
         );
  OAI211XLTS U880 ( .A0(n3571), .A1(n647), .B0(n1658), .C0(n1659), .Y(n2643)
         );
  OAI211XLTS U881 ( .A0(n3568), .A1(n646), .B0(n1628), .C0(n1629), .Y(n2658)
         );
  OAI211XLTS U882 ( .A0(n3567), .A1(n645), .B0(n1626), .C0(n1627), .Y(n2659)
         );
  OAI211XLTS U883 ( .A0(n3566), .A1(n644), .B0(n1618), .C0(n1619), .Y(n2663)
         );
  OAI211XLTS U884 ( .A0(n3564), .A1(n643), .B0(n1598), .C0(n1599), .Y(n2673)
         );
  OAI211XLTS U885 ( .A0(n3571), .A1(n636), .B0(n1656), .C0(n1657), .Y(n2644)
         );
  OAI211XLTS U886 ( .A0(n3571), .A1(n635), .B0(n1654), .C0(n1655), .Y(n2645)
         );
  OAI211XLTS U887 ( .A0(n3571), .A1(n634), .B0(n1652), .C0(n1653), .Y(n2646)
         );
  OAI211XLTS U888 ( .A0(n3570), .A1(n633), .B0(n1650), .C0(n1651), .Y(n2647)
         );
  OAI211XLTS U889 ( .A0(n3570), .A1(n632), .B0(n1648), .C0(n1649), .Y(n2648)
         );
  OAI211XLTS U890 ( .A0(n3570), .A1(n631), .B0(n1646), .C0(n1647), .Y(n2649)
         );
  OAI211XLTS U891 ( .A0(n3570), .A1(n630), .B0(n1644), .C0(n1645), .Y(n2650)
         );
  OAI211XLTS U892 ( .A0(n3569), .A1(n629), .B0(n1642), .C0(n1643), .Y(n2651)
         );
  OAI211XLTS U893 ( .A0(n3569), .A1(n628), .B0(n1640), .C0(n1641), .Y(n2652)
         );
  OAI211XLTS U894 ( .A0(n3569), .A1(n627), .B0(n1638), .C0(n1639), .Y(n2653)
         );
  OAI211XLTS U895 ( .A0(n3569), .A1(n626), .B0(n1636), .C0(n1637), .Y(n2654)
         );
  OAI211XLTS U896 ( .A0(n3568), .A1(n625), .B0(n1634), .C0(n1635), .Y(n2655)
         );
  OAI211XLTS U897 ( .A0(n3568), .A1(n624), .B0(n1632), .C0(n1633), .Y(n2656)
         );
  OAI211XLTS U898 ( .A0(n3568), .A1(n623), .B0(n1630), .C0(n1631), .Y(n2657)
         );
  OAI211XLTS U899 ( .A0(n3567), .A1(n622), .B0(n1624), .C0(n1625), .Y(n2660)
         );
  OAI211XLTS U900 ( .A0(n3567), .A1(n621), .B0(n1622), .C0(n1623), .Y(n2661)
         );
  OAI211XLTS U901 ( .A0(n3566), .A1(n620), .B0(n1620), .C0(n1621), .Y(n2662)
         );
  OAI211XLTS U902 ( .A0(n3566), .A1(n619), .B0(n1616), .C0(n1617), .Y(n2664)
         );
  OAI211XLTS U903 ( .A0(n3566), .A1(n618), .B0(n1614), .C0(n1615), .Y(n2665)
         );
  OAI211XLTS U904 ( .A0(n3565), .A1(n617), .B0(n1612), .C0(n1613), .Y(n2666)
         );
  OAI211XLTS U905 ( .A0(n3565), .A1(n616), .B0(n1610), .C0(n1611), .Y(n2667)
         );
  OAI211XLTS U906 ( .A0(n3565), .A1(n615), .B0(n1608), .C0(n1609), .Y(n2668)
         );
  OAI211XLTS U907 ( .A0(n3565), .A1(n614), .B0(n1606), .C0(n1607), .Y(n2669)
         );
  OAI211XLTS U908 ( .A0(n3564), .A1(n613), .B0(n1604), .C0(n1605), .Y(n2670)
         );
  OAI211XLTS U909 ( .A0(n3564), .A1(n612), .B0(n1602), .C0(n1603), .Y(n2671)
         );
  OAI211XLTS U910 ( .A0(n3564), .A1(n611), .B0(n1600), .C0(n1601), .Y(n2672)
         );
  OAI211XLTS U911 ( .A0(n3240), .A1(n870), .B0(n1394), .C0(n1395), .Y(n2775)
         );
  OAI211XLTS U912 ( .A0(n3239), .A1(n869), .B0(n1384), .C0(n1385), .Y(n2780)
         );
  OAI211XLTS U913 ( .A0(n3239), .A1(n868), .B0(n1380), .C0(n1381), .Y(n2782)
         );
  OAI211XLTS U914 ( .A0(n3238), .A1(n867), .B0(n1378), .C0(n1379), .Y(n2783)
         );
  OAI211XLTS U915 ( .A0(n3236), .A1(n866), .B0(n1360), .C0(n1361), .Y(n2792)
         );
  OAI211XLTS U916 ( .A0(n3235), .A1(n865), .B0(n1356), .C0(n1357), .Y(n2794)
         );
  OAI211XLTS U917 ( .A0(n3235), .A1(n864), .B0(n1350), .C0(n1351), .Y(n2797)
         );
  OAI211XLTS U918 ( .A0(n3234), .A1(n863), .B0(n1344), .C0(n1345), .Y(n2800)
         );
  OAI211XLTS U919 ( .A0(n3241), .A1(n856), .B0(n1402), .C0(n1403), .Y(n2771)
         );
  OAI211XLTS U920 ( .A0(n3241), .A1(n855), .B0(n1400), .C0(n1401), .Y(n2772)
         );
  OAI211XLTS U921 ( .A0(n3241), .A1(n854), .B0(n1398), .C0(n1399), .Y(n2773)
         );
  OAI211XLTS U922 ( .A0(n3241), .A1(n853), .B0(n1396), .C0(n1397), .Y(n2774)
         );
  OAI211XLTS U923 ( .A0(n3240), .A1(n852), .B0(n1392), .C0(n1393), .Y(n2776)
         );
  OAI211XLTS U924 ( .A0(n3240), .A1(n851), .B0(n1390), .C0(n1391), .Y(n2777)
         );
  OAI211XLTS U925 ( .A0(n3240), .A1(n850), .B0(n1388), .C0(n1389), .Y(n2778)
         );
  OAI211XLTS U926 ( .A0(n3239), .A1(n849), .B0(n1386), .C0(n1387), .Y(n2779)
         );
  OAI211XLTS U927 ( .A0(n3239), .A1(n848), .B0(n1382), .C0(n1383), .Y(n2781)
         );
  OAI211XLTS U928 ( .A0(n3238), .A1(n847), .B0(n1376), .C0(n1377), .Y(n2784)
         );
  OAI211XLTS U929 ( .A0(n3238), .A1(n846), .B0(n1374), .C0(n1375), .Y(n2785)
         );
  OAI211XLTS U930 ( .A0(n3238), .A1(n845), .B0(n1372), .C0(n1373), .Y(n2786)
         );
  OAI211XLTS U931 ( .A0(n3237), .A1(n844), .B0(n1370), .C0(n1371), .Y(n2787)
         );
  OAI211XLTS U932 ( .A0(n3237), .A1(n843), .B0(n1368), .C0(n1369), .Y(n2788)
         );
  OAI211XLTS U933 ( .A0(n3237), .A1(n842), .B0(n1366), .C0(n1367), .Y(n2789)
         );
  OAI211XLTS U934 ( .A0(n3236), .A1(n841), .B0(n1364), .C0(n1365), .Y(n2790)
         );
  OAI211XLTS U935 ( .A0(n3236), .A1(n840), .B0(n1362), .C0(n1363), .Y(n2791)
         );
  OAI211XLTS U936 ( .A0(n3236), .A1(n839), .B0(n1358), .C0(n1359), .Y(n2793)
         );
  OAI211XLTS U937 ( .A0(n3235), .A1(n838), .B0(n1354), .C0(n1355), .Y(n2795)
         );
  OAI211XLTS U938 ( .A0(n3235), .A1(n837), .B0(n1352), .C0(n1353), .Y(n2796)
         );
  OAI211XLTS U939 ( .A0(n3234), .A1(n836), .B0(n1348), .C0(n1349), .Y(n2798)
         );
  OAI211XLTS U940 ( .A0(n3234), .A1(n835), .B0(n1346), .C0(n1347), .Y(n2799)
         );
  OAI211XLTS U941 ( .A0(n3234), .A1(n834), .B0(n1342), .C0(n1343), .Y(n2801)
         );
  OAI211XLTS U942 ( .A0(n3233), .A1(n797), .B0(n1340), .C0(n1341), .Y(n2802)
         );
  OAI211XLTS U943 ( .A0(n3563), .A1(n654), .B0(n1189), .C0(n1190), .Y(n2868)
         );
  OAI211XLTS U944 ( .A0(n3563), .A1(n657), .B0(n1195), .C0(n1196), .Y(n2865)
         );
  OAI211XLTS U945 ( .A0(n3563), .A1(n656), .B0(n1193), .C0(n1194), .Y(n2866)
         );
  OAI211XLTS U946 ( .A0(n3567), .A1(n652), .B0(n1181), .C0(n1182), .Y(n2870)
         );
  OAI211XLTS U947 ( .A0(n3572), .A1(n640), .B0(n1924), .C0(n1925), .Y(n2531)
         );
  OAI211XLTS U948 ( .A0(n3572), .A1(n639), .B0(n1922), .C0(n1923), .Y(n2532)
         );
  OAI211XLTS U949 ( .A0(n3572), .A1(n638), .B0(n1920), .C0(n1921), .Y(n2533)
         );
  OAI211XLTS U950 ( .A0(n3572), .A1(n637), .B0(n1918), .C0(n1919), .Y(n2534)
         );
  OAI211XLTS U951 ( .A0(n3233), .A1(n889), .B0(n1253), .C0(n1254), .Y(n2844)
         );
  OAI211XLTS U952 ( .A0(n3233), .A1(n892), .B0(n1259), .C0(n1260), .Y(n2841)
         );
  OAI211XLTS U953 ( .A0(n3233), .A1(n891), .B0(n1257), .C0(n1258), .Y(n2842)
         );
  OAI211XLTS U954 ( .A0(n3237), .A1(n887), .B0(n1245), .C0(n1246), .Y(n2846)
         );
  OAI211XLTS U955 ( .A0(n3242), .A1(n860), .B0(n2018), .C0(n2019), .Y(n2475)
         );
  OAI211XLTS U956 ( .A0(n3242), .A1(n859), .B0(n2016), .C0(n2017), .Y(n2476)
         );
  OAI211XLTS U957 ( .A0(n3242), .A1(n858), .B0(n2014), .C0(n2015), .Y(n2477)
         );
  OAI211XLTS U958 ( .A0(n3242), .A1(n857), .B0(n2012), .C0(n2013), .Y(n2478)
         );
  OAI211XLTS U959 ( .A0(n4026), .A1(n3423), .B0(n1222), .C0(n1223), .Y(n2855)
         );
  OAI211XLTS U960 ( .A0(n4023), .A1(n3423), .B0(n1220), .C0(n1221), .Y(n2856)
         );
  OAI211XLTS U961 ( .A0(n4020), .A1(n3423), .B0(n1218), .C0(n1219), .Y(n2857)
         );
  OAI211XLTS U962 ( .A0(n4017), .A1(n3423), .B0(n1214), .C0(n1215), .Y(n2858)
         );
  OAI211XLTS U963 ( .A0(n4029), .A1(n3422), .B0(n1224), .C0(n1225), .Y(n2854)
         );
  OAI211XLTS U964 ( .A0(n4032), .A1(n3422), .B0(n1226), .C0(n1227), .Y(n2853)
         );
  OAI211XLTS U965 ( .A0(n4135), .A1(n3370), .B0(n1240), .C0(n1241), .Y(n2848)
         );
  OAI211XLTS U966 ( .A0(n4138), .A1(n3370), .B0(n1242), .C0(n1243), .Y(n2847)
         );
  OAI211XLTS U967 ( .A0(n4126), .A1(n3371), .B0(n1234), .C0(n1235), .Y(n2851)
         );
  OAI211XLTS U968 ( .A0(n4123), .A1(n3371), .B0(n1229), .C0(n1230), .Y(n2852)
         );
  OAI211XLTS U969 ( .A0(n4132), .A1(n3371), .B0(n1238), .C0(n1239), .Y(n2849)
         );
  OAI211XLTS U970 ( .A0(n4129), .A1(n3371), .B0(n1236), .C0(n1237), .Y(n2850)
         );
  OAI211XLTS U971 ( .A0(n1127), .A1(n932), .B0(n1661), .C0(n1662), .Y(n2642)
         );
  INVXLTS U972 ( .A(n1128), .Y(n1127) );
  OAI211XLTS U973 ( .A0(n3243), .A1(n872), .B0(n2020), .C0(n2021), .Y(n2474)
         );
  INVXLTS U974 ( .A(n3244), .Y(n3243) );
  OAI211XLTS U975 ( .A0(n3573), .A1(n641), .B0(n1926), .C0(n1927), .Y(n2530)
         );
  INVXLTS U976 ( .A(n3574), .Y(n3573) );
  OAI211XLTS U977 ( .A0(n3708), .A1(n882), .B0(n1158), .C0(n1159), .Y(n2879)
         );
  OAI211XLTS U978 ( .A0(n3708), .A1(n881), .B0(n1154), .C0(n1155), .Y(n2881)
         );
  OAI211XLTS U979 ( .A0(n3717), .A1(n833), .B0(n1876), .C0(n1877), .Y(n2557)
         );
  OAI211XLTS U980 ( .A0(n3709), .A1(n885), .B0(n1162), .C0(n1163), .Y(n2877)
         );
  OAI211XLTS U981 ( .A0(n3708), .A1(n884), .B0(n1160), .C0(n1161), .Y(n2878)
         );
  OAI211XLTS U982 ( .A0(n3708), .A1(n883), .B0(n1156), .C0(n1157), .Y(n2880)
         );
  OAI211XLTS U983 ( .A0(n3713), .A1(n880), .B0(n1147), .C0(n1148), .Y(n2882)
         );
  OAI211XLTS U984 ( .A0(n3716), .A1(n829), .B0(n1787), .C0(n1788), .Y(n2579)
         );
  OAI211XLTS U985 ( .A0(n3716), .A1(n828), .B0(n1785), .C0(n1786), .Y(n2580)
         );
  OAI211XLTS U986 ( .A0(n3715), .A1(n827), .B0(n1783), .C0(n1784), .Y(n2581)
         );
  OAI211XLTS U987 ( .A0(n3715), .A1(n826), .B0(n1781), .C0(n1782), .Y(n2582)
         );
  OAI211XLTS U988 ( .A0(n3715), .A1(n825), .B0(n1779), .C0(n1780), .Y(n2583)
         );
  OAI211XLTS U989 ( .A0(n3715), .A1(n824), .B0(n1777), .C0(n1778), .Y(n2584)
         );
  OAI211XLTS U990 ( .A0(n3714), .A1(n823), .B0(n1775), .C0(n1776), .Y(n2585)
         );
  OAI211XLTS U991 ( .A0(n3714), .A1(n822), .B0(n1773), .C0(n1774), .Y(n2586)
         );
  OAI211XLTS U992 ( .A0(n3714), .A1(n821), .B0(n1771), .C0(n1772), .Y(n2587)
         );
  OAI211XLTS U993 ( .A0(n3714), .A1(n820), .B0(n1769), .C0(n1770), .Y(n2588)
         );
  OAI211XLTS U994 ( .A0(n3720), .A1(n819), .B0(n1767), .C0(n1768), .Y(n2589)
         );
  OAI211XLTS U995 ( .A0(n3721), .A1(n818), .B0(n1765), .C0(n1766), .Y(n2590)
         );
  OAI211XLTS U996 ( .A0(n3718), .A1(n817), .B0(n1763), .C0(n1764), .Y(n2591)
         );
  OAI211XLTS U997 ( .A0(n1146), .A1(n816), .B0(n1761), .C0(n1762), .Y(n2592)
         );
  OAI211XLTS U998 ( .A0(n3713), .A1(n815), .B0(n1759), .C0(n1760), .Y(n2593)
         );
  OAI211XLTS U999 ( .A0(n3713), .A1(n814), .B0(n1757), .C0(n1758), .Y(n2594)
         );
  OAI211XLTS U1000 ( .A0(n3713), .A1(n813), .B0(n1755), .C0(n1756), .Y(n2595)
         );
  OAI211XLTS U1001 ( .A0(n3712), .A1(n812), .B0(n1753), .C0(n1754), .Y(n2596)
         );
  OAI211XLTS U1002 ( .A0(n3712), .A1(n811), .B0(n1751), .C0(n1752), .Y(n2597)
         );
  OAI211XLTS U1003 ( .A0(n3712), .A1(n810), .B0(n1749), .C0(n1750), .Y(n2598)
         );
  OAI211XLTS U1004 ( .A0(n3712), .A1(n809), .B0(n1747), .C0(n1748), .Y(n2599)
         );
  OAI211XLTS U1005 ( .A0(n3711), .A1(n808), .B0(n1745), .C0(n1746), .Y(n2600)
         );
  OAI211XLTS U1006 ( .A0(n3711), .A1(n807), .B0(n1743), .C0(n1744), .Y(n2601)
         );
  OAI211XLTS U1007 ( .A0(n3711), .A1(n806), .B0(n1741), .C0(n1742), .Y(n2602)
         );
  OAI211XLTS U1008 ( .A0(n3711), .A1(n805), .B0(n1739), .C0(n1740), .Y(n2603)
         );
  OAI211XLTS U1009 ( .A0(n3710), .A1(n804), .B0(n1737), .C0(n1738), .Y(n2604)
         );
  OAI211XLTS U1010 ( .A0(n3710), .A1(n803), .B0(n1735), .C0(n1736), .Y(n2605)
         );
  OAI211XLTS U1011 ( .A0(n3710), .A1(n802), .B0(n1733), .C0(n1734), .Y(n2606)
         );
  OAI211XLTS U1012 ( .A0(n3710), .A1(n801), .B0(n1731), .C0(n1732), .Y(n2607)
         );
  OAI211XLTS U1013 ( .A0(n3709), .A1(n800), .B0(n1729), .C0(n1730), .Y(n2608)
         );
  OAI211XLTS U1014 ( .A0(n3709), .A1(n799), .B0(n1727), .C0(n1728), .Y(n2609)
         );
  OAI211XLTS U1015 ( .A0(n3709), .A1(n798), .B0(n1725), .C0(n1726), .Y(n2610)
         );
  OAI211XLTS U1016 ( .A0(n3716), .A1(n862), .B0(n1866), .C0(n1867), .Y(n2562)
         );
  OAI211XLTS U1017 ( .A0(n3717), .A1(n832), .B0(n1872), .C0(n1873), .Y(n2559)
         );
  OAI211XLTS U1018 ( .A0(n3717), .A1(n831), .B0(n1870), .C0(n1871), .Y(n2560)
         );
  OAI211XLTS U1019 ( .A0(n3716), .A1(n830), .B0(n1868), .C0(n1869), .Y(n2561)
         );
  OAI211XLTS U1020 ( .A0(n3717), .A1(n796), .B0(n1874), .C0(n1875), .Y(n2558)
         );
  AOI32XLTS U1021 ( .A0(n23), .A1(n1847), .A2(n1848), .B0(n3819), .B1(n751), 
        .Y(n2565) );
  AOI32XLTS U1022 ( .A0(n162), .A1(n1861), .A2(n1862), .B0(n3897), .B1(n886), 
        .Y(n2563) );
  AOI21XLTS U1023 ( .A0(readIn_NORTH), .A1(n1863), .B0(n1864), .Y(n1862) );
  AOI32XLTS U1024 ( .A0(n130), .A1(n1817), .A2(n1818), .B0(n1153), .B1(n649), 
        .Y(n2569) );
  NAND4XLTS U1025 ( .A(n429), .B(n2962), .C(n2), .D(n523), .Y(n2071) );
  NAND4XLTS U1026 ( .A(n423), .B(n432), .C(n1029), .D(n426), .Y(n2070) );
  NAND2X1TS U1027 ( .A(n10), .B(n173), .Y(n2024) );
  NAND2X1TS U1028 ( .A(n166), .B(n165), .Y(n1141) );
  NOR2X1TS U1029 ( .A(n1141), .B(n8), .Y(n2096) );
  NAND3X1TS U1030 ( .A(n168), .B(n160), .C(n459), .Y(n2081) );
  NAND3X1TS U1031 ( .A(n12), .B(n160), .C(n8), .Y(n2083) );
  NAND3X1TS U1032 ( .A(n11), .B(n440), .C(n125), .Y(n2080) );
  NAND3X1TS U1033 ( .A(n125), .B(n430), .C(n8), .Y(n2082) );
  NAND3XLTS U1034 ( .A(n435), .B(n432), .C(n422), .Y(n2072) );
  NAND4XLTS U1035 ( .A(selectBit_WEST), .B(n435), .C(n1130), .D(n2), .Y(n2073)
         );
  NAND4XLTS U1036 ( .A(readReady), .B(n435), .C(n2), .D(n1084), .Y(n2074) );
  AND3XLTS U1037 ( .A(n2962), .B(n450), .C(n435), .Y(n2064) );
  CLKBUFX2TS U1038 ( .A(n3887), .Y(n3878) );
  CLKBUFX2TS U1039 ( .A(n3776), .Y(n3767) );
  CLKBUFX2TS U1040 ( .A(n769), .Y(n3884) );
  CLKBUFX2TS U1041 ( .A(n3885), .Y(n3883) );
  CLKBUFX2TS U1042 ( .A(n3885), .Y(n3882) );
  CLKBUFX2TS U1043 ( .A(n3886), .Y(n3881) );
  CLKBUFX2TS U1044 ( .A(n3886), .Y(n3880) );
  CLKBUFX2TS U1045 ( .A(n3887), .Y(n3879) );
  CLKBUFX2TS U1046 ( .A(n3779), .Y(n3773) );
  CLKBUFX2TS U1047 ( .A(n3774), .Y(n3772) );
  CLKBUFX2TS U1048 ( .A(n3774), .Y(n3771) );
  CLKBUFX2TS U1049 ( .A(n3775), .Y(n3770) );
  CLKBUFX2TS U1050 ( .A(n3775), .Y(n3769) );
  CLKBUFX2TS U1051 ( .A(n3776), .Y(n3768) );
  CLKBUFX2TS U1052 ( .A(n3748), .Y(n3740) );
  CLKBUFX2TS U1053 ( .A(n3748), .Y(n3741) );
  CLKBUFX2TS U1054 ( .A(n3747), .Y(n3742) );
  CLKBUFX2TS U1055 ( .A(n3747), .Y(n3743) );
  CLKBUFX2TS U1056 ( .A(n3746), .Y(n3744) );
  CLKBUFX2TS U1057 ( .A(n3929), .Y(n3920) );
  CLKBUFX2TS U1058 ( .A(n3834), .Y(n3824) );
  CLKBUFX2TS U1059 ( .A(n3928), .Y(n3923) );
  CLKBUFX2TS U1060 ( .A(n3834), .Y(n3829) );
  CLKBUFX2TS U1061 ( .A(n3834), .Y(n3832) );
  CLKBUFX2TS U1062 ( .A(n3833), .Y(n3830) );
  CLKBUFX2TS U1063 ( .A(n775), .Y(n3827) );
  CLKBUFX2TS U1064 ( .A(n3926), .Y(n3925) );
  CLKBUFX2TS U1065 ( .A(n3926), .Y(n3924) );
  CLKBUFX2TS U1066 ( .A(n3928), .Y(n3922) );
  CLKBUFX2TS U1067 ( .A(n3929), .Y(n3921) );
  CLKBUFX2TS U1068 ( .A(n3833), .Y(n3831) );
  CLKBUFX2TS U1069 ( .A(n3834), .Y(n3828) );
  CLKBUFX2TS U1070 ( .A(n775), .Y(n3826) );
  CLKBUFX2TS U1071 ( .A(n3833), .Y(n3825) );
  CLKBUFX2TS U1072 ( .A(n3751), .Y(n3746) );
  CLKBUFX2TS U1073 ( .A(n3750), .Y(n3748) );
  CLKBUFX2TS U1074 ( .A(n3750), .Y(n3747) );
  CLKBUFX2TS U1075 ( .A(n769), .Y(n3885) );
  CLKBUFX2TS U1076 ( .A(n3889), .Y(n3886) );
  CLKBUFX2TS U1077 ( .A(n3889), .Y(n3887) );
  CLKBUFX2TS U1078 ( .A(n3932), .Y(n3926) );
  CLKBUFX2TS U1079 ( .A(n3932), .Y(n3927) );
  CLKBUFX2TS U1080 ( .A(n3931), .Y(n3928) );
  CLKBUFX2TS U1081 ( .A(n224), .Y(n3833) );
  CLKBUFX2TS U1082 ( .A(n224), .Y(n3834) );
  CLKBUFX2TS U1083 ( .A(n3931), .Y(n3929) );
  CLKBUFX2TS U1084 ( .A(n3779), .Y(n3774) );
  CLKBUFX2TS U1085 ( .A(n3778), .Y(n3775) );
  CLKBUFX2TS U1086 ( .A(n3778), .Y(n3776) );
  CLKBUFX2TS U1087 ( .A(n3508), .Y(n3495) );
  CLKBUFX2TS U1088 ( .A(n3508), .Y(n3496) );
  CLKBUFX2TS U1089 ( .A(n3506), .Y(n3500) );
  CLKBUFX2TS U1090 ( .A(n3506), .Y(n3499) );
  CLKBUFX2TS U1091 ( .A(n3507), .Y(n3498) );
  CLKBUFX2TS U1092 ( .A(n3507), .Y(n3497) );
  CLKBUFX2TS U1093 ( .A(n3592), .Y(n3578) );
  CLKBUFX2TS U1094 ( .A(n2366), .Y(n1244) );
  CLKBUFX2TS U1095 ( .A(n3888), .Y(n3877) );
  CLKBUFX2TS U1096 ( .A(n3889), .Y(n3888) );
  CLKBUFX2TS U1097 ( .A(n3777), .Y(n3766) );
  CLKBUFX2TS U1098 ( .A(n3778), .Y(n3777) );
  CLKBUFX2TS U1099 ( .A(n3592), .Y(n3579) );
  CLKBUFX2TS U1100 ( .A(n2366), .Y(n1660) );
  CLKBUFX2TS U1101 ( .A(n3761), .Y(n3758) );
  CLKBUFX2TS U1102 ( .A(n3763), .Y(n3757) );
  CLKBUFX2TS U1103 ( .A(n3764), .Y(n3756) );
  CLKBUFX2TS U1104 ( .A(n3762), .Y(n3755) );
  CLKBUFX2TS U1105 ( .A(n3762), .Y(n3754) );
  CLKBUFX2TS U1106 ( .A(n3762), .Y(n3753) );
  CLKBUFX2TS U1107 ( .A(n2155), .Y(n1823) );
  CLKBUFX2TS U1108 ( .A(n2155), .Y(n1806) );
  CLKBUFX2TS U1109 ( .A(n2359), .Y(n1803) );
  CLKBUFX2TS U1110 ( .A(n2033), .Y(n1916) );
  CLKBUFX2TS U1111 ( .A(n2057), .Y(n1891) );
  CLKBUFX2TS U1112 ( .A(n2057), .Y(n1845) );
  CLKBUFX2TS U1113 ( .A(n2359), .Y(n1797) );
  CLKBUFX2TS U1114 ( .A(n3227), .Y(n3213) );
  CLKBUFX2TS U1115 ( .A(n3557), .Y(n3543) );
  CLKBUFX2TS U1116 ( .A(n3227), .Y(n3214) );
  CLKBUFX2TS U1117 ( .A(n3223), .Y(n3221) );
  CLKBUFX2TS U1118 ( .A(n3224), .Y(n3220) );
  CLKBUFX2TS U1119 ( .A(n3225), .Y(n3218) );
  CLKBUFX2TS U1120 ( .A(n3225), .Y(n3217) );
  CLKBUFX2TS U1121 ( .A(n3224), .Y(n3219) );
  CLKBUFX2TS U1122 ( .A(n3226), .Y(n3216) );
  CLKBUFX2TS U1123 ( .A(n3226), .Y(n3215) );
  CLKBUFX2TS U1124 ( .A(n3552), .Y(n3549) );
  CLKBUFX2TS U1125 ( .A(n3553), .Y(n3548) );
  CLKBUFX2TS U1126 ( .A(n3553), .Y(n3547) );
  CLKBUFX2TS U1127 ( .A(n3554), .Y(n3546) );
  CLKBUFX2TS U1128 ( .A(n3554), .Y(n3545) );
  CLKBUFX2TS U1129 ( .A(n3556), .Y(n3544) );
  CLKBUFX2TS U1130 ( .A(n3788), .Y(n3786) );
  CLKBUFX2TS U1131 ( .A(n3789), .Y(n3784) );
  CLKBUFX2TS U1132 ( .A(n3789), .Y(n3785) );
  CLKBUFX2TS U1133 ( .A(n3790), .Y(n3783) );
  CLKBUFX2TS U1134 ( .A(n3792), .Y(n3780) );
  CLKBUFX2TS U1135 ( .A(n3790), .Y(n3782) );
  CLKBUFX2TS U1136 ( .A(n3791), .Y(n3781) );
  CLKBUFX2TS U1137 ( .A(n3475), .Y(n3461) );
  CLKBUFX2TS U1138 ( .A(n3475), .Y(n3462) );
  CLKBUFX2TS U1139 ( .A(n3358), .Y(n3344) );
  CLKBUFX2TS U1140 ( .A(n3358), .Y(n3345) );
  CLKBUFX2TS U1141 ( .A(n3749), .Y(n3739) );
  CLKBUFX2TS U1142 ( .A(n3750), .Y(n3749) );
  CLKBUFX2TS U1143 ( .A(n3357), .Y(n3346) );
  CLKBUFX2TS U1144 ( .A(n3874), .Y(n3865) );
  CLKBUFX2TS U1145 ( .A(n3874), .Y(n3866) );
  CLKBUFX2TS U1146 ( .A(n3873), .Y(n3867) );
  CLKBUFX2TS U1147 ( .A(n3873), .Y(n3868) );
  CLKBUFX2TS U1148 ( .A(n3872), .Y(n3869) );
  CLKBUFX2TS U1149 ( .A(n3875), .Y(n3870) );
  CLKBUFX2TS U1150 ( .A(n3872), .Y(n3871) );
  CLKBUFX2TS U1151 ( .A(n3470), .Y(n3467) );
  CLKBUFX2TS U1152 ( .A(n3473), .Y(n3465) );
  CLKBUFX2TS U1153 ( .A(n3473), .Y(n3466) );
  CLKBUFX2TS U1154 ( .A(n3474), .Y(n3464) );
  CLKBUFX2TS U1155 ( .A(n3356), .Y(n3349) );
  CLKBUFX2TS U1156 ( .A(n3356), .Y(n3348) );
  CLKBUFX2TS U1157 ( .A(n3354), .Y(n3351) );
  CLKBUFX2TS U1158 ( .A(n3360), .Y(n3350) );
  CLKBUFX2TS U1159 ( .A(n3357), .Y(n3347) );
  CLKBUFX2TS U1160 ( .A(n3470), .Y(n3468) );
  CLKBUFX2TS U1161 ( .A(n3354), .Y(n3352) );
  CLKBUFX2TS U1162 ( .A(n3525), .Y(n3512) );
  CLKBUFX2TS U1163 ( .A(n3761), .Y(n3759) );
  CLKBUFX2TS U1164 ( .A(n3525), .Y(n3513) );
  CLKBUFX2TS U1165 ( .A(n3805), .Y(n3796) );
  CLKBUFX2TS U1166 ( .A(n3223), .Y(n3222) );
  CLKBUFX2TS U1167 ( .A(n3808), .Y(n3802) );
  CLKBUFX2TS U1168 ( .A(n3806), .Y(n3801) );
  CLKBUFX2TS U1169 ( .A(n3804), .Y(n3799) );
  CLKBUFX2TS U1170 ( .A(n3804), .Y(n3798) );
  CLKBUFX2TS U1171 ( .A(n3805), .Y(n3797) );
  CLKBUFX2TS U1172 ( .A(n3552), .Y(n3550) );
  CLKBUFX2TS U1173 ( .A(n3589), .Y(n3580) );
  CLKBUFX2TS U1174 ( .A(n3589), .Y(n3581) );
  CLKBUFX2TS U1175 ( .A(n3588), .Y(n3582) );
  CLKBUFX2TS U1176 ( .A(n3588), .Y(n3583) );
  CLKBUFX2TS U1177 ( .A(n3587), .Y(n3584) );
  CLKBUFX2TS U1178 ( .A(n3587), .Y(n3585) );
  CLKBUFX2TS U1179 ( .A(n3527), .Y(n3521) );
  CLKBUFX2TS U1180 ( .A(n3523), .Y(n3520) );
  CLKBUFX2TS U1181 ( .A(n3522), .Y(n3519) );
  CLKBUFX2TS U1182 ( .A(n3522), .Y(n3518) );
  CLKBUFX2TS U1183 ( .A(n3523), .Y(n3516) );
  CLKBUFX2TS U1184 ( .A(n3523), .Y(n3517) );
  CLKBUFX2TS U1185 ( .A(n3524), .Y(n3515) );
  CLKBUFX2TS U1186 ( .A(n3524), .Y(n3514) );
  CLKBUFX2TS U1187 ( .A(n3930), .Y(n3919) );
  CLKBUFX2TS U1188 ( .A(n3931), .Y(n3930) );
  CLKBUFX2TS U1189 ( .A(n3835), .Y(n3823) );
  CLKBUFX2TS U1190 ( .A(n775), .Y(n3835) );
  CLKBUFX2TS U1191 ( .A(n3918), .Y(n3908) );
  CLKBUFX2TS U1192 ( .A(n3916), .Y(n3909) );
  CLKBUFX2TS U1193 ( .A(n3917), .Y(n3905) );
  CLKBUFX2TS U1194 ( .A(n3917), .Y(n3906) );
  CLKBUFX2TS U1195 ( .A(n3916), .Y(n3907) );
  CLKBUFX2TS U1196 ( .A(n3915), .Y(n3910) );
  CLKBUFX2TS U1197 ( .A(n3915), .Y(n3911) );
  CLKBUFX2TS U1198 ( .A(n3914), .Y(n3912) );
  CLKBUFX2TS U1199 ( .A(n3914), .Y(n3913) );
  CLKBUFX2TS U1200 ( .A(n3788), .Y(n3787) );
  INVX2TS U1201 ( .A(n4504), .Y(n4502) );
  CLKBUFX2TS U1202 ( .A(n3847), .Y(n3836) );
  CLKBUFX2TS U1203 ( .A(n3847), .Y(n3837) );
  CLKBUFX2TS U1204 ( .A(n3844), .Y(n3843) );
  CLKBUFX2TS U1205 ( .A(n3846), .Y(n3838) );
  CLKBUFX2TS U1206 ( .A(n3845), .Y(n3840) );
  CLKBUFX2TS U1207 ( .A(n3846), .Y(n3839) );
  CLKBUFX2TS U1208 ( .A(n3844), .Y(n3842) );
  CLKBUFX2TS U1209 ( .A(n3845), .Y(n3841) );
  INVX2TS U1210 ( .A(n4504), .Y(n4503) );
  CLKBUFX2TS U1211 ( .A(n3429), .Y(n3424) );
  CLKBUFX2TS U1212 ( .A(n3429), .Y(n3425) );
  CLKBUFX2TS U1213 ( .A(n3429), .Y(n3426) );
  CLKBUFX2TS U1214 ( .A(n3558), .Y(n3557) );
  CLKBUFX2TS U1215 ( .A(n3558), .Y(n3555) );
  CLKBUFX2TS U1216 ( .A(n3558), .Y(n3556) );
  CLKBUFX2TS U1217 ( .A(n3876), .Y(n3874) );
  CLKBUFX2TS U1218 ( .A(n3876), .Y(n3873) );
  CLKBUFX2TS U1219 ( .A(n771), .Y(n3872) );
  CLKBUFX2TS U1220 ( .A(n3477), .Y(n3470) );
  CLKBUFX2TS U1221 ( .A(n3477), .Y(n3471) );
  CLKBUFX2TS U1222 ( .A(n3807), .Y(n3804) );
  CLKBUFX2TS U1223 ( .A(n3477), .Y(n3472) );
  CLKBUFX2TS U1224 ( .A(n3808), .Y(n3803) );
  CLKBUFX2TS U1225 ( .A(n3476), .Y(n3473) );
  CLKBUFX2TS U1226 ( .A(n3807), .Y(n3805) );
  CLKBUFX2TS U1227 ( .A(n3476), .Y(n3474) );
  CLKBUFX2TS U1228 ( .A(n3526), .Y(n3525) );
  CLKBUFX2TS U1229 ( .A(n3593), .Y(n3591) );
  CLKBUFX2TS U1230 ( .A(n3510), .Y(n3503) );
  CLKBUFX2TS U1231 ( .A(n3594), .Y(n3589) );
  CLKBUFX2TS U1232 ( .A(n3594), .Y(n3588) );
  CLKBUFX2TS U1233 ( .A(n3594), .Y(n3587) );
  CLKBUFX2TS U1234 ( .A(n3764), .Y(n3762) );
  CLKBUFX2TS U1235 ( .A(n3765), .Y(n3761) );
  CLKBUFX2TS U1236 ( .A(n3593), .Y(n3592) );
  CLKBUFX2TS U1237 ( .A(n3765), .Y(n3760) );
  CLKBUFX2TS U1238 ( .A(n3228), .Y(n3225) );
  CLKBUFX2TS U1239 ( .A(n3229), .Y(n3224) );
  CLKBUFX2TS U1240 ( .A(n3228), .Y(n3226) );
  CLKBUFX2TS U1241 ( .A(n3228), .Y(n3227) );
  CLKBUFX2TS U1242 ( .A(n2372), .Y(n2155) );
  CLKBUFX2TS U1243 ( .A(n3359), .Y(n3356) );
  CLKBUFX2TS U1244 ( .A(n2380), .Y(n2057) );
  CLKBUFX2TS U1245 ( .A(n2372), .Y(n2359) );
  CLKBUFX2TS U1246 ( .A(n3360), .Y(n3355) );
  CLKBUFX2TS U1247 ( .A(n3359), .Y(n3357) );
  CLKBUFX2TS U1248 ( .A(n2372), .Y(n2366) );
  CLKBUFX2TS U1249 ( .A(n3360), .Y(n3354) );
  CLKBUFX2TS U1250 ( .A(n3509), .Y(n3508) );
  CLKBUFX2TS U1251 ( .A(n3510), .Y(n3504) );
  CLKBUFX2TS U1252 ( .A(n3527), .Y(n3522) );
  CLKBUFX2TS U1253 ( .A(n3509), .Y(n3506) );
  CLKBUFX2TS U1254 ( .A(n3510), .Y(n3505) );
  CLKBUFX2TS U1255 ( .A(n3527), .Y(n3523) );
  CLKBUFX2TS U1256 ( .A(n3526), .Y(n3524) );
  CLKBUFX2TS U1257 ( .A(n3509), .Y(n3507) );
  CLKBUFX2TS U1258 ( .A(n3794), .Y(n3788) );
  CLKBUFX2TS U1259 ( .A(n3794), .Y(n3789) );
  CLKBUFX2TS U1260 ( .A(n3794), .Y(n3790) );
  CLKBUFX2TS U1261 ( .A(n3793), .Y(n3791) );
  CLKBUFX2TS U1262 ( .A(n3476), .Y(n3475) );
  CLKBUFX2TS U1263 ( .A(n3359), .Y(n3358) );
  CLKBUFX2TS U1264 ( .A(n3918), .Y(n3917) );
  CLKBUFX2TS U1265 ( .A(n767), .Y(n3916) );
  CLKBUFX2TS U1266 ( .A(n3918), .Y(n3915) );
  CLKBUFX2TS U1267 ( .A(n3918), .Y(n3914) );
  CLKBUFX2TS U1268 ( .A(n3559), .Y(n3553) );
  CLKBUFX2TS U1269 ( .A(n3559), .Y(n3554) );
  CLKBUFX2TS U1270 ( .A(n209), .Y(n3779) );
  CLKBUFX2TS U1271 ( .A(n209), .Y(n3778) );
  CLKBUFX2TS U1272 ( .A(n784), .Y(n3750) );
  CLKBUFX2TS U1273 ( .A(n766), .Y(n3932) );
  CLKBUFX2TS U1274 ( .A(n766), .Y(n3931) );
  CLKBUFX2TS U1275 ( .A(n769), .Y(n3889) );
  CLKBUFX2TS U1276 ( .A(n3114), .Y(n3026) );
  CLKBUFX2TS U1277 ( .A(n3410), .Y(n3396) );
  CLKBUFX2TS U1278 ( .A(n3114), .Y(n3027) );
  CLKBUFX2TS U1279 ( .A(n3410), .Y(n3397) );
  CLKBUFX2TS U1280 ( .A(n3087), .Y(n3082) );
  CLKBUFX2TS U1281 ( .A(n3100), .Y(n3069) );
  CLKBUFX2TS U1282 ( .A(n3100), .Y(n3060) );
  CLKBUFX2TS U1283 ( .A(n3103), .Y(n3049) );
  CLKBUFX2TS U1284 ( .A(n3112), .Y(n3037) );
  CLKBUFX2TS U1285 ( .A(n3112), .Y(n3028) );
  CLKBUFX2TS U1286 ( .A(n3103), .Y(n3044) );
  CLKBUFX2TS U1287 ( .A(n3654), .Y(n3649) );
  CLKBUFX2TS U1288 ( .A(n3654), .Y(n3648) );
  CLKBUFX2TS U1289 ( .A(n3655), .Y(n3647) );
  CLKBUFX2TS U1290 ( .A(n3655), .Y(n3646) );
  CLKBUFX2TS U1291 ( .A(n3656), .Y(n3645) );
  CLKBUFX2TS U1292 ( .A(n3656), .Y(n3644) );
  CLKBUFX2TS U1293 ( .A(n3657), .Y(n3643) );
  CLKBUFX2TS U1294 ( .A(n3653), .Y(n3650) );
  CLKBUFX2TS U1295 ( .A(n3407), .Y(n3403) );
  CLKBUFX2TS U1296 ( .A(n3407), .Y(n3402) );
  CLKBUFX2TS U1297 ( .A(n3406), .Y(n3404) );
  CLKBUFX2TS U1298 ( .A(n3408), .Y(n3401) );
  CLKBUFX2TS U1299 ( .A(n3408), .Y(n3400) );
  CLKBUFX2TS U1300 ( .A(n3409), .Y(n3398) );
  CLKBUFX2TS U1301 ( .A(n3409), .Y(n3399) );
  CLKBUFX2TS U1302 ( .A(n3444), .Y(n3430) );
  CLKBUFX2TS U1303 ( .A(n3260), .Y(n3249) );
  CLKBUFX2TS U1304 ( .A(n3259), .Y(n3251) );
  CLKBUFX2TS U1305 ( .A(n3257), .Y(n3255) );
  CLKBUFX2TS U1306 ( .A(n3258), .Y(n3253) );
  CLKBUFX2TS U1307 ( .A(n3258), .Y(n3254) );
  CLKBUFX2TS U1308 ( .A(n3259), .Y(n3252) );
  CLKBUFX2TS U1309 ( .A(n3260), .Y(n3250) );
  CLKBUFX2TS U1310 ( .A(n3261), .Y(n3248) );
  CLKBUFX2TS U1311 ( .A(n3441), .Y(n3437) );
  CLKBUFX2TS U1312 ( .A(n3442), .Y(n3436) );
  CLKBUFX2TS U1313 ( .A(n3442), .Y(n3435) );
  CLKBUFX2TS U1314 ( .A(n3443), .Y(n3434) );
  CLKBUFX2TS U1315 ( .A(n3443), .Y(n3433) );
  CLKBUFX2TS U1316 ( .A(n3445), .Y(n3432) );
  CLKBUFX2TS U1317 ( .A(n3445), .Y(n3431) );
  CLKBUFX2TS U1318 ( .A(n3763), .Y(n3752) );
  CLKBUFX2TS U1319 ( .A(n3764), .Y(n3763) );
  INVX2TS U1320 ( .A(n3637), .Y(n3636) );
  INVX2TS U1321 ( .A(n3639), .Y(n3634) );
  INVX2TS U1322 ( .A(n3638), .Y(n3635) );
  CLKBUFX2TS U1323 ( .A(n3821), .Y(n3810) );
  CLKBUFX2TS U1324 ( .A(n3821), .Y(n3809) );
  CLKBUFX2TS U1325 ( .A(n3819), .Y(n3814) );
  CLKBUFX2TS U1326 ( .A(n3818), .Y(n3816) );
  CLKBUFX2TS U1327 ( .A(n3820), .Y(n3812) );
  CLKBUFX2TS U1328 ( .A(n206), .Y(n3817) );
  CLKBUFX2TS U1329 ( .A(n3818), .Y(n3815) );
  CLKBUFX2TS U1330 ( .A(n3819), .Y(n3813) );
  CLKBUFX2TS U1331 ( .A(n3820), .Y(n3811) );
  CLKBUFX2TS U1332 ( .A(n3902), .Y(n3890) );
  CLKBUFX2TS U1333 ( .A(n3705), .Y(n3691) );
  CLKBUFX2TS U1334 ( .A(n3653), .Y(n3651) );
  CLKBUFX2TS U1335 ( .A(n3707), .Y(n3697) );
  CLKBUFX2TS U1336 ( .A(n3703), .Y(n3696) );
  CLKBUFX2TS U1337 ( .A(n3703), .Y(n3695) );
  CLKBUFX2TS U1338 ( .A(n3704), .Y(n3694) );
  CLKBUFX2TS U1339 ( .A(n3704), .Y(n3693) );
  CLKBUFX2TS U1340 ( .A(n3705), .Y(n3692) );
  CLKBUFX2TS U1341 ( .A(n3701), .Y(n3698) );
  CLKBUFX2TS U1342 ( .A(n3899), .Y(n3895) );
  CLKBUFX2TS U1343 ( .A(n3899), .Y(n3894) );
  CLKBUFX2TS U1344 ( .A(n3900), .Y(n3893) );
  CLKBUFX2TS U1345 ( .A(n3898), .Y(n3896) );
  CLKBUFX2TS U1346 ( .A(n3902), .Y(n3891) );
  CLKBUFX2TS U1347 ( .A(n3900), .Y(n3892) );
  CLKBUFX2TS U1348 ( .A(n3023), .Y(n2979) );
  CLKBUFX2TS U1349 ( .A(n3023), .Y(n2985) );
  CLKBUFX2TS U1350 ( .A(n3022), .Y(n2986) );
  CLKBUFX2TS U1351 ( .A(n3195), .Y(n3138) );
  CLKBUFX2TS U1352 ( .A(n3674), .Y(n3661) );
  CLKBUFX2TS U1353 ( .A(n3674), .Y(n3660) );
  CLKBUFX2TS U1354 ( .A(n3019), .Y(n3014) );
  CLKBUFX2TS U1355 ( .A(n3021), .Y(n3004) );
  CLKBUFX2TS U1356 ( .A(n3018), .Y(n3016) );
  CLKBUFX2TS U1357 ( .A(n3018), .Y(n3015) );
  CLKBUFX2TS U1358 ( .A(n3021), .Y(n2996) );
  CLKBUFX2TS U1359 ( .A(n3022), .Y(n2992) );
  CLKBUFX2TS U1360 ( .A(n3441), .Y(n3438) );
  CLKBUFX2TS U1361 ( .A(n3257), .Y(n3256) );
  CLKBUFX2TS U1362 ( .A(n3673), .Y(n3662) );
  CLKBUFX2TS U1363 ( .A(n3358), .Y(n3353) );
  CLKBUFX2TS U1364 ( .A(n3875), .Y(n3864) );
  CLKBUFX2TS U1365 ( .A(n3876), .Y(n3875) );
  CLKBUFX2TS U1366 ( .A(n3593), .Y(n3586) );
  CLKBUFX2TS U1367 ( .A(n3701), .Y(n3699) );
  CLKBUFX2TS U1368 ( .A(n3184), .Y(n3172) );
  CLKBUFX2TS U1369 ( .A(n3184), .Y(n3161) );
  CLKBUFX2TS U1370 ( .A(n3193), .Y(n3157) );
  CLKBUFX2TS U1371 ( .A(n3193), .Y(n3148) );
  CLKBUFX2TS U1372 ( .A(n3194), .Y(n3143) );
  CLKBUFX2TS U1373 ( .A(n3194), .Y(n3147) );
  CLKBUFX2TS U1374 ( .A(n3198), .Y(n3140) );
  CLKBUFX2TS U1375 ( .A(n3670), .Y(n3669) );
  CLKBUFX2TS U1376 ( .A(n3670), .Y(n3668) );
  CLKBUFX2TS U1377 ( .A(n3671), .Y(n3667) );
  CLKBUFX2TS U1378 ( .A(n3671), .Y(n3666) );
  CLKBUFX2TS U1379 ( .A(n3672), .Y(n3665) );
  CLKBUFX2TS U1380 ( .A(n3672), .Y(n3664) );
  CLKBUFX2TS U1381 ( .A(n3673), .Y(n3663) );
  CLKBUFX2TS U1382 ( .A(n3198), .Y(n3139) );
  CLKBUFX2TS U1383 ( .A(n3860), .Y(n3856) );
  CLKBUFX2TS U1384 ( .A(n3862), .Y(n3850) );
  CLKBUFX2TS U1385 ( .A(n3859), .Y(n3857) );
  CLKBUFX2TS U1386 ( .A(n3860), .Y(n3855) );
  CLKBUFX2TS U1387 ( .A(n3861), .Y(n3854) );
  CLKBUFX2TS U1388 ( .A(n3861), .Y(n3853) );
  CLKBUFX2TS U1389 ( .A(n3862), .Y(n3852) );
  CLKBUFX2TS U1390 ( .A(n3862), .Y(n3851) );
  CLKBUFX2TS U1391 ( .A(n3806), .Y(n3795) );
  CLKBUFX2TS U1392 ( .A(n3807), .Y(n3806) );
  CLKBUFX2TS U1393 ( .A(n3898), .Y(n3897) );
  CLKBUFX2TS U1394 ( .A(n3859), .Y(n3858) );
  INVX2TS U1395 ( .A(n3427), .Y(n3414) );
  INVX2TS U1396 ( .A(n3427), .Y(n3415) );
  INVX2TS U1397 ( .A(n3427), .Y(n3413) );
  INVX2TS U1398 ( .A(n3428), .Y(n3416) );
  INVX2TS U1399 ( .A(n3428), .Y(n3417) );
  INVX2TS U1400 ( .A(n3427), .Y(n3418) );
  INVX2TS U1401 ( .A(n3428), .Y(n3419) );
  INVX2TS U1402 ( .A(n3428), .Y(n3420) );
  INVX2TS U1403 ( .A(n3575), .Y(n3570) );
  INVX2TS U1404 ( .A(n3576), .Y(n3569) );
  INVX2TS U1405 ( .A(n3577), .Y(n3568) );
  INVX2TS U1406 ( .A(n3575), .Y(n3562) );
  INVX2TS U1407 ( .A(n3575), .Y(n3563) );
  INVX2TS U1408 ( .A(n3574), .Y(n3567) );
  INVX2TS U1409 ( .A(n3574), .Y(n3566) );
  INVX2TS U1410 ( .A(n3574), .Y(n3565) );
  INVX2TS U1411 ( .A(n3575), .Y(n3564) );
  INVX2TS U1412 ( .A(n529), .Y(n1126) );
  INVX2TS U1413 ( .A(n1129), .Y(n1125) );
  INVX2TS U1414 ( .A(n1133), .Y(n1124) );
  INVX2TS U1415 ( .A(n1153), .Y(n1123) );
  INVX2TS U1416 ( .A(n3576), .Y(n3560) );
  INVX2TS U1417 ( .A(n3576), .Y(n3561) );
  CLKBUFX2TS U1418 ( .A(reset), .Y(n4504) );
  CLKBUFX2TS U1419 ( .A(n3848), .Y(n3847) );
  CLKBUFX2TS U1420 ( .A(n3849), .Y(n3846) );
  CLKBUFX2TS U1421 ( .A(n3849), .Y(n3844) );
  CLKBUFX2TS U1422 ( .A(n3849), .Y(n3845) );
  CLKBUFX2TS U1423 ( .A(n3605), .Y(n3596) );
  CLKBUFX2TS U1424 ( .A(n3605), .Y(n3597) );
  CLKBUFX2TS U1425 ( .A(n3458), .Y(n3447) );
  CLKBUFX2TS U1426 ( .A(n3455), .Y(n3451) );
  CLKBUFX2TS U1427 ( .A(n3454), .Y(n3452) );
  CLKBUFX2TS U1428 ( .A(n3456), .Y(n3448) );
  CLKBUFX2TS U1429 ( .A(n3455), .Y(n3450) );
  CLKBUFX2TS U1430 ( .A(n3456), .Y(n3449) );
  CLKBUFX2TS U1431 ( .A(n3454), .Y(n3453) );
  CLKBUFX2TS U1432 ( .A(n3603), .Y(n3601) );
  CLKBUFX2TS U1433 ( .A(n3603), .Y(n3600) );
  CLKBUFX2TS U1434 ( .A(n3604), .Y(n3599) );
  CLKBUFX2TS U1435 ( .A(n3604), .Y(n3598) );
  CLKBUFX2TS U1436 ( .A(n3687), .Y(n3678) );
  CLKBUFX2TS U1437 ( .A(n3687), .Y(n3679) );
  CLKBUFX2TS U1438 ( .A(n3686), .Y(n3680) );
  CLKBUFX2TS U1439 ( .A(n3686), .Y(n3681) );
  CLKBUFX2TS U1440 ( .A(n3683), .Y(n3682) );
  CLKBUFX2TS U1441 ( .A(n3540), .Y(n3529) );
  CLKBUFX2TS U1442 ( .A(n3538), .Y(n3530) );
  CLKBUFX2TS U1443 ( .A(n3538), .Y(n3531) );
  CLKBUFX2TS U1444 ( .A(n3537), .Y(n3532) );
  CLKBUFX2TS U1445 ( .A(n3537), .Y(n3533) );
  CLKBUFX2TS U1446 ( .A(n3536), .Y(n3535) );
  CLKBUFX2TS U1447 ( .A(n3536), .Y(n3534) );
  CLKBUFX2TS U1448 ( .A(n529), .Y(n1128) );
  CLKBUFX2TS U1449 ( .A(n3642), .Y(n3639) );
  CLKBUFX2TS U1450 ( .A(n3642), .Y(n3638) );
  CLKBUFX2TS U1451 ( .A(n3642), .Y(n3637) );
  CLKBUFX2TS U1452 ( .A(n3494), .Y(n3491) );
  CLKBUFX2TS U1453 ( .A(n3494), .Y(n3489) );
  CLKBUFX2TS U1454 ( .A(n3494), .Y(n3490) );
  CLKBUFX2TS U1455 ( .A(n3377), .Y(n3372) );
  CLKBUFX2TS U1456 ( .A(n3377), .Y(n3373) );
  CLKBUFX2TS U1457 ( .A(n3377), .Y(n3374) );
  CLKBUFX2TS U1458 ( .A(n229), .Y(n3808) );
  CLKBUFX2TS U1459 ( .A(n229), .Y(n3807) );
  CLKBUFX2TS U1460 ( .A(n1183), .Y(n3558) );
  CLKBUFX2TS U1461 ( .A(n3706), .Y(n3703) );
  CLKBUFX2TS U1462 ( .A(n3706), .Y(n3704) );
  CLKBUFX2TS U1463 ( .A(n3706), .Y(n3705) );
  CLKBUFX2TS U1464 ( .A(n3819), .Y(n3818) );
  CLKBUFX2TS U1465 ( .A(n3196), .Y(n3195) );
  CLKBUFX2TS U1466 ( .A(n3136), .Y(n3100) );
  CLKBUFX2TS U1467 ( .A(n3197), .Y(n3184) );
  CLKBUFX2TS U1468 ( .A(n3197), .Y(n3193) );
  CLKBUFX2TS U1469 ( .A(n3121), .Y(n3112) );
  CLKBUFX2TS U1470 ( .A(n3136), .Y(n3103) );
  CLKBUFX2TS U1471 ( .A(n3197), .Y(n3194) );
  CLKBUFX2TS U1472 ( .A(n3659), .Y(n3654) );
  CLKBUFX2TS U1473 ( .A(n3676), .Y(n3670) );
  CLKBUFX2TS U1474 ( .A(n3659), .Y(n3655) );
  CLKBUFX2TS U1475 ( .A(n3658), .Y(n3656) );
  CLKBUFX2TS U1476 ( .A(n3676), .Y(n3671) );
  CLKBUFX2TS U1477 ( .A(n3658), .Y(n3657) );
  CLKBUFX2TS U1478 ( .A(n3675), .Y(n3672) );
  CLKBUFX2TS U1479 ( .A(n3675), .Y(n3673) );
  CLKBUFX2TS U1480 ( .A(n3121), .Y(n3114) );
  CLKBUFX2TS U1481 ( .A(n3659), .Y(n3653) );
  CLKBUFX2TS U1482 ( .A(n3136), .Y(n3087) );
  CLKBUFX2TS U1483 ( .A(n3675), .Y(n3674) );
  CLKBUFX2TS U1484 ( .A(n3904), .Y(n3899) );
  CLKBUFX2TS U1485 ( .A(n3412), .Y(n3407) );
  CLKBUFX2TS U1486 ( .A(n3411), .Y(n3410) );
  CLKBUFX2TS U1487 ( .A(n3904), .Y(n3898) );
  CLKBUFX2TS U1488 ( .A(n3863), .Y(n3859) );
  CLKBUFX2TS U1489 ( .A(n3863), .Y(n3860) );
  CLKBUFX2TS U1490 ( .A(n3412), .Y(n3408) );
  CLKBUFX2TS U1491 ( .A(n3863), .Y(n3861) );
  CLKBUFX2TS U1492 ( .A(n773), .Y(n3862) );
  CLKBUFX2TS U1493 ( .A(n3025), .Y(n3018) );
  CLKBUFX2TS U1494 ( .A(n3025), .Y(n3019) );
  CLKBUFX2TS U1495 ( .A(n3024), .Y(n3021) );
  CLKBUFX2TS U1496 ( .A(n3024), .Y(n3022) );
  CLKBUFX2TS U1497 ( .A(n3264), .Y(n3258) );
  CLKBUFX2TS U1498 ( .A(n3264), .Y(n3259) );
  CLKBUFX2TS U1499 ( .A(n3263), .Y(n3260) );
  CLKBUFX2TS U1500 ( .A(n3263), .Y(n3261) );
  CLKBUFX2TS U1501 ( .A(n3411), .Y(n3409) );
  CLKBUFX2TS U1502 ( .A(n3025), .Y(n3017) );
  CLKBUFX2TS U1503 ( .A(n3903), .Y(n3901) );
  CLKBUFX2TS U1504 ( .A(n3903), .Y(n3902) );
  CLKBUFX2TS U1505 ( .A(n3904), .Y(n3900) );
  CLKBUFX2TS U1506 ( .A(n3263), .Y(n3262) );
  CLKBUFX2TS U1507 ( .A(n3446), .Y(n3442) );
  CLKBUFX2TS U1508 ( .A(n3446), .Y(n3443) );
  CLKBUFX2TS U1509 ( .A(n3445), .Y(n3444) );
  CLKBUFX2TS U1510 ( .A(n3446), .Y(n3441) );
  CLKBUFX2TS U1511 ( .A(n3412), .Y(n3406) );
  CLKBUFX2TS U1512 ( .A(n3024), .Y(n3023) );
  CLKBUFX2TS U1513 ( .A(n3264), .Y(n3257) );
  CLKBUFX2TS U1514 ( .A(n3511), .Y(n3502) );
  CLKBUFX2TS U1515 ( .A(n1186), .Y(n3511) );
  CLKBUFX2TS U1516 ( .A(n3707), .Y(n3702) );
  CLKBUFX2TS U1517 ( .A(n3707), .Y(n3701) );
  CLKBUFX2TS U1518 ( .A(n3822), .Y(n3819) );
  CLKBUFX2TS U1519 ( .A(n3822), .Y(n3820) );
  CLKBUFX2TS U1520 ( .A(n1185), .Y(n3528) );
  CLKBUFX2TS U1521 ( .A(n1186), .Y(n3509) );
  CLKBUFX2TS U1522 ( .A(n1265), .Y(n2372) );
  CLKBUFX2TS U1523 ( .A(n1231), .Y(n3360) );
  CLKBUFX2TS U1524 ( .A(n1231), .Y(n3359) );
  CLKBUFX2TS U1525 ( .A(n767), .Y(n3918) );
  CLKBUFX2TS U1526 ( .A(n780), .Y(n3793) );
  CLKBUFX2TS U1527 ( .A(n780), .Y(n3794) );
  CLKBUFX2TS U1528 ( .A(n771), .Y(n3876) );
  CLKBUFX2TS U1529 ( .A(n1169), .Y(n3593) );
  CLKBUFX2TS U1530 ( .A(n1185), .Y(n3526) );
  CLKBUFX2TS U1531 ( .A(n1169), .Y(n3594) );
  CLKBUFX2TS U1532 ( .A(n1185), .Y(n3527) );
  CLKBUFX2TS U1533 ( .A(n218), .Y(n3764) );
  CLKBUFX2TS U1534 ( .A(n3624), .Y(n3609) );
  CLKBUFX2TS U1535 ( .A(n3624), .Y(n3610) );
  CLKBUFX2TS U1536 ( .A(n3623), .Y(n3611) );
  CLKBUFX2TS U1537 ( .A(n3623), .Y(n3612) );
  CLKBUFX2TS U1538 ( .A(n3622), .Y(n3613) );
  CLKBUFX2TS U1539 ( .A(n3622), .Y(n3614) );
  CLKBUFX2TS U1540 ( .A(n3393), .Y(n3379) );
  CLKBUFX2TS U1541 ( .A(n3393), .Y(n3380) );
  CLKBUFX2TS U1542 ( .A(n3389), .Y(n3387) );
  CLKBUFX2TS U1543 ( .A(n3390), .Y(n3386) );
  CLKBUFX2TS U1544 ( .A(n3390), .Y(n3385) );
  CLKBUFX2TS U1545 ( .A(n3391), .Y(n3384) );
  CLKBUFX2TS U1546 ( .A(n3391), .Y(n3383) );
  CLKBUFX2TS U1547 ( .A(n3392), .Y(n3381) );
  CLKBUFX2TS U1548 ( .A(n3392), .Y(n3382) );
  CLKBUFX2TS U1549 ( .A(n1183), .Y(n3559) );
  INVX2TS U1550 ( .A(n212), .Y(n769) );
  CLKBUFX2TS U1551 ( .A(n526), .Y(n3427) );
  CLKBUFX2TS U1552 ( .A(n526), .Y(n3428) );
  CLKBUFX2TS U1553 ( .A(n526), .Y(n3429) );
  CLKBUFX2TS U1554 ( .A(n3654), .Y(n3652) );
  CLKBUFX2TS U1555 ( .A(n3621), .Y(n3615) );
  CLKBUFX2TS U1556 ( .A(n3621), .Y(n3616) );
  CLKBUFX2TS U1557 ( .A(n3620), .Y(n3617) );
  CLKBUFX2TS U1558 ( .A(n3440), .Y(n3439) );
  CLKBUFX2TS U1559 ( .A(n3620), .Y(n3618) );
  CLKBUFX2TS U1560 ( .A(n3706), .Y(n3700) );
  CLKBUFX2TS U1561 ( .A(n3198), .Y(n3179) );
  INVX2TS U1562 ( .A(n3376), .Y(n3365) );
  INVX2TS U1563 ( .A(n3375), .Y(n3361) );
  INVX2TS U1564 ( .A(n3375), .Y(n3363) );
  INVX2TS U1565 ( .A(n3376), .Y(n3367) );
  INVX2TS U1566 ( .A(n3376), .Y(n3362) );
  INVX2TS U1567 ( .A(n3375), .Y(n3364) );
  INVX2TS U1568 ( .A(n3375), .Y(n3366) );
  INVX2TS U1569 ( .A(n3376), .Y(n3368) );
  CLKBUFX2TS U1570 ( .A(n3493), .Y(n3492) );
  INVX2TS U1571 ( .A(n3494), .Y(n3479) );
  INVX2TS U1572 ( .A(n3492), .Y(n3480) );
  INVX2TS U1573 ( .A(n3493), .Y(n3481) );
  INVX2TS U1574 ( .A(n3493), .Y(n3482) );
  INVX2TS U1575 ( .A(n3492), .Y(n3484) );
  INVX2TS U1576 ( .A(n3493), .Y(n3485) );
  INVX2TS U1577 ( .A(n3492), .Y(n3483) );
  CLKBUFX2TS U1578 ( .A(n1213), .Y(n1133) );
  CLKBUFX2TS U1579 ( .A(n1213), .Y(n1129) );
  CLKBUFX2TS U1580 ( .A(n1213), .Y(n1153) );
  INVX2TS U1581 ( .A(n1197), .Y(n1117) );
  CLKBUFX2TS U1582 ( .A(n1180), .Y(n1197) );
  INVX2TS U1583 ( .A(n1197), .Y(n1118) );
  CLKBUFX2TS U1584 ( .A(n3577), .Y(n3576) );
  INVX2TS U1585 ( .A(n530), .Y(n3572) );
  INVX2TS U1586 ( .A(n530), .Y(n3571) );
  INVX2TS U1587 ( .A(n3246), .Y(n3240) );
  INVX2TS U1588 ( .A(n3247), .Y(n3239) );
  INVX2TS U1589 ( .A(n3245), .Y(n3238) );
  INVX2TS U1590 ( .A(n3245), .Y(n3232) );
  INVX2TS U1591 ( .A(n3244), .Y(n3237) );
  INVX2TS U1592 ( .A(n3244), .Y(n3236) );
  INVX2TS U1593 ( .A(n3244), .Y(n3235) );
  INVX2TS U1594 ( .A(n3245), .Y(n3234) );
  INVX2TS U1595 ( .A(n3245), .Y(n3233) );
  INVX2TS U1596 ( .A(n3246), .Y(n3230) );
  INVX2TS U1597 ( .A(n3246), .Y(n3231) );
  INVX2TS U1598 ( .A(n1197), .Y(n1119) );
  INVX2TS U1599 ( .A(n1180), .Y(n1122) );
  CLKBUFX2TS U1600 ( .A(n1213), .Y(n1180) );
  INVX2TS U1601 ( .A(n1180), .Y(n1121) );
  INVX2TS U1602 ( .A(n1180), .Y(n1120) );
  CLKBUFX2TS U1603 ( .A(n3608), .Y(n3603) );
  CLKBUFX2TS U1604 ( .A(n3608), .Y(n3602) );
  CLKBUFX2TS U1605 ( .A(n3607), .Y(n3604) );
  CLKBUFX2TS U1606 ( .A(n3607), .Y(n3605) );
  CLKBUFX2TS U1607 ( .A(n3689), .Y(n3687) );
  CLKBUFX2TS U1608 ( .A(n3689), .Y(n3686) );
  CLKBUFX2TS U1609 ( .A(n3690), .Y(n3685) );
  CLKBUFX2TS U1610 ( .A(n3690), .Y(n3684) );
  CLKBUFX2TS U1611 ( .A(n3690), .Y(n3683) );
  CLKBUFX2TS U1612 ( .A(n3542), .Y(n3536) );
  CLKBUFX2TS U1613 ( .A(n3541), .Y(n3540) );
  CLKBUFX2TS U1614 ( .A(n3541), .Y(n3539) );
  CLKBUFX2TS U1615 ( .A(n3542), .Y(n3538) );
  CLKBUFX2TS U1616 ( .A(n3542), .Y(n3537) );
  CLKBUFX2TS U1617 ( .A(n3459), .Y(n3458) );
  CLKBUFX2TS U1618 ( .A(n3459), .Y(n3457) );
  CLKBUFX2TS U1619 ( .A(n3460), .Y(n3455) );
  CLKBUFX2TS U1620 ( .A(n3460), .Y(n3456) );
  CLKBUFX2TS U1621 ( .A(n3460), .Y(n3454) );
  CLKBUFX2TS U1622 ( .A(n774), .Y(n3848) );
  CLKBUFX2TS U1623 ( .A(n774), .Y(n3849) );
  CLKBUFX2TS U1624 ( .A(n2952), .Y(n2909) );
  CLKBUFX2TS U1625 ( .A(n3340), .Y(n3267) );
  CLKBUFX2TS U1626 ( .A(n2952), .Y(n2907) );
  CLKBUFX2TS U1627 ( .A(n3340), .Y(n3266) );
  CLKBUFX2TS U1628 ( .A(n3339), .Y(n3268) );
  CLKBUFX2TS U1629 ( .A(n3337), .Y(n3335) );
  CLKBUFX2TS U1630 ( .A(n2950), .Y(n2913) );
  CLKBUFX2TS U1631 ( .A(n2950), .Y(n2914) );
  CLKBUFX2TS U1632 ( .A(n2974), .Y(n2923) );
  CLKBUFX2TS U1633 ( .A(n2950), .Y(n2925) );
  CLKBUFX2TS U1634 ( .A(n3339), .Y(n3269) );
  INVX2TS U1635 ( .A(n1112), .Y(n1100) );
  INVX2TS U1636 ( .A(n1112), .Y(n1101) );
  INVX2TS U1637 ( .A(n1116), .Y(n1110) );
  INVX2TS U1638 ( .A(n1111), .Y(n1109) );
  INVX2TS U1639 ( .A(n1115), .Y(n1108) );
  INVX2TS U1640 ( .A(n1115), .Y(n1107) );
  INVX2TS U1641 ( .A(n1112), .Y(n1106) );
  INVX2TS U1642 ( .A(n1111), .Y(n1104) );
  INVX2TS U1643 ( .A(n1111), .Y(n1103) );
  INVX2TS U1644 ( .A(n1111), .Y(n1105) );
  INVX2TS U1645 ( .A(n1112), .Y(n1102) );
  CLKBUFX2TS U1646 ( .A(n3606), .Y(n3595) );
  CLKBUFX2TS U1647 ( .A(n3607), .Y(n3606) );
  CLKBUFX2TS U1648 ( .A(n3688), .Y(n3677) );
  CLKBUFX2TS U1649 ( .A(n3689), .Y(n3688) );
  CLKBUFX2TS U1650 ( .A(n1074), .Y(n1073) );
  CLKBUFX2TS U1651 ( .A(n1078), .Y(n1065) );
  CLKBUFX2TS U1652 ( .A(n1077), .Y(n1066) );
  CLKBUFX2TS U1653 ( .A(n1077), .Y(n1067) );
  CLKBUFX2TS U1654 ( .A(n1076), .Y(n1068) );
  CLKBUFX2TS U1655 ( .A(n1076), .Y(n1069) );
  CLKBUFX2TS U1656 ( .A(n1074), .Y(n1072) );
  CLKBUFX2TS U1657 ( .A(n1075), .Y(n1070) );
  CLKBUFX2TS U1658 ( .A(n1075), .Y(n1071) );
  CLKBUFX2TS U1659 ( .A(n3210), .Y(n3200) );
  CLKBUFX2TS U1660 ( .A(n3209), .Y(n3202) );
  CLKBUFX2TS U1661 ( .A(n3210), .Y(n3201) );
  CLKBUFX2TS U1662 ( .A(n3208), .Y(n3204) );
  CLKBUFX2TS U1663 ( .A(n3209), .Y(n3203) );
  CLKBUFX2TS U1664 ( .A(n1097), .Y(n1083) );
  CLKBUFX2TS U1665 ( .A(n1097), .Y(n1082) );
  CLKBUFX2TS U1666 ( .A(n3207), .Y(n3206) );
  CLKBUFX2TS U1667 ( .A(n3207), .Y(n3205) );
  CLKBUFX2TS U1668 ( .A(n1061), .Y(n1050) );
  CLKBUFX2TS U1669 ( .A(n1093), .Y(n1092) );
  CLKBUFX2TS U1670 ( .A(n1093), .Y(n1091) );
  CLKBUFX2TS U1671 ( .A(n1094), .Y(n1090) );
  CLKBUFX2TS U1672 ( .A(n1095), .Y(n1088) );
  CLKBUFX2TS U1673 ( .A(n1094), .Y(n1089) );
  CLKBUFX2TS U1674 ( .A(n1096), .Y(n1085) );
  CLKBUFX2TS U1675 ( .A(n1095), .Y(n1087) );
  CLKBUFX2TS U1676 ( .A(n1096), .Y(n1086) );
  CLKBUFX2TS U1677 ( .A(n3720), .Y(n3708) );
  CLKBUFX2TS U1678 ( .A(n3719), .Y(n3715) );
  CLKBUFX2TS U1679 ( .A(n3719), .Y(n3714) );
  CLKBUFX2TS U1680 ( .A(n3720), .Y(n3713) );
  CLKBUFX2TS U1681 ( .A(n3721), .Y(n3712) );
  CLKBUFX2TS U1682 ( .A(n3721), .Y(n3711) );
  CLKBUFX2TS U1683 ( .A(n3722), .Y(n3710) );
  CLKBUFX2TS U1684 ( .A(n3722), .Y(n3709) );
  CLKBUFX2TS U1685 ( .A(n1057), .Y(n1056) );
  CLKBUFX2TS U1686 ( .A(n1057), .Y(n1055) );
  CLKBUFX2TS U1687 ( .A(n1058), .Y(n1054) );
  CLKBUFX2TS U1688 ( .A(n1061), .Y(n1051) );
  CLKBUFX2TS U1689 ( .A(n1060), .Y(n1053) );
  CLKBUFX2TS U1690 ( .A(n1060), .Y(n1052) );
  INVX2TS U1691 ( .A(n1044), .Y(n1043) );
  INVX2TS U1692 ( .A(n1045), .Y(n1042) );
  INVX2TS U1693 ( .A(n1046), .Y(n1041) );
  CLKBUFX2TS U1694 ( .A(n1002), .Y(n989) );
  CLKBUFX2TS U1695 ( .A(n2163), .Y(n990) );
  CLKBUFX2TS U1696 ( .A(n1001), .Y(n991) );
  CLKBUFX2TS U1697 ( .A(n1001), .Y(n992) );
  CLKBUFX2TS U1698 ( .A(n1003), .Y(n993) );
  CLKBUFX2TS U1699 ( .A(n1000), .Y(n994) );
  CLKBUFX2TS U1700 ( .A(n999), .Y(n998) );
  CLKBUFX2TS U1701 ( .A(n1000), .Y(n995) );
  CLKBUFX2TS U1702 ( .A(n999), .Y(n997) );
  CLKBUFX2TS U1703 ( .A(n1144), .Y(n3725) );
  CLKBUFX2TS U1704 ( .A(n1144), .Y(n3726) );
  CLKBUFX2TS U1705 ( .A(n986), .Y(n968) );
  CLKBUFX2TS U1706 ( .A(n3736), .Y(n3727) );
  CLKBUFX2TS U1707 ( .A(n3736), .Y(n3728) );
  CLKBUFX2TS U1708 ( .A(n984), .Y(n971) );
  CLKBUFX2TS U1709 ( .A(n3736), .Y(n3729) );
  CLKBUFX2TS U1710 ( .A(n984), .Y(n973) );
  CLKBUFX2TS U1711 ( .A(n3736), .Y(n3730) );
  CLKBUFX2TS U1712 ( .A(n983), .Y(n974) );
  CLKBUFX2TS U1713 ( .A(n3734), .Y(n3733) );
  CLKBUFX2TS U1714 ( .A(n978), .Y(n977) );
  CLKBUFX2TS U1715 ( .A(n3735), .Y(n3731) );
  CLKBUFX2TS U1716 ( .A(n983), .Y(n975) );
  CLKBUFX2TS U1717 ( .A(n3735), .Y(n3732) );
  CLKBUFX2TS U1718 ( .A(n978), .Y(n976) );
  CLKBUFX2TS U1719 ( .A(n964), .Y(n785) );
  CLKBUFX2TS U1720 ( .A(n964), .Y(n786) );
  CLKBUFX2TS U1721 ( .A(n963), .Y(n787) );
  CLKBUFX2TS U1722 ( .A(n965), .Y(n899) );
  CLKBUFX2TS U1723 ( .A(n963), .Y(n900) );
  CLKBUFX2TS U1724 ( .A(n962), .Y(n935) );
  CLKBUFX2TS U1725 ( .A(n961), .Y(n959) );
  CLKBUFX2TS U1726 ( .A(n962), .Y(n937) );
  CLKBUFX2TS U1727 ( .A(n961), .Y(n938) );
  CLKBUFX2TS U1728 ( .A(n547), .Y(n535) );
  CLKBUFX2TS U1729 ( .A(n561), .Y(n549) );
  CLKBUFX2TS U1730 ( .A(n547), .Y(n536) );
  CLKBUFX2TS U1731 ( .A(n561), .Y(n550) );
  CLKBUFX2TS U1732 ( .A(n546), .Y(n537) );
  CLKBUFX2TS U1733 ( .A(n560), .Y(n551) );
  CLKBUFX2TS U1734 ( .A(n548), .Y(n538) );
  CLKBUFX2TS U1735 ( .A(n562), .Y(n552) );
  CLKBUFX2TS U1736 ( .A(n546), .Y(n539) );
  CLKBUFX2TS U1737 ( .A(n560), .Y(n553) );
  CLKBUFX2TS U1738 ( .A(n545), .Y(n540) );
  CLKBUFX2TS U1739 ( .A(n559), .Y(n554) );
  CLKBUFX2TS U1740 ( .A(n544), .Y(n543) );
  CLKBUFX2TS U1741 ( .A(n558), .Y(n557) );
  CLKBUFX2TS U1742 ( .A(n545), .Y(n541) );
  CLKBUFX2TS U1743 ( .A(n559), .Y(n555) );
  CLKBUFX2TS U1744 ( .A(n544), .Y(n542) );
  CLKBUFX2TS U1745 ( .A(n558), .Y(n556) );
  CLKBUFX2TS U1746 ( .A(n1030), .Y(n1019) );
  CLKBUFX2TS U1747 ( .A(n2160), .Y(n1020) );
  CLKBUFX2TS U1748 ( .A(n778), .Y(n755) );
  CLKBUFX2TS U1749 ( .A(n1030), .Y(n1021) );
  CLKBUFX2TS U1750 ( .A(n778), .Y(n756) );
  CLKBUFX2TS U1751 ( .A(n1030), .Y(n1022) );
  CLKBUFX2TS U1752 ( .A(n776), .Y(n763) );
  CLKBUFX2TS U1753 ( .A(n1028), .Y(n1023) );
  CLKBUFX2TS U1754 ( .A(n772), .Y(n770) );
  CLKBUFX2TS U1755 ( .A(n1027), .Y(n1026) );
  CLKBUFX2TS U1756 ( .A(n776), .Y(n765) );
  CLKBUFX2TS U1757 ( .A(n1028), .Y(n1024) );
  CLKBUFX2TS U1758 ( .A(n772), .Y(n768) );
  CLKBUFX2TS U1759 ( .A(n1027), .Y(n1025) );
  CLKBUFX2TS U1760 ( .A(n1015), .Y(n1004) );
  CLKBUFX2TS U1761 ( .A(n1013), .Y(n1005) );
  CLKBUFX2TS U1762 ( .A(n1013), .Y(n1006) );
  CLKBUFX2TS U1763 ( .A(n1012), .Y(n1007) );
  CLKBUFX2TS U1764 ( .A(n1011), .Y(n1010) );
  CLKBUFX2TS U1765 ( .A(n1012), .Y(n1008) );
  CLKBUFX2TS U1766 ( .A(n1011), .Y(n1009) );
  NOR2BX1TS U1767 ( .AN(n132), .B(n1827), .Y(n1186) );
  NOR2BX1TS U1768 ( .AN(n1846), .B(n1853), .Y(n1231) );
  NAND2X1TS U1769 ( .A(n942), .B(n1846), .Y(n1800) );
  AND3X2TS U1770 ( .A(n447), .B(n1827), .C(n132), .Y(n1185) );
  INVX2TS U1771 ( .A(n1827), .Y(n945) );
  AND2X2TS U1772 ( .A(n1821), .B(n130), .Y(n1169) );
  INVX2TS U1773 ( .A(n215), .Y(n771) );
  CLKBUFX2TS U1774 ( .A(n1149), .Y(n3706) );
  CLKBUFX2TS U1775 ( .A(n3622), .Y(n3624) );
  CLKBUFX2TS U1776 ( .A(n3621), .Y(n3623) );
  CLKBUFX2TS U1777 ( .A(n3625), .Y(n3622) );
  CLKBUFX2TS U1778 ( .A(n3625), .Y(n3620) );
  CLKBUFX2TS U1779 ( .A(n3625), .Y(n3621) );
  CLKBUFX2TS U1780 ( .A(n3395), .Y(n3389) );
  CLKBUFX2TS U1781 ( .A(n1249), .Y(n3198) );
  CLKBUFX2TS U1782 ( .A(n3394), .Y(n3393) );
  CLKBUFX2TS U1783 ( .A(n3395), .Y(n3390) );
  CLKBUFX2TS U1784 ( .A(n3394), .Y(n3391) );
  CLKBUFX2TS U1785 ( .A(n3394), .Y(n3392) );
  CLKBUFX2TS U1786 ( .A(n3446), .Y(n3440) );
  CLKBUFX2TS U1787 ( .A(n1151), .Y(n3676) );
  CLKBUFX2TS U1788 ( .A(n1152), .Y(n3658) );
  CLKBUFX2TS U1789 ( .A(n1152), .Y(n3659) );
  CLKBUFX2TS U1790 ( .A(n1151), .Y(n3675) );
  CLKBUFX2TS U1791 ( .A(n1202), .Y(n3445) );
  CLKBUFX2TS U1792 ( .A(n1202), .Y(n3446) );
  CLKBUFX2TS U1793 ( .A(n1249), .Y(n3196) );
  CLKBUFX2TS U1794 ( .A(n1249), .Y(n3197) );
  CLKBUFX2TS U1795 ( .A(n1263), .Y(n3025) );
  CLKBUFX2TS U1796 ( .A(n1233), .Y(n3263) );
  CLKBUFX2TS U1797 ( .A(n1263), .Y(n3024) );
  CLKBUFX2TS U1798 ( .A(n1233), .Y(n3264) );
  CLKBUFX2TS U1799 ( .A(n4), .Y(n3903) );
  CLKBUFX2TS U1800 ( .A(n4), .Y(n3904) );
  CLKBUFX2TS U1801 ( .A(n773), .Y(n3863) );
  CLKBUFX2TS U1802 ( .A(n1250), .Y(n3121) );
  CLKBUFX2TS U1803 ( .A(n1250), .Y(n3136) );
  CLKBUFX2TS U1804 ( .A(n1216), .Y(n3411) );
  CLKBUFX2TS U1805 ( .A(n1216), .Y(n3412) );
  INVX2TS U1806 ( .A(n2989), .Y(n969) );
  INVX2TS U1807 ( .A(n1812), .Y(n946) );
  CLKBUFX2TS U1808 ( .A(n777), .Y(n3822) );
  CLKBUFX2TS U1809 ( .A(n528), .Y(n3493) );
  CLKBUFX2TS U1810 ( .A(n527), .Y(n3641) );
  CLKBUFX2TS U1811 ( .A(n527), .Y(n3640) );
  CLKBUFX2TS U1812 ( .A(n3378), .Y(n3375) );
  CLKBUFX2TS U1813 ( .A(n3378), .Y(n3376) );
  INVX2TS U1814 ( .A(n1811), .Y(n949) );
  CLKBUFX2TS U1815 ( .A(n527), .Y(n3642) );
  CLKBUFX2TS U1816 ( .A(n528), .Y(n3494) );
  CLKBUFX2TS U1817 ( .A(n3378), .Y(n3377) );
  CLKBUFX2TS U1818 ( .A(n3621), .Y(n3619) );
  CLKBUFX2TS U1819 ( .A(n3247), .Y(n3246) );
  CLKBUFX2TS U1820 ( .A(n530), .Y(n3577) );
  CLKBUFX2TS U1821 ( .A(n529), .Y(n1213) );
  INVX2TS U1822 ( .A(n531), .Y(n3242) );
  INVX2TS U1823 ( .A(n531), .Y(n3241) );
  CLKBUFX2TS U1824 ( .A(n1048), .Y(n1044) );
  CLKBUFX2TS U1825 ( .A(n1048), .Y(n1045) );
  CLKBUFX2TS U1826 ( .A(n1048), .Y(n1046) );
  CLKBUFX2TS U1827 ( .A(n3723), .Y(n3719) );
  CLKBUFX2TS U1828 ( .A(n3723), .Y(n3720) );
  CLKBUFX2TS U1829 ( .A(n3723), .Y(n3721) );
  CLKBUFX2TS U1830 ( .A(n1248), .Y(n3207) );
  CLKBUFX2TS U1831 ( .A(n3212), .Y(n3210) );
  CLKBUFX2TS U1832 ( .A(n1248), .Y(n3208) );
  CLKBUFX2TS U1833 ( .A(n3212), .Y(n3209) );
  CLKBUFX2TS U1834 ( .A(n1098), .Y(n1097) );
  CLKBUFX2TS U1835 ( .A(n1079), .Y(n1078) );
  CLKBUFX2TS U1836 ( .A(n1064), .Y(n1057) );
  CLKBUFX2TS U1837 ( .A(n1099), .Y(n1093) );
  CLKBUFX2TS U1838 ( .A(n1064), .Y(n1058) );
  CLKBUFX2TS U1839 ( .A(n1079), .Y(n1077) );
  CLKBUFX2TS U1840 ( .A(n1064), .Y(n1059) );
  CLKBUFX2TS U1841 ( .A(n1080), .Y(n1076) );
  CLKBUFX2TS U1842 ( .A(n1099), .Y(n1094) );
  CLKBUFX2TS U1843 ( .A(n1063), .Y(n1061) );
  CLKBUFX2TS U1844 ( .A(n1080), .Y(n1074) );
  CLKBUFX2TS U1845 ( .A(n1098), .Y(n1095) );
  CLKBUFX2TS U1846 ( .A(n1063), .Y(n1060) );
  CLKBUFX2TS U1847 ( .A(n1098), .Y(n1096) );
  CLKBUFX2TS U1848 ( .A(n1080), .Y(n1075) );
  CLKBUFX2TS U1849 ( .A(n3343), .Y(n3337) );
  CLKBUFX2TS U1850 ( .A(n2961), .Y(n2950) );
  CLKBUFX2TS U1851 ( .A(n2974), .Y(n2945) );
  CLKBUFX2TS U1852 ( .A(n2974), .Y(n2938) );
  CLKBUFX2TS U1853 ( .A(n3342), .Y(n3339) );
  CLKBUFX2TS U1854 ( .A(n3343), .Y(n3338) );
  CLKBUFX2TS U1855 ( .A(n3343), .Y(n3336) );
  CLKBUFX2TS U1856 ( .A(n2961), .Y(n2952) );
  CLKBUFX2TS U1857 ( .A(n3342), .Y(n3340) );
  CLKBUFX2TS U1858 ( .A(n3724), .Y(n3722) );
  CLKBUFX2TS U1859 ( .A(n1168), .Y(n3608) );
  CLKBUFX2TS U1860 ( .A(n1168), .Y(n3607) );
  CLKBUFX2TS U1861 ( .A(n1150), .Y(n3690) );
  CLKBUFX2TS U1862 ( .A(n1150), .Y(n3689) );
  CLKBUFX2TS U1863 ( .A(n1184), .Y(n3541) );
  CLKBUFX2TS U1864 ( .A(n1184), .Y(n3542) );
  CLKBUFX2TS U1865 ( .A(n1201), .Y(n3459) );
  CLKBUFX2TS U1866 ( .A(n1201), .Y(n3460) );
  CLKBUFX2TS U1867 ( .A(n2959), .Y(n2895) );
  CLKBUFX2TS U1868 ( .A(n2961), .Y(n2959) );
  CLKBUFX2TS U1869 ( .A(n3341), .Y(n3265) );
  CLKBUFX2TS U1870 ( .A(n3342), .Y(n3341) );
  CLKBUFX2TS U1871 ( .A(n1115), .Y(n1113) );
  CLKBUFX2TS U1872 ( .A(n1115), .Y(n1114) );
  CLKBUFX2TS U1873 ( .A(n3211), .Y(n3199) );
  CLKBUFX2TS U1874 ( .A(n3212), .Y(n3211) );
  INVX2TS U1875 ( .A(n1975), .Y(n774) );
  CLKBUFX2TS U1876 ( .A(n4172), .Y(n4174) );
  CLKBUFX2TS U1877 ( .A(n4175), .Y(n4177) );
  CLKBUFX2TS U1878 ( .A(n1062), .Y(n1049) );
  CLKBUFX2TS U1879 ( .A(n1063), .Y(n1062) );
  CLKBUFX2TS U1880 ( .A(n3718), .Y(n3716) );
  CLKBUFX2TS U1881 ( .A(n3718), .Y(n3717) );
  INVX2TS U1882 ( .A(n1047), .Y(n1033) );
  INVX2TS U1883 ( .A(n532), .Y(n1034) );
  INVX2TS U1884 ( .A(n1047), .Y(n1035) );
  INVX2TS U1885 ( .A(n1046), .Y(n1036) );
  INVX2TS U1886 ( .A(n1048), .Y(n1037) );
  INVX2TS U1887 ( .A(n1047), .Y(n1038) );
  INVX2TS U1888 ( .A(n1047), .Y(n1039) );
  INVX2TS U1889 ( .A(n532), .Y(n1040) );
  CLKBUFX2TS U1890 ( .A(n987), .Y(n986) );
  CLKBUFX2TS U1891 ( .A(n3738), .Y(n3737) );
  CLKBUFX2TS U1892 ( .A(n987), .Y(n985) );
  CLKBUFX2TS U1893 ( .A(n1003), .Y(n1001) );
  CLKBUFX2TS U1894 ( .A(n1144), .Y(n3736) );
  CLKBUFX2TS U1895 ( .A(n988), .Y(n984) );
  CLKBUFX2TS U1896 ( .A(n3738), .Y(n3734) );
  CLKBUFX2TS U1897 ( .A(n988), .Y(n983) );
  CLKBUFX2TS U1898 ( .A(n1003), .Y(n1000) );
  CLKBUFX2TS U1899 ( .A(n3738), .Y(n3735) );
  CLKBUFX2TS U1900 ( .A(n988), .Y(n978) );
  CLKBUFX2TS U1901 ( .A(n1003), .Y(n999) );
  CLKBUFX2TS U1902 ( .A(n548), .Y(n547) );
  CLKBUFX2TS U1903 ( .A(n562), .Y(n561) );
  CLKBUFX2TS U1904 ( .A(n782), .Y(n779) );
  CLKBUFX2TS U1905 ( .A(n965), .Y(n964) );
  CLKBUFX2TS U1906 ( .A(n1016), .Y(n1015) );
  CLKBUFX2TS U1907 ( .A(n2169), .Y(n546) );
  CLKBUFX2TS U1908 ( .A(n2167), .Y(n560) );
  CLKBUFX2TS U1909 ( .A(n2165), .Y(n963) );
  CLKBUFX2TS U1910 ( .A(n1016), .Y(n1014) );
  CLKBUFX2TS U1911 ( .A(n783), .Y(n778) );
  CLKBUFX2TS U1912 ( .A(n1017), .Y(n1013) );
  CLKBUFX2TS U1913 ( .A(n1032), .Y(n1030) );
  CLKBUFX2TS U1914 ( .A(n548), .Y(n545) );
  CLKBUFX2TS U1915 ( .A(n562), .Y(n559) );
  CLKBUFX2TS U1916 ( .A(n783), .Y(n776) );
  CLKBUFX2TS U1917 ( .A(n965), .Y(n962) );
  CLKBUFX2TS U1918 ( .A(n1017), .Y(n1012) );
  CLKBUFX2TS U1919 ( .A(n1032), .Y(n1028) );
  CLKBUFX2TS U1920 ( .A(n548), .Y(n544) );
  CLKBUFX2TS U1921 ( .A(n562), .Y(n558) );
  CLKBUFX2TS U1922 ( .A(n783), .Y(n772) );
  CLKBUFX2TS U1923 ( .A(n965), .Y(n961) );
  CLKBUFX2TS U1924 ( .A(n1017), .Y(n1011) );
  CLKBUFX2TS U1925 ( .A(n1032), .Y(n1027) );
  CLKBUFX2TS U1926 ( .A(n2163), .Y(n1002) );
  CLKBUFX2TS U1927 ( .A(n4175), .Y(n4176) );
  CLKBUFX2TS U1928 ( .A(n4172), .Y(n4173) );
  CLKBUFX2TS U1929 ( .A(n781), .Y(n710) );
  CLKBUFX2TS U1930 ( .A(n782), .Y(n781) );
  CLKBUFX2TS U1931 ( .A(n1031), .Y(n1018) );
  CLKBUFX2TS U1932 ( .A(n2160), .Y(n1031) );
  INVX2TS U1933 ( .A(n4150), .Y(n4147) );
  OAI21X1TS U1934 ( .A0(n127), .A1(n3003), .B0(n2971), .Y(n2989) );
  OAI211X1TS U1935 ( .A0(n954), .A1(n956), .B0(n1859), .C0(n1986), .Y(n1836)
         );
  OAI21X1TS U1936 ( .A0(n951), .A1(n2009), .B0(n1986), .Y(n1850) );
  NOR2X1TS U1937 ( .A(n954), .B(n956), .Y(n2009) );
  NAND2X1TS U1938 ( .A(n127), .B(n3003), .Y(n2971) );
  AND3X2TS U1939 ( .A(n1894), .B(n947), .C(n957), .Y(n1821) );
  INVX2TS U1940 ( .A(n1842), .Y(n944) );
  NAND2X1TS U1941 ( .A(n969), .B(n2972), .Y(n2973) );
  NAND2BX1TS U1942 ( .AN(n2971), .B(n2972), .Y(n2970) );
  INVX2TS U1943 ( .A(n2011), .Y(n956) );
  OA22X1TS U1944 ( .A0(n1820), .A1(n233), .B0(n1879), .B1(n1917), .Y(n529) );
  CLKBUFX2TS U1945 ( .A(n1167), .Y(n3625) );
  CLKBUFX2TS U1946 ( .A(n1217), .Y(n3394) );
  OAI22X1TS U1947 ( .A0(n1135), .A1(n148), .B0(n1134), .B1(n9), .Y(n2887) );
  NAND2X1TS U1948 ( .A(n2010), .B(n2011), .Y(n1853) );
  NAND2X1TS U1949 ( .A(n960), .B(n1878), .Y(n1975) );
  CLKBUFX2TS U1950 ( .A(n531), .Y(n3247) );
  INVX2TS U1951 ( .A(n2054), .Y(n940) );
  NOR2BX1TS U1952 ( .AN(n1907), .B(n170), .Y(n1168) );
  NOR2BX1TS U1953 ( .AN(n1878), .B(n1879), .Y(n1150) );
  NOR2BX1TS U1954 ( .AN(n1878), .B(n1930), .Y(n1184) );
  NOR2BX1TS U1955 ( .AN(n1907), .B(n143), .Y(n1201) );
  NOR2BX1TS U1956 ( .AN(n140), .B(n233), .Y(n1907) );
  CLKBUFX2TS U1957 ( .A(n1146), .Y(n3723) );
  CLKBUFX2TS U1958 ( .A(destinationAddressIn_SOUTH[7]), .Y(n4175) );
  CLKBUFX2TS U1959 ( .A(destinationAddressIn_SOUTH[6]), .Y(n4172) );
  CLKBUFX2TS U1960 ( .A(n2087), .Y(n1081) );
  CLKBUFX2TS U1961 ( .A(n3724), .Y(n3718) );
  CLKBUFX2TS U1962 ( .A(n1146), .Y(n3724) );
  CLKBUFX2TS U1963 ( .A(n1116), .Y(n1115) );
  CLKBUFX2TS U1964 ( .A(n1248), .Y(n3212) );
  CLKBUFX2TS U1965 ( .A(n1264), .Y(n2974) );
  CLKBUFX2TS U1966 ( .A(n1232), .Y(n3343) );
  CLKBUFX2TS U1967 ( .A(n1264), .Y(n2961) );
  CLKBUFX2TS U1968 ( .A(n1232), .Y(n3342) );
  CLKBUFX2TS U1969 ( .A(n2087), .Y(n1079) );
  CLKBUFX2TS U1970 ( .A(n2100), .Y(n1064) );
  CLKBUFX2TS U1971 ( .A(n2086), .Y(n1099) );
  CLKBUFX2TS U1972 ( .A(n2100), .Y(n1063) );
  CLKBUFX2TS U1973 ( .A(n2086), .Y(n1098) );
  CLKBUFX2TS U1974 ( .A(n2087), .Y(n1080) );
  INVX2TS U1975 ( .A(n2010), .Y(n950) );
  INVX2TS U1976 ( .A(n1852), .Y(n943) );
  CLKBUFX2TS U1977 ( .A(n532), .Y(n1047) );
  CLKBUFX2TS U1978 ( .A(n532), .Y(n1048) );
  INVX2TS U1979 ( .A(n4143), .Y(n4141) );
  CLKBUFX2TS U1980 ( .A(n1144), .Y(n3738) );
  CLKBUFX2TS U1981 ( .A(n2164), .Y(n987) );
  CLKBUFX2TS U1982 ( .A(n2164), .Y(n988) );
  CLKBUFX2TS U1983 ( .A(n2163), .Y(n1003) );
  CLKBUFX2TS U1984 ( .A(n2166), .Y(n782) );
  CLKBUFX2TS U1985 ( .A(n2161), .Y(n1016) );
  CLKBUFX2TS U1986 ( .A(n2167), .Y(n562) );
  CLKBUFX2TS U1987 ( .A(n2166), .Y(n783) );
  CLKBUFX2TS U1988 ( .A(n2165), .Y(n965) );
  CLKBUFX2TS U1989 ( .A(n2161), .Y(n1017) );
  CLKBUFX2TS U1990 ( .A(n2160), .Y(n1032) );
  CLKBUFX2TS U1991 ( .A(n2169), .Y(n548) );
  CLKBUFX2TS U1992 ( .A(n4057), .Y(n4058) );
  CLKBUFX2TS U1993 ( .A(dataIn_NORTH[31]), .Y(n4119) );
  CLKBUFX2TS U1994 ( .A(n4089), .Y(n4090) );
  CLKBUFX2TS U1995 ( .A(n4087), .Y(n4088) );
  CLKBUFX2TS U1996 ( .A(n4079), .Y(n4080) );
  CLKBUFX2TS U1997 ( .A(dataIn_NORTH[1]), .Y(n4059) );
  CLKBUFX2TS U1998 ( .A(n4117), .Y(n4118) );
  CLKBUFX2TS U1999 ( .A(n4115), .Y(n4116) );
  CLKBUFX2TS U2000 ( .A(n4113), .Y(n4114) );
  CLKBUFX2TS U2001 ( .A(dataIn_NORTH[27]), .Y(n4111) );
  CLKBUFX2TS U2002 ( .A(n4109), .Y(n4110) );
  CLKBUFX2TS U2003 ( .A(n4107), .Y(n4108) );
  CLKBUFX2TS U2004 ( .A(n4105), .Y(n4106) );
  CLKBUFX2TS U2005 ( .A(n4103), .Y(n4104) );
  CLKBUFX2TS U2006 ( .A(n4101), .Y(n4102) );
  CLKBUFX2TS U2007 ( .A(n4099), .Y(n4100) );
  CLKBUFX2TS U2008 ( .A(n4097), .Y(n4098) );
  CLKBUFX2TS U2009 ( .A(n4095), .Y(n4096) );
  CLKBUFX2TS U2010 ( .A(n4093), .Y(n4094) );
  CLKBUFX2TS U2011 ( .A(n4091), .Y(n4092) );
  CLKBUFX2TS U2012 ( .A(n4085), .Y(n4086) );
  CLKBUFX2TS U2013 ( .A(n4083), .Y(n4084) );
  CLKBUFX2TS U2014 ( .A(n4081), .Y(n4082) );
  CLKBUFX2TS U2015 ( .A(n4077), .Y(n4078) );
  CLKBUFX2TS U2016 ( .A(dataIn_NORTH[9]), .Y(n4075) );
  CLKBUFX2TS U2017 ( .A(n4073), .Y(n4074) );
  CLKBUFX2TS U2018 ( .A(n4071), .Y(n4072) );
  CLKBUFX2TS U2019 ( .A(n4069), .Y(n4070) );
  CLKBUFX2TS U2020 ( .A(dataIn_NORTH[5]), .Y(n4067) );
  CLKBUFX2TS U2021 ( .A(n4065), .Y(n4066) );
  CLKBUFX2TS U2022 ( .A(n4063), .Y(n4064) );
  CLKBUFX2TS U2023 ( .A(n4061), .Y(n4062) );
  INVX2TS U2024 ( .A(n3992), .Y(n3990) );
  INVX2TS U2025 ( .A(n3989), .Y(n3987) );
  INVX2TS U2026 ( .A(n3986), .Y(n3984) );
  INVX2TS U2027 ( .A(n3983), .Y(n3981) );
  INVX2TS U2028 ( .A(n3980), .Y(n3978) );
  INVX2TS U2029 ( .A(n3977), .Y(n3975) );
  INVX2TS U2030 ( .A(n3950), .Y(n3948) );
  INVX2TS U2031 ( .A(n3947), .Y(n3945) );
  INVX2TS U2032 ( .A(n3944), .Y(n3942) );
  INVX2TS U2033 ( .A(n3941), .Y(n3939) );
  INVX2TS U2034 ( .A(n3938), .Y(n3936) );
  INVX2TS U2035 ( .A(n3935), .Y(n3933) );
  INVX2TS U2036 ( .A(n4384), .Y(n4382) );
  INVX2TS U2037 ( .A(n4378), .Y(n4376) );
  INVX2TS U2038 ( .A(n4375), .Y(n4373) );
  INVX2TS U2039 ( .A(n4372), .Y(n4370) );
  INVX2TS U2040 ( .A(n4369), .Y(n4367) );
  INVX2TS U2041 ( .A(n4366), .Y(n4364) );
  INVX2TS U2042 ( .A(n4363), .Y(n4361) );
  INVX2TS U2043 ( .A(n4348), .Y(n4346) );
  INVX2TS U2044 ( .A(n4333), .Y(n4331) );
  INVX2TS U2045 ( .A(n4321), .Y(n4319) );
  INVX2TS U2046 ( .A(n4315), .Y(n4313) );
  INVX2TS U2047 ( .A(n4309), .Y(n4307) );
  INVX2TS U2048 ( .A(n4306), .Y(n4304) );
  INVX2TS U2049 ( .A(n4300), .Y(n4298) );
  INVX2TS U2050 ( .A(n4387), .Y(n4385) );
  INVX2TS U2051 ( .A(n4381), .Y(n4379) );
  INVX2TS U2052 ( .A(n4360), .Y(n4358) );
  INVX2TS U2053 ( .A(n4357), .Y(n4355) );
  INVX2TS U2054 ( .A(n4354), .Y(n4352) );
  INVX2TS U2055 ( .A(n4351), .Y(n4349) );
  INVX2TS U2056 ( .A(n4342), .Y(n4340) );
  INVX2TS U2057 ( .A(n4330), .Y(n4328) );
  INVX2TS U2058 ( .A(n4327), .Y(n4325) );
  INVX2TS U2059 ( .A(n4324), .Y(n4322) );
  INVX2TS U2060 ( .A(n4318), .Y(n4316) );
  INVX2TS U2061 ( .A(n4312), .Y(n4310) );
  INVX2TS U2062 ( .A(n4297), .Y(n4295) );
  INVX2TS U2063 ( .A(n4294), .Y(n4292) );
  INVX2TS U2064 ( .A(n4345), .Y(n4343) );
  INVX2TS U2065 ( .A(n4339), .Y(n4337) );
  INVX2TS U2066 ( .A(n4336), .Y(n4334) );
  INVX2TS U2067 ( .A(n4303), .Y(n4301) );
  INVX2TS U2068 ( .A(n4029), .Y(n4027) );
  INVX2TS U2069 ( .A(n4020), .Y(n4018) );
  INVX2TS U2070 ( .A(n4017), .Y(n4015) );
  INVX2TS U2071 ( .A(n4032), .Y(n4030) );
  INVX2TS U2072 ( .A(n4026), .Y(n4024) );
  INVX2TS U2073 ( .A(n4023), .Y(n4021) );
  CLKBUFX2TS U2074 ( .A(destinationAddressIn_NORTH[5]), .Y(n4043) );
  CLKBUFX2TS U2075 ( .A(n4041), .Y(n4042) );
  CLKBUFX2TS U2076 ( .A(destinationAddressIn_NORTH[3]), .Y(n4039) );
  CLKBUFX2TS U2077 ( .A(n4037), .Y(n4038) );
  CLKBUFX2TS U2078 ( .A(n4035), .Y(n4036) );
  CLKBUFX2TS U2079 ( .A(destinationAddressIn_NORTH[0]), .Y(n4033) );
  INVX2TS U2080 ( .A(n4138), .Y(n4136) );
  INVX2TS U2081 ( .A(n4132), .Y(n4130) );
  INVX2TS U2082 ( .A(n4135), .Y(n4133) );
  INVX2TS U2083 ( .A(n4129), .Y(n4127) );
  INVX2TS U2084 ( .A(n4126), .Y(n4124) );
  INVX2TS U2085 ( .A(n4123), .Y(n4121) );
  CLKBUFX2TS U2086 ( .A(requesterAddressIn_NORTH[5]), .Y(n4055) );
  CLKBUFX2TS U2087 ( .A(n4053), .Y(n4054) );
  CLKBUFX2TS U2088 ( .A(n4051), .Y(n4052) );
  CLKBUFX2TS U2089 ( .A(n4049), .Y(n4050) );
  CLKBUFX2TS U2090 ( .A(n4047), .Y(n4048) );
  CLKBUFX2TS U2091 ( .A(n4045), .Y(n4046) );
  INVX2TS U2092 ( .A(n4198), .Y(n4196) );
  INVX2TS U2093 ( .A(n4291), .Y(n4289) );
  INVX2TS U2094 ( .A(n4246), .Y(n4244) );
  INVX2TS U2095 ( .A(n4243), .Y(n4241) );
  INVX2TS U2096 ( .A(n4231), .Y(n4229) );
  INVX2TS U2097 ( .A(n4201), .Y(n4199) );
  INVX2TS U2098 ( .A(n4288), .Y(n4286) );
  INVX2TS U2099 ( .A(n4285), .Y(n4283) );
  INVX2TS U2100 ( .A(n4282), .Y(n4280) );
  INVX2TS U2101 ( .A(n4279), .Y(n4277) );
  INVX2TS U2102 ( .A(n4276), .Y(n4274) );
  INVX2TS U2103 ( .A(n4273), .Y(n4271) );
  INVX2TS U2104 ( .A(n4270), .Y(n4268) );
  INVX2TS U2105 ( .A(n4267), .Y(n4265) );
  INVX2TS U2106 ( .A(n4264), .Y(n4262) );
  INVX2TS U2107 ( .A(n4261), .Y(n4259) );
  INVX2TS U2108 ( .A(n4258), .Y(n4256) );
  INVX2TS U2109 ( .A(n4255), .Y(n4253) );
  INVX2TS U2110 ( .A(n4252), .Y(n4250) );
  INVX2TS U2111 ( .A(n4249), .Y(n4247) );
  INVX2TS U2112 ( .A(n4240), .Y(n4238) );
  INVX2TS U2113 ( .A(n4237), .Y(n4235) );
  INVX2TS U2114 ( .A(n4234), .Y(n4232) );
  INVX2TS U2115 ( .A(n4228), .Y(n4226) );
  INVX2TS U2116 ( .A(n4225), .Y(n4223) );
  INVX2TS U2117 ( .A(n4222), .Y(n4220) );
  INVX2TS U2118 ( .A(n4219), .Y(n4217) );
  INVX2TS U2119 ( .A(n4216), .Y(n4214) );
  INVX2TS U2120 ( .A(n4213), .Y(n4211) );
  INVX2TS U2121 ( .A(n4210), .Y(n4208) );
  INVX2TS U2122 ( .A(n4207), .Y(n4205) );
  INVX2TS U2123 ( .A(n4204), .Y(n4202) );
  INVX2TS U2124 ( .A(n4143), .Y(n4142) );
  INVX2TS U2125 ( .A(n4390), .Y(n4388) );
  INVX2TS U2126 ( .A(n4483), .Y(n4481) );
  INVX2TS U2127 ( .A(n4438), .Y(n4436) );
  INVX2TS U2128 ( .A(n4435), .Y(n4433) );
  INVX2TS U2129 ( .A(n4423), .Y(n4421) );
  INVX2TS U2130 ( .A(n4393), .Y(n4391) );
  INVX2TS U2131 ( .A(n4480), .Y(n4478) );
  INVX2TS U2132 ( .A(n4477), .Y(n4475) );
  INVX2TS U2133 ( .A(n4474), .Y(n4472) );
  INVX2TS U2134 ( .A(n4471), .Y(n4469) );
  INVX2TS U2135 ( .A(n4468), .Y(n4466) );
  INVX2TS U2136 ( .A(n4465), .Y(n4463) );
  INVX2TS U2137 ( .A(n4462), .Y(n4460) );
  INVX2TS U2138 ( .A(n4459), .Y(n4457) );
  INVX2TS U2139 ( .A(n4456), .Y(n4454) );
  INVX2TS U2140 ( .A(n4453), .Y(n4451) );
  INVX2TS U2141 ( .A(n4450), .Y(n4448) );
  INVX2TS U2142 ( .A(n4447), .Y(n4445) );
  INVX2TS U2143 ( .A(n4444), .Y(n4442) );
  INVX2TS U2144 ( .A(n4441), .Y(n4439) );
  INVX2TS U2145 ( .A(n4432), .Y(n4430) );
  INVX2TS U2146 ( .A(n4429), .Y(n4427) );
  INVX2TS U2147 ( .A(n4426), .Y(n4424) );
  INVX2TS U2148 ( .A(n4420), .Y(n4418) );
  INVX2TS U2149 ( .A(n4417), .Y(n4415) );
  INVX2TS U2150 ( .A(n4414), .Y(n4412) );
  INVX2TS U2151 ( .A(n4411), .Y(n4409) );
  INVX2TS U2152 ( .A(n4408), .Y(n4406) );
  INVX2TS U2153 ( .A(n4405), .Y(n4403) );
  INVX2TS U2154 ( .A(n4402), .Y(n4400) );
  INVX2TS U2155 ( .A(n4399), .Y(n4397) );
  INVX2TS U2156 ( .A(n4396), .Y(n4394) );
  CLKBUFX2TS U2157 ( .A(n3), .Y(n4139) );
  CLKBUFX2TS U2158 ( .A(n4012), .Y(n4013) );
  CLKBUFX2TS U2159 ( .A(n4009), .Y(n4010) );
  CLKBUFX2TS U2160 ( .A(n3999), .Y(n4000) );
  CLKBUFX2TS U2161 ( .A(destinationAddressIn_WEST[10]), .Y(n4004) );
  CLKBUFX2TS U2162 ( .A(n3993), .Y(n3994) );
  CLKBUFX2TS U2163 ( .A(n4006), .Y(n4007) );
  CLKBUFX2TS U2164 ( .A(destinationAddressIn_WEST[9]), .Y(n4002) );
  CLKBUFX2TS U2165 ( .A(n3996), .Y(n3997) );
  CLKBUFX2TS U2166 ( .A(n4193), .Y(n4194) );
  CLKBUFX2TS U2167 ( .A(n4187), .Y(n4188) );
  CLKBUFX2TS U2168 ( .A(n4181), .Y(n4182) );
  CLKBUFX2TS U2169 ( .A(n4190), .Y(n4191) );
  CLKBUFX2TS U2170 ( .A(n4184), .Y(n4185) );
  CLKBUFX2TS U2171 ( .A(n4178), .Y(n4179) );
  CLKBUFX2TS U2172 ( .A(n4151), .Y(n4152) );
  CLKBUFX2TS U2173 ( .A(n4151), .Y(n4153) );
  CLKBUFX2TS U2174 ( .A(n4193), .Y(n4195) );
  CLKBUFX2TS U2175 ( .A(n4190), .Y(n4192) );
  CLKBUFX2TS U2176 ( .A(n4178), .Y(n4180) );
  CLKBUFX2TS U2177 ( .A(n4184), .Y(n4186) );
  CLKBUFX2TS U2178 ( .A(n4187), .Y(n4189) );
  CLKBUFX2TS U2179 ( .A(n4181), .Y(n4183) );
  CLKBUFX2TS U2180 ( .A(destinationAddressIn_NORTH[5]), .Y(n4044) );
  CLKBUFX2TS U2181 ( .A(destinationAddressIn_NORTH[3]), .Y(n4040) );
  CLKBUFX2TS U2182 ( .A(destinationAddressIn_NORTH[0]), .Y(n4034) );
  CLKBUFX2TS U2183 ( .A(dataIn_NORTH[27]), .Y(n4112) );
  CLKBUFX2TS U2184 ( .A(dataIn_NORTH[9]), .Y(n4076) );
  CLKBUFX2TS U2185 ( .A(dataIn_NORTH[5]), .Y(n4068) );
  CLKBUFX2TS U2186 ( .A(dataIn_NORTH[31]), .Y(n4120) );
  CLKBUFX2TS U2187 ( .A(dataIn_NORTH[1]), .Y(n4060) );
  CLKBUFX2TS U2188 ( .A(n3), .Y(n4140) );
  CLKBUFX2TS U2189 ( .A(n4012), .Y(n4014) );
  CLKBUFX2TS U2190 ( .A(n4006), .Y(n4008) );
  CLKBUFX2TS U2191 ( .A(destinationAddressIn_WEST[9]), .Y(n4003) );
  CLKBUFX2TS U2192 ( .A(n3996), .Y(n3998) );
  CLKBUFX2TS U2193 ( .A(n4009), .Y(n4011) );
  CLKBUFX2TS U2194 ( .A(destinationAddressIn_WEST[10]), .Y(n4005) );
  CLKBUFX2TS U2195 ( .A(n3999), .Y(n4001) );
  CLKBUFX2TS U2196 ( .A(n3993), .Y(n3995) );
  CLKBUFX2TS U2197 ( .A(requesterAddressIn_NORTH[5]), .Y(n4056) );
  CLKBUFX2TS U2198 ( .A(n4150), .Y(n4149) );
  INVX2TS U2199 ( .A(n4171), .Y(n4169) );
  INVX2TS U2200 ( .A(n4168), .Y(n4166) );
  INVX2TS U2201 ( .A(n4165), .Y(n4163) );
  INVX2TS U2202 ( .A(n4162), .Y(n4160) );
  INVX2TS U2203 ( .A(n4159), .Y(n4157) );
  INVX2TS U2204 ( .A(n4156), .Y(n4154) );
  INVX2TS U2205 ( .A(n4501), .Y(n4499) );
  INVX2TS U2206 ( .A(n4498), .Y(n4496) );
  INVX2TS U2207 ( .A(n4495), .Y(n4493) );
  INVX2TS U2208 ( .A(n4492), .Y(n4490) );
  INVX2TS U2209 ( .A(n4489), .Y(n4487) );
  INVX2TS U2210 ( .A(n4486), .Y(n4484) );
  INVX2TS U2211 ( .A(n4480), .Y(n4479) );
  INVX2TS U2212 ( .A(n4474), .Y(n4473) );
  INVX2TS U2213 ( .A(n4471), .Y(n4470) );
  INVX2TS U2214 ( .A(n4468), .Y(n4467) );
  INVX2TS U2215 ( .A(n4465), .Y(n4464) );
  INVX2TS U2216 ( .A(n4462), .Y(n4461) );
  INVX2TS U2217 ( .A(n4459), .Y(n4458) );
  INVX2TS U2218 ( .A(n4444), .Y(n4443) );
  INVX2TS U2219 ( .A(n4429), .Y(n4428) );
  INVX2TS U2220 ( .A(n4417), .Y(n4416) );
  INVX2TS U2221 ( .A(n4411), .Y(n4410) );
  INVX2TS U2222 ( .A(n4405), .Y(n4404) );
  INVX2TS U2223 ( .A(n4402), .Y(n4401) );
  INVX2TS U2224 ( .A(n4396), .Y(n4395) );
  INVX2TS U2225 ( .A(n4483), .Y(n4482) );
  INVX2TS U2226 ( .A(n4477), .Y(n4476) );
  INVX2TS U2227 ( .A(n4456), .Y(n4455) );
  INVX2TS U2228 ( .A(n4453), .Y(n4452) );
  INVX2TS U2229 ( .A(n4450), .Y(n4449) );
  INVX2TS U2230 ( .A(n4447), .Y(n4446) );
  INVX2TS U2231 ( .A(n4438), .Y(n4437) );
  INVX2TS U2232 ( .A(n4426), .Y(n4425) );
  INVX2TS U2233 ( .A(n4423), .Y(n4422) );
  INVX2TS U2234 ( .A(n4420), .Y(n4419) );
  INVX2TS U2235 ( .A(n4414), .Y(n4413) );
  INVX2TS U2236 ( .A(n4408), .Y(n4407) );
  INVX2TS U2237 ( .A(n4393), .Y(n4392) );
  INVX2TS U2238 ( .A(n4390), .Y(n4389) );
  INVX2TS U2239 ( .A(n4441), .Y(n4440) );
  INVX2TS U2240 ( .A(n4435), .Y(n4434) );
  INVX2TS U2241 ( .A(n4432), .Y(n4431) );
  INVX2TS U2242 ( .A(n4399), .Y(n4398) );
  INVX2TS U2243 ( .A(n4146), .Y(n4144) );
  INVX2TS U2244 ( .A(n3974), .Y(n3972) );
  INVX2TS U2245 ( .A(n3968), .Y(n3966) );
  INVX2TS U2246 ( .A(n3962), .Y(n3960) );
  INVX2TS U2247 ( .A(n3956), .Y(n3954) );
  INVX2TS U2248 ( .A(n3971), .Y(n3969) );
  INVX2TS U2249 ( .A(n3965), .Y(n3963) );
  INVX2TS U2250 ( .A(n3959), .Y(n3957) );
  INVX2TS U2251 ( .A(n3953), .Y(n3951) );
  INVX2TS U2252 ( .A(n4294), .Y(n4293) );
  INVX2TS U2253 ( .A(n4387), .Y(n4386) );
  INVX2TS U2254 ( .A(n4342), .Y(n4341) );
  INVX2TS U2255 ( .A(n4339), .Y(n4338) );
  INVX2TS U2256 ( .A(n4327), .Y(n4326) );
  INVX2TS U2257 ( .A(n4297), .Y(n4296) );
  INVX2TS U2258 ( .A(n4384), .Y(n4383) );
  INVX2TS U2259 ( .A(n4381), .Y(n4380) );
  INVX2TS U2260 ( .A(n4378), .Y(n4377) );
  INVX2TS U2261 ( .A(n4375), .Y(n4374) );
  INVX2TS U2262 ( .A(n4372), .Y(n4371) );
  INVX2TS U2263 ( .A(n4369), .Y(n4368) );
  INVX2TS U2264 ( .A(n4366), .Y(n4365) );
  INVX2TS U2265 ( .A(n4363), .Y(n4362) );
  INVX2TS U2266 ( .A(n4360), .Y(n4359) );
  INVX2TS U2267 ( .A(n4357), .Y(n4356) );
  INVX2TS U2268 ( .A(n4354), .Y(n4353) );
  INVX2TS U2269 ( .A(n4351), .Y(n4350) );
  INVX2TS U2270 ( .A(n4348), .Y(n4347) );
  INVX2TS U2271 ( .A(n4345), .Y(n4344) );
  INVX2TS U2272 ( .A(n4336), .Y(n4335) );
  INVX2TS U2273 ( .A(n4333), .Y(n4332) );
  INVX2TS U2274 ( .A(n4330), .Y(n4329) );
  INVX2TS U2275 ( .A(n4324), .Y(n4323) );
  INVX2TS U2276 ( .A(n4321), .Y(n4320) );
  INVX2TS U2277 ( .A(n4318), .Y(n4317) );
  INVX2TS U2278 ( .A(n4315), .Y(n4314) );
  INVX2TS U2279 ( .A(n4312), .Y(n4311) );
  INVX2TS U2280 ( .A(n4309), .Y(n4308) );
  INVX2TS U2281 ( .A(n4306), .Y(n4305) );
  INVX2TS U2282 ( .A(n4303), .Y(n4302) );
  INVX2TS U2283 ( .A(n4300), .Y(n4299) );
  INVX2TS U2284 ( .A(n4498), .Y(n4497) );
  INVX2TS U2285 ( .A(n4489), .Y(n4488) );
  INVX2TS U2286 ( .A(n4486), .Y(n4485) );
  INVX2TS U2287 ( .A(n4501), .Y(n4500) );
  INVX2TS U2288 ( .A(n4495), .Y(n4494) );
  INVX2TS U2289 ( .A(n4492), .Y(n4491) );
  INVX2TS U2290 ( .A(n4171), .Y(n4170) );
  INVX2TS U2291 ( .A(n4168), .Y(n4167) );
  INVX2TS U2292 ( .A(n4165), .Y(n4164) );
  INVX2TS U2293 ( .A(n4162), .Y(n4161) );
  INVX2TS U2294 ( .A(n4159), .Y(n4158) );
  INVX2TS U2295 ( .A(n4156), .Y(n4155) );
  INVX2TS U2296 ( .A(n4146), .Y(n4145) );
  INVX2TS U2297 ( .A(n3971), .Y(n3970) );
  INVX2TS U2298 ( .A(n3968), .Y(n3967) );
  INVX2TS U2299 ( .A(n3962), .Y(n3961) );
  INVX2TS U2300 ( .A(n3959), .Y(n3958) );
  INVX2TS U2301 ( .A(n3953), .Y(n3952) );
  INVX2TS U2302 ( .A(n3974), .Y(n3973) );
  INVX2TS U2303 ( .A(n3965), .Y(n3964) );
  INVX2TS U2304 ( .A(n3956), .Y(n3955) );
  INVX2TS U2305 ( .A(n4032), .Y(n4031) );
  INVX2TS U2306 ( .A(n4026), .Y(n4025) );
  INVX2TS U2307 ( .A(n4029), .Y(n4028) );
  INVX2TS U2308 ( .A(n4023), .Y(n4022) );
  INVX2TS U2309 ( .A(n4020), .Y(n4019) );
  INVX2TS U2310 ( .A(n4017), .Y(n4016) );
  INVX2TS U2311 ( .A(n3992), .Y(n3991) );
  INVX2TS U2312 ( .A(n3986), .Y(n3985) );
  INVX2TS U2313 ( .A(n3983), .Y(n3982) );
  INVX2TS U2314 ( .A(n3980), .Y(n3979) );
  INVX2TS U2315 ( .A(n3989), .Y(n3988) );
  INVX2TS U2316 ( .A(n3977), .Y(n3976) );
  INVX2TS U2317 ( .A(n4291), .Y(n4290) );
  INVX2TS U2318 ( .A(n4288), .Y(n4287) );
  INVX2TS U2319 ( .A(n4285), .Y(n4284) );
  INVX2TS U2320 ( .A(n4276), .Y(n4275) );
  INVX2TS U2321 ( .A(n4273), .Y(n4272) );
  INVX2TS U2322 ( .A(n4270), .Y(n4269) );
  INVX2TS U2323 ( .A(n4264), .Y(n4263) );
  INVX2TS U2324 ( .A(n4261), .Y(n4260) );
  INVX2TS U2325 ( .A(n4255), .Y(n4254) );
  INVX2TS U2326 ( .A(n4252), .Y(n4251) );
  INVX2TS U2327 ( .A(n4249), .Y(n4248) );
  INVX2TS U2328 ( .A(n4246), .Y(n4245) );
  INVX2TS U2329 ( .A(n4243), .Y(n4242) );
  INVX2TS U2330 ( .A(n4240), .Y(n4239) );
  INVX2TS U2331 ( .A(n4237), .Y(n4236) );
  INVX2TS U2332 ( .A(n4234), .Y(n4233) );
  INVX2TS U2333 ( .A(n4231), .Y(n4230) );
  INVX2TS U2334 ( .A(n4228), .Y(n4227) );
  INVX2TS U2335 ( .A(n4222), .Y(n4221) );
  INVX2TS U2336 ( .A(n4219), .Y(n4218) );
  INVX2TS U2337 ( .A(n4216), .Y(n4215) );
  INVX2TS U2338 ( .A(n4210), .Y(n4209) );
  INVX2TS U2339 ( .A(n4207), .Y(n4206) );
  INVX2TS U2340 ( .A(n4282), .Y(n4281) );
  INVX2TS U2341 ( .A(n4279), .Y(n4278) );
  INVX2TS U2342 ( .A(n4267), .Y(n4266) );
  INVX2TS U2343 ( .A(n4258), .Y(n4257) );
  INVX2TS U2344 ( .A(n4225), .Y(n4224) );
  INVX2TS U2345 ( .A(n4213), .Y(n4212) );
  INVX2TS U2346 ( .A(n4204), .Y(n4203) );
  INVX2TS U2347 ( .A(n4201), .Y(n4200) );
  INVX2TS U2348 ( .A(n4198), .Y(n4197) );
  INVX2TS U2349 ( .A(n3950), .Y(n3949) );
  INVX2TS U2350 ( .A(n3947), .Y(n3946) );
  INVX2TS U2351 ( .A(n3944), .Y(n3943) );
  INVX2TS U2352 ( .A(n3941), .Y(n3940) );
  INVX2TS U2353 ( .A(n3938), .Y(n3937) );
  INVX2TS U2354 ( .A(n3935), .Y(n3934) );
  INVX2TS U2355 ( .A(n4138), .Y(n4137) );
  INVX2TS U2356 ( .A(n4135), .Y(n4134) );
  INVX2TS U2357 ( .A(n4132), .Y(n4131) );
  INVX2TS U2358 ( .A(n4129), .Y(n4128) );
  INVX2TS U2359 ( .A(n4126), .Y(n4125) );
  INVX2TS U2360 ( .A(n4123), .Y(n4122) );
  INVX2TS U2361 ( .A(n2991), .Y(n758) );
  INVX2TS U2362 ( .A(n1140), .Y(n757) );
  INVX2TS U2363 ( .A(n2097), .Y(n762) );
  AOI222XLTS U2364 ( .A0(n4139), .A1(n3426), .B0(n4145), .B1(n3405), .C0(n4153), .C1(n3388), .Y(n1799) );
  AOI222XLTS U2365 ( .A0(n4152), .A1(n3463), .B0(n4145), .B1(n3438), .C0(n4140), .C1(n3491), .Y(n1796) );
  XNOR2X1TS U2366 ( .A(n2967), .B(n2969), .Y(n1136) );
  OAI2BB1X1TS U2367 ( .A0N(n2973), .A1N(n2976), .B0(n2977), .Y(n2967) );
  XOR2X1TS U2368 ( .A(n124), .B(n2970), .Y(n2969) );
  OAI21X1TS U2369 ( .A0(n2973), .A1(n2976), .B0(n173), .Y(n2977) );
  XNOR2X1TS U2370 ( .A(n2981), .B(n439), .Y(n1132) );
  NAND2X1TS U2371 ( .A(n2982), .B(n2972), .Y(n2981) );
  XNOR2X1TS U2372 ( .A(n2983), .B(n2976), .Y(n1135) );
  XOR2X1TS U2373 ( .A(n2973), .B(n6), .Y(n2983) );
  OAI21X1TS U2374 ( .A0(n170), .A1(n1889), .B0(n1890), .Y(n1146) );
  NAND3X1TS U2375 ( .A(n2982), .B(n424), .C(n2972), .Y(n2976) );
  OAI21X1TS U2376 ( .A0(n9), .A1(n2061), .B0(n139), .Y(n2060) );
  OAI211X1TS U2377 ( .A0(n757), .A1(n969), .B0(n1138), .C0(n2982), .Y(n2995)
         );
  INVX2TS U2378 ( .A(n2999), .Y(n970) );
  XOR2X1TS U2379 ( .A(n12), .B(n1135), .Y(n2978) );
  OAI221XLTS U2380 ( .A0(n213), .A1(n204), .B0(n3232), .B1(n898), .C0(n1804), 
        .Y(n2572) );
  AOI222XLTS U2381 ( .A0(n4144), .A1(n3085), .B0(n4140), .B1(n3196), .C0(n4153), .C1(n3222), .Y(n1804) );
  OAI221XLTS U2382 ( .A0(n219), .A1(n203), .B0(n1119), .B1(n749), .C0(n1791), 
        .Y(n2577) );
  AOI222XLTS U2383 ( .A0(n4152), .A1(n3615), .B0(n4140), .B1(n3590), .C0(n4144), .C1(n3745), .Y(n1791) );
  OAI221XLTS U2384 ( .A0(n1805), .A1(n204), .B0(n149), .B1(n747), .C0(n1807), 
        .Y(n2571) );
  OAI221XLTS U2385 ( .A0(n225), .A1(n982), .B0(n1801), .B1(n660), .C0(n1802), 
        .Y(n2573) );
  AOI222XLTS U2386 ( .A0(n4152), .A1(n3346), .B0(n4140), .B1(n3256), .C0(n4144), .C1(n3374), .Y(n1802) );
  INVX2TS U2387 ( .A(n2007), .Y(n952) );
  AOI32X1TS U2388 ( .A0(n1142), .A1(n757), .A2(n1138), .B0(n2988), .B1(n2971), 
        .Y(n2987) );
  NOR2X1TS U2389 ( .A(n1888), .B(n232), .Y(n1878) );
  NAND2X1TS U2390 ( .A(n439), .B(n144), .Y(n1917) );
  INVX2TS U2391 ( .A(n1888), .Y(n958) );
  NOR2BX1TS U2392 ( .AN(n1878), .B(n164), .Y(n1248) );
  NOR2BX1TS U2393 ( .AN(n1907), .B(n2024), .Y(n1264) );
  NOR2BX1TS U2394 ( .AN(n1907), .B(n1985), .Y(n1232) );
  INVX2TS U2395 ( .A(n2065), .Y(n1116) );
  NAND4X1TS U2396 ( .A(n2072), .B(n2070), .C(n939), .D(n2960), .Y(n2065) );
  AND3X2TS U2397 ( .A(n2073), .B(n2071), .C(n2074), .Y(n2960) );
  NOR2X1TS U2398 ( .A(n2070), .B(n172), .Y(n2100) );
  NOR2X1TS U2399 ( .A(n2071), .B(n171), .Y(n2087) );
  NOR2X1TS U2400 ( .A(n2073), .B(n171), .Y(n2086) );
  INVX2TS U2401 ( .A(n2085), .Y(n659) );
  AOI221X1TS U2402 ( .A0(n3), .A1(n1093), .B0(writeIn_SOUTH), .B1(n1081), .C0(
        n2088), .Y(n2085) );
  INVX2TS U2403 ( .A(writeIn_EAST), .Y(n4146) );
  INVX2TS U2404 ( .A(n171), .Y(n939) );
  OR2X2TS U2405 ( .A(n2072), .B(n172), .Y(n532) );
  OAI221XLTS U2406 ( .A0(n4149), .A1(n2072), .B0(n4143), .B1(n2073), .C0(n2074), .Y(n2068) );
  NOR2BX1TS U2407 ( .AN(n241), .B(n2082), .Y(n2167) );
  NOR2BX1TS U2408 ( .AN(n242), .B(n2083), .Y(n2166) );
  NOR2BX1TS U2409 ( .AN(n153), .B(n2081), .Y(n2165) );
  NOR2BX1TS U2410 ( .AN(n154), .B(n2097), .Y(n2161) );
  NOR2BX1TS U2411 ( .AN(n240), .B(n2080), .Y(n2160) );
  OAI22X1TS U2412 ( .A0(n647), .A1(n1002), .B0(n829), .B1(n987), .Y(n2956) );
  OAI22X1TS U2413 ( .A0(n636), .A1(n1002), .B0(n828), .B1(n987), .Y(n2947) );
  OAI22X1TS U2414 ( .A0(n635), .A1(n1002), .B0(n827), .B1(n988), .Y(n2937) );
  OAI22X1TS U2415 ( .A0(n634), .A1(n1000), .B0(n826), .B1(n2164), .Y(n2931) );
  OAI22X1TS U2416 ( .A0(n633), .A1(n989), .B0(n825), .B1(n968), .Y(n2920) );
  OAI22X1TS U2417 ( .A0(n632), .A1(n989), .B0(n824), .B1(n968), .Y(n2911) );
  OAI22X1TS U2418 ( .A0(n631), .A1(n989), .B0(n823), .B1(n968), .Y(n2898) );
  OAI22X1TS U2419 ( .A0(n630), .A1(n989), .B0(n822), .B1(n968), .Y(n2891) );
  OAI22X1TS U2420 ( .A0(n629), .A1(n990), .B0(n821), .B1(n986), .Y(n2392) );
  OAI22X1TS U2421 ( .A0(n628), .A1(n990), .B0(n820), .B1(n983), .Y(n2384) );
  OAI22X1TS U2422 ( .A0(n627), .A1(n990), .B0(n819), .B1(n978), .Y(n2376) );
  OAI22X1TS U2423 ( .A0(n626), .A1(n990), .B0(n818), .B1(n984), .Y(n2368) );
  OAI22X1TS U2424 ( .A0(n625), .A1(n991), .B0(n817), .B1(n985), .Y(n2360) );
  OAI22X1TS U2425 ( .A0(n624), .A1(n991), .B0(n816), .B1(n985), .Y(n2353) );
  OAI22X1TS U2426 ( .A0(n623), .A1(n991), .B0(n815), .B1(n985), .Y(n2347) );
  OAI22X1TS U2427 ( .A0(n646), .A1(n991), .B0(n814), .B1(n986), .Y(n2341) );
  OAI22X1TS U2428 ( .A0(n645), .A1(n992), .B0(n813), .B1(n985), .Y(n2335) );
  OAI22X1TS U2429 ( .A0(n622), .A1(n992), .B0(n812), .B1(n983), .Y(n2329) );
  OAI22X1TS U2430 ( .A0(n621), .A1(n992), .B0(n811), .B1(n978), .Y(n2323) );
  OAI22X1TS U2431 ( .A0(n620), .A1(n992), .B0(n810), .B1(n984), .Y(n2317) );
  OAI22X1TS U2432 ( .A0(n644), .A1(n1001), .B0(n809), .B1(n971), .Y(n2311) );
  OAI22X1TS U2433 ( .A0(n619), .A1(n999), .B0(n808), .B1(n971), .Y(n2305) );
  OAI22X1TS U2434 ( .A0(n618), .A1(n1001), .B0(n807), .B1(n971), .Y(n2299) );
  OAI22X1TS U2435 ( .A0(n617), .A1(n1000), .B0(n806), .B1(n971), .Y(n2293) );
  OAI22X1TS U2436 ( .A0(n616), .A1(n993), .B0(n805), .B1(n973), .Y(n2282) );
  OAI22X1TS U2437 ( .A0(n615), .A1(n993), .B0(n804), .B1(n973), .Y(n2276) );
  OAI22X1TS U2438 ( .A0(n614), .A1(n993), .B0(n803), .B1(n973), .Y(n2270) );
  OAI22X1TS U2439 ( .A0(n613), .A1(n993), .B0(n802), .B1(n973), .Y(n2264) );
  OAI22X1TS U2440 ( .A0(n612), .A1(n994), .B0(n801), .B1(n974), .Y(n2258) );
  OAI22X1TS U2441 ( .A0(n611), .A1(n994), .B0(n800), .B1(n974), .Y(n2252) );
  OAI22X1TS U2442 ( .A0(n643), .A1(n994), .B0(n799), .B1(n974), .Y(n2246) );
  OAI22X1TS U2443 ( .A0(n967), .A1(n994), .B0(n798), .B1(n974), .Y(n2240) );
  OAI22X1TS U2444 ( .A0(n657), .A1(n995), .B0(n885), .B1(n975), .Y(n2234) );
  OAI22X1TS U2445 ( .A0(n656), .A1(n995), .B0(n884), .B1(n975), .Y(n2228) );
  OAI22X1TS U2446 ( .A0(n654), .A1(n995), .B0(n883), .B1(n975), .Y(n2216) );
  OAI22X1TS U2447 ( .A0(n653), .A1(n997), .B0(n881), .B1(n976), .Y(n2210) );
  OAI22X1TS U2448 ( .A0(n642), .A1(n997), .B0(n833), .B1(n976), .Y(n2198) );
  OAI22X1TS U2449 ( .A0(n641), .A1(n997), .B0(n796), .B1(n976), .Y(n2192) );
  OAI22X1TS U2450 ( .A0(n640), .A1(n998), .B0(n832), .B1(n977), .Y(n2186) );
  OAI22X1TS U2451 ( .A0(n639), .A1(n998), .B0(n831), .B1(n977), .Y(n2180) );
  OAI22X1TS U2452 ( .A0(n638), .A1(n998), .B0(n830), .B1(n977), .Y(n2174) );
  OAI22X1TS U2453 ( .A0(n637), .A1(n998), .B0(n862), .B1(n977), .Y(n2162) );
  OAI22X1TS U2454 ( .A0(n655), .A1(n995), .B0(n882), .B1(n975), .Y(n2222) );
  OAI22X1TS U2455 ( .A0(n652), .A1(n997), .B0(n880), .B1(n976), .Y(n2204) );
  OAI22X1TS U2456 ( .A0(n981), .A1(n2070), .B0(n431), .B1(n2071), .Y(n2069) );
  NOR2X1TS U2457 ( .A(n2074), .B(n172), .Y(n2169) );
  NAND2X1TS U2458 ( .A(n223), .B(n154), .Y(n1144) );
  NAND2X1TS U2459 ( .A(n238), .B(n241), .Y(n2164) );
  NAND2X1TS U2460 ( .A(n235), .B(n242), .Y(n2163) );
  INVX2TS U2461 ( .A(requesterAddressIn_WEST[3]), .Y(n4026) );
  INVX2TS U2462 ( .A(requesterAddressIn_WEST[2]), .Y(n4023) );
  INVX2TS U2463 ( .A(requesterAddressIn_WEST[1]), .Y(n4020) );
  INVX2TS U2464 ( .A(requesterAddressIn_WEST[0]), .Y(n4017) );
  INVX2TS U2465 ( .A(requesterAddressIn_WEST[5]), .Y(n4032) );
  INVX2TS U2466 ( .A(requesterAddressIn_WEST[4]), .Y(n4029) );
  INVX2TS U2467 ( .A(requesterAddressIn_EAST[4]), .Y(n4135) );
  INVX2TS U2468 ( .A(requesterAddressIn_EAST[1]), .Y(n4126) );
  INVX2TS U2469 ( .A(requesterAddressIn_EAST[0]), .Y(n4123) );
  INVX2TS U2470 ( .A(requesterAddressIn_EAST[5]), .Y(n4138) );
  INVX2TS U2471 ( .A(requesterAddressIn_EAST[3]), .Y(n4132) );
  INVX2TS U2472 ( .A(requesterAddressIn_EAST[2]), .Y(n4129) );
  INVX2TS U2473 ( .A(destinationAddressIn_EAST[2]), .Y(n3941) );
  INVX2TS U2474 ( .A(destinationAddressIn_EAST[5]), .Y(n3950) );
  INVX2TS U2475 ( .A(destinationAddressIn_EAST[4]), .Y(n3947) );
  INVX2TS U2476 ( .A(destinationAddressIn_EAST[3]), .Y(n3944) );
  INVX2TS U2477 ( .A(destinationAddressIn_EAST[1]), .Y(n3938) );
  INVX2TS U2478 ( .A(destinationAddressIn_EAST[0]), .Y(n3935) );
  INVX2TS U2479 ( .A(destinationAddressIn_WEST[5]), .Y(n3992) );
  INVX2TS U2480 ( .A(destinationAddressIn_WEST[4]), .Y(n3989) );
  INVX2TS U2481 ( .A(destinationAddressIn_WEST[3]), .Y(n3986) );
  INVX2TS U2482 ( .A(destinationAddressIn_WEST[2]), .Y(n3983) );
  INVX2TS U2483 ( .A(destinationAddressIn_WEST[1]), .Y(n3980) );
  INVX2TS U2484 ( .A(destinationAddressIn_WEST[0]), .Y(n3977) );
  INVX2TS U2485 ( .A(dataIn_WEST[30]), .Y(n4288) );
  INVX2TS U2486 ( .A(dataIn_WEST[28]), .Y(n4282) );
  INVX2TS U2487 ( .A(dataIn_WEST[27]), .Y(n4279) );
  INVX2TS U2488 ( .A(dataIn_WEST[26]), .Y(n4276) );
  INVX2TS U2489 ( .A(dataIn_WEST[25]), .Y(n4273) );
  INVX2TS U2490 ( .A(dataIn_WEST[24]), .Y(n4270) );
  INVX2TS U2491 ( .A(dataIn_WEST[23]), .Y(n4267) );
  INVX2TS U2492 ( .A(dataIn_WEST[18]), .Y(n4252) );
  INVX2TS U2493 ( .A(dataIn_WEST[13]), .Y(n4237) );
  INVX2TS U2494 ( .A(dataIn_WEST[9]), .Y(n4225) );
  INVX2TS U2495 ( .A(dataIn_WEST[7]), .Y(n4219) );
  INVX2TS U2496 ( .A(dataIn_WEST[5]), .Y(n4213) );
  INVX2TS U2497 ( .A(dataIn_WEST[4]), .Y(n4210) );
  INVX2TS U2498 ( .A(dataIn_WEST[2]), .Y(n4204) );
  INVX2TS U2499 ( .A(dataIn_WEST[31]), .Y(n4291) );
  INVX2TS U2500 ( .A(dataIn_WEST[29]), .Y(n4285) );
  INVX2TS U2501 ( .A(dataIn_WEST[22]), .Y(n4264) );
  INVX2TS U2502 ( .A(dataIn_WEST[21]), .Y(n4261) );
  INVX2TS U2503 ( .A(dataIn_WEST[20]), .Y(n4258) );
  INVX2TS U2504 ( .A(dataIn_WEST[19]), .Y(n4255) );
  INVX2TS U2505 ( .A(dataIn_WEST[16]), .Y(n4246) );
  INVX2TS U2506 ( .A(dataIn_WEST[12]), .Y(n4234) );
  INVX2TS U2507 ( .A(dataIn_WEST[11]), .Y(n4231) );
  INVX2TS U2508 ( .A(dataIn_WEST[10]), .Y(n4228) );
  INVX2TS U2509 ( .A(dataIn_WEST[8]), .Y(n4222) );
  INVX2TS U2510 ( .A(dataIn_WEST[6]), .Y(n4216) );
  INVX2TS U2511 ( .A(dataIn_WEST[1]), .Y(n4201) );
  INVX2TS U2512 ( .A(dataIn_WEST[0]), .Y(n4198) );
  INVX2TS U2513 ( .A(dataIn_WEST[17]), .Y(n4249) );
  INVX2TS U2514 ( .A(dataIn_WEST[15]), .Y(n4243) );
  INVX2TS U2515 ( .A(dataIn_WEST[14]), .Y(n4240) );
  INVX2TS U2516 ( .A(dataIn_WEST[3]), .Y(n4207) );
  INVX2TS U2517 ( .A(readIn_WEST), .Y(n4143) );
  INVX2TS U2518 ( .A(destinationAddressIn_EAST[13]), .Y(n3974) );
  INVX2TS U2519 ( .A(destinationAddressIn_EAST[11]), .Y(n3968) );
  INVX2TS U2520 ( .A(destinationAddressIn_EAST[9]), .Y(n3962) );
  INVX2TS U2521 ( .A(destinationAddressIn_EAST[7]), .Y(n3956) );
  INVX2TS U2522 ( .A(destinationAddressIn_EAST[12]), .Y(n3971) );
  INVX2TS U2523 ( .A(destinationAddressIn_EAST[10]), .Y(n3965) );
  INVX2TS U2524 ( .A(destinationAddressIn_EAST[8]), .Y(n3959) );
  INVX2TS U2525 ( .A(destinationAddressIn_EAST[6]), .Y(n3953) );
  INVX2TS U2526 ( .A(dataIn_EAST[30]), .Y(n4384) );
  INVX2TS U2527 ( .A(dataIn_EAST[28]), .Y(n4378) );
  INVX2TS U2528 ( .A(dataIn_EAST[27]), .Y(n4375) );
  INVX2TS U2529 ( .A(dataIn_EAST[26]), .Y(n4372) );
  INVX2TS U2530 ( .A(dataIn_EAST[25]), .Y(n4369) );
  INVX2TS U2531 ( .A(dataIn_EAST[24]), .Y(n4366) );
  INVX2TS U2532 ( .A(dataIn_EAST[23]), .Y(n4363) );
  INVX2TS U2533 ( .A(dataIn_EAST[18]), .Y(n4348) );
  INVX2TS U2534 ( .A(dataIn_EAST[13]), .Y(n4333) );
  INVX2TS U2535 ( .A(dataIn_EAST[9]), .Y(n4321) );
  INVX2TS U2536 ( .A(dataIn_EAST[7]), .Y(n4315) );
  INVX2TS U2537 ( .A(dataIn_EAST[5]), .Y(n4309) );
  INVX2TS U2538 ( .A(dataIn_EAST[4]), .Y(n4306) );
  INVX2TS U2539 ( .A(dataIn_EAST[2]), .Y(n4300) );
  INVX2TS U2540 ( .A(dataIn_EAST[31]), .Y(n4387) );
  INVX2TS U2541 ( .A(dataIn_EAST[29]), .Y(n4381) );
  INVX2TS U2542 ( .A(dataIn_EAST[22]), .Y(n4360) );
  INVX2TS U2543 ( .A(dataIn_EAST[21]), .Y(n4357) );
  INVX2TS U2544 ( .A(dataIn_EAST[20]), .Y(n4354) );
  INVX2TS U2545 ( .A(dataIn_EAST[19]), .Y(n4351) );
  INVX2TS U2546 ( .A(dataIn_EAST[16]), .Y(n4342) );
  INVX2TS U2547 ( .A(dataIn_EAST[12]), .Y(n4330) );
  INVX2TS U2548 ( .A(dataIn_EAST[11]), .Y(n4327) );
  INVX2TS U2549 ( .A(dataIn_EAST[10]), .Y(n4324) );
  INVX2TS U2550 ( .A(dataIn_EAST[8]), .Y(n4318) );
  INVX2TS U2551 ( .A(dataIn_EAST[6]), .Y(n4312) );
  INVX2TS U2552 ( .A(dataIn_EAST[1]), .Y(n4297) );
  INVX2TS U2553 ( .A(dataIn_EAST[0]), .Y(n4294) );
  INVX2TS U2554 ( .A(dataIn_EAST[17]), .Y(n4345) );
  INVX2TS U2555 ( .A(dataIn_EAST[15]), .Y(n4339) );
  INVX2TS U2556 ( .A(dataIn_EAST[14]), .Y(n4336) );
  INVX2TS U2557 ( .A(dataIn_EAST[3]), .Y(n4303) );
  INVX2TS U2558 ( .A(requesterAddressIn_SOUTH[4]), .Y(n4498) );
  INVX2TS U2559 ( .A(requesterAddressIn_SOUTH[1]), .Y(n4489) );
  INVX2TS U2560 ( .A(requesterAddressIn_SOUTH[0]), .Y(n4486) );
  INVX2TS U2561 ( .A(requesterAddressIn_SOUTH[5]), .Y(n4501) );
  INVX2TS U2562 ( .A(requesterAddressIn_SOUTH[3]), .Y(n4495) );
  INVX2TS U2563 ( .A(requesterAddressIn_SOUTH[2]), .Y(n4492) );
  INVX2TS U2564 ( .A(destinationAddressIn_SOUTH[5]), .Y(n4171) );
  INVX2TS U2565 ( .A(destinationAddressIn_SOUTH[4]), .Y(n4168) );
  INVX2TS U2566 ( .A(destinationAddressIn_SOUTH[3]), .Y(n4165) );
  INVX2TS U2567 ( .A(destinationAddressIn_SOUTH[2]), .Y(n4162) );
  INVX2TS U2568 ( .A(destinationAddressIn_SOUTH[1]), .Y(n4159) );
  INVX2TS U2569 ( .A(destinationAddressIn_SOUTH[0]), .Y(n4156) );
  INVX2TS U2570 ( .A(dataIn_SOUTH[30]), .Y(n4480) );
  INVX2TS U2571 ( .A(dataIn_SOUTH[28]), .Y(n4474) );
  INVX2TS U2572 ( .A(dataIn_SOUTH[27]), .Y(n4471) );
  INVX2TS U2573 ( .A(dataIn_SOUTH[26]), .Y(n4468) );
  INVX2TS U2574 ( .A(dataIn_SOUTH[25]), .Y(n4465) );
  INVX2TS U2575 ( .A(dataIn_SOUTH[24]), .Y(n4462) );
  INVX2TS U2576 ( .A(dataIn_SOUTH[23]), .Y(n4459) );
  INVX2TS U2577 ( .A(dataIn_SOUTH[18]), .Y(n4444) );
  INVX2TS U2578 ( .A(dataIn_SOUTH[13]), .Y(n4429) );
  INVX2TS U2579 ( .A(dataIn_SOUTH[9]), .Y(n4417) );
  INVX2TS U2580 ( .A(dataIn_SOUTH[7]), .Y(n4411) );
  INVX2TS U2581 ( .A(dataIn_SOUTH[5]), .Y(n4405) );
  INVX2TS U2582 ( .A(dataIn_SOUTH[4]), .Y(n4402) );
  INVX2TS U2583 ( .A(dataIn_SOUTH[2]), .Y(n4396) );
  INVX2TS U2584 ( .A(dataIn_SOUTH[31]), .Y(n4483) );
  INVX2TS U2585 ( .A(dataIn_SOUTH[29]), .Y(n4477) );
  INVX2TS U2586 ( .A(dataIn_SOUTH[22]), .Y(n4456) );
  INVX2TS U2587 ( .A(dataIn_SOUTH[21]), .Y(n4453) );
  INVX2TS U2588 ( .A(dataIn_SOUTH[20]), .Y(n4450) );
  INVX2TS U2589 ( .A(dataIn_SOUTH[19]), .Y(n4447) );
  INVX2TS U2590 ( .A(dataIn_SOUTH[16]), .Y(n4438) );
  INVX2TS U2591 ( .A(dataIn_SOUTH[12]), .Y(n4426) );
  INVX2TS U2592 ( .A(dataIn_SOUTH[11]), .Y(n4423) );
  INVX2TS U2593 ( .A(dataIn_SOUTH[10]), .Y(n4420) );
  INVX2TS U2594 ( .A(dataIn_SOUTH[8]), .Y(n4414) );
  INVX2TS U2595 ( .A(dataIn_SOUTH[6]), .Y(n4408) );
  INVX2TS U2596 ( .A(dataIn_SOUTH[1]), .Y(n4393) );
  INVX2TS U2597 ( .A(dataIn_SOUTH[0]), .Y(n4390) );
  INVX2TS U2598 ( .A(dataIn_SOUTH[17]), .Y(n4441) );
  INVX2TS U2599 ( .A(dataIn_SOUTH[15]), .Y(n4435) );
  INVX2TS U2600 ( .A(dataIn_SOUTH[14]), .Y(n4432) );
  INVX2TS U2601 ( .A(dataIn_SOUTH[3]), .Y(n4399) );
  CLKBUFX2TS U2602 ( .A(destinationAddressIn_WEST[13]), .Y(n4012) );
  CLKBUFX2TS U2603 ( .A(destinationAddressIn_WEST[11]), .Y(n4006) );
  CLKBUFX2TS U2604 ( .A(destinationAddressIn_WEST[7]), .Y(n3996) );
  CLKBUFX2TS U2605 ( .A(destinationAddressIn_WEST[12]), .Y(n4009) );
  CLKBUFX2TS U2606 ( .A(destinationAddressIn_WEST[8]), .Y(n3999) );
  CLKBUFX2TS U2607 ( .A(destinationAddressIn_WEST[6]), .Y(n3993) );
  CLKBUFX2TS U2608 ( .A(writeIn_SOUTH), .Y(n4151) );
  CLKBUFX2TS U2609 ( .A(requesterAddressIn_NORTH[4]), .Y(n4053) );
  CLKBUFX2TS U2610 ( .A(requesterAddressIn_NORTH[1]), .Y(n4047) );
  CLKBUFX2TS U2611 ( .A(requesterAddressIn_NORTH[0]), .Y(n4045) );
  CLKBUFX2TS U2612 ( .A(requesterAddressIn_NORTH[3]), .Y(n4051) );
  CLKBUFX2TS U2613 ( .A(requesterAddressIn_NORTH[2]), .Y(n4049) );
  CLKBUFX2TS U2614 ( .A(destinationAddressIn_NORTH[4]), .Y(n4041) );
  CLKBUFX2TS U2615 ( .A(destinationAddressIn_NORTH[2]), .Y(n4037) );
  CLKBUFX2TS U2616 ( .A(destinationAddressIn_NORTH[1]), .Y(n4035) );
  CLKBUFX2TS U2617 ( .A(dataIn_NORTH[30]), .Y(n4117) );
  CLKBUFX2TS U2618 ( .A(dataIn_NORTH[28]), .Y(n4113) );
  CLKBUFX2TS U2619 ( .A(dataIn_NORTH[26]), .Y(n4109) );
  CLKBUFX2TS U2620 ( .A(dataIn_NORTH[25]), .Y(n4107) );
  CLKBUFX2TS U2621 ( .A(dataIn_NORTH[24]), .Y(n4105) );
  CLKBUFX2TS U2622 ( .A(dataIn_NORTH[23]), .Y(n4103) );
  CLKBUFX2TS U2623 ( .A(dataIn_NORTH[18]), .Y(n4093) );
  CLKBUFX2TS U2624 ( .A(dataIn_NORTH[13]), .Y(n4083) );
  CLKBUFX2TS U2625 ( .A(dataIn_NORTH[7]), .Y(n4071) );
  CLKBUFX2TS U2626 ( .A(dataIn_NORTH[4]), .Y(n4065) );
  CLKBUFX2TS U2627 ( .A(dataIn_NORTH[2]), .Y(n4061) );
  CLKBUFX2TS U2628 ( .A(dataIn_NORTH[29]), .Y(n4115) );
  CLKBUFX2TS U2629 ( .A(dataIn_NORTH[22]), .Y(n4101) );
  CLKBUFX2TS U2630 ( .A(dataIn_NORTH[21]), .Y(n4099) );
  CLKBUFX2TS U2631 ( .A(dataIn_NORTH[20]), .Y(n4097) );
  CLKBUFX2TS U2632 ( .A(dataIn_NORTH[19]), .Y(n4095) );
  CLKBUFX2TS U2633 ( .A(dataIn_NORTH[16]), .Y(n4089) );
  CLKBUFX2TS U2634 ( .A(dataIn_NORTH[12]), .Y(n4081) );
  CLKBUFX2TS U2635 ( .A(dataIn_NORTH[11]), .Y(n4079) );
  CLKBUFX2TS U2636 ( .A(dataIn_NORTH[10]), .Y(n4077) );
  CLKBUFX2TS U2637 ( .A(dataIn_NORTH[8]), .Y(n4073) );
  CLKBUFX2TS U2638 ( .A(dataIn_NORTH[6]), .Y(n4069) );
  CLKBUFX2TS U2639 ( .A(dataIn_NORTH[0]), .Y(n4057) );
  CLKBUFX2TS U2640 ( .A(dataIn_NORTH[17]), .Y(n4091) );
  CLKBUFX2TS U2641 ( .A(destinationAddressIn_SOUTH[13]), .Y(n4193) );
  CLKBUFX2TS U2642 ( .A(destinationAddressIn_SOUTH[11]), .Y(n4187) );
  CLKBUFX2TS U2643 ( .A(destinationAddressIn_SOUTH[9]), .Y(n4181) );
  CLKBUFX2TS U2644 ( .A(destinationAddressIn_SOUTH[12]), .Y(n4190) );
  CLKBUFX2TS U2645 ( .A(destinationAddressIn_SOUTH[10]), .Y(n4184) );
  CLKBUFX2TS U2646 ( .A(destinationAddressIn_SOUTH[8]), .Y(n4178) );
  CLKBUFX2TS U2647 ( .A(dataIn_NORTH[15]), .Y(n4087) );
  CLKBUFX2TS U2648 ( .A(dataIn_NORTH[14]), .Y(n4085) );
  CLKBUFX2TS U2649 ( .A(dataIn_NORTH[3]), .Y(n4063) );
  INVX2TS U2650 ( .A(readIn_EAST), .Y(n4150) );
  AOI21X1TS U2651 ( .A0(n242), .A1(n1137), .B0(n7), .Y(n2885) );
  NAND3BX1TS U2652 ( .AN(n1138), .B(n1139), .C(n1140), .Y(n1137) );
  XNOR2X1TS U2653 ( .A(n1141), .B(n1142), .Y(n1139) );
  OAI21X1TS U2654 ( .A0(n168), .A1(n1143), .B0(n3734), .Y(n2884) );
  XOR2X1TS U2655 ( .A(n12), .B(n533), .Y(n3001) );
  NAND2X1TS U2656 ( .A(n424), .B(n430), .Y(n2991) );
  OAI22X1TS U2657 ( .A0(n747), .A1(n2081), .B0(n750), .B1(n2082), .Y(n2095) );
  OAI22X1TS U2658 ( .A0(n221), .A1(n748), .B0(n749), .B1(n2083), .Y(n2094) );
  INVX2TS U2659 ( .A(n2079), .Y(n753) );
  NOR2X1TS U2660 ( .A(n1141), .B(n440), .Y(n2084) );
  XOR2X1TS U2661 ( .A(n441), .B(n168), .Y(n1142) );
  INVX2TS U2662 ( .A(n1985), .Y(n960) );
  OAI22X1TS U2663 ( .A0(n660), .A1(n2097), .B0(n898), .B1(n2080), .Y(n2092) );
  OAI22X1TS U2664 ( .A0(n221), .A1(n648), .B0(n2079), .B1(n650), .Y(n2078) );
  OAI22X1TS U2665 ( .A0(n2080), .A1(n651), .B0(n2081), .B1(n886), .Y(n2077) );
  INVX2TS U2666 ( .A(n2080), .Y(n754) );
  INVX2TS U2667 ( .A(n2083), .Y(n760) );
  NOR2X1TS U2668 ( .A(n533), .B(n127), .Y(n2056) );
  AOI222XLTS U2669 ( .A0(n4007), .A1(n3424), .B0(n3967), .B1(n3407), .C0(n4189), .C1(n1217), .Y(n1981) );
  AOI222XLTS U2670 ( .A0(n3994), .A1(n3426), .B0(n3952), .B1(n3405), .C0(n4174), .C1(n3388), .Y(n1976) );
  AOI222XLTS U2671 ( .A0(n4010), .A1(n3424), .B0(n3970), .B1(n3408), .C0(n4192), .C1(n1217), .Y(n1982) );
  AOI222XLTS U2672 ( .A0(n4002), .A1(n3425), .B0(n3961), .B1(n3407), .C0(n4183), .C1(n3389), .Y(n1979) );
  AOI222XLTS U2673 ( .A0(n4000), .A1(n3425), .B0(n3958), .B1(n3405), .C0(n4180), .C1(n3388), .Y(n1978) );
  AOI222XLTS U2674 ( .A0(n4013), .A1(n3424), .B0(n3973), .B1(n3411), .C0(n4195), .C1(n3394), .Y(n1983) );
  AOI222XLTS U2675 ( .A0(n4004), .A1(n3425), .B0(n3964), .B1(n3408), .C0(n4186), .C1(n3395), .Y(n1980) );
  AOI222XLTS U2676 ( .A0(n3997), .A1(n3426), .B0(n3955), .B1(n3405), .C0(n4177), .C1(n3388), .Y(n1977) );
  AOI222XLTS U2677 ( .A0(n4191), .A1(n3461), .B0(n3970), .B1(n3439), .C0(n4011), .C1(n3489), .Y(n1959) );
  AOI222XLTS U2678 ( .A0(n4188), .A1(n3461), .B0(n3967), .B1(n3439), .C0(n4008), .C1(n3489), .Y(n1958) );
  AOI222XLTS U2679 ( .A0(n4185), .A1(n3461), .B0(n3964), .B1(n3439), .C0(n4005), .C1(n3490), .Y(n1957) );
  AOI222XLTS U2680 ( .A0(n4179), .A1(n3462), .B0(n3958), .B1(n3438), .C0(n4001), .C1(n3490), .Y(n1955) );
  AOI222XLTS U2681 ( .A0(n4176), .A1(n3462), .B0(n3955), .B1(n3438), .C0(n3998), .C1(n3491), .Y(n1954) );
  AOI222XLTS U2682 ( .A0(n4173), .A1(n3462), .B0(n3952), .B1(n3438), .C0(n3995), .C1(n3491), .Y(n1953) );
  AOI222XLTS U2683 ( .A0(n4194), .A1(n3461), .B0(n3973), .B1(n3445), .C0(n4014), .C1(n3489), .Y(n1960) );
  AOI222XLTS U2684 ( .A0(n4182), .A1(n3462), .B0(n3961), .B1(n3439), .C0(n4003), .C1(n3490), .Y(n1956) );
  NOR2X1TS U2685 ( .A(n427), .B(n425), .Y(n2962) );
  OAI2BB2XLTS U2686 ( .B0(n10), .B1(n147), .A0N(n170), .A1N(n147), .Y(n2063)
         );
  XOR2X1TS U2687 ( .A(n166), .B(n1132), .Y(n2980) );
  OAI32X1TS U2688 ( .A0(n2964), .A1(n2965), .A2(n148), .B0(n171), .B1(n764), 
        .Y(N4718) );
  XOR2X1TS U2689 ( .A(n1136), .B(n440), .Y(n2965) );
  NAND2X1TS U2690 ( .A(n2978), .B(n2980), .Y(n2964) );
  OAI221XLTS U2691 ( .A0(n228), .A1(n187), .B0(n205), .B1(n966), .C0(n2053), 
        .Y(n2451) );
  AOI222XLTS U2692 ( .A0(n4013), .A1(n2979), .B0(n3972), .B1(n2389), .C0(n4195), .C1(n524), .Y(n2053) );
  OAI221XLTS U2693 ( .A0(n214), .A1(n186), .B0(n3230), .B1(n934), .C0(n2032), 
        .Y(n2465) );
  OAI221XLTS U2694 ( .A0(n212), .A1(n192), .B0(n3230), .B1(n795), .C0(n2031), 
        .Y(n2466) );
  AOI222XLTS U2695 ( .A0(n3969), .A1(n3100), .B0(n4011), .B1(n3138), .C0(
        destinationAddressIn_SOUTH[12]), .C1(n3229), .Y(n2031) );
  OAI221XLTS U2696 ( .A0(n213), .A1(n188), .B0(n3230), .B1(n794), .C0(n2030), 
        .Y(n2467) );
  AOI222XLTS U2697 ( .A0(n3966), .A1(n3103), .B0(n4008), .B1(n3138), .C0(
        destinationAddressIn_SOUTH[11]), .C1(n3224), .Y(n2030) );
  OAI221XLTS U2698 ( .A0(n214), .A1(n194), .B0(n3230), .B1(n793), .C0(n2029), 
        .Y(n2468) );
  AOI222XLTS U2699 ( .A0(n3963), .A1(n3100), .B0(n4005), .B1(n3138), .C0(
        destinationAddressIn_SOUTH[10]), .C1(n3226), .Y(n2029) );
  OAI221XLTS U2700 ( .A0(n212), .A1(n190), .B0(n3231), .B1(n792), .C0(n2028), 
        .Y(n2469) );
  AOI222XLTS U2701 ( .A0(n3960), .A1(n3103), .B0(n4003), .B1(n3195), .C0(
        destinationAddressIn_SOUTH[9]), .C1(n3227), .Y(n2028) );
  OAI221XLTS U2702 ( .A0(n213), .A1(n196), .B0(n3231), .B1(n791), .C0(n2027), 
        .Y(n2470) );
  AOI222XLTS U2703 ( .A0(n3957), .A1(n3085), .B0(n4001), .B1(n3184), .C0(
        destinationAddressIn_SOUTH[8]), .C1(n3222), .Y(n2027) );
  OAI221XLTS U2704 ( .A0(n214), .A1(n181), .B0(n3231), .B1(n790), .C0(n2026), 
        .Y(n2471) );
  AOI222XLTS U2705 ( .A0(n3954), .A1(n3085), .B0(n3998), .B1(n3193), .C0(n4175), .C1(n3222), .Y(n2026) );
  OAI221XLTS U2706 ( .A0(n212), .A1(n184), .B0(n3231), .B1(n789), .C0(n2025), 
        .Y(n2472) );
  AOI222XLTS U2707 ( .A0(n3951), .A1(n3085), .B0(n3995), .B1(n3195), .C0(n4172), .C1(n3222), .Y(n2025) );
  OAI221XLTS U2708 ( .A0(n220), .A1(n193), .B0(n1117), .B1(n604), .C0(n1914), 
        .Y(n2536) );
  AOI222XLTS U2709 ( .A0(n4191), .A1(n3616), .B0(n4011), .B1(n3588), .C0(n3969), .C1(n3749), .Y(n1914) );
  OAI221XLTS U2710 ( .A0(n1790), .A1(n195), .B0(n1117), .B1(n603), .C0(n1912), 
        .Y(n2538) );
  AOI222XLTS U2711 ( .A0(n4185), .A1(n3615), .B0(n4005), .B1(n3587), .C0(n3963), .C1(n3749), .Y(n1912) );
  OAI221XLTS U2712 ( .A0(n220), .A1(n191), .B0(n1118), .B1(n602), .C0(n1911), 
        .Y(n2539) );
  AOI222XLTS U2713 ( .A0(n4182), .A1(n3616), .B0(n4003), .B1(n3591), .C0(n3960), .C1(n3750), .Y(n1911) );
  OAI221XLTS U2714 ( .A0(n1790), .A1(n184), .B0(n1118), .B1(n601), .C0(n1908), 
        .Y(n2542) );
  AOI222XLTS U2715 ( .A0(n4173), .A1(n3615), .B0(n3995), .B1(n3589), .C0(n3951), .C1(n3745), .Y(n1908) );
  OAI221XLTS U2716 ( .A0(n220), .A1(n186), .B0(n1117), .B1(n598), .C0(n1915), 
        .Y(n2535) );
  AOI222XLTS U2717 ( .A0(n4194), .A1(n3615), .B0(n4014), .B1(n3591), .C0(n3972), .C1(n784), .Y(n1915) );
  OAI221XLTS U2718 ( .A0(n1790), .A1(n189), .B0(n1117), .B1(n597), .C0(n1913), 
        .Y(n2537) );
  AOI222XLTS U2719 ( .A0(n4188), .A1(n3617), .B0(n4008), .B1(n1169), .C0(n3966), .C1(n3746), .Y(n1913) );
  OAI221XLTS U2720 ( .A0(n220), .A1(n196), .B0(n1118), .B1(n596), .C0(n1910), 
        .Y(n2540) );
  AOI222XLTS U2721 ( .A0(n4179), .A1(n3616), .B0(n4001), .B1(n3588), .C0(n3957), .C1(n3745), .Y(n1910) );
  OAI221XLTS U2722 ( .A0(n219), .A1(n181), .B0(n1118), .B1(n595), .C0(n1909), 
        .Y(n2541) );
  AOI222XLTS U2723 ( .A0(n4176), .A1(n3616), .B0(n3998), .B1(n3590), .C0(n3954), .C1(n3745), .Y(n1909) );
  OAI221XLTS U2724 ( .A0(n227), .A1(n192), .B0(n205), .B1(n577), .C0(n2052), 
        .Y(n2452) );
  AOI222XLTS U2725 ( .A0(n4010), .A1(n2979), .B0(n3969), .B1(n2389), .C0(n4192), .C1(n1808), .Y(n2052) );
  OAI221XLTS U2726 ( .A0(n228), .A1(n197), .B0(n149), .B1(n576), .C0(n2048), 
        .Y(n2456) );
  OAI221XLTS U2727 ( .A0(n227), .A1(n194), .B0(n128), .B1(n574), .C0(n2050), 
        .Y(n2454) );
  AOI222XLTS U2728 ( .A0(n4004), .A1(n2979), .B0(n3963), .B1(n2389), .C0(n4186), .C1(n1808), .Y(n2050) );
  OAI221XLTS U2729 ( .A0(n228), .A1(n185), .B0(n149), .B1(n573), .C0(n2046), 
        .Y(n2458) );
  OAI221XLTS U2730 ( .A0(n227), .A1(n188), .B0(n128), .B1(n569), .C0(n2051), 
        .Y(n2453) );
  AOI222XLTS U2731 ( .A0(n4007), .A1(n2979), .B0(n3966), .B1(n2372), .C0(n4189), .C1(n524), .Y(n2051) );
  OAI221XLTS U2732 ( .A0(n228), .A1(n191), .B0(n149), .B1(n568), .C0(n2049), 
        .Y(n2455) );
  AOI222XLTS U2733 ( .A0(n4002), .A1(n2985), .B0(n3960), .B1(n2389), .C0(n4183), .C1(n524), .Y(n2049) );
  OAI221XLTS U2734 ( .A0(n227), .A1(n182), .B0(n205), .B1(n567), .C0(n2047), 
        .Y(n2457) );
  OAI221XLTS U2735 ( .A0(n226), .A1(n187), .B0(n207), .B1(n575), .C0(n2006), 
        .Y(n2479) );
  AOI222XLTS U2736 ( .A0(n4194), .A1(n3344), .B0(n4014), .B1(n3260), .C0(n3972), .C1(n3372), .Y(n2006) );
  OAI221XLTS U2737 ( .A0(n1800), .A1(n189), .B0(n208), .B1(n572), .C0(n2004), 
        .Y(n2481) );
  AOI222XLTS U2738 ( .A0(n4188), .A1(n3344), .B0(n4008), .B1(n3258), .C0(n3966), .C1(n3372), .Y(n2004) );
  OAI221XLTS U2739 ( .A0(n226), .A1(n191), .B0(n207), .B1(n571), .C0(n2002), 
        .Y(n2483) );
  AOI222XLTS U2740 ( .A0(n4182), .A1(n3345), .B0(n4003), .B1(n3259), .C0(n3960), .C1(n3373), .Y(n2002) );
  OAI221XLTS U2741 ( .A0(n225), .A1(n181), .B0(n208), .B1(n570), .C0(n2000), 
        .Y(n2485) );
  AOI222XLTS U2742 ( .A0(n4176), .A1(n3345), .B0(n3998), .B1(n3256), .C0(n3954), .C1(n3374), .Y(n2000) );
  OAI221XLTS U2743 ( .A0(n226), .A1(n192), .B0(n207), .B1(n566), .C0(n2005), 
        .Y(n2480) );
  AOI222XLTS U2744 ( .A0(n4191), .A1(n3344), .B0(n4011), .B1(n3261), .C0(n3969), .C1(n3372), .Y(n2005) );
  OAI221XLTS U2745 ( .A0(n1800), .A1(n194), .B0(n208), .B1(n565), .C0(n2003), 
        .Y(n2482) );
  AOI222XLTS U2746 ( .A0(n4185), .A1(n3344), .B0(n4005), .B1(n3262), .C0(n3963), .C1(n3373), .Y(n2003) );
  OAI221XLTS U2747 ( .A0(n226), .A1(n197), .B0(n207), .B1(n564), .C0(n2001), 
        .Y(n2484) );
  AOI222XLTS U2748 ( .A0(n4179), .A1(n3345), .B0(n4001), .B1(n3256), .C0(n3957), .C1(n3373), .Y(n2001) );
  OAI221XLTS U2749 ( .A0(n1800), .A1(n185), .B0(n208), .B1(n563), .C0(n1999), 
        .Y(n2486) );
  AOI222XLTS U2750 ( .A0(n4173), .A1(n3345), .B0(n3995), .B1(n3256), .C0(n3951), .C1(n3374), .Y(n1999) );
  OAI221XLTS U2751 ( .A0(n211), .A1(n187), .B0(n3560), .B1(n588), .C0(n1938), 
        .Y(n2521) );
  AOI222XLTS U2752 ( .A0(n4013), .A1(n3509), .B0(n3973), .B1(n3524), .C0(n4195), .C1(n3555), .Y(n1938) );
  OAI221XLTS U2753 ( .A0(n1792), .A1(n193), .B0(n3560), .B1(n587), .C0(n1937), 
        .Y(n2522) );
  AOI222XLTS U2754 ( .A0(n4010), .A1(n3501), .B0(n3970), .B1(n3526), .C0(n4192), .C1(n3551), .Y(n1937) );
  OAI221XLTS U2755 ( .A0(n210), .A1(n188), .B0(n3560), .B1(n586), .C0(n1936), 
        .Y(n2523) );
  AOI222XLTS U2756 ( .A0(n4007), .A1(n3501), .B0(n3967), .B1(n1185), .C0(n4189), .C1(n3551), .Y(n1936) );
  OAI221XLTS U2757 ( .A0(n211), .A1(n195), .B0(n3560), .B1(n585), .C0(n1935), 
        .Y(n2524) );
  AOI222XLTS U2758 ( .A0(n4004), .A1(n3501), .B0(n3964), .B1(n3527), .C0(n4186), .C1(n3551), .Y(n1935) );
  OAI221XLTS U2759 ( .A0(n1792), .A1(n190), .B0(n3561), .B1(n584), .C0(n1934), 
        .Y(n2525) );
  AOI222XLTS U2760 ( .A0(n4002), .A1(n3501), .B0(n3961), .B1(n3528), .C0(n4183), .C1(n3551), .Y(n1934) );
  OAI221XLTS U2761 ( .A0(n210), .A1(n196), .B0(n3561), .B1(n583), .C0(n1933), 
        .Y(n2526) );
  AOI222XLTS U2762 ( .A0(n4000), .A1(n3503), .B0(n3958), .B1(n3528), .C0(n4180), .C1(n3550), .Y(n1933) );
  OAI221XLTS U2763 ( .A0(n211), .A1(n182), .B0(n3561), .B1(n582), .C0(n1932), 
        .Y(n2527) );
  AOI222XLTS U2764 ( .A0(n3997), .A1(n3503), .B0(n3955), .B1(n3526), .C0(n4177), .C1(n3550), .Y(n1932) );
  OAI221XLTS U2765 ( .A0(n211), .A1(n184), .B0(n3561), .B1(n581), .C0(n1931), 
        .Y(n2528) );
  AOI222XLTS U2766 ( .A0(n3994), .A1(n3503), .B0(n3952), .B1(n3522), .C0(n4174), .C1(n3550), .Y(n1931) );
  OAI221XLTS U2767 ( .A0(n210), .A1(n203), .B0(n3562), .B1(n658), .C0(n1793), 
        .Y(n2576) );
  AOI222XLTS U2768 ( .A0(n4139), .A1(n3502), .B0(n4145), .B1(n3512), .C0(n4152), .C1(n3550), .Y(n1793) );
  OAI221XLTS U2769 ( .A0(n3638), .A1(n191), .B0(n3723), .B1(n897), .C0(n1883), 
        .Y(n2553) );
  AOI222XLTS U2770 ( .A0(n4002), .A1(n3652), .B0(n3961), .B1(n3661), .C0(n4183), .C1(n3700), .Y(n1883) );
  OAI221XLTS U2771 ( .A0(n3637), .A1(n189), .B0(n3722), .B1(n896), .C0(n1885), 
        .Y(n2551) );
  AOI222XLTS U2772 ( .A0(n4007), .A1(n3652), .B0(n3967), .B1(n3660), .C0(n4189), .C1(n3700), .Y(n1885) );
  OAI221XLTS U2773 ( .A0(n3638), .A1(n197), .B0(n3721), .B1(n895), .C0(n1882), 
        .Y(n2554) );
  AOI222XLTS U2774 ( .A0(n4000), .A1(n3651), .B0(n3958), .B1(n3661), .C0(n4180), .C1(n3699), .Y(n1882) );
  OAI221XLTS U2775 ( .A0(n3639), .A1(n181), .B0(n3718), .B1(n894), .C0(n1881), 
        .Y(n2555) );
  AOI222XLTS U2776 ( .A0(n3997), .A1(n3651), .B0(n3955), .B1(n3661), .C0(n4177), .C1(n3699), .Y(n1881) );
  OAI221XLTS U2777 ( .A0(n3639), .A1(n185), .B0(n3724), .B1(n893), .C0(n1880), 
        .Y(n2556) );
  AOI222XLTS U2778 ( .A0(n3994), .A1(n3651), .B0(n3952), .B1(n3661), .C0(n4174), .C1(n3699), .Y(n1880) );
  OAI221XLTS U2779 ( .A0(n3639), .A1(n204), .B0(n3724), .B1(n879), .C0(n1789), 
        .Y(n2578) );
  AOI222XLTS U2780 ( .A0(n4139), .A1(n3651), .B0(n4145), .B1(n3662), .C0(n4153), .C1(n3699), .Y(n1789) );
  OAI221XLTS U2781 ( .A0(n3638), .A1(n194), .B0(n3722), .B1(n871), .C0(n1884), 
        .Y(n2552) );
  AOI222XLTS U2782 ( .A0(n4004), .A1(n3652), .B0(n3964), .B1(n3660), .C0(n4186), .C1(n3700), .Y(n1884) );
  OAI221XLTS U2783 ( .A0(n3637), .A1(n192), .B0(n3720), .B1(n933), .C0(n1886), 
        .Y(n2550) );
  AOI222XLTS U2784 ( .A0(n4010), .A1(n3652), .B0(n3970), .B1(n3660), .C0(n4192), .C1(n3700), .Y(n1886) );
  OAI221XLTS U2785 ( .A0(n3637), .A1(n186), .B0(n3719), .B1(n788), .C0(n1887), 
        .Y(n2549) );
  AOI222XLTS U2786 ( .A0(n4013), .A1(n3658), .B0(n3973), .B1(n3660), .C0(n4195), .C1(n1149), .Y(n1887) );
  AOI22X1TS U2787 ( .A0(n3027), .A1(n4136), .B0(n3878), .B1(n4055), .Y(n1259)
         );
  AOI222XLTS U2788 ( .A0(n3214), .A1(n4500), .B0(n3205), .B1(n119), .C0(n3197), 
        .C1(n4031), .Y(n1260) );
  AOI22X1TS U2789 ( .A0(n3026), .A1(n4133), .B0(n3878), .B1(n4054), .Y(n1257)
         );
  AOI222XLTS U2790 ( .A0(n3213), .A1(n4497), .B0(n3205), .B1(n114), .C0(n3194), 
        .C1(n4028), .Y(n1258) );
  AOI22X1TS U2791 ( .A0(n3026), .A1(n4130), .B0(n3877), .B1(n4052), .Y(n1255)
         );
  AOI222XLTS U2792 ( .A0(n3213), .A1(n4494), .B0(n3210), .B1(n109), .C0(n3196), 
        .C1(n4025), .Y(n1256) );
  AOI22X1TS U2793 ( .A0(n3026), .A1(n4127), .B0(n3877), .B1(n4050), .Y(n1253)
         );
  AOI222XLTS U2794 ( .A0(n3213), .A1(n4491), .B0(n3209), .B1(n104), .C0(n3184), 
        .C1(n4022), .Y(n1254) );
  AOI22X1TS U2795 ( .A0(n3026), .A1(n4124), .B0(n3877), .B1(n4048), .Y(n1251)
         );
  AOI222XLTS U2796 ( .A0(n3213), .A1(n4488), .B0(n3210), .B1(n35), .C0(n3193), 
        .C1(n4019), .Y(n1252) );
  AOI22X1TS U2797 ( .A0(n3027), .A1(n4121), .B0(n3877), .B1(n4046), .Y(n1245)
         );
  AOI222XLTS U2798 ( .A0(n3214), .A1(n4485), .B0(n3205), .B1(n30), .C0(n3196), 
        .C1(n4016), .Y(n1246) );
  AOI22X1TS U2799 ( .A0(n3496), .A1(n4030), .B0(n3767), .B1(n4055), .Y(n1195)
         );
  AOI222XLTS U2800 ( .A0(n1183), .A1(n4499), .B0(n3534), .B1(n120), .C0(n3513), 
        .C1(n4137), .Y(n1196) );
  AOI22X1TS U2801 ( .A0(n3495), .A1(n4027), .B0(n3767), .B1(n4054), .Y(n1193)
         );
  AOI222XLTS U2802 ( .A0(n3543), .A1(n4496), .B0(n3534), .B1(n115), .C0(n3513), 
        .C1(n4134), .Y(n1194) );
  AOI22X1TS U2803 ( .A0(n3495), .A1(n4024), .B0(n3766), .B1(n4052), .Y(n1191)
         );
  AOI222XLTS U2804 ( .A0(n3543), .A1(n4493), .B0(n3533), .B1(n110), .C0(n3512), 
        .C1(n4131), .Y(n1192) );
  AOI22X1TS U2805 ( .A0(n3495), .A1(n4021), .B0(n3766), .B1(n4050), .Y(n1189)
         );
  AOI222XLTS U2806 ( .A0(n3543), .A1(n4490), .B0(n3533), .B1(n105), .C0(n3512), 
        .C1(n4128), .Y(n1190) );
  AOI22X1TS U2807 ( .A0(n3495), .A1(n4018), .B0(n3766), .B1(n4048), .Y(n1187)
         );
  AOI222XLTS U2808 ( .A0(n3543), .A1(n4487), .B0(n3533), .B1(n100), .C0(n3512), 
        .C1(n4125), .Y(n1188) );
  AOI22X1TS U2809 ( .A0(n3496), .A1(n4015), .B0(n3766), .B1(n4046), .Y(n1181)
         );
  AOI222XLTS U2810 ( .A0(n1183), .A1(n4484), .B0(n3534), .B1(n31), .C0(n3513), 
        .C1(n4122), .Y(n1182) );
  AOI222XLTS U2811 ( .A0(n4293), .A1(n3739), .B0(n512), .B1(n3606), .C0(n4197), 
        .C1(n3580), .Y(n1662) );
  AOI222XLTS U2812 ( .A0(n4166), .A1(n3221), .B0(n3206), .B1(n116), .C0(n3988), 
        .C1(n3198), .Y(n2021) );
  AOI22X1TS U2813 ( .A0(n3948), .A1(n3404), .B0(n4169), .B1(n3387), .Y(n1973)
         );
  AOI222XLTS U2814 ( .A0(n3848), .A1(n120), .B0(n4044), .B1(n3864), .C0(n63), 
        .C1(n3860), .Y(n1974) );
  AOI22X1TS U2815 ( .A0(n3945), .A1(n3404), .B0(n4166), .B1(n3387), .Y(n1971)
         );
  AOI222XLTS U2816 ( .A0(n3837), .A1(n115), .B0(n4041), .B1(n3864), .C0(n64), 
        .C1(n3858), .Y(n1972) );
  AOI22X1TS U2817 ( .A0(n3942), .A1(n3404), .B0(n4163), .B1(n3387), .Y(n1969)
         );
  AOI222XLTS U2818 ( .A0(n3837), .A1(n110), .B0(n4040), .B1(n3864), .C0(n65), 
        .C1(n3857), .Y(n1970) );
  AOI22X1TS U2819 ( .A0(n3936), .A1(n3403), .B0(n4157), .B1(n3391), .Y(n1965)
         );
  AOI222XLTS U2820 ( .A0(n3836), .A1(n100), .B0(n4035), .B1(n3865), .C0(n66), 
        .C1(n3857), .Y(n1966) );
  AOI22X1TS U2821 ( .A0(n3933), .A1(n3403), .B0(n4154), .B1(n3393), .Y(n1963)
         );
  AOI222XLTS U2822 ( .A0(n3837), .A1(n31), .B0(n4034), .B1(n3865), .C0(n67), 
        .C1(n3857), .Y(n1964) );
  AOI22X1TS U2823 ( .A0(n3939), .A1(n3404), .B0(n4160), .B1(n3387), .Y(n1967)
         );
  AOI222XLTS U2824 ( .A0(n3837), .A1(n105), .B0(n4037), .B1(n3864), .C0(n92), 
        .C1(n3857), .Y(n1968) );
  AOI22X1TS U2825 ( .A0(n3596), .A1(n32), .B0(n3578), .B1(n4015), .Y(n1165) );
  AOI222XLTS U2826 ( .A0(\requesterAddressbuffer[6][0] ), .A1(n1153), .B0(
        n3625), .B1(n4485), .C0(n3760), .C1(n4045), .Y(n1166) );
  AOI22X1TS U2827 ( .A0(n3596), .A1(n121), .B0(n3579), .B1(n4030), .Y(n1178)
         );
  AOI222XLTS U2828 ( .A0(\requesterAddressbuffer[6][5] ), .A1(n1129), .B0(
        n3618), .B1(n4500), .C0(n3760), .C1(n4056), .Y(n1179) );
  AOI22X1TS U2829 ( .A0(n3596), .A1(n116), .B0(n3578), .B1(n4027), .Y(n1176)
         );
  AOI222XLTS U2830 ( .A0(\requesterAddressbuffer[6][4] ), .A1(n1197), .B0(
        n3619), .B1(n4497), .C0(n3759), .C1(requesterAddressIn_NORTH[4]), .Y(
        n1177) );
  AOI22X1TS U2831 ( .A0(n3595), .A1(n111), .B0(n3578), .B1(n4024), .Y(n1174)
         );
  AOI222XLTS U2832 ( .A0(\requesterAddressbuffer[6][3] ), .A1(n1129), .B0(
        n3619), .B1(n4494), .C0(n3759), .C1(requesterAddressIn_NORTH[3]), .Y(
        n1175) );
  AOI22X1TS U2833 ( .A0(n3595), .A1(n106), .B0(n3578), .B1(n4021), .Y(n1172)
         );
  AOI222XLTS U2834 ( .A0(\requesterAddressbuffer[6][2] ), .A1(n529), .B0(n3619), .B1(n4491), .C0(n3759), .C1(requesterAddressIn_NORTH[2]), .Y(n1173) );
  AOI22X1TS U2835 ( .A0(n3595), .A1(n102), .B0(n3579), .B1(n4018), .Y(n1170)
         );
  AOI222XLTS U2836 ( .A0(\requesterAddressbuffer[6][1] ), .A1(n1128), .B0(
        n3619), .B1(n4488), .C0(n3759), .C1(n4047), .Y(n1171) );
  AOI22X1TS U2837 ( .A0(n3597), .A1(n117), .B0(n3987), .B1(n3592), .Y(n1903)
         );
  AOI222XLTS U2838 ( .A0(n3126), .A1(n1153), .B0(n4167), .B1(n3618), .C0(n4042), .C1(n3761), .Y(n1904) );
  AOI22X1TS U2839 ( .A0(n3595), .A1(n120), .B0(n3990), .B1(n3579), .Y(n1905)
         );
  AOI222XLTS U2840 ( .A0(n3124), .A1(n1128), .B0(n4170), .B1(n3617), .C0(n4043), .C1(n3765), .Y(n1906) );
  AOI22X1TS U2841 ( .A0(n3597), .A1(n112), .B0(n3984), .B1(n3591), .Y(n1901)
         );
  AOI222XLTS U2842 ( .A0(n3129), .A1(n1133), .B0(n4164), .B1(n3618), .C0(n4039), .C1(n3761), .Y(n1902) );
  AOI22X1TS U2843 ( .A0(n3597), .A1(n105), .B0(n3981), .B1(n3579), .Y(n1899)
         );
  AOI222XLTS U2844 ( .A0(n3131), .A1(n1133), .B0(n4161), .B1(n3618), .C0(n4038), .C1(n3765), .Y(n1900) );
  AOI22X1TS U2845 ( .A0(n3596), .A1(n102), .B0(n3978), .B1(n3591), .Y(n1897)
         );
  AOI222XLTS U2846 ( .A0(n3133), .A1(n1133), .B0(n4158), .B1(n3617), .C0(n4036), .C1(n3760), .Y(n1898) );
  AOI22X1TS U2847 ( .A0(n3597), .A1(n33), .B0(n3975), .B1(n3594), .Y(n1895) );
  AOI222XLTS U2848 ( .A0(n3135), .A1(n1129), .B0(n4155), .B1(n3617), .C0(n4033), .C1(n3760), .Y(n1896) );
  AOI22X1TS U2849 ( .A0(n3396), .A1(n4130), .B0(n3379), .B1(n4493), .Y(n1222)
         );
  AOI222XLTS U2850 ( .A0(n3847), .A1(n109), .B0(n3875), .B1(n4052), .C0(
        \requesterAddressbuffer[3][3] ), .C1(n3860), .Y(n1223) );
  AOI22X1TS U2851 ( .A0(n3396), .A1(n4127), .B0(n3379), .B1(n4490), .Y(n1220)
         );
  AOI222XLTS U2852 ( .A0(n3845), .A1(n104), .B0(n3874), .B1(n4050), .C0(
        \requesterAddressbuffer[3][2] ), .C1(n3861), .Y(n1221) );
  AOI22X1TS U2853 ( .A0(n3396), .A1(n4124), .B0(n3379), .B1(n4487), .Y(n1218)
         );
  AOI222XLTS U2854 ( .A0(n3848), .A1(n35), .B0(n3873), .B1(n4048), .C0(
        \requesterAddressbuffer[3][1] ), .C1(n3850), .Y(n1219) );
  AOI22X1TS U2855 ( .A0(n3397), .A1(n4121), .B0(n3380), .B1(n4484), .Y(n1214)
         );
  AOI222XLTS U2856 ( .A0(n3836), .A1(n30), .B0(n3874), .B1(n4046), .C0(
        \requesterAddressbuffer[3][0] ), .C1(n3852), .Y(n1215) );
  AOI22X1TS U2857 ( .A0(n3459), .A1(n112), .B0(n3430), .B1(n4130), .Y(n1207)
         );
  AOI222XLTS U2858 ( .A0(n3034), .A1(n3780), .B0(n3469), .B1(n4494), .C0(n3795), .C1(n4051), .Y(n1208) );
  AOI22X1TS U2859 ( .A0(n3460), .A1(n107), .B0(n3430), .B1(n4127), .Y(n1205)
         );
  AOI222XLTS U2860 ( .A0(n3032), .A1(n3792), .B0(n3469), .B1(n4491), .C0(n3795), .C1(n4049), .Y(n1206) );
  AOI22X1TS U2861 ( .A0(n3459), .A1(n35), .B0(n3430), .B1(n4124), .Y(n1203) );
  AOI222XLTS U2862 ( .A0(n3033), .A1(n3792), .B0(n3469), .B1(n4488), .C0(n3795), .C1(n4047), .Y(n1204) );
  AOI22X1TS U2863 ( .A0(n3447), .A1(n30), .B0(n3441), .B1(n4121), .Y(n1198) );
  AOI222XLTS U2864 ( .A0(n3035), .A1(n3788), .B0(n3469), .B1(n4485), .C0(n3795), .C1(n4045), .Y(n1199) );
  AOI22X1TS U2865 ( .A0(n3265), .A1(n100), .B0(n3263), .B1(n4018), .Y(n1234)
         );
  AOI222XLTS U2866 ( .A0(\requesterAddressbuffer[2][1] ), .A1(n3820), .B0(
        n3353), .B1(n4488), .C0(n3823), .C1(n4047), .Y(n1235) );
  AOI22X1TS U2867 ( .A0(n3266), .A1(n33), .B0(n3260), .B1(n4015), .Y(n1229) );
  AOI222XLTS U2868 ( .A0(\requesterAddressbuffer[2][0] ), .A1(n3821), .B0(
        n3353), .B1(n4485), .C0(n3823), .C1(requesterAddressIn_NORTH[0]), .Y(
        n1230) );
  AOI22X1TS U2869 ( .A0(n3265), .A1(n109), .B0(n3262), .B1(n4024), .Y(n1238)
         );
  AOI222XLTS U2870 ( .A0(\requesterAddressbuffer[2][3] ), .A1(n206), .B0(n3353), .B1(n4494), .C0(n3823), .C1(n4051), .Y(n1239) );
  AOI22X1TS U2871 ( .A0(n3265), .A1(n104), .B0(n3259), .B1(n4021), .Y(n1236)
         );
  AOI222XLTS U2872 ( .A0(\requesterAddressbuffer[2][2] ), .A1(n3820), .B0(
        n3353), .B1(n4491), .C0(n3823), .C1(n4049), .Y(n1237) );
  AOI22X1TS U2873 ( .A0(n3396), .A1(n4133), .B0(n3379), .B1(n4496), .Y(n1224)
         );
  AOI222XLTS U2874 ( .A0(n3836), .A1(n114), .B0(n3876), .B1(n4054), .C0(
        \requesterAddressbuffer[3][4] ), .C1(n3859), .Y(n1225) );
  AOI22X1TS U2875 ( .A0(n3397), .A1(n4136), .B0(n3380), .B1(n4499), .Y(n1226)
         );
  AOI222XLTS U2876 ( .A0(n3836), .A1(n119), .B0(n3875), .B1(n4055), .C0(
        \requesterAddressbuffer[3][5] ), .C1(n3850), .Y(n1227) );
  AOI22X1TS U2877 ( .A0(n3447), .A1(n122), .B0(n3440), .B1(n4136), .Y(n1211)
         );
  AOI222XLTS U2878 ( .A0(n3030), .A1(n3780), .B0(n3468), .B1(n4500), .C0(n3796), .C1(n4056), .Y(n1212) );
  AOI22X1TS U2879 ( .A0(n3447), .A1(n117), .B0(n3430), .B1(n4133), .Y(n1209)
         );
  AOI222XLTS U2880 ( .A0(n3031), .A1(n3780), .B0(n3475), .B1(n4497), .C0(n3796), .C1(n4053), .Y(n1210) );
  AOI22X1TS U2881 ( .A0(n3266), .A1(n114), .B0(n3261), .B1(n4027), .Y(n1240)
         );
  AOI222XLTS U2882 ( .A0(\requesterAddressbuffer[2][4] ), .A1(n777), .B0(n3358), .B1(n4497), .C0(n3824), .C1(n4053), .Y(n1241) );
  AOI22X1TS U2883 ( .A0(n3266), .A1(n119), .B0(n3258), .B1(n4030), .Y(n1242)
         );
  AOI222XLTS U2884 ( .A0(\requesterAddressbuffer[2][5] ), .A1(n777), .B0(n3352), .B1(n4500), .C0(n3824), .C1(n4056), .Y(n1243) );
  AOI22X1TS U2885 ( .A0(n2907), .A1(n120), .B0(n1660), .B1(n4136), .Y(n1274)
         );
  AOI222XLTS U2886 ( .A0(\requesterAddressbuffer[0][5] ), .A1(n3891), .B0(
        n3024), .B1(n4031), .C0(n3920), .C1(n4056), .Y(n1275) );
  AOI22X1TS U2887 ( .A0(n2895), .A1(n110), .B0(n1244), .B1(n4130), .Y(n1270)
         );
  AOI222XLTS U2888 ( .A0(\requesterAddressbuffer[0][3] ), .A1(n3901), .B0(
        n3025), .B1(n4025), .C0(n3919), .C1(n4051), .Y(n1271) );
  AOI22X1TS U2889 ( .A0(n2907), .A1(n115), .B0(n1244), .B1(n4133), .Y(n1272)
         );
  AOI222XLTS U2890 ( .A0(\requesterAddressbuffer[0][4] ), .A1(n3891), .B0(
        n3017), .B1(n4028), .C0(n3920), .C1(n4053), .Y(n1273) );
  AOI22X1TS U2891 ( .A0(n2895), .A1(n105), .B0(n1244), .B1(n4127), .Y(n1268)
         );
  AOI222XLTS U2892 ( .A0(\requesterAddressbuffer[0][2] ), .A1(n3891), .B0(
        n3021), .B1(n4022), .C0(n3919), .C1(n4049), .Y(n1269) );
  AOI22X1TS U2893 ( .A0(n2895), .A1(n101), .B0(n1244), .B1(n4124), .Y(n1266)
         );
  AOI222XLTS U2894 ( .A0(\requesterAddressbuffer[0][1] ), .A1(n3890), .B0(
        n3023), .B1(n4019), .C0(n3919), .C1(requesterAddressIn_NORTH[1]), .Y(
        n1267) );
  AOI22X1TS U2895 ( .A0(n2907), .A1(n31), .B0(n1660), .B1(n4121), .Y(n1261) );
  AOI222XLTS U2896 ( .A0(\requesterAddressbuffer[0][0] ), .A1(n3892), .B0(
        n3023), .B1(n4016), .C0(n3919), .C1(n4045), .Y(n1262) );
  AOI22X1TS U2897 ( .A0(n4030), .A1(n3643), .B0(n4055), .B1(n3635), .Y(n1162)
         );
  AOI222XLTS U2898 ( .A0(n4499), .A1(n3692), .B0(n121), .B1(n3682), .C0(n4137), 
        .C1(n3663), .Y(n1163) );
  AOI22X1TS U2899 ( .A0(n4027), .A1(n3655), .B0(n4054), .B1(n3635), .Y(n1160)
         );
  AOI222XLTS U2900 ( .A0(n4496), .A1(n3691), .B0(n116), .B1(n3682), .C0(n4134), 
        .C1(n3663), .Y(n1161) );
  AOI22X1TS U2901 ( .A0(n4021), .A1(n3657), .B0(n4050), .B1(n3636), .Y(n1156)
         );
  AOI222XLTS U2902 ( .A0(n4490), .A1(n3691), .B0(n106), .B1(n3688), .C0(n4128), 
        .C1(n3663), .Y(n1157) );
  AOI22X1TS U2903 ( .A0(n4024), .A1(n3655), .B0(n4052), .B1(n3636), .Y(n1158)
         );
  AOI222XLTS U2904 ( .A0(n4493), .A1(n3691), .B0(n111), .B1(n3683), .C0(n4131), 
        .C1(n3662), .Y(n1159) );
  AOI22X1TS U2905 ( .A0(n4018), .A1(n3656), .B0(n4048), .B1(n3636), .Y(n1154)
         );
  AOI222XLTS U2906 ( .A0(n4487), .A1(n3691), .B0(n102), .B1(n3688), .C0(n4125), 
        .C1(n3662), .Y(n1155) );
  AOI22X1TS U2907 ( .A0(n4015), .A1(n3646), .B0(n4046), .B1(n3636), .Y(n1147)
         );
  AOI22X1TS U2908 ( .A0(n3975), .A1(n3649), .B0(n4033), .B1(n3627), .Y(n1866)
         );
  AOI222XLTS U2909 ( .A0(n4154), .A1(n3702), .B0(n32), .B1(n3678), .C0(n3934), 
        .C1(n3674), .Y(n1867) );
  AOI22X1TS U2910 ( .A0(n3990), .A1(n3650), .B0(n4043), .B1(n3626), .Y(n1876)
         );
  AOI222XLTS U2911 ( .A0(n4169), .A1(n3698), .B0(n122), .B1(n3677), .C0(n3949), 
        .C1(n3662), .Y(n1877) );
  AOI22X1TS U2912 ( .A0(n3984), .A1(n3650), .B0(n4039), .B1(n3626), .Y(n1872)
         );
  AOI222XLTS U2913 ( .A0(n4163), .A1(n3698), .B0(n112), .B1(n3677), .C0(n3943), 
        .C1(n3675), .Y(n1873) );
  AOI22X1TS U2914 ( .A0(n3981), .A1(n3650), .B0(n4038), .B1(n3626), .Y(n1870)
         );
  AOI222XLTS U2915 ( .A0(n4160), .A1(n3698), .B0(n107), .B1(n3677), .C0(n3940), 
        .C1(n3671), .Y(n1871) );
  AOI22X1TS U2916 ( .A0(n3978), .A1(n3649), .B0(n4036), .B1(n3627), .Y(n1868)
         );
  AOI222XLTS U2917 ( .A0(n4157), .A1(n3703), .B0(n101), .B1(n3678), .C0(n3937), 
        .C1(n3674), .Y(n1869) );
  AOI22X1TS U2918 ( .A0(n4289), .A1(n3649), .B0(n4119), .B1(n3627), .Y(n1787)
         );
  AOI22X1TS U2919 ( .A0(n4286), .A1(n3649), .B0(n4118), .B1(n3627), .Y(n1785)
         );
  AOI22X1TS U2920 ( .A0(n4283), .A1(n3648), .B0(n4116), .B1(n3628), .Y(n1783)
         );
  AOI22X1TS U2921 ( .A0(n4280), .A1(n3648), .B0(n4114), .B1(n3628), .Y(n1781)
         );
  AOI22X1TS U2922 ( .A0(n4277), .A1(n3648), .B0(n4111), .B1(n3628), .Y(n1779)
         );
  AOI22X1TS U2923 ( .A0(n4274), .A1(n3648), .B0(n4110), .B1(n3628), .Y(n1777)
         );
  AOI22X1TS U2924 ( .A0(n4271), .A1(n3647), .B0(n4108), .B1(n3629), .Y(n1775)
         );
  AOI22X1TS U2925 ( .A0(n4268), .A1(n3647), .B0(n4106), .B1(n3629), .Y(n1773)
         );
  AOI22X1TS U2926 ( .A0(n4265), .A1(n3647), .B0(n4104), .B1(n3629), .Y(n1771)
         );
  AOI22X1TS U2927 ( .A0(n4262), .A1(n3647), .B0(n4102), .B1(n3629), .Y(n1769)
         );
  AOI22X1TS U2928 ( .A0(n4259), .A1(n3646), .B0(n4100), .B1(n3630), .Y(n1767)
         );
  AOI22X1TS U2929 ( .A0(n4256), .A1(n3646), .B0(n4098), .B1(n3630), .Y(n1765)
         );
  AOI22X1TS U2930 ( .A0(n4253), .A1(n3646), .B0(n4096), .B1(n3630), .Y(n1763)
         );
  AOI22X1TS U2931 ( .A0(n4250), .A1(n3645), .B0(n4094), .B1(n3630), .Y(n1761)
         );
  AOI22X1TS U2932 ( .A0(n4247), .A1(n3645), .B0(n4092), .B1(n3631), .Y(n1759)
         );
  AOI22X1TS U2933 ( .A0(n4244), .A1(n3645), .B0(n4090), .B1(n3631), .Y(n1757)
         );
  AOI22X1TS U2934 ( .A0(n4241), .A1(n3645), .B0(n4088), .B1(n3631), .Y(n1755)
         );
  AOI22X1TS U2935 ( .A0(n4238), .A1(n3644), .B0(n4086), .B1(n3631), .Y(n1753)
         );
  AOI22X1TS U2936 ( .A0(n4235), .A1(n3644), .B0(n4084), .B1(n3632), .Y(n1751)
         );
  AOI22X1TS U2937 ( .A0(n4232), .A1(n3644), .B0(n4082), .B1(n3632), .Y(n1749)
         );
  AOI22X1TS U2938 ( .A0(n4229), .A1(n3644), .B0(n4080), .B1(n3632), .Y(n1747)
         );
  AOI22X1TS U2939 ( .A0(n4226), .A1(n3657), .B0(n4078), .B1(n3632), .Y(n1745)
         );
  AOI22X1TS U2940 ( .A0(n4223), .A1(n3654), .B0(n4075), .B1(n3633), .Y(n1743)
         );
  AOI22X1TS U2941 ( .A0(n4220), .A1(n3659), .B0(n4074), .B1(n3633), .Y(n1741)
         );
  AOI22X1TS U2942 ( .A0(n4217), .A1(n1152), .B0(n4072), .B1(n3633), .Y(n1739)
         );
  AOI22X1TS U2943 ( .A0(n4214), .A1(n3658), .B0(n4070), .B1(n3633), .Y(n1737)
         );
  AOI22X1TS U2944 ( .A0(n4211), .A1(n3657), .B0(n4067), .B1(n3634), .Y(n1735)
         );
  AOI22X1TS U2945 ( .A0(n4208), .A1(n3656), .B0(n4066), .B1(n3634), .Y(n1733)
         );
  AOI22X1TS U2946 ( .A0(n4205), .A1(n3653), .B0(n4064), .B1(n3634), .Y(n1731)
         );
  AOI22X1TS U2947 ( .A0(n4202), .A1(n3643), .B0(n4062), .B1(n3634), .Y(n1729)
         );
  AOI22X1TS U2948 ( .A0(n4199), .A1(n3643), .B0(n4059), .B1(n3635), .Y(n1727)
         );
  AOI22X1TS U2949 ( .A0(n4196), .A1(n3643), .B0(n4058), .B1(n3635), .Y(n1725)
         );
  AOI22X1TS U2950 ( .A0(n3987), .A1(n3650), .B0(n4042), .B1(n3626), .Y(n1874)
         );
  AOI222XLTS U2951 ( .A0(n4166), .A1(n3698), .B0(n117), .B1(n3677), .C0(n3946), 
        .C1(n3676), .Y(n1875) );
  AOI22X1TS U2952 ( .A0(n2895), .A1(n122), .B0(n3948), .B1(n1916), .Y(n2044)
         );
  AOI222XLTS U2953 ( .A0(n36), .A1(n3890), .B0(n3991), .B1(n2986), .C0(n4044), 
        .C1(n3932), .Y(n2045) );
  AOI22X1TS U2954 ( .A0(n2909), .A1(n109), .B0(n3942), .B1(n1916), .Y(n2040)
         );
  AOI222XLTS U2955 ( .A0(n37), .A1(n3896), .B0(n3985), .B1(n3022), .C0(n4040), 
        .C1(n3932), .Y(n2041) );
  AOI22X1TS U2956 ( .A0(n2909), .A1(n107), .B0(n3939), .B1(n1916), .Y(n2038)
         );
  AOI222XLTS U2957 ( .A0(n38), .A1(n3896), .B0(n3982), .B1(n3017), .C0(n4037), 
        .C1(n3931), .Y(n2039) );
  AOI22X1TS U2958 ( .A0(n2907), .A1(n35), .B0(n3936), .B1(n2366), .Y(n2036) );
  AOI222XLTS U2959 ( .A0(n39), .A1(n3896), .B0(n3979), .B1(n3017), .C0(n4035), 
        .C1(n3928), .Y(n2037) );
  AOI22X1TS U2960 ( .A0(n458), .A1(n2925), .B0(n4385), .B1(n2057), .Y(n1338)
         );
  AOI222XLTS U2961 ( .A0(n40), .A1(n3895), .B0(n4290), .B1(n3017), .C0(n4120), 
        .C1(n3930), .Y(n1339) );
  AOI22X1TS U2962 ( .A0(n461), .A1(n2913), .B0(n4382), .B1(n2155), .Y(n1336)
         );
  AOI222XLTS U2963 ( .A0(n41), .A1(n3895), .B0(n4287), .B1(n3018), .C0(n4117), 
        .C1(n766), .Y(n1337) );
  AOI22X1TS U2964 ( .A0(n463), .A1(n2913), .B0(n4379), .B1(n2057), .Y(n1334)
         );
  AOI222XLTS U2965 ( .A0(n42), .A1(n3895), .B0(n4284), .B1(n3016), .C0(n4115), 
        .C1(n3925), .Y(n1335) );
  AOI22X1TS U2966 ( .A0(n469), .A1(n2938), .B0(n4370), .B1(n2359), .Y(n1328)
         );
  AOI222XLTS U2967 ( .A0(n43), .A1(n3895), .B0(n4275), .B1(n3016), .C0(n4109), 
        .C1(n3925), .Y(n1329) );
  AOI22X1TS U2968 ( .A0(n471), .A1(n2913), .B0(n4367), .B1(n1891), .Y(n1326)
         );
  AOI222XLTS U2969 ( .A0(n44), .A1(n3894), .B0(n4272), .B1(n3015), .C0(n4107), 
        .C1(n3924), .Y(n1327) );
  AOI22X1TS U2970 ( .A0(n473), .A1(n2914), .B0(n4364), .B1(n1891), .Y(n1324)
         );
  AOI222XLTS U2971 ( .A0(n45), .A1(n3894), .B0(n4269), .B1(n3015), .C0(n4105), 
        .C1(n3924), .Y(n1325) );
  AOI22X1TS U2972 ( .A0(n477), .A1(n2914), .B0(n4358), .B1(n1891), .Y(n1320)
         );
  AOI222XLTS U2973 ( .A0(n46), .A1(n3894), .B0(n4263), .B1(n3015), .C0(n4101), 
        .C1(n3924), .Y(n1321) );
  AOI22X1TS U2974 ( .A0(n479), .A1(n2945), .B0(n4355), .B1(n1845), .Y(n1318)
         );
  AOI222XLTS U2975 ( .A0(n47), .A1(n3894), .B0(n4260), .B1(n3019), .C0(n4099), 
        .C1(n3927), .Y(n1319) );
  AOI22X1TS U2976 ( .A0(n483), .A1(n2952), .B0(n4349), .B1(n1845), .Y(n1314)
         );
  AOI222XLTS U2977 ( .A0(n48), .A1(n3893), .B0(n4254), .B1(n3018), .C0(n4095), 
        .C1(n3927), .Y(n1315) );
  AOI22X1TS U2978 ( .A0(n485), .A1(n2945), .B0(n4346), .B1(n1823), .Y(n1312)
         );
  AOI222XLTS U2979 ( .A0(n49), .A1(n3893), .B0(n4251), .B1(n3014), .C0(n4093), 
        .C1(n3926), .Y(n1313) );
  AOI22X1TS U2980 ( .A0(n487), .A1(n2961), .B0(n4343), .B1(n1823), .Y(n1310)
         );
  AOI222XLTS U2981 ( .A0(n50), .A1(n3893), .B0(n4248), .B1(n3014), .C0(n4091), 
        .C1(n3927), .Y(n1311) );
  AOI22X1TS U2982 ( .A0(n489), .A1(n2945), .B0(n4340), .B1(n1823), .Y(n1308)
         );
  AOI222XLTS U2983 ( .A0(n51), .A1(n3893), .B0(n4245), .B1(n3014), .C0(n4089), 
        .C1(n3928), .Y(n1309) );
  AOI22X1TS U2984 ( .A0(n491), .A1(n2938), .B0(n4337), .B1(n1823), .Y(n1306)
         );
  AOI222XLTS U2985 ( .A0(n52), .A1(n3892), .B0(n4242), .B1(n3014), .C0(n4087), 
        .C1(n3929), .Y(n1307) );
  AOI22X1TS U2986 ( .A0(n493), .A1(n2945), .B0(n4334), .B1(n1806), .Y(n1304)
         );
  AOI222XLTS U2987 ( .A0(n53), .A1(n3892), .B0(n4239), .B1(n3004), .C0(n4085), 
        .C1(n3926), .Y(n1305) );
  AOI22X1TS U2988 ( .A0(n495), .A1(n2959), .B0(n4331), .B1(n1806), .Y(n1302)
         );
  AOI222XLTS U2989 ( .A0(n54), .A1(n3892), .B0(n4236), .B1(n3004), .C0(n4083), 
        .C1(n3923), .Y(n1303) );
  AOI22X1TS U2990 ( .A0(n497), .A1(n2938), .B0(n4328), .B1(n1806), .Y(n1300)
         );
  AOI222XLTS U2991 ( .A0(n55), .A1(n3901), .B0(n4233), .B1(n3004), .C0(n4081), 
        .C1(n3923), .Y(n1301) );
  AOI22X1TS U2992 ( .A0(n499), .A1(n2974), .B0(n4325), .B1(n1806), .Y(n1298)
         );
  AOI222XLTS U2993 ( .A0(n56), .A1(n3902), .B0(n4230), .B1(n3004), .C0(n4079), 
        .C1(n3923), .Y(n1299) );
  AOI22X1TS U2994 ( .A0(n501), .A1(n2925), .B0(n4322), .B1(n1803), .Y(n1296)
         );
  AOI222XLTS U2995 ( .A0(n57), .A1(n3898), .B0(n4227), .B1(n2996), .C0(n4077), 
        .C1(n3923), .Y(n1297) );
  AOI22X1TS U2996 ( .A0(n505), .A1(n2952), .B0(n4316), .B1(n1803), .Y(n1292)
         );
  AOI222XLTS U2997 ( .A0(n58), .A1(n3899), .B0(n4221), .B1(n2996), .C0(n4073), 
        .C1(n3922), .Y(n1293) );
  AOI22X1TS U2998 ( .A0(n452), .A1(n2959), .B0(n4313), .B1(n1803), .Y(n1290)
         );
  AOI222XLTS U2999 ( .A0(n59), .A1(n3901), .B0(n4218), .B1(n2996), .C0(n4071), 
        .C1(n3922), .Y(n1291) );
  AOI22X1TS U3000 ( .A0(n507), .A1(n2923), .B0(n4310), .B1(n1803), .Y(n1288)
         );
  AOI222XLTS U3001 ( .A0(n60), .A1(n3901), .B0(n4215), .B1(n3021), .C0(n4069), 
        .C1(n3922), .Y(n1289) );
  AOI22X1TS U3002 ( .A0(n454), .A1(n2923), .B0(n4304), .B1(n1797), .Y(n1284)
         );
  AOI222XLTS U3003 ( .A0(n61), .A1(n3904), .B0(n4209), .B1(n2992), .C0(n4065), 
        .C1(n3921), .Y(n1285) );
  AOI22X1TS U3004 ( .A0(n511), .A1(n2925), .B0(n4301), .B1(n1797), .Y(n1282)
         );
  AOI222XLTS U3005 ( .A0(n62), .A1(n3891), .B0(n4206), .B1(n2992), .C0(n4063), 
        .C1(n3921), .Y(n1283) );
  AOI22X1TS U3006 ( .A0(n2909), .A1(n114), .B0(n3945), .B1(n1916), .Y(n2042)
         );
  AOI222XLTS U3007 ( .A0(n90), .A1(n3897), .B0(n3988), .B1(n3022), .C0(n4041), 
        .C1(n766), .Y(n2043) );
  AOI22X1TS U3008 ( .A0(n2909), .A1(n30), .B0(n3933), .B1(n2359), .Y(n2034) );
  AOI222XLTS U3009 ( .A0(n91), .A1(n3896), .B0(n3976), .B1(n3019), .C0(n4034), 
        .C1(n3929), .Y(n2035) );
  AOI22X1TS U3010 ( .A0(n465), .A1(n2913), .B0(n4376), .B1(n2366), .Y(n1332)
         );
  AOI222XLTS U3011 ( .A0(n3900), .A1(n677), .B0(n4281), .B1(n3016), .C0(n4113), 
        .C1(n3925), .Y(n1333) );
  AOI22X1TS U3012 ( .A0(n467), .A1(n2914), .B0(n4373), .B1(n2155), .Y(n1330)
         );
  AOI222XLTS U3013 ( .A0(n3902), .A1(n676), .B0(n4278), .B1(n3016), .C0(n4112), 
        .C1(n3925), .Y(n1331) );
  AOI22X1TS U3014 ( .A0(n475), .A1(n2914), .B0(n4361), .B1(n1891), .Y(n1322)
         );
  AOI222XLTS U3015 ( .A0(n3900), .A1(n675), .B0(n4266), .B1(n3015), .C0(n4103), 
        .C1(n3924), .Y(n1323) );
  AOI22X1TS U3016 ( .A0(n481), .A1(n2950), .B0(n4352), .B1(n1845), .Y(n1316)
         );
  AOI222XLTS U3017 ( .A0(n3890), .A1(n674), .B0(n4257), .B1(n3019), .C0(n4097), 
        .C1(n3927), .Y(n1317) );
  AOI22X1TS U3018 ( .A0(n503), .A1(n2959), .B0(n4319), .B1(n1845), .Y(n1294)
         );
  AOI222XLTS U3019 ( .A0(n3890), .A1(n673), .B0(n4224), .B1(n2996), .C0(n4076), 
        .C1(n3922), .Y(n1295) );
  AOI22X1TS U3020 ( .A0(n509), .A1(n2938), .B0(n4307), .B1(n1797), .Y(n1286)
         );
  AOI222XLTS U3021 ( .A0(n3903), .A1(n672), .B0(n4212), .B1(n2992), .C0(n4068), 
        .C1(n3921), .Y(n1287) );
  AOI22X1TS U3022 ( .A0(n456), .A1(n2923), .B0(n4298), .B1(n1797), .Y(n1280)
         );
  AOI222XLTS U3023 ( .A0(n3898), .A1(n671), .B0(n4203), .B1(n2992), .C0(n4061), 
        .C1(n3921), .Y(n1281) );
  AOI22X1TS U3024 ( .A0(n515), .A1(n2923), .B0(n4295), .B1(n1660), .Y(n1278)
         );
  AOI222XLTS U3025 ( .A0(n3903), .A1(n670), .B0(n4200), .B1(n2986), .C0(n4060), 
        .C1(n3920), .Y(n1279) );
  AOI22X1TS U3026 ( .A0(n513), .A1(n2925), .B0(n4292), .B1(n1660), .Y(n1276)
         );
  AOI222XLTS U3027 ( .A0(n3899), .A1(n669), .B0(n4197), .B1(n2986), .C0(n4057), 
        .C1(n3920), .Y(n1277) );
  AOI22X1TS U3028 ( .A0(n4196), .A1(n3496), .B0(n4058), .B1(n3767), .Y(n1596)
         );
  AOI222XLTS U3029 ( .A0(n4388), .A1(n3557), .B0(n513), .B1(n3538), .C0(n4293), 
        .C1(n3514), .Y(n1597) );
  AOI22X1TS U3030 ( .A0(n4373), .A1(n3060), .B0(n4111), .B1(n3888), .Y(n1394)
         );
  AOI222XLTS U3031 ( .A0(n4469), .A1(n1247), .B0(n466), .B1(n3199), .C0(n4278), 
        .C1(n3161), .Y(n1395) );
  AOI22X1TS U3032 ( .A0(n4358), .A1(n3049), .B0(n4102), .B1(n3884), .Y(n1384)
         );
  AOI222XLTS U3033 ( .A0(n4454), .A1(n3220), .B0(n476), .B1(n3202), .C0(n4263), 
        .C1(n3157), .Y(n1385) );
  AOI22X1TS U3034 ( .A0(n4352), .A1(n3044), .B0(n4098), .B1(n3883), .Y(n1380)
         );
  AOI222XLTS U3035 ( .A0(n4448), .A1(n3219), .B0(n480), .B1(n3202), .C0(n4257), 
        .C1(n3157), .Y(n1381) );
  AOI22X1TS U3036 ( .A0(n4349), .A1(n3044), .B0(n4096), .B1(n3883), .Y(n1378)
         );
  AOI222XLTS U3037 ( .A0(n4445), .A1(n3219), .B0(n482), .B1(n3203), .C0(n4254), 
        .C1(n3148), .Y(n1379) );
  AOI22X1TS U3038 ( .A0(n4322), .A1(n3121), .B0(n4078), .B1(n3881), .Y(n1360)
         );
  AOI222XLTS U3039 ( .A0(n4418), .A1(n3216), .B0(n500), .B1(n3207), .C0(n4227), 
        .C1(n3143), .Y(n1361) );
  AOI22X1TS U3040 ( .A0(n4316), .A1(n3136), .B0(n4074), .B1(n3880), .Y(n1356)
         );
  AOI222XLTS U3041 ( .A0(n4412), .A1(n3216), .B0(n504), .B1(n3207), .C0(n4221), 
        .C1(n3140), .Y(n1357) );
  AOI22X1TS U3042 ( .A0(n4307), .A1(n1250), .B0(n4067), .B1(n3879), .Y(n1350)
         );
  AOI222XLTS U3043 ( .A0(n4403), .A1(n3215), .B0(n508), .B1(n3204), .C0(n4212), 
        .C1(n3140), .Y(n1351) );
  AOI22X1TS U3044 ( .A0(n4298), .A1(n3112), .B0(n4062), .B1(n3879), .Y(n1344)
         );
  AOI222XLTS U3045 ( .A0(n4394), .A1(n3215), .B0(n455), .B1(n3204), .C0(n4203), 
        .C1(n3139), .Y(n1345) );
  AOI22X1TS U3046 ( .A0(n3948), .A1(n3082), .B0(n4043), .B1(n3888), .Y(n2022)
         );
  AOI222XLTS U3047 ( .A0(n4169), .A1(n3221), .B0(n3208), .B1(n121), .C0(n3991), 
        .C1(n3194), .Y(n2023) );
  AOI22X1TS U3048 ( .A0(n3942), .A1(n3082), .B0(n4039), .B1(n3887), .Y(n2018)
         );
  AOI222XLTS U3049 ( .A0(n4163), .A1(n3221), .B0(n3206), .B1(n111), .C0(n3985), 
        .C1(n3179), .Y(n2019) );
  AOI22X1TS U3050 ( .A0(n3939), .A1(n3082), .B0(n4038), .B1(n3885), .Y(n2016)
         );
  AOI222XLTS U3051 ( .A0(n4160), .A1(n3221), .B0(n3206), .B1(n106), .C0(n3982), 
        .C1(n3179), .Y(n2017) );
  AOI22X1TS U3052 ( .A0(n3936), .A1(n3069), .B0(n4036), .B1(n3889), .Y(n2014)
         );
  AOI222XLTS U3053 ( .A0(n4157), .A1(n3227), .B0(n3206), .B1(n101), .C0(n3979), 
        .C1(n3179), .Y(n2015) );
  AOI22X1TS U3054 ( .A0(n3933), .A1(n3069), .B0(n4033), .B1(n3886), .Y(n2012)
         );
  AOI222XLTS U3055 ( .A0(n4154), .A1(n3228), .B0(n3205), .B1(n32), .C0(n3976), 
        .C1(n3179), .Y(n2013) );
  AOI22X1TS U3056 ( .A0(n4385), .A1(n3069), .B0(n4119), .B1(n3886), .Y(n1402)
         );
  AOI222XLTS U3057 ( .A0(n4481), .A1(n1247), .B0(n457), .B1(n3200), .C0(n4290), 
        .C1(n3172), .Y(n1403) );
  AOI22X1TS U3058 ( .A0(n4382), .A1(n3069), .B0(n4118), .B1(n3887), .Y(n1400)
         );
  AOI222XLTS U3059 ( .A0(n4478), .A1(n3226), .B0(n460), .B1(n3199), .C0(n4287), 
        .C1(n3172), .Y(n1401) );
  AOI22X1TS U3060 ( .A0(n4379), .A1(n3060), .B0(n4116), .B1(n769), .Y(n1398)
         );
  AOI222XLTS U3061 ( .A0(n4475), .A1(n3229), .B0(n462), .B1(n3200), .C0(n4284), 
        .C1(n3172), .Y(n1399) );
  AOI22X1TS U3062 ( .A0(n4376), .A1(n3060), .B0(n4114), .B1(n3888), .Y(n1396)
         );
  AOI222XLTS U3063 ( .A0(n4472), .A1(n3224), .B0(n464), .B1(n3199), .C0(n4281), 
        .C1(n3172), .Y(n1397) );
  AOI22X1TS U3064 ( .A0(n4370), .A1(n3060), .B0(n4110), .B1(n14), .Y(n1392) );
  AOI222XLTS U3065 ( .A0(n4466), .A1(n3225), .B0(n468), .B1(n3201), .C0(n4275), 
        .C1(n3161), .Y(n1393) );
  AOI22X1TS U3066 ( .A0(n4367), .A1(n3049), .B0(n4108), .B1(n3884), .Y(n1390)
         );
  AOI222XLTS U3067 ( .A0(n4463), .A1(n3220), .B0(n470), .B1(n3201), .C0(n4272), 
        .C1(n3161), .Y(n1391) );
  AOI22X1TS U3068 ( .A0(n4364), .A1(n3049), .B0(n4106), .B1(n3884), .Y(n1388)
         );
  AOI222XLTS U3069 ( .A0(n4460), .A1(n3220), .B0(n472), .B1(n3200), .C0(n4269), 
        .C1(n3161), .Y(n1389) );
  AOI22X1TS U3070 ( .A0(n4361), .A1(n3049), .B0(n4104), .B1(n3884), .Y(n1386)
         );
  AOI222XLTS U3071 ( .A0(n4457), .A1(n3220), .B0(n474), .B1(n3202), .C0(n4266), 
        .C1(n3157), .Y(n1387) );
  AOI22X1TS U3072 ( .A0(n4355), .A1(n3044), .B0(n4100), .B1(n3883), .Y(n1382)
         );
  AOI222XLTS U3073 ( .A0(n4451), .A1(n3219), .B0(n478), .B1(n3200), .C0(n4260), 
        .C1(n3157), .Y(n1383) );
  AOI22X1TS U3074 ( .A0(n4346), .A1(n3037), .B0(n4094), .B1(n3883), .Y(n1376)
         );
  AOI222XLTS U3075 ( .A0(n4442), .A1(n3218), .B0(n484), .B1(n3201), .C0(n4251), 
        .C1(n3148), .Y(n1377) );
  AOI22X1TS U3076 ( .A0(n4343), .A1(n3037), .B0(n4092), .B1(n3882), .Y(n1374)
         );
  AOI222XLTS U3077 ( .A0(n4439), .A1(n3218), .B0(n486), .B1(n3203), .C0(n4248), 
        .C1(n3148), .Y(n1375) );
  AOI22X1TS U3078 ( .A0(n4340), .A1(n3037), .B0(n4090), .B1(n3882), .Y(n1372)
         );
  AOI222XLTS U3079 ( .A0(n4436), .A1(n3218), .B0(n488), .B1(n3199), .C0(n4245), 
        .C1(n3148), .Y(n1373) );
  AOI22X1TS U3080 ( .A0(n4337), .A1(n3037), .B0(n4088), .B1(n3882), .Y(n1370)
         );
  AOI222XLTS U3081 ( .A0(n4433), .A1(n3218), .B0(n490), .B1(n3202), .C0(n4242), 
        .C1(n3147), .Y(n1371) );
  AOI22X1TS U3082 ( .A0(n4334), .A1(n3028), .B0(n4086), .B1(n3882), .Y(n1368)
         );
  AOI222XLTS U3083 ( .A0(n4430), .A1(n3217), .B0(n492), .B1(n3201), .C0(n4239), 
        .C1(n3147), .Y(n1369) );
  AOI22X1TS U3084 ( .A0(n4331), .A1(n3028), .B0(n4084), .B1(n3881), .Y(n1366)
         );
  AOI222XLTS U3085 ( .A0(n4427), .A1(n3217), .B0(n494), .B1(n3211), .C0(n4236), 
        .C1(n3147), .Y(n1367) );
  AOI22X1TS U3086 ( .A0(n4328), .A1(n3028), .B0(n4082), .B1(n3881), .Y(n1364)
         );
  AOI222XLTS U3087 ( .A0(n4424), .A1(n3217), .B0(n496), .B1(n3203), .C0(n4233), 
        .C1(n3143), .Y(n1365) );
  AOI22X1TS U3088 ( .A0(n4325), .A1(n3028), .B0(n4080), .B1(n3881), .Y(n1362)
         );
  AOI222XLTS U3089 ( .A0(n4421), .A1(n3217), .B0(n498), .B1(n3208), .C0(n4230), 
        .C1(n3143), .Y(n1363) );
  AOI22X1TS U3090 ( .A0(n4319), .A1(n3044), .B0(n4075), .B1(n3880), .Y(n1358)
         );
  AOI222XLTS U3091 ( .A0(n4415), .A1(n3219), .B0(n502), .B1(n3211), .C0(n4224), 
        .C1(n3143), .Y(n1359) );
  AOI22X1TS U3092 ( .A0(n4313), .A1(n3112), .B0(n4072), .B1(n3880), .Y(n1354)
         );
  AOI222XLTS U3093 ( .A0(n4409), .A1(n3216), .B0(n451), .B1(n3212), .C0(n4218), 
        .C1(n3140), .Y(n1355) );
  AOI22X1TS U3094 ( .A0(n4310), .A1(n3114), .B0(n4070), .B1(n3880), .Y(n1352)
         );
  AOI222XLTS U3095 ( .A0(n4406), .A1(n3216), .B0(n506), .B1(n1248), .C0(n4215), 
        .C1(n3147), .Y(n1353) );
  AOI22X1TS U3096 ( .A0(n4304), .A1(n1250), .B0(n4066), .B1(n3879), .Y(n1348)
         );
  AOI222XLTS U3097 ( .A0(n4400), .A1(n3215), .B0(n453), .B1(n3204), .C0(n4209), 
        .C1(n3140), .Y(n1349) );
  AOI22X1TS U3098 ( .A0(n4301), .A1(n3114), .B0(n4064), .B1(n3879), .Y(n1346)
         );
  AOI222XLTS U3099 ( .A0(n4397), .A1(n3215), .B0(n510), .B1(n3208), .C0(n4206), 
        .C1(n3139), .Y(n1347) );
  AOI22X1TS U3100 ( .A0(n4295), .A1(n3027), .B0(n4059), .B1(n3878), .Y(n1342)
         );
  AOI222XLTS U3101 ( .A0(n4391), .A1(n3214), .B0(n514), .B1(n3204), .C0(n4200), 
        .C1(n3139), .Y(n1343) );
  AOI22X1TS U3102 ( .A0(n4292), .A1(n3027), .B0(n4058), .B1(n3878), .Y(n1340)
         );
  AOI222XLTS U3103 ( .A0(n4388), .A1(n3214), .B0(n513), .B1(n3203), .C0(n4197), 
        .C1(n3139), .Y(n1341) );
  AOI22X1TS U3104 ( .A0(n4289), .A1(n3504), .B0(n4119), .B1(n3776), .Y(n1658)
         );
  AOI222XLTS U3105 ( .A0(n4481), .A1(n3548), .B0(n458), .B1(n3529), .C0(n4386), 
        .C1(n3521), .Y(n1659) );
  AOI22X1TS U3106 ( .A0(n4244), .A1(n3500), .B0(n4090), .B1(n3771), .Y(n1628)
         );
  AOI222XLTS U3107 ( .A0(n4436), .A1(n3555), .B0(n489), .B1(n3536), .C0(n4341), 
        .C1(n3518), .Y(n1629) );
  AOI22X1TS U3108 ( .A0(n4241), .A1(n3500), .B0(n4088), .B1(n3771), .Y(n1626)
         );
  AOI222XLTS U3109 ( .A0(n4433), .A1(n3555), .B0(n491), .B1(n3539), .C0(n4338), 
        .C1(n3517), .Y(n1627) );
  AOI22X1TS U3110 ( .A0(n4229), .A1(n3499), .B0(n4080), .B1(n3770), .Y(n1618)
         );
  AOI222XLTS U3111 ( .A0(n4421), .A1(n3555), .B0(n499), .B1(n3531), .C0(n4326), 
        .C1(n3516), .Y(n1619) );
  AOI22X1TS U3112 ( .A0(n4199), .A1(n3496), .B0(n4059), .B1(n3767), .Y(n1598)
         );
  AOI222XLTS U3113 ( .A0(n4391), .A1(n3559), .B0(n515), .B1(n3532), .C0(n4296), 
        .C1(n3514), .Y(n1599) );
  AOI22X1TS U3114 ( .A0(n3990), .A1(n3510), .B0(n4043), .B1(n3779), .Y(n1928)
         );
  AOI222XLTS U3115 ( .A0(n4169), .A1(n3549), .B0(n3533), .B1(n122), .C0(n3949), 
        .C1(n3513), .Y(n1929) );
  AOI22X1TS U3116 ( .A0(n3984), .A1(n3511), .B0(n4039), .B1(n3778), .Y(n1924)
         );
  AOI222XLTS U3117 ( .A0(n4163), .A1(n3549), .B0(n3535), .B1(n112), .C0(n3943), 
        .C1(n3528), .Y(n1925) );
  AOI22X1TS U3118 ( .A0(n3981), .A1(n1186), .B0(n4038), .B1(n3775), .Y(n1922)
         );
  AOI222XLTS U3119 ( .A0(n4160), .A1(n3549), .B0(n3535), .B1(n107), .C0(n3940), 
        .C1(n3522), .Y(n1923) );
  AOI22X1TS U3120 ( .A0(n3978), .A1(n3511), .B0(n4036), .B1(n3776), .Y(n1920)
         );
  AOI222XLTS U3121 ( .A0(n4157), .A1(n3548), .B0(n3535), .B1(n102), .C0(n3937), 
        .C1(n3523), .Y(n1921) );
  AOI22X1TS U3122 ( .A0(n3975), .A1(n3511), .B0(n4033), .B1(n3774), .Y(n1918)
         );
  AOI222XLTS U3123 ( .A0(n4154), .A1(n3548), .B0(n3534), .B1(n33), .C0(n3934), 
        .C1(n3525), .Y(n1919) );
  AOI22X1TS U3124 ( .A0(n4286), .A1(n3507), .B0(n4118), .B1(n3777), .Y(n1656)
         );
  AOI222XLTS U3125 ( .A0(n4478), .A1(n3548), .B0(n461), .B1(n3536), .C0(n4383), 
        .C1(n3521), .Y(n1657) );
  AOI22X1TS U3126 ( .A0(n4283), .A1(n3508), .B0(n4116), .B1(n3777), .Y(n1654)
         );
  AOI222XLTS U3127 ( .A0(n4475), .A1(n3547), .B0(n463), .B1(n3529), .C0(n4380), 
        .C1(n3521), .Y(n1655) );
  AOI22X1TS U3128 ( .A0(n4280), .A1(n3508), .B0(n4114), .B1(n3779), .Y(n1652)
         );
  AOI222XLTS U3129 ( .A0(n4472), .A1(n3547), .B0(n465), .B1(n3541), .C0(n4377), 
        .C1(n3521), .Y(n1653) );
  AOI22X1TS U3130 ( .A0(n4277), .A1(n3504), .B0(n4111), .B1(n3777), .Y(n1650)
         );
  AOI222XLTS U3131 ( .A0(n4469), .A1(n3547), .B0(n467), .B1(n3541), .C0(n4374), 
        .C1(n3520), .Y(n1651) );
  AOI22X1TS U3132 ( .A0(n4274), .A1(n3506), .B0(n4110), .B1(n3775), .Y(n1648)
         );
  AOI222XLTS U3133 ( .A0(n4466), .A1(n3547), .B0(n469), .B1(n3540), .C0(n4371), 
        .C1(n3520), .Y(n1649) );
  AOI22X1TS U3134 ( .A0(n4271), .A1(n3505), .B0(n4108), .B1(n3773), .Y(n1646)
         );
  AOI222XLTS U3135 ( .A0(n4463), .A1(n3546), .B0(n471), .B1(n3540), .C0(n4368), 
        .C1(n3520), .Y(n1647) );
  AOI22X1TS U3136 ( .A0(n4268), .A1(n3505), .B0(n4106), .B1(n3773), .Y(n1644)
         );
  AOI222XLTS U3137 ( .A0(n4460), .A1(n3546), .B0(n473), .B1(n3529), .C0(n4365), 
        .C1(n3520), .Y(n1645) );
  AOI22X1TS U3138 ( .A0(n4265), .A1(n3506), .B0(n4104), .B1(n3773), .Y(n1642)
         );
  AOI222XLTS U3139 ( .A0(n4457), .A1(n3546), .B0(n475), .B1(n3539), .C0(n4362), 
        .C1(n3519), .Y(n1643) );
  AOI22X1TS U3140 ( .A0(n4262), .A1(n3507), .B0(n4102), .B1(n3773), .Y(n1640)
         );
  AOI222XLTS U3141 ( .A0(n4454), .A1(n3546), .B0(n477), .B1(n3539), .C0(n4359), 
        .C1(n3519), .Y(n1641) );
  AOI22X1TS U3142 ( .A0(n4259), .A1(n3505), .B0(n4100), .B1(n3772), .Y(n1638)
         );
  AOI222XLTS U3143 ( .A0(n4451), .A1(n3545), .B0(n479), .B1(n3529), .C0(n4356), 
        .C1(n3519), .Y(n1639) );
  AOI22X1TS U3144 ( .A0(n4256), .A1(n3504), .B0(n4098), .B1(n3772), .Y(n1636)
         );
  AOI222XLTS U3145 ( .A0(n4448), .A1(n3545), .B0(n481), .B1(n3540), .C0(n4353), 
        .C1(n3519), .Y(n1637) );
  AOI22X1TS U3146 ( .A0(n4253), .A1(n3505), .B0(n4096), .B1(n3772), .Y(n1634)
         );
  AOI222XLTS U3147 ( .A0(n4445), .A1(n3545), .B0(n483), .B1(n3537), .C0(n4350), 
        .C1(n3518), .Y(n1635) );
  AOI22X1TS U3148 ( .A0(n4250), .A1(n3500), .B0(n4094), .B1(n3772), .Y(n1632)
         );
  AOI222XLTS U3149 ( .A0(n4442), .A1(n3556), .B0(n485), .B1(n3538), .C0(n4347), 
        .C1(n3518), .Y(n1633) );
  AOI22X1TS U3150 ( .A0(n4247), .A1(n3500), .B0(n4092), .B1(n3771), .Y(n1630)
         );
  AOI222XLTS U3151 ( .A0(n4439), .A1(n3557), .B0(n487), .B1(n3539), .C0(n4344), 
        .C1(n3518), .Y(n1631) );
  AOI22X1TS U3152 ( .A0(n4238), .A1(n3499), .B0(n4086), .B1(n3771), .Y(n1624)
         );
  AOI222XLTS U3153 ( .A0(n4430), .A1(n3554), .B0(n493), .B1(n3537), .C0(n4335), 
        .C1(n3517), .Y(n1625) );
  AOI22X1TS U3154 ( .A0(n4235), .A1(n3499), .B0(n4084), .B1(n3770), .Y(n1622)
         );
  AOI222XLTS U3155 ( .A0(n4427), .A1(n3556), .B0(n495), .B1(n3530), .C0(n4332), 
        .C1(n3517), .Y(n1623) );
  AOI22X1TS U3156 ( .A0(n4232), .A1(n3499), .B0(n4082), .B1(n3770), .Y(n1620)
         );
  AOI222XLTS U3157 ( .A0(n4424), .A1(n3557), .B0(n497), .B1(n3542), .C0(n4329), 
        .C1(n3516), .Y(n1621) );
  AOI22X1TS U3158 ( .A0(n4226), .A1(n3498), .B0(n4078), .B1(n3770), .Y(n1616)
         );
  AOI222XLTS U3159 ( .A0(n4418), .A1(n3556), .B0(n501), .B1(n3531), .C0(n4323), 
        .C1(n3516), .Y(n1617) );
  AOI22X1TS U3160 ( .A0(n4223), .A1(n3504), .B0(n4075), .B1(n3769), .Y(n1614)
         );
  AOI222XLTS U3161 ( .A0(n4415), .A1(n3545), .B0(n503), .B1(n3530), .C0(n4320), 
        .C1(n3516), .Y(n1615) );
  AOI22X1TS U3162 ( .A0(n4220), .A1(n3498), .B0(n4074), .B1(n3769), .Y(n1612)
         );
  AOI222XLTS U3163 ( .A0(n4412), .A1(n3553), .B0(n505), .B1(n3531), .C0(n4317), 
        .C1(n3515), .Y(n1613) );
  AOI22X1TS U3164 ( .A0(n4217), .A1(n3498), .B0(n4072), .B1(n3769), .Y(n1610)
         );
  AOI222XLTS U3165 ( .A0(n4409), .A1(n3554), .B0(n452), .B1(n3530), .C0(n4314), 
        .C1(n3515), .Y(n1611) );
  AOI22X1TS U3166 ( .A0(n4214), .A1(n3498), .B0(n4070), .B1(n3769), .Y(n1608)
         );
  AOI222XLTS U3167 ( .A0(n4406), .A1(n3553), .B0(n507), .B1(n3530), .C0(n4311), 
        .C1(n3517), .Y(n1609) );
  AOI22X1TS U3168 ( .A0(n4211), .A1(n3497), .B0(n4067), .B1(n3768), .Y(n1606)
         );
  AOI222XLTS U3169 ( .A0(n4403), .A1(n3544), .B0(n509), .B1(n3532), .C0(n4308), 
        .C1(n3515), .Y(n1607) );
  AOI22X1TS U3170 ( .A0(n4208), .A1(n3497), .B0(n4066), .B1(n3768), .Y(n1604)
         );
  AOI222XLTS U3171 ( .A0(n4400), .A1(n3544), .B0(n454), .B1(n3532), .C0(n4305), 
        .C1(n3515), .Y(n1605) );
  AOI22X1TS U3172 ( .A0(n4205), .A1(n3497), .B0(n4064), .B1(n3768), .Y(n1602)
         );
  AOI222XLTS U3173 ( .A0(n4397), .A1(n3544), .B0(n511), .B1(n3531), .C0(n4302), 
        .C1(n3514), .Y(n1603) );
  AOI22X1TS U3174 ( .A0(n4202), .A1(n3497), .B0(n4062), .B1(n3768), .Y(n1600)
         );
  AOI222XLTS U3175 ( .A0(n4394), .A1(n3544), .B0(n456), .B1(n3532), .C0(n4299), 
        .C1(n3514), .Y(n1601) );
  AOI22X1TS U3176 ( .A0(n4385), .A1(n3403), .B0(n4481), .B1(n3392), .Y(n1530)
         );
  AOI222XLTS U3177 ( .A0(n457), .A1(n3843), .B0(n4120), .B1(n3865), .C0(n68), 
        .C1(n3856), .Y(n1531) );
  AOI22X1TS U3178 ( .A0(n4382), .A1(n3403), .B0(n4478), .B1(n3392), .Y(n1528)
         );
  AOI222XLTS U3179 ( .A0(n460), .A1(n3849), .B0(n4117), .B1(n3865), .C0(n69), 
        .C1(n3856), .Y(n1529) );
  AOI22X1TS U3180 ( .A0(n4379), .A1(n3402), .B0(n4475), .B1(n3390), .Y(n1526)
         );
  AOI222XLTS U3181 ( .A0(n462), .A1(n3848), .B0(n4115), .B1(n3866), .C0(n70), 
        .C1(n3856), .Y(n1527) );
  AOI22X1TS U3182 ( .A0(n4376), .A1(n3402), .B0(n4472), .B1(n3390), .Y(n1524)
         );
  AOI222XLTS U3183 ( .A0(n464), .A1(n774), .B0(n4113), .B1(n3866), .C0(n71), 
        .C1(n3856), .Y(n1525) );
  AOI22X1TS U3184 ( .A0(n4373), .A1(n3402), .B0(n4469), .B1(n3391), .Y(n1522)
         );
  AOI222XLTS U3185 ( .A0(n466), .A1(n3846), .B0(n4112), .B1(n3866), .C0(n72), 
        .C1(n3855), .Y(n1523) );
  AOI22X1TS U3186 ( .A0(n4370), .A1(n3402), .B0(n4466), .B1(n3393), .Y(n1520)
         );
  AOI222XLTS U3187 ( .A0(n468), .A1(n3840), .B0(n4109), .B1(n3866), .C0(n73), 
        .C1(n3855), .Y(n1521) );
  AOI22X1TS U3188 ( .A0(n4364), .A1(n3401), .B0(n4460), .B1(n3386), .Y(n1516)
         );
  AOI222XLTS U3189 ( .A0(n472), .A1(n3846), .B0(n4105), .B1(n3867), .C0(n74), 
        .C1(n3855), .Y(n1517) );
  AOI22X1TS U3190 ( .A0(n4358), .A1(n3401), .B0(n4454), .B1(n3386), .Y(n1512)
         );
  AOI222XLTS U3191 ( .A0(n476), .A1(n3844), .B0(n4101), .B1(n3867), .C0(n75), 
        .C1(n3854), .Y(n1513) );
  AOI22X1TS U3192 ( .A0(n4355), .A1(n3400), .B0(n4451), .B1(n3385), .Y(n1510)
         );
  AOI222XLTS U3193 ( .A0(n478), .A1(n3838), .B0(n4099), .B1(n3868), .C0(n76), 
        .C1(n3854), .Y(n1511) );
  AOI22X1TS U3194 ( .A0(n4349), .A1(n3400), .B0(n4445), .B1(n3385), .Y(n1506)
         );
  AOI222XLTS U3195 ( .A0(n482), .A1(n3838), .B0(n4095), .B1(n3868), .C0(n77), 
        .C1(n3853), .Y(n1507) );
  AOI22X1TS U3196 ( .A0(n4343), .A1(n3411), .B0(n4439), .B1(n3384), .Y(n1502)
         );
  AOI222XLTS U3197 ( .A0(n486), .A1(n3838), .B0(n4091), .B1(n3869), .C0(n78), 
        .C1(n3853), .Y(n1503) );
  AOI22X1TS U3198 ( .A0(n4340), .A1(n3410), .B0(n4436), .B1(n3384), .Y(n1500)
         );
  AOI222XLTS U3199 ( .A0(n488), .A1(n3839), .B0(n4089), .B1(n3869), .C0(n79), 
        .C1(n3853), .Y(n1501) );
  AOI22X1TS U3200 ( .A0(n4334), .A1(n3412), .B0(n4430), .B1(n3383), .Y(n1496)
         );
  AOI222XLTS U3201 ( .A0(n492), .A1(n3839), .B0(n4085), .B1(n3869), .C0(n80), 
        .C1(n3852), .Y(n1497) );
  AOI22X1TS U3202 ( .A0(n4328), .A1(n1216), .B0(n4424), .B1(n3383), .Y(n1492)
         );
  AOI222XLTS U3203 ( .A0(n496), .A1(n3840), .B0(n4081), .B1(n3870), .C0(n81), 
        .C1(n3858), .Y(n1493) );
  AOI22X1TS U3204 ( .A0(n4325), .A1(n3410), .B0(n4421), .B1(n3383), .Y(n1490)
         );
  AOI222XLTS U3205 ( .A0(n498), .A1(n3840), .B0(n4079), .B1(n3870), .C0(n82), 
        .C1(n3858), .Y(n1491) );
  AOI22X1TS U3206 ( .A0(n4322), .A1(n3399), .B0(n4418), .B1(n3382), .Y(n1488)
         );
  AOI222XLTS U3207 ( .A0(n500), .A1(n3843), .B0(n4077), .B1(n3870), .C0(n83), 
        .C1(n3862), .Y(n1489) );
  AOI22X1TS U3208 ( .A0(n4319), .A1(n3400), .B0(n4415), .B1(n3385), .Y(n1486)
         );
  AOI222XLTS U3209 ( .A0(n502), .A1(n3841), .B0(n4076), .B1(n3872), .C0(n84), 
        .C1(n3863), .Y(n1487) );
  AOI22X1TS U3210 ( .A0(n4316), .A1(n3399), .B0(n4412), .B1(n3382), .Y(n1484)
         );
  AOI222XLTS U3211 ( .A0(n504), .A1(n3841), .B0(n4073), .B1(n771), .C0(n85), 
        .C1(n3851), .Y(n1485) );
  AOI22X1TS U3212 ( .A0(n4310), .A1(n3399), .B0(n4406), .B1(n3382), .Y(n1480)
         );
  AOI222XLTS U3213 ( .A0(n506), .A1(n3842), .B0(n4069), .B1(n771), .C0(n86), 
        .C1(n3851), .Y(n1481) );
  AOI22X1TS U3214 ( .A0(n4301), .A1(n3398), .B0(n4397), .B1(n3381), .Y(n1474)
         );
  AOI222XLTS U3215 ( .A0(n510), .A1(n3843), .B0(n4063), .B1(n3871), .C0(n87), 
        .C1(n3851), .Y(n1475) );
  AOI22X1TS U3216 ( .A0(n4295), .A1(n3397), .B0(n4391), .B1(n3380), .Y(n1470)
         );
  AOI222XLTS U3217 ( .A0(n514), .A1(n3842), .B0(n4060), .B1(n3873), .C0(n88), 
        .C1(n3850), .Y(n1471) );
  AOI22X1TS U3218 ( .A0(n4292), .A1(n3397), .B0(n4388), .B1(n3380), .Y(n1468)
         );
  AOI222XLTS U3219 ( .A0(n512), .A1(n3843), .B0(n4057), .B1(n15), .C0(n89), 
        .C1(n3850), .Y(n1469) );
  AOI22X1TS U3220 ( .A0(n4367), .A1(n3401), .B0(n4463), .B1(n3386), .Y(n1518)
         );
  AOI222XLTS U3221 ( .A0(n470), .A1(n3847), .B0(n4107), .B1(n3867), .C0(n93), 
        .C1(n3855), .Y(n1519) );
  AOI22X1TS U3222 ( .A0(n4361), .A1(n3401), .B0(n4457), .B1(n3386), .Y(n1514)
         );
  AOI222XLTS U3223 ( .A0(n474), .A1(n774), .B0(n4103), .B1(n3867), .C0(n94), 
        .C1(n3854), .Y(n1515) );
  AOI22X1TS U3224 ( .A0(n4352), .A1(n3400), .B0(n4448), .B1(n3385), .Y(n1508)
         );
  AOI222XLTS U3225 ( .A0(n480), .A1(n3838), .B0(n4097), .B1(n3868), .C0(n95), 
        .C1(n3854), .Y(n1509) );
  AOI22X1TS U3226 ( .A0(n4346), .A1(n3409), .B0(n4442), .B1(n3384), .Y(n1504)
         );
  AOI222XLTS U3227 ( .A0(n484), .A1(n3839), .B0(n4093), .B1(n3868), .C0(n96), 
        .C1(n3853), .Y(n1505) );
  AOI22X1TS U3228 ( .A0(n4337), .A1(n3409), .B0(n4433), .B1(n3384), .Y(n1498)
         );
  AOI222XLTS U3229 ( .A0(n490), .A1(n3840), .B0(n4087), .B1(n3869), .C0(n97), 
        .C1(n3852), .Y(n1499) );
  AOI22X1TS U3230 ( .A0(n4331), .A1(n1216), .B0(n4427), .B1(n3383), .Y(n1494)
         );
  AOI222XLTS U3231 ( .A0(n494), .A1(n3839), .B0(n4083), .B1(n3870), .C0(n98), 
        .C1(n3852), .Y(n1495) );
  AOI22X1TS U3232 ( .A0(n4307), .A1(n3398), .B0(n4403), .B1(n3381), .Y(n1478)
         );
  AOI222XLTS U3233 ( .A0(n508), .A1(n3841), .B0(n4068), .B1(n3871), .C0(n99), 
        .C1(n3851), .Y(n1479) );
  AOI22X1TS U3234 ( .A0(n4304), .A1(n3398), .B0(n4400), .B1(n3381), .Y(n1476)
         );
  AOI222XLTS U3235 ( .A0(n453), .A1(n3842), .B0(n4065), .B1(n3871), .C0(n3861), 
        .C1(n679), .Y(n1477) );
  AOI22X1TS U3236 ( .A0(n4298), .A1(n3398), .B0(n4394), .B1(n3381), .Y(n1472)
         );
  AOI222XLTS U3237 ( .A0(n455), .A1(n3842), .B0(n4061), .B1(n3871), .C0(n3859), 
        .C1(n678), .Y(n1473) );
  AOI22X1TS U3238 ( .A0(n4313), .A1(n3399), .B0(n4409), .B1(n3382), .Y(n1482)
         );
  AOI222XLTS U3239 ( .A0(n451), .A1(n3841), .B0(n4071), .B1(n3872), .C0(n773), 
        .C1(n661), .Y(n1483) );
  AOI22X1TS U3240 ( .A0(n3458), .A1(n121), .B0(n3948), .B1(n3437), .Y(n1951)
         );
  AOI222XLTS U3241 ( .A0(n3123), .A1(n3792), .B0(n4170), .B1(n3463), .C0(n4044), .C1(n3806), .Y(n1952) );
  AOI22X1TS U3242 ( .A0(n3454), .A1(n116), .B0(n3945), .B1(n3437), .Y(n1949)
         );
  AOI222XLTS U3243 ( .A0(n3125), .A1(n3787), .B0(n4167), .B1(n3468), .C0(
        destinationAddressIn_NORTH[4]), .C1(n3805), .Y(n1950) );
  AOI22X1TS U3244 ( .A0(n3455), .A1(n111), .B0(n3942), .B1(n3437), .Y(n1947)
         );
  AOI222XLTS U3245 ( .A0(n3127), .A1(n3786), .B0(n4164), .B1(n3468), .C0(n4040), .C1(n3803), .Y(n1948) );
  AOI22X1TS U3246 ( .A0(n3456), .A1(n106), .B0(n3939), .B1(n3437), .Y(n1945)
         );
  AOI222XLTS U3247 ( .A0(n3130), .A1(n3786), .B0(n4161), .B1(n3468), .C0(
        destinationAddressIn_NORTH[2]), .C1(n3804), .Y(n1946) );
  AOI22X1TS U3248 ( .A0(n3447), .A1(n101), .B0(n3936), .B1(n3436), .Y(n1943)
         );
  AOI222XLTS U3249 ( .A0(n3132), .A1(n3786), .B0(n4158), .B1(n3467), .C0(
        destinationAddressIn_NORTH[1]), .C1(n3808), .Y(n1944) );
  AOI22X1TS U3250 ( .A0(n3458), .A1(n32), .B0(n3933), .B1(n3436), .Y(n1941) );
  AOI222XLTS U3251 ( .A0(n3134), .A1(n3786), .B0(n4155), .B1(n3467), .C0(n4034), .C1(n3806), .Y(n1942) );
  AOI22X1TS U3252 ( .A0(n460), .A1(n3457), .B0(n4382), .B1(n3436), .Y(n1592)
         );
  AOI222XLTS U3253 ( .A0(n3040), .A1(n3785), .B0(n4479), .B1(n3467), .C0(
        dataIn_NORTH[30]), .C1(n3808), .Y(n1593) );
  AOI22X1TS U3254 ( .A0(n464), .A1(n3457), .B0(n4376), .B1(n3435), .Y(n1588)
         );
  AOI222XLTS U3255 ( .A0(n3045), .A1(n3785), .B0(n4473), .B1(n3471), .C0(
        dataIn_NORTH[28]), .C1(n3802), .Y(n1589) );
  AOI22X1TS U3256 ( .A0(n466), .A1(n3457), .B0(n4373), .B1(n3435), .Y(n1586)
         );
  AOI222XLTS U3257 ( .A0(n3048), .A1(n3784), .B0(n4470), .B1(n3477), .C0(n4112), .C1(n3802), .Y(n1587) );
  AOI22X1TS U3258 ( .A0(n468), .A1(n3450), .B0(n4370), .B1(n3435), .Y(n1584)
         );
  AOI222XLTS U3259 ( .A0(n3051), .A1(n3784), .B0(n4467), .B1(n3474), .C0(
        dataIn_NORTH[26]), .C1(n3802), .Y(n1585) );
  AOI22X1TS U3260 ( .A0(n470), .A1(n3457), .B0(n4367), .B1(n3434), .Y(n1582)
         );
  AOI222XLTS U3261 ( .A0(n3053), .A1(n3784), .B0(n4464), .B1(n3471), .C0(
        dataIn_NORTH[25]), .C1(n3801), .Y(n1583) );
  AOI22X1TS U3262 ( .A0(n472), .A1(n3454), .B0(n4364), .B1(n3434), .Y(n1580)
         );
  AOI222XLTS U3263 ( .A0(n3055), .A1(n3784), .B0(n4461), .B1(n3471), .C0(
        dataIn_NORTH[24]), .C1(n3801), .Y(n1581) );
  AOI22X1TS U3264 ( .A0(n474), .A1(n3455), .B0(n4361), .B1(n3434), .Y(n1578)
         );
  AOI222XLTS U3265 ( .A0(n3058), .A1(n3783), .B0(n4458), .B1(n3473), .C0(
        dataIn_NORTH[23]), .C1(n3801), .Y(n1579) );
  AOI22X1TS U3266 ( .A0(n484), .A1(n3449), .B0(n4346), .B1(n3444), .Y(n1568)
         );
  AOI222XLTS U3267 ( .A0(n3071), .A1(n3782), .B0(n4443), .B1(n3472), .C0(
        dataIn_NORTH[18]), .C1(n3800), .Y(n1569) );
  AOI22X1TS U3268 ( .A0(n494), .A1(n3449), .B0(n4331), .B1(n3442), .Y(n1558)
         );
  AOI222XLTS U3269 ( .A0(n3084), .A1(n3791), .B0(n4428), .B1(n3466), .C0(
        dataIn_NORTH[13]), .C1(n3799), .Y(n1559) );
  AOI22X1TS U3270 ( .A0(n502), .A1(n3451), .B0(n4319), .B1(n3433), .Y(n1550)
         );
  AOI222XLTS U3271 ( .A0(n3095), .A1(n3791), .B0(n4416), .B1(n3465), .C0(n4076), .C1(n3798), .Y(n1551) );
  AOI22X1TS U3272 ( .A0(n451), .A1(n3451), .B0(n4313), .B1(n3432), .Y(n1546)
         );
  AOI222XLTS U3273 ( .A0(n3099), .A1(n3788), .B0(n4410), .B1(n3465), .C0(
        dataIn_NORTH[7]), .C1(n3798), .Y(n1547) );
  AOI22X1TS U3274 ( .A0(n508), .A1(n3451), .B0(n4307), .B1(n3431), .Y(n1542)
         );
  AOI222XLTS U3275 ( .A0(n3106), .A1(n3789), .B0(n4404), .B1(n3464), .C0(n4068), .C1(n3797), .Y(n1543) );
  AOI22X1TS U3276 ( .A0(n453), .A1(n3452), .B0(n4304), .B1(n3431), .Y(n1540)
         );
  AOI222XLTS U3277 ( .A0(n3108), .A1(n3781), .B0(n4401), .B1(n3464), .C0(
        dataIn_NORTH[4]), .C1(n3797), .Y(n1541) );
  AOI22X1TS U3278 ( .A0(n455), .A1(n3452), .B0(n4298), .B1(n3431), .Y(n1536)
         );
  AOI222XLTS U3279 ( .A0(n3115), .A1(n3781), .B0(n4395), .B1(n3464), .C0(
        dataIn_NORTH[2]), .C1(n3797), .Y(n1537) );
  AOI22X1TS U3280 ( .A0(n457), .A1(n3453), .B0(n4385), .B1(n3436), .Y(n1594)
         );
  AOI222XLTS U3281 ( .A0(n3036), .A1(n3785), .B0(n4482), .B1(n3467), .C0(n4120), .C1(n3807), .Y(n1595) );
  AOI22X1TS U3282 ( .A0(n462), .A1(n3458), .B0(n4379), .B1(n3435), .Y(n1590)
         );
  AOI222XLTS U3283 ( .A0(n3042), .A1(n3785), .B0(n4476), .B1(n3470), .C0(
        dataIn_NORTH[29]), .C1(n3802), .Y(n1591) );
  AOI22X1TS U3284 ( .A0(n476), .A1(n3456), .B0(n4358), .B1(n3434), .Y(n1576)
         );
  AOI222XLTS U3285 ( .A0(n3061), .A1(n3783), .B0(n4455), .B1(n3476), .C0(
        dataIn_NORTH[22]), .C1(n3801), .Y(n1577) );
  AOI22X1TS U3286 ( .A0(n478), .A1(n3448), .B0(n4355), .B1(n3433), .Y(n1574)
         );
  AOI222XLTS U3287 ( .A0(n3063), .A1(n3783), .B0(n4452), .B1(n3472), .C0(
        dataIn_NORTH[21]), .C1(n3800), .Y(n1575) );
  AOI22X1TS U3288 ( .A0(n480), .A1(n3448), .B0(n4352), .B1(n3433), .Y(n1572)
         );
  AOI222XLTS U3289 ( .A0(n3066), .A1(n3783), .B0(n4449), .B1(n3472), .C0(
        dataIn_NORTH[20]), .C1(n3800), .Y(n1573) );
  AOI22X1TS U3290 ( .A0(n482), .A1(n3448), .B0(n4349), .B1(n3433), .Y(n1570)
         );
  AOI222XLTS U3291 ( .A0(n3068), .A1(n3782), .B0(n4446), .B1(n3474), .C0(
        dataIn_NORTH[19]), .C1(n3800), .Y(n1571) );
  AOI22X1TS U3292 ( .A0(n488), .A1(n3449), .B0(n4340), .B1(n3440), .Y(n1564)
         );
  AOI222XLTS U3293 ( .A0(n3076), .A1(n3782), .B0(n4437), .B1(n3472), .C0(
        dataIn_NORTH[16]), .C1(n3803), .Y(n1565) );
  AOI22X1TS U3294 ( .A0(n496), .A1(n3450), .B0(n4328), .B1(n3443), .Y(n1556)
         );
  AOI222XLTS U3295 ( .A0(n3088), .A1(n3789), .B0(n4425), .B1(n3466), .C0(
        dataIn_NORTH[12]), .C1(n3799), .Y(n1557) );
  AOI22X1TS U3296 ( .A0(n498), .A1(n3450), .B0(n4325), .B1(n3440), .Y(n1554)
         );
  AOI222XLTS U3297 ( .A0(n3090), .A1(n780), .B0(n4422), .B1(n3466), .C0(
        dataIn_NORTH[11]), .C1(n3799), .Y(n1555) );
  AOI22X1TS U3298 ( .A0(n500), .A1(n3453), .B0(n4322), .B1(n3432), .Y(n1552)
         );
  AOI222XLTS U3299 ( .A0(n3093), .A1(n780), .B0(n4419), .B1(n3465), .C0(
        dataIn_NORTH[10]), .C1(n3799), .Y(n1553) );
  AOI22X1TS U3300 ( .A0(n504), .A1(n3451), .B0(n4316), .B1(n3432), .Y(n1548)
         );
  AOI222XLTS U3301 ( .A0(n3097), .A1(n3794), .B0(n4413), .B1(n3465), .C0(
        dataIn_NORTH[8]), .C1(n3798), .Y(n1549) );
  AOI22X1TS U3302 ( .A0(n506), .A1(n3452), .B0(n4310), .B1(n3432), .Y(n1544)
         );
  AOI222XLTS U3303 ( .A0(n3104), .A1(n3791), .B0(n4407), .B1(n3470), .C0(
        dataIn_NORTH[6]), .C1(n3798), .Y(n1545) );
  AOI22X1TS U3304 ( .A0(n514), .A1(n3452), .B0(n4295), .B1(n3444), .Y(n1534)
         );
  AOI222XLTS U3305 ( .A0(n3117), .A1(n3781), .B0(n4392), .B1(n3463), .C0(n4060), .C1(n3796), .Y(n1535) );
  AOI22X1TS U3306 ( .A0(n512), .A1(n3453), .B0(n4292), .B1(n3441), .Y(n1532)
         );
  AOI222XLTS U3307 ( .A0(n3120), .A1(n3780), .B0(n4389), .B1(n3463), .C0(
        dataIn_NORTH[0]), .C1(n3796), .Y(n1533) );
  AOI22X1TS U3308 ( .A0(n486), .A1(n3448), .B0(n4343), .B1(n3442), .Y(n1566)
         );
  AOI222XLTS U3309 ( .A0(n3073), .A1(n3782), .B0(n4440), .B1(n3471), .C0(
        dataIn_NORTH[17]), .C1(n3803), .Y(n1567) );
  AOI22X1TS U3310 ( .A0(n490), .A1(n3450), .B0(n4337), .B1(n3443), .Y(n1562)
         );
  AOI222XLTS U3311 ( .A0(n3078), .A1(n3790), .B0(n4434), .B1(n3473), .C0(
        dataIn_NORTH[15]), .C1(n3804), .Y(n1563) );
  AOI22X1TS U3312 ( .A0(n492), .A1(n3449), .B0(n4334), .B1(n3444), .Y(n1560)
         );
  AOI222XLTS U3313 ( .A0(n3080), .A1(n3790), .B0(n4431), .B1(n3466), .C0(
        dataIn_NORTH[14]), .C1(n3805), .Y(n1561) );
  AOI22X1TS U3314 ( .A0(n510), .A1(n3453), .B0(n4301), .B1(n3431), .Y(n1538)
         );
  AOI222XLTS U3315 ( .A0(n3111), .A1(n3781), .B0(n4398), .B1(n3464), .C0(
        dataIn_NORTH[3]), .C1(n3797), .Y(n1539) );
  AOI22X1TS U3316 ( .A0(n4391), .A1(n3609), .B0(n4059), .B1(n3756), .Y(n1663)
         );
  AOI222XLTS U3317 ( .A0(n4296), .A1(n3739), .B0(n515), .B1(n3608), .C0(n4200), 
        .C1(n3590), .Y(n1664) );
  AOI22X1TS U3318 ( .A0(n4394), .A1(n3609), .B0(n4062), .B1(n3758), .Y(n1665)
         );
  AOI222XLTS U3319 ( .A0(n4299), .A1(n3739), .B0(n456), .B1(n3608), .C0(n4203), 
        .C1(n3590), .Y(n1666) );
  AOI22X1TS U3320 ( .A0(n4397), .A1(n3609), .B0(n4064), .B1(n3758), .Y(n1667)
         );
  AOI222XLTS U3321 ( .A0(n4302), .A1(n3739), .B0(n511), .B1(n3605), .C0(n4206), 
        .C1(n3580), .Y(n1668) );
  AOI22X1TS U3322 ( .A0(n4400), .A1(n3610), .B0(n4066), .B1(n3757), .Y(n1669)
         );
  AOI222XLTS U3323 ( .A0(n4305), .A1(n3740), .B0(n454), .B1(n3607), .C0(n4209), 
        .C1(n3580), .Y(n1670) );
  AOI22X1TS U3324 ( .A0(n4403), .A1(n3610), .B0(n4067), .B1(n3758), .Y(n1671)
         );
  AOI222XLTS U3325 ( .A0(n4308), .A1(n3740), .B0(n509), .B1(n3602), .C0(n4212), 
        .C1(n3580), .Y(n1672) );
  AOI22X1TS U3326 ( .A0(n4406), .A1(n3610), .B0(n4070), .B1(n3758), .Y(n1673)
         );
  AOI222XLTS U3327 ( .A0(n4311), .A1(n3740), .B0(n507), .B1(n3606), .C0(n4215), 
        .C1(n3582), .Y(n1674) );
  AOI22X1TS U3328 ( .A0(n4409), .A1(n3610), .B0(n4072), .B1(n3763), .Y(n1675)
         );
  AOI222XLTS U3329 ( .A0(n4314), .A1(n3740), .B0(n452), .B1(n3602), .C0(n4218), 
        .C1(n3581), .Y(n1676) );
  AOI22X1TS U3330 ( .A0(n4412), .A1(n3622), .B0(n4074), .B1(n3763), .Y(n1677)
         );
  AOI222XLTS U3331 ( .A0(n4317), .A1(n3741), .B0(n505), .B1(n3604), .C0(n4221), 
        .C1(n3581), .Y(n1678) );
  AOI22X1TS U3332 ( .A0(n4415), .A1(n3620), .B0(n4075), .B1(n3757), .Y(n1679)
         );
  AOI222XLTS U3333 ( .A0(n4320), .A1(n3741), .B0(n503), .B1(n3603), .C0(n4224), 
        .C1(n3581), .Y(n1680) );
  AOI22X1TS U3334 ( .A0(n4418), .A1(n3624), .B0(n4078), .B1(n3764), .Y(n1681)
         );
  AOI222XLTS U3335 ( .A0(n4323), .A1(n3741), .B0(n501), .B1(n3606), .C0(n4227), 
        .C1(n3581), .Y(n1682) );
  AOI22X1TS U3336 ( .A0(n4421), .A1(n3623), .B0(n4080), .B1(n3757), .Y(n1683)
         );
  AOI222XLTS U3337 ( .A0(n4326), .A1(n3741), .B0(n499), .B1(n3602), .C0(n4230), 
        .C1(n3582), .Y(n1684) );
  AOI22X1TS U3338 ( .A0(n4424), .A1(n1167), .B0(n4082), .B1(n3757), .Y(n1685)
         );
  AOI222XLTS U3339 ( .A0(n4329), .A1(n3742), .B0(n497), .B1(n3602), .C0(n4233), 
        .C1(n3582), .Y(n1686) );
  AOI22X1TS U3340 ( .A0(n4427), .A1(n3624), .B0(n4084), .B1(n3756), .Y(n1687)
         );
  AOI222XLTS U3341 ( .A0(n4332), .A1(n3742), .B0(n495), .B1(n3601), .C0(n4236), 
        .C1(n3582), .Y(n1688) );
  AOI22X1TS U3342 ( .A0(n4430), .A1(n3623), .B0(n4086), .B1(n3762), .Y(n1689)
         );
  AOI222XLTS U3343 ( .A0(n4335), .A1(n3742), .B0(n493), .B1(n3601), .C0(n4239), 
        .C1(n3583), .Y(n1690) );
  AOI22X1TS U3344 ( .A0(n4433), .A1(n1167), .B0(n4088), .B1(n3754), .Y(n1691)
         );
  AOI222XLTS U3345 ( .A0(n4338), .A1(n3742), .B0(n491), .B1(n3604), .C0(n4242), 
        .C1(n3583), .Y(n1692) );
  AOI22X1TS U3346 ( .A0(n4436), .A1(n3611), .B0(n4090), .B1(n3755), .Y(n1693)
         );
  AOI222XLTS U3347 ( .A0(n4341), .A1(n3743), .B0(n489), .B1(n3601), .C0(n4245), 
        .C1(n3583), .Y(n1694) );
  AOI22X1TS U3348 ( .A0(n4439), .A1(n3611), .B0(n4092), .B1(n3752), .Y(n1695)
         );
  AOI222XLTS U3349 ( .A0(n4344), .A1(n3743), .B0(n487), .B1(n3600), .C0(n4248), 
        .C1(n3583), .Y(n1696) );
  AOI22X1TS U3350 ( .A0(n4442), .A1(n3611), .B0(n4094), .B1(n3756), .Y(n1697)
         );
  AOI222XLTS U3351 ( .A0(n4347), .A1(n3743), .B0(n485), .B1(n3601), .C0(n4251), 
        .C1(n3584), .Y(n1698) );
  AOI22X1TS U3352 ( .A0(n4445), .A1(n3611), .B0(n4096), .B1(n3754), .Y(n1699)
         );
  AOI222XLTS U3353 ( .A0(n4350), .A1(n3743), .B0(n483), .B1(n3600), .C0(n4254), 
        .C1(n3584), .Y(n1700) );
  AOI22X1TS U3354 ( .A0(n4448), .A1(n3612), .B0(n4098), .B1(n3756), .Y(n1701)
         );
  AOI222XLTS U3355 ( .A0(n4353), .A1(n3751), .B0(n481), .B1(n3600), .C0(n4257), 
        .C1(n3584), .Y(n1702) );
  AOI22X1TS U3356 ( .A0(n4451), .A1(n3612), .B0(n4100), .B1(n3755), .Y(n1703)
         );
  AOI222XLTS U3357 ( .A0(n4356), .A1(n3749), .B0(n479), .B1(n3600), .C0(n4260), 
        .C1(n3584), .Y(n1704) );
  AOI22X1TS U3358 ( .A0(n4454), .A1(n3612), .B0(n4102), .B1(n3753), .Y(n1705)
         );
  AOI222XLTS U3359 ( .A0(n4359), .A1(n3747), .B0(n477), .B1(n3599), .C0(n4263), 
        .C1(n3585), .Y(n1706) );
  AOI22X1TS U3360 ( .A0(n4457), .A1(n3612), .B0(n4104), .B1(n3755), .Y(n1707)
         );
  AOI222XLTS U3361 ( .A0(n4362), .A1(n784), .B0(n475), .B1(n3599), .C0(n4266), 
        .C1(n3585), .Y(n1708) );
  AOI22X1TS U3362 ( .A0(n4460), .A1(n3613), .B0(n4106), .B1(n3755), .Y(n1709)
         );
  AOI222XLTS U3363 ( .A0(n4365), .A1(n3751), .B0(n473), .B1(n3599), .C0(n4269), 
        .C1(n3585), .Y(n1710) );
  AOI22X1TS U3364 ( .A0(n4463), .A1(n3613), .B0(n4108), .B1(n3753), .Y(n1711)
         );
  AOI222XLTS U3365 ( .A0(n4368), .A1(n3748), .B0(n471), .B1(n3598), .C0(n4272), 
        .C1(n3585), .Y(n1712) );
  AOI22X1TS U3366 ( .A0(n4466), .A1(n3613), .B0(n4110), .B1(n3754), .Y(n1713)
         );
  AOI222XLTS U3367 ( .A0(n4371), .A1(n3747), .B0(n469), .B1(n3603), .C0(n4275), 
        .C1(n3586), .Y(n1714) );
  AOI22X1TS U3368 ( .A0(n4469), .A1(n3613), .B0(n4111), .B1(n3754), .Y(n1715)
         );
  AOI222XLTS U3369 ( .A0(n4374), .A1(n3748), .B0(n467), .B1(n3599), .C0(n4278), 
        .C1(n3586), .Y(n1716) );
  AOI22X1TS U3370 ( .A0(n4472), .A1(n3614), .B0(n4114), .B1(n3752), .Y(n1717)
         );
  AOI222XLTS U3371 ( .A0(n4377), .A1(n3744), .B0(n465), .B1(n3598), .C0(n4281), 
        .C1(n3586), .Y(n1718) );
  AOI22X1TS U3372 ( .A0(n4475), .A1(n3614), .B0(n4116), .B1(n3752), .Y(n1719)
         );
  AOI222XLTS U3373 ( .A0(n4380), .A1(n3744), .B0(n463), .B1(n3598), .C0(n4284), 
        .C1(n3586), .Y(n1720) );
  AOI22X1TS U3374 ( .A0(n4478), .A1(n3614), .B0(n4118), .B1(n3753), .Y(n1721)
         );
  AOI222XLTS U3375 ( .A0(n4383), .A1(n3744), .B0(n461), .B1(n3598), .C0(n4287), 
        .C1(n3592), .Y(n1722) );
  AOI22X1TS U3376 ( .A0(n4481), .A1(n3614), .B0(n4119), .B1(n3752), .Y(n1723)
         );
  AOI222XLTS U3377 ( .A0(n4386), .A1(n3744), .B0(n458), .B1(n3605), .C0(n4290), 
        .C1(n1169), .Y(n1724) );
  AOI22X1TS U3378 ( .A0(n3945), .A1(n3082), .B0(n4042), .B1(n3885), .Y(n2020)
         );
  AOI22X1TS U3379 ( .A0(n3267), .A1(n104), .B0(n3981), .B1(n3255), .Y(n1991)
         );
  AOI222XLTS U3380 ( .A0(n3818), .A1(n746), .B0(n4161), .B1(n3352), .C0(n4037), 
        .C1(n3832), .Y(n1992) );
  AOI22X1TS U3381 ( .A0(n460), .A1(n3268), .B0(n4286), .B1(n3254), .Y(n1464)
         );
  AOI222XLTS U3382 ( .A0(n3817), .A1(n745), .B0(n4479), .B1(n3351), .C0(n4117), 
        .C1(n3831), .Y(n1465) );
  AOI22X1TS U3383 ( .A0(n462), .A1(n3268), .B0(n4283), .B1(n3253), .Y(n1462)
         );
  AOI222XLTS U3384 ( .A0(n3814), .A1(n744), .B0(n4476), .B1(n3355), .C0(n4115), 
        .C1(n3830), .Y(n1463) );
  AOI22X1TS U3385 ( .A0(n464), .A1(n3268), .B0(n4280), .B1(n3253), .Y(n1460)
         );
  AOI222XLTS U3386 ( .A0(n3816), .A1(n743), .B0(n4473), .B1(n3356), .C0(n4113), 
        .C1(n3830), .Y(n1461) );
  AOI22X1TS U3387 ( .A0(n468), .A1(n3335), .B0(n4274), .B1(n3253), .Y(n1456)
         );
  AOI222XLTS U3388 ( .A0(n3816), .A1(n742), .B0(n4467), .B1(n3360), .C0(n4109), 
        .C1(n3830), .Y(n1457) );
  AOI22X1TS U3389 ( .A0(n470), .A1(n3268), .B0(n4271), .B1(n3252), .Y(n1454)
         );
  AOI222XLTS U3390 ( .A0(n3816), .A1(n741), .B0(n4464), .B1(n3355), .C0(n4107), 
        .C1(n3835), .Y(n1455) );
  AOI22X1TS U3391 ( .A0(n474), .A1(n3269), .B0(n4265), .B1(n3252), .Y(n1450)
         );
  AOI222XLTS U3392 ( .A0(n3815), .A1(n740), .B0(n4458), .B1(n3357), .C0(n4103), 
        .C1(n3835), .Y(n1451) );
  AOI22X1TS U3393 ( .A0(n478), .A1(n3338), .B0(n4259), .B1(n3251), .Y(n1446)
         );
  AOI222XLTS U3394 ( .A0(n3815), .A1(n739), .B0(n4452), .B1(n3350), .C0(n4099), 
        .C1(n3829), .Y(n1447) );
  AOI22X1TS U3395 ( .A0(n480), .A1(n3338), .B0(n4256), .B1(n3251), .Y(n1444)
         );
  AOI222XLTS U3396 ( .A0(n3814), .A1(n738), .B0(n4449), .B1(n3350), .C0(n4097), 
        .C1(n3829), .Y(n1445) );
  AOI22X1TS U3397 ( .A0(n482), .A1(n3338), .B0(n4253), .B1(n3251), .Y(n1442)
         );
  AOI222XLTS U3398 ( .A0(n3814), .A1(n737), .B0(n4446), .B1(n3350), .C0(n4095), 
        .C1(n3829), .Y(n1443) );
  AOI22X1TS U3399 ( .A0(n484), .A1(n3339), .B0(n4250), .B1(n3250), .Y(n1440)
         );
  AOI222XLTS U3400 ( .A0(n3814), .A1(n736), .B0(n4443), .B1(n3357), .C0(n4093), 
        .C1(n3829), .Y(n1441) );
  AOI22X1TS U3401 ( .A0(n486), .A1(n3341), .B0(n4247), .B1(n3250), .Y(n1438)
         );
  AOI222XLTS U3402 ( .A0(n3813), .A1(n735), .B0(n4440), .B1(n3354), .C0(n4091), 
        .C1(n3828), .Y(n1439) );
  AOI22X1TS U3403 ( .A0(n490), .A1(n3335), .B0(n4241), .B1(n3250), .Y(n1434)
         );
  AOI222XLTS U3404 ( .A0(n3813), .A1(n734), .B0(n4434), .B1(n3355), .C0(n4087), 
        .C1(n3828), .Y(n1435) );
  AOI22X1TS U3405 ( .A0(n492), .A1(n3338), .B0(n4238), .B1(n3249), .Y(n1432)
         );
  AOI222XLTS U3406 ( .A0(n3813), .A1(n733), .B0(n4431), .B1(n3349), .C0(n4085), 
        .C1(n3828), .Y(n1433) );
  AOI22X1TS U3407 ( .A0(n494), .A1(n3340), .B0(n4235), .B1(n3249), .Y(n1430)
         );
  AOI222XLTS U3408 ( .A0(n3812), .A1(n732), .B0(n4428), .B1(n3349), .C0(n4083), 
        .C1(n3827), .Y(n1431) );
  AOI22X1TS U3409 ( .A0(n496), .A1(n3335), .B0(n4232), .B1(n3249), .Y(n1428)
         );
  AOI222XLTS U3410 ( .A0(n3812), .A1(n731), .B0(n4425), .B1(n3349), .C0(n4081), 
        .C1(n3827), .Y(n1429) );
  AOI22X1TS U3411 ( .A0(n498), .A1(n3335), .B0(n4229), .B1(n3249), .Y(n1426)
         );
  AOI222XLTS U3412 ( .A0(n3812), .A1(n730), .B0(n4422), .B1(n3349), .C0(n4079), 
        .C1(n3827), .Y(n1427) );
  AOI22X1TS U3413 ( .A0(n502), .A1(n3337), .B0(n4223), .B1(n3251), .Y(n1422)
         );
  AOI222XLTS U3414 ( .A0(n3811), .A1(n729), .B0(n4416), .B1(n3348), .C0(n4076), 
        .C1(n3826), .Y(n1423) );
  AOI22X1TS U3415 ( .A0(n504), .A1(n3337), .B0(n4220), .B1(n3248), .Y(n1420)
         );
  AOI222XLTS U3416 ( .A0(n3811), .A1(n728), .B0(n4413), .B1(n3348), .C0(n4073), 
        .C1(n3826), .Y(n1421) );
  AOI22X1TS U3417 ( .A0(n451), .A1(n3337), .B0(n4217), .B1(n3248), .Y(n1418)
         );
  AOI222XLTS U3418 ( .A0(n3811), .A1(n727), .B0(n4410), .B1(n3348), .C0(n4071), 
        .C1(n3826), .Y(n1419) );
  AOI22X1TS U3419 ( .A0(n508), .A1(n3342), .B0(n4211), .B1(n3261), .Y(n1414)
         );
  AOI222XLTS U3420 ( .A0(n3810), .A1(n726), .B0(n4404), .B1(n3347), .C0(n4068), 
        .C1(n3825), .Y(n1415) );
  AOI22X1TS U3421 ( .A0(n453), .A1(n3336), .B0(n4208), .B1(n3264), .Y(n1412)
         );
  AOI222XLTS U3422 ( .A0(n3810), .A1(n725), .B0(n4401), .B1(n3347), .C0(n4065), 
        .C1(n3825), .Y(n1413) );
  AOI22X1TS U3423 ( .A0(n510), .A1(n3341), .B0(n4205), .B1(n3257), .Y(n1410)
         );
  AOI222XLTS U3424 ( .A0(n3810), .A1(n724), .B0(n4398), .B1(n3347), .C0(n4063), 
        .C1(n3825), .Y(n1411) );
  AOI22X1TS U3425 ( .A0(n3265), .A1(n119), .B0(n3990), .B1(n3255), .Y(n1997)
         );
  AOI222XLTS U3426 ( .A0(n3809), .A1(n695), .B0(n4170), .B1(n3346), .C0(n4044), 
        .C1(n3832), .Y(n1998) );
  AOI22X1TS U3427 ( .A0(n3267), .A1(n115), .B0(n3987), .B1(n3255), .Y(n1995)
         );
  AOI222XLTS U3428 ( .A0(n3817), .A1(n694), .B0(n4167), .B1(n3352), .C0(n4041), 
        .C1(n3832), .Y(n1996) );
  AOI22X1TS U3429 ( .A0(n3267), .A1(n110), .B0(n3984), .B1(n3255), .Y(n1993)
         );
  AOI222XLTS U3430 ( .A0(n3818), .A1(n693), .B0(n4164), .B1(n3352), .C0(n4040), 
        .C1(n3832), .Y(n1994) );
  AOI22X1TS U3431 ( .A0(n3266), .A1(n100), .B0(n3978), .B1(n3254), .Y(n1989)
         );
  AOI222XLTS U3432 ( .A0(n3822), .A1(n692), .B0(n4158), .B1(n3351), .C0(n4035), 
        .C1(n3831), .Y(n1990) );
  AOI22X1TS U3433 ( .A0(n3267), .A1(n31), .B0(n3975), .B1(n3254), .Y(n1987) );
  AOI222XLTS U3434 ( .A0(n3817), .A1(n691), .B0(n4155), .B1(n3351), .C0(n4034), 
        .C1(n3831), .Y(n1988) );
  AOI22X1TS U3435 ( .A0(n466), .A1(n3269), .B0(n4277), .B1(n3253), .Y(n1458)
         );
  AOI222XLTS U3436 ( .A0(n3816), .A1(n690), .B0(n4470), .B1(n3359), .C0(n4112), 
        .C1(n3830), .Y(n1459) );
  AOI22X1TS U3437 ( .A0(n500), .A1(n3336), .B0(n4226), .B1(n3248), .Y(n1424)
         );
  AOI222XLTS U3438 ( .A0(n3812), .A1(n689), .B0(n4419), .B1(n3348), .C0(n4077), 
        .C1(n3827), .Y(n1425) );
  AOI22X1TS U3439 ( .A0(n514), .A1(n3336), .B0(n4199), .B1(n3262), .Y(n1406)
         );
  AOI222XLTS U3440 ( .A0(n3809), .A1(n688), .B0(n4392), .B1(n3346), .C0(n4060), 
        .C1(n3824), .Y(n1407) );
  AOI22X1TS U3441 ( .A0(n457), .A1(n3340), .B0(n4289), .B1(n3254), .Y(n1466)
         );
  AOI222XLTS U3442 ( .A0(n3817), .A1(n668), .B0(n4482), .B1(n3351), .C0(n4120), 
        .C1(n3831), .Y(n1467) );
  AOI22X1TS U3443 ( .A0(n472), .A1(n3269), .B0(n4268), .B1(n3252), .Y(n1452)
         );
  AOI222XLTS U3444 ( .A0(n3815), .A1(n667), .B0(n4461), .B1(n3354), .C0(n4105), 
        .C1(n3835), .Y(n1453) );
  AOI22X1TS U3445 ( .A0(n476), .A1(n3269), .B0(n4262), .B1(n3252), .Y(n1448)
         );
  AOI222XLTS U3446 ( .A0(n3815), .A1(n666), .B0(n4455), .B1(n3355), .C0(n4101), 
        .C1(n3833), .Y(n1449) );
  AOI22X1TS U3447 ( .A0(n488), .A1(n3339), .B0(n4244), .B1(n3250), .Y(n1436)
         );
  AOI222XLTS U3448 ( .A0(n3813), .A1(n665), .B0(n4437), .B1(n3356), .C0(n4089), 
        .C1(n3828), .Y(n1437) );
  AOI22X1TS U3449 ( .A0(n506), .A1(n3336), .B0(n4214), .B1(n3248), .Y(n1416)
         );
  AOI222XLTS U3450 ( .A0(n3811), .A1(n664), .B0(n4407), .B1(n3350), .C0(n4069), 
        .C1(n3826), .Y(n1417) );
  AOI22X1TS U3451 ( .A0(n455), .A1(n3343), .B0(n4202), .B1(n1233), .Y(n1408)
         );
  AOI222XLTS U3452 ( .A0(n3810), .A1(n663), .B0(n4395), .B1(n3347), .C0(n4061), 
        .C1(n3825), .Y(n1409) );
  AOI22X1TS U3453 ( .A0(n512), .A1(n3341), .B0(n4196), .B1(n3262), .Y(n1404)
         );
  AOI222XLTS U3454 ( .A0(n3809), .A1(n662), .B0(n4389), .B1(n3346), .C0(n4057), 
        .C1(n3824), .Y(n1405) );
  AOI22X1TS U3455 ( .A0(n3987), .A1(n3503), .B0(n4042), .B1(n3774), .Y(n1926)
         );
  AOI222XLTS U3456 ( .A0(n4166), .A1(n3549), .B0(n3535), .B1(n117), .C0(n3946), 
        .C1(n3528), .Y(n1927) );
  AOI22X1TS U3457 ( .A0(n4388), .A1(n3609), .B0(n4058), .B1(n3753), .Y(n1661)
         );
  NOR2BX1TS U3458 ( .AN(n3000), .B(n432), .Y(n2997) );
  XOR2X1TS U3459 ( .A(n1130), .B(selectBit_WEST), .Y(n2998) );
  OAI33XLTS U3460 ( .A0(n4150), .A1(n129), .A2(n161), .B0(n996), .B1(n156), 
        .B2(n1837), .Y(n1834) );
  NAND2X1TS U3461 ( .A(readReady), .B(n534), .Y(n1888) );
  OAI22X1TS U3462 ( .A0(n148), .A1(n1136), .B0(n10), .B1(n1134), .Y(n2886) );
  INVX2TS U3463 ( .A(n4149), .Y(n4148) );
  OAI22X1TS U3464 ( .A0(n1132), .A1(n148), .B0(n439), .B1(n1134), .Y(n2888) );
  INVX2TS U3465 ( .A(readReady), .Y(n1130) );
  INVX2TS U3466 ( .A(selectBit_WEST), .Y(n1084) );
  NAND2X1TS U3467 ( .A(n4141), .B(n940), .Y(n1861) );
  OAI33XLTS U3468 ( .A0(n4150), .A1(n940), .A2(n161), .B0(n431), .B1(n950), 
        .B2(n1865), .Y(n1864) );
  NAND2X1TS U3469 ( .A(readIn_SOUTH), .B(n1822), .Y(n1817) );
  AOI222XLTS U3470 ( .A0(n4147), .A1(n1819), .B0(readIn_NORTH), .B1(n1820), 
        .C0(n4142), .C1(n1821), .Y(n1818) );
  NAND2BX1TS U3471 ( .AN(n1853), .B(readIn_SOUTH), .Y(n1847) );
  AOI21X1TS U3472 ( .A0(n4142), .A1(n943), .B0(n1849), .Y(n1848) );
  OAI221XLTS U3473 ( .A0(n4146), .A1(n2072), .B0(n203), .B1(n2070), .C0(n126), 
        .Y(n2089) );
  AOI221X1TS U3474 ( .A0(n1033), .A1(n4383), .B0(n1058), .B1(dataIn_NORTH[30]), 
        .C0(n2949), .Y(n2942) );
  OAI22X1TS U3475 ( .A0(n3182), .A1(n1110), .B0(n717), .B1(n3725), .Y(n2949)
         );
  AOI221X1TS U3476 ( .A0(n1033), .A1(n4380), .B0(n1060), .B1(dataIn_NORTH[29]), 
        .C0(n2940), .Y(n2934) );
  OAI22X1TS U3477 ( .A0(n3173), .A1(n1110), .B0(n716), .B1(n3725), .Y(n2940)
         );
  AOI221X1TS U3478 ( .A0(n1033), .A1(n4377), .B0(n1060), .B1(dataIn_NORTH[28]), 
        .C0(n2932), .Y(n2927) );
  OAI22X1TS U3479 ( .A0(n3164), .A1(n1110), .B0(n715), .B1(n3725), .Y(n2932)
         );
  AOI221X1TS U3480 ( .A0(n1034), .A1(n4374), .B0(n1059), .B1(dataIn_NORTH[27]), 
        .C0(n2922), .Y(n2917) );
  OAI22X1TS U3481 ( .A0(n3155), .A1(n1110), .B0(n714), .B1(n3726), .Y(n2922)
         );
  AOI221X1TS U3482 ( .A0(n1034), .A1(n4371), .B0(n1058), .B1(dataIn_NORTH[26]), 
        .C0(n2915), .Y(n2906) );
  OAI22X1TS U3483 ( .A0(n3146), .A1(n1109), .B0(n713), .B1(n3726), .Y(n2915)
         );
  AOI221X1TS U3484 ( .A0(n1034), .A1(n4368), .B0(n1059), .B1(dataIn_NORTH[25]), 
        .C0(n2904), .Y(n2894) );
  OAI22X1TS U3485 ( .A0(n3137), .A1(n1109), .B0(n686), .B1(n3726), .Y(n2904)
         );
  AOI221X1TS U3486 ( .A0(n1034), .A1(n4365), .B0(n1064), .B1(dataIn_NORTH[24]), 
        .C0(n2892), .Y(n2395) );
  OAI22X1TS U3487 ( .A0(n3128), .A1(n1109), .B0(n712), .B1(n3726), .Y(n2892)
         );
  AOI221X1TS U3488 ( .A0(n1035), .A1(n4362), .B0(n1056), .B1(dataIn_NORTH[23]), 
        .C0(n2393), .Y(n2387) );
  OAI22X1TS U3489 ( .A0(n3119), .A1(n1109), .B0(n685), .B1(n3737), .Y(n2393)
         );
  AOI221X1TS U3490 ( .A0(n1035), .A1(n4359), .B0(n1056), .B1(dataIn_NORTH[22]), 
        .C0(n2385), .Y(n2381) );
  OAI22X1TS U3491 ( .A0(n3110), .A1(n1108), .B0(n711), .B1(n3737), .Y(n2385)
         );
  AOI221X1TS U3492 ( .A0(n1035), .A1(n4356), .B0(n1056), .B1(dataIn_NORTH[21]), 
        .C0(n2377), .Y(n2373) );
  OAI22X1TS U3493 ( .A0(n3101), .A1(n1108), .B0(n709), .B1(n3734), .Y(n2377)
         );
  AOI221X1TS U3494 ( .A0(n1035), .A1(n4353), .B0(n1056), .B1(dataIn_NORTH[20]), 
        .C0(n2369), .Y(n2364) );
  OAI22X1TS U3495 ( .A0(n3092), .A1(n1108), .B0(n684), .B1(n3734), .Y(n2369)
         );
  AOI221X1TS U3496 ( .A0(n1036), .A1(n4350), .B0(n1055), .B1(dataIn_NORTH[19]), 
        .C0(n2362), .Y(n2356) );
  OAI22X1TS U3497 ( .A0(n3083), .A1(n1108), .B0(n708), .B1(n3737), .Y(n2362)
         );
  AOI221X1TS U3498 ( .A0(n1036), .A1(n4347), .B0(n1055), .B1(dataIn_NORTH[18]), 
        .C0(n2354), .Y(n2350) );
  OAI22X1TS U3499 ( .A0(n3074), .A1(n1107), .B0(n683), .B1(n3737), .Y(n2354)
         );
  AOI221X1TS U3500 ( .A0(n1036), .A1(n4344), .B0(n1055), .B1(dataIn_NORTH[17]), 
        .C0(n2348), .Y(n2344) );
  OAI22X1TS U3501 ( .A0(n3065), .A1(n1107), .B0(n707), .B1(n3735), .Y(n2348)
         );
  AOI221X1TS U3502 ( .A0(n1036), .A1(n4341), .B0(n1055), .B1(dataIn_NORTH[16]), 
        .C0(n2342), .Y(n2338) );
  OAI22X1TS U3503 ( .A0(n3056), .A1(n1107), .B0(n706), .B1(n3738), .Y(n2342)
         );
  AOI221X1TS U3504 ( .A0(n1037), .A1(n4338), .B0(n1054), .B1(dataIn_NORTH[15]), 
        .C0(n2336), .Y(n2332) );
  OAI22X1TS U3505 ( .A0(n3047), .A1(n1107), .B0(n682), .B1(n3727), .Y(n2336)
         );
  AOI221X1TS U3506 ( .A0(n1037), .A1(n4335), .B0(n1054), .B1(dataIn_NORTH[14]), 
        .C0(n2330), .Y(n2326) );
  OAI22X1TS U3507 ( .A0(n3038), .A1(n1106), .B0(n705), .B1(n3727), .Y(n2330)
         );
  AOI221X1TS U3508 ( .A0(n1037), .A1(n4332), .B0(n1054), .B1(dataIn_NORTH[13]), 
        .C0(n2324), .Y(n2320) );
  OAI22X1TS U3509 ( .A0(n3029), .A1(n1106), .B0(n681), .B1(n3727), .Y(n2324)
         );
  AOI221X1TS U3510 ( .A0(n1037), .A1(n4329), .B0(n1054), .B1(dataIn_NORTH[12]), 
        .C0(n2318), .Y(n2314) );
  OAI22X1TS U3511 ( .A0(n3020), .A1(n1106), .B0(n704), .B1(n3727), .Y(n2318)
         );
  AOI221X1TS U3512 ( .A0(n1038), .A1(n4326), .B0(n1058), .B1(dataIn_NORTH[11]), 
        .C0(n2312), .Y(n2308) );
  OAI22X1TS U3513 ( .A0(n3011), .A1(n1106), .B0(n703), .B1(n3728), .Y(n2312)
         );
  AOI221X1TS U3514 ( .A0(n1038), .A1(n4323), .B0(n1061), .B1(dataIn_NORTH[10]), 
        .C0(n2306), .Y(n2302) );
  OAI22X1TS U3515 ( .A0(n3002), .A1(n1105), .B0(n702), .B1(n3728), .Y(n2306)
         );
  AOI221X1TS U3516 ( .A0(n1038), .A1(n4320), .B0(n1062), .B1(dataIn_NORTH[9]), 
        .C0(n2300), .Y(n2296) );
  OAI22X1TS U3517 ( .A0(n2993), .A1(n1105), .B0(n701), .B1(n3728), .Y(n2300)
         );
  AOI221X1TS U3518 ( .A0(n1038), .A1(n4317), .B0(n2100), .B1(dataIn_NORTH[8]), 
        .C0(n2294), .Y(n2290) );
  OAI22X1TS U3519 ( .A0(n2984), .A1(n1105), .B0(n700), .B1(n3728), .Y(n2294)
         );
  AOI221X1TS U3520 ( .A0(n1039), .A1(n4311), .B0(n1059), .B1(dataIn_NORTH[6]), 
        .C0(n2277), .Y(n2273) );
  OAI22X1TS U3521 ( .A0(n2966), .A1(n1104), .B0(n699), .B1(n3729), .Y(n2277)
         );
  AOI221X1TS U3522 ( .A0(n1039), .A1(n4308), .B0(n1061), .B1(dataIn_NORTH[5]), 
        .C0(n2271), .Y(n2267) );
  OAI22X1TS U3523 ( .A0(n2957), .A1(n1104), .B0(n680), .B1(n3729), .Y(n2271)
         );
  AOI221X1TS U3524 ( .A0(n1040), .A1(n4302), .B0(n1057), .B1(dataIn_NORTH[3]), 
        .C0(n2259), .Y(n2255) );
  OAI22X1TS U3525 ( .A0(n2939), .A1(n1103), .B0(n698), .B1(n3730), .Y(n2259)
         );
  AOI221X1TS U3526 ( .A0(n1040), .A1(n4296), .B0(n1059), .B1(dataIn_NORTH[1]), 
        .C0(n2247), .Y(n2243) );
  OAI22X1TS U3527 ( .A0(n2921), .A1(n1103), .B0(n697), .B1(n3730), .Y(n2247)
         );
  AOI221X1TS U3528 ( .A0(n1040), .A1(n4293), .B0(n1062), .B1(dataIn_NORTH[0]), 
        .C0(n2241), .Y(n2237) );
  OAI22X1TS U3529 ( .A0(n2912), .A1(n1103), .B0(n696), .B1(n3730), .Y(n2241)
         );
  AOI221X1TS U3530 ( .A0(n1042), .A1(n3949), .B0(n1052), .B1(
        destinationAddressIn_NORTH[5]), .C0(n2199), .Y(n2195) );
  OAI22X1TS U3531 ( .A0(n2899), .A1(n1102), .B0(n723), .B1(n3732), .Y(n2199)
         );
  AOI221X1TS U3532 ( .A0(n1042), .A1(n3946), .B0(n1052), .B1(
        destinationAddressIn_NORTH[4]), .C0(n2193), .Y(n2189) );
  OAI22X1TS U3533 ( .A0(n2890), .A1(n1102), .B0(n722), .B1(n3732), .Y(n2193)
         );
  AOI221X1TS U3534 ( .A0(n1043), .A1(n3943), .B0(n1051), .B1(
        destinationAddressIn_NORTH[3]), .C0(n2187), .Y(n2183) );
  OAI22X1TS U3535 ( .A0(n2388), .A1(n1105), .B0(n721), .B1(n3733), .Y(n2187)
         );
  AOI221X1TS U3536 ( .A0(n1043), .A1(n3940), .B0(n1051), .B1(
        destinationAddressIn_NORTH[2]), .C0(n2181), .Y(n2177) );
  OAI22X1TS U3537 ( .A0(n2379), .A1(n1102), .B0(n687), .B1(n3733), .Y(n2181)
         );
  AOI221X1TS U3538 ( .A0(n1043), .A1(n3934), .B0(n1051), .B1(
        destinationAddressIn_NORTH[0]), .C0(n2168), .Y(n2157) );
  OAI22X1TS U3539 ( .A0(n2361), .A1(n1102), .B0(n719), .B1(n3733), .Y(n2168)
         );
  AOI221X1TS U3540 ( .A0(n1039), .A1(n4314), .B0(n1062), .B1(dataIn_NORTH[7]), 
        .C0(n2287), .Y(n2279) );
  OAI22X1TS U3541 ( .A0(n2975), .A1(n1104), .B0(n2968), .B1(n3729), .Y(n2287)
         );
  AOI221X1TS U3542 ( .A0(n1039), .A1(n4305), .B0(n2100), .B1(dataIn_NORTH[4]), 
        .C0(n2265), .Y(n2261) );
  OAI22X1TS U3543 ( .A0(n2948), .A1(n1104), .B0(n2944), .B1(n3729), .Y(n2265)
         );
  AOI221X1TS U3544 ( .A0(n1040), .A1(n4299), .B0(n1063), .B1(dataIn_NORTH[2]), 
        .C0(n2253), .Y(n2249) );
  OAI22X1TS U3545 ( .A0(n2930), .A1(n1103), .B0(n2924), .B1(n3730), .Y(n2253)
         );
  AOI221X1TS U3546 ( .A0(n1033), .A1(n4386), .B0(n1057), .B1(dataIn_NORTH[31]), 
        .C0(n2958), .Y(n2953) );
  OAI22X1TS U3547 ( .A0(n3191), .A1(n1101), .B0(n718), .B1(n3725), .Y(n2958)
         );
  AOI221X1TS U3548 ( .A0(n1041), .A1(n4137), .B0(n1053), .B1(
        requesterAddressIn_NORTH[5]), .C0(n2235), .Y(n2231) );
  OAI22X1TS U3549 ( .A0(n1101), .A1(n2903), .B0(n877), .B1(n3731), .Y(n2235)
         );
  AOI221X1TS U3550 ( .A0(n1041), .A1(n4134), .B0(n1053), .B1(
        requesterAddressIn_NORTH[4]), .C0(n2229), .Y(n2225) );
  OAI22X1TS U3551 ( .A0(n1101), .A1(n2902), .B0(n878), .B1(n3731), .Y(n2229)
         );
  AOI221X1TS U3552 ( .A0(n1041), .A1(n4128), .B0(n1053), .B1(
        requesterAddressIn_NORTH[2]), .C0(n2217), .Y(n2213) );
  OAI22X1TS U3553 ( .A0(n1100), .A1(n2901), .B0(n875), .B1(n3731), .Y(n2217)
         );
  AOI221X1TS U3554 ( .A0(n1042), .A1(n4125), .B0(n1052), .B1(
        requesterAddressIn_NORTH[1]), .C0(n2211), .Y(n2207) );
  OAI22X1TS U3555 ( .A0(n1100), .A1(n2900), .B0(n874), .B1(n3732), .Y(n2211)
         );
  AOI221X1TS U3556 ( .A0(n1043), .A1(n3937), .B0(n1051), .B1(
        destinationAddressIn_NORTH[1]), .C0(n2175), .Y(n2171) );
  OAI22X1TS U3557 ( .A0(n2370), .A1(n1101), .B0(n720), .B1(n3733), .Y(n2175)
         );
  AOI221X1TS U3558 ( .A0(n1041), .A1(n4131), .B0(n1053), .B1(
        requesterAddressIn_NORTH[3]), .C0(n2223), .Y(n2219) );
  OAI22X1TS U3559 ( .A0(n1100), .A1(n2283), .B0(n876), .B1(n3731), .Y(n2223)
         );
  AOI221X1TS U3560 ( .A0(n1042), .A1(n4122), .B0(n1052), .B1(
        requesterAddressIn_NORTH[0]), .C0(n2205), .Y(n2201) );
  OAI22X1TS U3561 ( .A0(n1100), .A1(n2284), .B0(n873), .B1(n3732), .Y(n2205)
         );
  NAND4X1TS U3562 ( .A(n2951), .B(n2953), .C(n2954), .D(n2955), .Y(n2397) );
  AOI221X1TS U3563 ( .A0(n1018), .A1(n3141), .B0(n1016), .B1(n668), .C0(n2956), 
        .Y(n2955) );
  AOI222XLTS U3564 ( .A0(n2165), .A1(n40), .B0(n710), .B1(n3039), .C0(n2167), 
        .C1(n3036), .Y(n2954) );
  AOI222XLTS U3565 ( .A0(n1065), .A1(n4482), .B0(n1085), .B1(n4289), .C0(n2169), .C1(cacheDataOut[31]), .Y(n2951) );
  NAND4X1TS U3566 ( .A(n2941), .B(n2942), .C(n2943), .D(n2946), .Y(n2398) );
  AOI221X1TS U3567 ( .A0(n1018), .A1(n3142), .B0(n1017), .B1(n745), .C0(n2947), 
        .Y(n2946) );
  AOI222XLTS U3568 ( .A0(n2165), .A1(n41), .B0(n710), .B1(n3041), .C0(n2167), 
        .C1(n3040), .Y(n2943) );
  AOI222XLTS U3569 ( .A0(n1065), .A1(n4479), .B0(n1094), .B1(n4286), .C0(n2169), .C1(cacheDataOut[30]), .Y(n2941) );
  NAND4X1TS U3570 ( .A(n2933), .B(n2934), .C(n2935), .D(n2936), .Y(n2399) );
  AOI221X1TS U3571 ( .A0(n1018), .A1(n3144), .B0(n1016), .B1(n744), .C0(n2937), 
        .Y(n2936) );
  AOI222XLTS U3572 ( .A0(n964), .A1(n42), .B0(n710), .B1(n3043), .C0(n561), 
        .C1(n3042), .Y(n2935) );
  AOI222XLTS U3573 ( .A0(n1065), .A1(n4476), .B0(n1094), .B1(n4283), .C0(n547), 
        .C1(cacheDataOut[29]), .Y(n2933) );
  NAND4X1TS U3574 ( .A(n2926), .B(n2927), .C(n2928), .D(n2929), .Y(n2400) );
  AOI221X1TS U3575 ( .A0(n1018), .A1(n3145), .B0(n2161), .B1(n743), .C0(n2931), 
        .Y(n2929) );
  AOI222XLTS U3576 ( .A0(n963), .A1(n677), .B0(n710), .B1(n3046), .C0(n560), 
        .C1(n3045), .Y(n2928) );
  AOI222XLTS U3577 ( .A0(n1065), .A1(n4473), .B0(n1098), .B1(n4280), .C0(n546), 
        .C1(cacheDataOut[28]), .Y(n2926) );
  NAND4X1TS U3578 ( .A(n2916), .B(n2917), .C(n2918), .D(n2919), .Y(n2401) );
  AOI221X1TS U3579 ( .A0(n1028), .A1(n3149), .B0(n1004), .B1(n690), .C0(n2920), 
        .Y(n2919) );
  AOI222XLTS U3580 ( .A0(n785), .A1(n676), .B0(n779), .B1(n3050), .C0(n549), 
        .C1(n3048), .Y(n2918) );
  AOI222XLTS U3581 ( .A0(n1078), .A1(n4470), .B0(n1097), .B1(n4277), .C0(n535), 
        .C1(cacheDataOut[27]), .Y(n2916) );
  NAND4X1TS U3582 ( .A(n2905), .B(n2906), .C(n2908), .D(n2910), .Y(n2402) );
  AOI221X1TS U3583 ( .A0(n1030), .A1(n3150), .B0(n1004), .B1(n742), .C0(n2911), 
        .Y(n2910) );
  AOI222XLTS U3584 ( .A0(n785), .A1(n43), .B0(n772), .B1(n3052), .C0(n549), 
        .C1(n3051), .Y(n2908) );
  AOI222XLTS U3585 ( .A0(n1074), .A1(n4467), .B0(n1099), .B1(n4274), .C0(n535), 
        .C1(cacheDataOut[26]), .Y(n2905) );
  NAND4X1TS U3586 ( .A(n2893), .B(n2894), .C(n2896), .D(n2897), .Y(n2403) );
  AOI221X1TS U3587 ( .A0(n1028), .A1(n3151), .B0(n1004), .B1(n741), .C0(n2898), 
        .Y(n2897) );
  AOI222XLTS U3588 ( .A0(n785), .A1(n44), .B0(n782), .B1(n3054), .C0(n549), 
        .C1(n3053), .Y(n2896) );
  AOI222XLTS U3589 ( .A0(n1075), .A1(n4464), .B0(n1095), .B1(n4271), .C0(n535), 
        .C1(cacheDataOut[25]), .Y(n2893) );
  NAND4X1TS U3590 ( .A(n2394), .B(n2395), .C(n2396), .D(n2449), .Y(n2404) );
  AOI221X1TS U3591 ( .A0(n2160), .A1(n3152), .B0(n1004), .B1(n667), .C0(n2891), 
        .Y(n2449) );
  AOI222XLTS U3592 ( .A0(n785), .A1(n45), .B0(n772), .B1(n3057), .C0(n549), 
        .C1(n3055), .Y(n2396) );
  AOI222XLTS U3593 ( .A0(n1078), .A1(n4461), .B0(n1096), .B1(n4268), .C0(n535), 
        .C1(cacheDataOut[24]), .Y(n2394) );
  NAND4X1TS U3594 ( .A(n2386), .B(n2387), .C(n2390), .D(n2391), .Y(n2405) );
  AOI221X1TS U3595 ( .A0(n1027), .A1(n3153), .B0(n1015), .B1(n740), .C0(n2392), 
        .Y(n2391) );
  AOI222XLTS U3596 ( .A0(n786), .A1(n675), .B0(n779), .B1(n3059), .C0(n550), 
        .C1(n3058), .Y(n2390) );
  AOI222XLTS U3597 ( .A0(n1076), .A1(n4458), .B0(n1097), .B1(n4265), .C0(n536), 
        .C1(cacheDataOut[23]), .Y(n2386) );
  NAND4X1TS U3598 ( .A(n2378), .B(n2381), .C(n2382), .D(n2383), .Y(n2406) );
  AOI221X1TS U3599 ( .A0(n1031), .A1(n3154), .B0(n1013), .B1(n666), .C0(n2384), 
        .Y(n2383) );
  AOI222XLTS U3600 ( .A0(n786), .A1(n46), .B0(n779), .B1(n3062), .C0(n550), 
        .C1(n3061), .Y(n2382) );
  AOI222XLTS U3601 ( .A0(n1075), .A1(n4455), .B0(n1096), .B1(n4262), .C0(n536), 
        .C1(cacheDataOut[22]), .Y(n2378) );
  NAND4X1TS U3602 ( .A(n2371), .B(n2373), .C(n2374), .D(n2375), .Y(n2407) );
  AOI221X1TS U3603 ( .A0(n1027), .A1(n3156), .B0(n1012), .B1(n739), .C0(n2376), 
        .Y(n2375) );
  AOI222XLTS U3604 ( .A0(n786), .A1(n47), .B0(n778), .B1(n3064), .C0(n550), 
        .C1(n3063), .Y(n2374) );
  AOI222XLTS U3605 ( .A0(n1078), .A1(n4452), .B0(n1093), .B1(n4259), .C0(n536), 
        .C1(cacheDataOut[21]), .Y(n2371) );
  NAND4X1TS U3606 ( .A(n2363), .B(n2364), .C(n2365), .D(n2367), .Y(n2408) );
  AOI221X1TS U3607 ( .A0(n1032), .A1(n3158), .B0(n1011), .B1(n738), .C0(n2368), 
        .Y(n2367) );
  AOI222XLTS U3608 ( .A0(n786), .A1(n674), .B0(n776), .B1(n3067), .C0(n550), 
        .C1(n3066), .Y(n2365) );
  AOI222XLTS U3609 ( .A0(n1077), .A1(n4449), .B0(n1099), .B1(n4256), .C0(n536), 
        .C1(cacheDataOut[20]), .Y(n2363) );
  NAND4X1TS U3610 ( .A(n2355), .B(n2356), .C(n2357), .D(n2358), .Y(n2409) );
  AOI221X1TS U3611 ( .A0(n1019), .A1(n3159), .B0(n1014), .B1(n737), .C0(n2360), 
        .Y(n2358) );
  AOI222XLTS U3612 ( .A0(n787), .A1(n48), .B0(n782), .B1(n3070), .C0(n551), 
        .C1(n3068), .Y(n2357) );
  AOI222XLTS U3613 ( .A0(n1079), .A1(n4446), .B0(n1095), .B1(n4253), .C0(n537), 
        .C1(cacheDataOut[19]), .Y(n2355) );
  NAND4X1TS U3614 ( .A(n2349), .B(n2350), .C(n2351), .D(n2352), .Y(n2410) );
  AOI221X1TS U3615 ( .A0(n1019), .A1(n3160), .B0(n1014), .B1(n736), .C0(n2353), 
        .Y(n2352) );
  AOI222XLTS U3616 ( .A0(n787), .A1(n49), .B0(n778), .B1(n3072), .C0(n551), 
        .C1(n3071), .Y(n2351) );
  AOI222XLTS U3617 ( .A0(n1076), .A1(n4443), .B0(n1092), .B1(n4250), .C0(n537), 
        .C1(cacheDataOut[18]), .Y(n2349) );
  NAND4X1TS U3618 ( .A(n2343), .B(n2344), .C(n2345), .D(n2346), .Y(n2411) );
  AOI221X1TS U3619 ( .A0(n1019), .A1(n3162), .B0(n1014), .B1(n735), .C0(n2347), 
        .Y(n2346) );
  AOI222XLTS U3620 ( .A0(n787), .A1(n50), .B0(n783), .B1(n3075), .C0(n551), 
        .C1(n3073), .Y(n2345) );
  AOI222XLTS U3621 ( .A0(n1079), .A1(n4440), .B0(n1092), .B1(n4247), .C0(n537), 
        .C1(cacheDataOut[17]), .Y(n2343) );
  NAND4X1TS U3622 ( .A(n2337), .B(n2338), .C(n2339), .D(n2340), .Y(n2412) );
  AOI221X1TS U3623 ( .A0(n1019), .A1(n3163), .B0(n1015), .B1(n665), .C0(n2341), 
        .Y(n2340) );
  AOI222XLTS U3624 ( .A0(n787), .A1(n51), .B0(n779), .B1(n3077), .C0(n551), 
        .C1(n3076), .Y(n2339) );
  AOI222XLTS U3625 ( .A0(n1074), .A1(n4437), .B0(n1092), .B1(n4244), .C0(n537), 
        .C1(cacheDataOut[16]), .Y(n2337) );
  NAND4X1TS U3626 ( .A(n2331), .B(n2332), .C(n2333), .D(n2334), .Y(n2413) );
  AOI221X1TS U3627 ( .A0(n1020), .A1(n3165), .B0(n1014), .B1(n734), .C0(n2335), 
        .Y(n2334) );
  AOI222XLTS U3628 ( .A0(n963), .A1(n52), .B0(n776), .B1(n3079), .C0(n560), 
        .C1(n3078), .Y(n2333) );
  AOI222XLTS U3629 ( .A0(n1066), .A1(n4434), .B0(n1092), .B1(n4241), .C0(n546), 
        .C1(cacheDataOut[15]), .Y(n2331) );
  NAND4X1TS U3630 ( .A(n2325), .B(n2326), .C(n2327), .D(n2328), .Y(n2414) );
  AOI221X1TS U3631 ( .A0(n1020), .A1(n3166), .B0(n1013), .B1(n733), .C0(n2329), 
        .Y(n2328) );
  AOI222XLTS U3632 ( .A0(n962), .A1(n53), .B0(n781), .B1(n3081), .C0(n559), 
        .C1(n3080), .Y(n2327) );
  AOI222XLTS U3633 ( .A0(n1066), .A1(n4431), .B0(n1091), .B1(n4238), .C0(n545), 
        .C1(cacheDataOut[14]), .Y(n2325) );
  NAND4X1TS U3634 ( .A(n2319), .B(n2320), .C(n2321), .D(n2322), .Y(n2415) );
  AOI221X1TS U3635 ( .A0(n1020), .A1(n3167), .B0(n1012), .B1(n732), .C0(n2323), 
        .Y(n2322) );
  AOI222XLTS U3636 ( .A0(n961), .A1(n54), .B0(n781), .B1(n3086), .C0(n558), 
        .C1(n3084), .Y(n2321) );
  AOI222XLTS U3637 ( .A0(n1066), .A1(n4428), .B0(n1091), .B1(n4235), .C0(n544), 
        .C1(cacheDataOut[13]), .Y(n2319) );
  NAND4X1TS U3638 ( .A(n2313), .B(n2314), .C(n2315), .D(n2316), .Y(n2416) );
  AOI221X1TS U3639 ( .A0(n1020), .A1(n3168), .B0(n1011), .B1(n731), .C0(n2317), 
        .Y(n2316) );
  AOI222XLTS U3640 ( .A0(n962), .A1(n55), .B0(n781), .B1(n3089), .C0(n559), 
        .C1(n3088), .Y(n2315) );
  AOI222XLTS U3641 ( .A0(n1066), .A1(n4425), .B0(n1091), .B1(n4232), .C0(n545), 
        .C1(cacheDataOut[12]), .Y(n2313) );
  NAND4X1TS U3642 ( .A(n2307), .B(n2308), .C(n2309), .D(n2310), .Y(n2417) );
  AOI221X1TS U3643 ( .A0(n1021), .A1(n3169), .B0(n1005), .B1(n730), .C0(n2311), 
        .Y(n2310) );
  AOI222XLTS U3644 ( .A0(n899), .A1(n56), .B0(n755), .B1(n3091), .C0(n552), 
        .C1(n3090), .Y(n2309) );
  AOI222XLTS U3645 ( .A0(n1067), .A1(n4422), .B0(n1091), .B1(n4229), .C0(n538), 
        .C1(cacheDataOut[11]), .Y(n2307) );
  NAND4X1TS U3646 ( .A(n2301), .B(n2302), .C(n2303), .D(n2304), .Y(n2418) );
  AOI221X1TS U3647 ( .A0(n1021), .A1(n3170), .B0(n1005), .B1(n689), .C0(n2305), 
        .Y(n2304) );
  AOI222XLTS U3648 ( .A0(n899), .A1(n57), .B0(n755), .B1(n3094), .C0(n552), 
        .C1(n3093), .Y(n2303) );
  AOI222XLTS U3649 ( .A0(n1067), .A1(n4419), .B0(n1090), .B1(n4226), .C0(n538), 
        .C1(cacheDataOut[10]), .Y(n2301) );
  NAND4X1TS U3650 ( .A(n2295), .B(n2296), .C(n2297), .D(n2298), .Y(n2419) );
  AOI221X1TS U3651 ( .A0(n1021), .A1(n3171), .B0(n1005), .B1(n729), .C0(n2299), 
        .Y(n2298) );
  AOI222XLTS U3652 ( .A0(n899), .A1(n673), .B0(n755), .B1(n3096), .C0(n552), 
        .C1(n3095), .Y(n2297) );
  AOI222XLTS U3653 ( .A0(n1067), .A1(n4416), .B0(n1090), .B1(n4223), .C0(n538), 
        .C1(cacheDataOut[9]), .Y(n2295) );
  NAND4X1TS U3654 ( .A(n2289), .B(n2290), .C(n2291), .D(n2292), .Y(n2420) );
  AOI221X1TS U3655 ( .A0(n1021), .A1(n3174), .B0(n1005), .B1(n728), .C0(n2293), 
        .Y(n2292) );
  AOI222XLTS U3656 ( .A0(n899), .A1(n58), .B0(n755), .B1(n3098), .C0(n552), 
        .C1(n3097), .Y(n2291) );
  AOI222XLTS U3657 ( .A0(n1067), .A1(n4413), .B0(n1090), .B1(n4220), .C0(n538), 
        .C1(cacheDataOut[8]), .Y(n2289) );
  NAND4X1TS U3658 ( .A(n2278), .B(n2279), .C(n2280), .D(n2281), .Y(n2421) );
  AOI221X1TS U3659 ( .A0(n1022), .A1(n3175), .B0(n1006), .B1(n727), .C0(n2282), 
        .Y(n2281) );
  AOI222XLTS U3660 ( .A0(n900), .A1(n59), .B0(n756), .B1(n3102), .C0(n553), 
        .C1(n3099), .Y(n2280) );
  AOI222XLTS U3661 ( .A0(n1068), .A1(n4410), .B0(n1090), .B1(n4217), .C0(n539), 
        .C1(cacheDataOut[7]), .Y(n2278) );
  NAND4X1TS U3662 ( .A(n2272), .B(n2273), .C(n2274), .D(n2275), .Y(n2422) );
  AOI221X1TS U3663 ( .A0(n1022), .A1(n3176), .B0(n1006), .B1(n664), .C0(n2276), 
        .Y(n2275) );
  AOI222XLTS U3664 ( .A0(n900), .A1(n60), .B0(n756), .B1(n3105), .C0(n553), 
        .C1(n3104), .Y(n2274) );
  AOI222XLTS U3665 ( .A0(n1068), .A1(n4407), .B0(n1089), .B1(n4214), .C0(n539), 
        .C1(cacheDataOut[6]), .Y(n2272) );
  NAND4X1TS U3666 ( .A(n2266), .B(n2267), .C(n2268), .D(n2269), .Y(n2423) );
  AOI221X1TS U3667 ( .A0(n1022), .A1(n3177), .B0(n1006), .B1(n726), .C0(n2270), 
        .Y(n2269) );
  AOI222XLTS U3668 ( .A0(n900), .A1(n672), .B0(n756), .B1(n3107), .C0(n553), 
        .C1(n3106), .Y(n2268) );
  AOI222XLTS U3669 ( .A0(n1068), .A1(n4404), .B0(n1089), .B1(n4211), .C0(n539), 
        .C1(cacheDataOut[5]), .Y(n2266) );
  NAND4X1TS U3670 ( .A(n2260), .B(n2261), .C(n2262), .D(n2263), .Y(n2424) );
  AOI221X1TS U3671 ( .A0(n1022), .A1(n3178), .B0(n1006), .B1(n725), .C0(n2264), 
        .Y(n2263) );
  AOI222XLTS U3672 ( .A0(n900), .A1(n61), .B0(n756), .B1(n3109), .C0(n553), 
        .C1(n3108), .Y(n2262) );
  AOI222XLTS U3673 ( .A0(n1068), .A1(n4401), .B0(n1089), .B1(n4208), .C0(n539), 
        .C1(cacheDataOut[4]), .Y(n2260) );
  NAND4X1TS U3674 ( .A(n2254), .B(n2255), .C(n2256), .D(n2257), .Y(n2425) );
  AOI221X1TS U3675 ( .A0(n1023), .A1(n3180), .B0(n1007), .B1(n724), .C0(n2258), 
        .Y(n2257) );
  AOI222XLTS U3676 ( .A0(n935), .A1(n62), .B0(n763), .B1(n3113), .C0(n554), 
        .C1(n3111), .Y(n2256) );
  AOI222XLTS U3677 ( .A0(n1069), .A1(n4398), .B0(n1088), .B1(n4205), .C0(n540), 
        .C1(cacheDataOut[3]), .Y(n2254) );
  NAND4X1TS U3678 ( .A(n2248), .B(n2249), .C(n2250), .D(n2251), .Y(n2426) );
  AOI221X1TS U3679 ( .A0(n1023), .A1(n3181), .B0(n1007), .B1(n663), .C0(n2252), 
        .Y(n2251) );
  AOI222XLTS U3680 ( .A0(n935), .A1(n671), .B0(n763), .B1(n3116), .C0(n554), 
        .C1(n3115), .Y(n2250) );
  AOI222XLTS U3681 ( .A0(n1069), .A1(n4395), .B0(n1088), .B1(n4202), .C0(n540), 
        .C1(cacheDataOut[2]), .Y(n2248) );
  NAND4X1TS U3682 ( .A(n2242), .B(n2243), .C(n2244), .D(n2245), .Y(n2427) );
  AOI221X1TS U3683 ( .A0(n1023), .A1(n3183), .B0(n1007), .B1(n688), .C0(n2246), 
        .Y(n2245) );
  AOI222XLTS U3684 ( .A0(n935), .A1(n670), .B0(n763), .B1(n3118), .C0(n554), 
        .C1(n3117), .Y(n2244) );
  AOI222XLTS U3685 ( .A0(n1069), .A1(n4392), .B0(n1088), .B1(n4199), .C0(n540), 
        .C1(cacheDataOut[1]), .Y(n2242) );
  NAND4X1TS U3686 ( .A(n2236), .B(n2237), .C(n2238), .D(n2239), .Y(n2428) );
  AOI221X1TS U3687 ( .A0(n1023), .A1(n3185), .B0(n1007), .B1(n662), .C0(n2240), 
        .Y(n2239) );
  AOI222XLTS U3688 ( .A0(n935), .A1(n669), .B0(n763), .B1(n3122), .C0(n554), 
        .C1(n3120), .Y(n2238) );
  AOI222XLTS U3689 ( .A0(n1069), .A1(n4389), .B0(n1088), .B1(n4196), .C0(n540), 
        .C1(cacheDataOut[0]), .Y(n2236) );
  NAND4X1TS U3690 ( .A(n2230), .B(n2231), .C(n2232), .D(n2233), .Y(n2429) );
  AOI221X1TS U3691 ( .A0(n1024), .A1(n3007), .B0(n1008), .B1(
        \requesterAddressbuffer[2][5] ), .C0(n2234), .Y(n2233) );
  AOI222XLTS U3692 ( .A0(n937), .A1(\requesterAddressbuffer[0][5] ), .B0(n765), 
        .B1(\requesterAddressbuffer[6][5] ), .C0(n555), .C1(n3030), .Y(n2232)
         );
  AOI222XLTS U3693 ( .A0(n1070), .A1(n4499), .B0(n1087), .B1(n4031), .C0(n541), 
        .C1(readRequesterAddress[5]), .Y(n2230) );
  NAND4X1TS U3694 ( .A(n2224), .B(n2225), .C(n2226), .D(n2227), .Y(n2430) );
  AOI221X1TS U3695 ( .A0(n1024), .A1(n3008), .B0(n1008), .B1(
        \requesterAddressbuffer[2][4] ), .C0(n2228), .Y(n2227) );
  AOI222XLTS U3696 ( .A0(n937), .A1(\requesterAddressbuffer[0][4] ), .B0(n765), 
        .B1(\requesterAddressbuffer[6][4] ), .C0(n555), .C1(n3031), .Y(n2226)
         );
  AOI222XLTS U3697 ( .A0(n1070), .A1(n4496), .B0(n1087), .B1(n4028), .C0(n541), 
        .C1(readRequesterAddress[4]), .Y(n2224) );
  NAND4X1TS U3698 ( .A(n2212), .B(n2213), .C(n2214), .D(n2215), .Y(n2432) );
  AOI221X1TS U3699 ( .A0(n1024), .A1(n3009), .B0(n1008), .B1(
        \requesterAddressbuffer[2][2] ), .C0(n2216), .Y(n2215) );
  AOI222XLTS U3700 ( .A0(n937), .A1(\requesterAddressbuffer[0][2] ), .B0(n765), 
        .B1(\requesterAddressbuffer[6][2] ), .C0(n555), .C1(n3032), .Y(n2214)
         );
  AOI222XLTS U3701 ( .A0(n1070), .A1(n4490), .B0(n1087), .B1(n4022), .C0(n541), 
        .C1(readRequesterAddress[2]), .Y(n2212) );
  NAND4X1TS U3702 ( .A(n2206), .B(n2207), .C(n2208), .D(n2209), .Y(n2433) );
  AOI221X1TS U3703 ( .A0(n1025), .A1(n3010), .B0(n1009), .B1(
        \requesterAddressbuffer[2][1] ), .C0(n2210), .Y(n2209) );
  AOI222XLTS U3704 ( .A0(n938), .A1(\requesterAddressbuffer[0][1] ), .B0(n768), 
        .B1(\requesterAddressbuffer[6][1] ), .C0(n556), .C1(n3033), .Y(n2208)
         );
  AOI222XLTS U3705 ( .A0(n1071), .A1(n4487), .B0(n1086), .B1(n4019), .C0(n542), 
        .C1(readRequesterAddress[1]), .Y(n2206) );
  NAND4X1TS U3706 ( .A(n2194), .B(n2195), .C(n2196), .D(n2197), .Y(n2435) );
  AOI221X1TS U3707 ( .A0(n1025), .A1(n3186), .B0(n1009), .B1(n695), .C0(n2198), 
        .Y(n2197) );
  AOI222XLTS U3708 ( .A0(n938), .A1(n36), .B0(n768), .B1(n3124), .C0(n556), 
        .C1(n3123), .Y(n2196) );
  AOI222XLTS U3709 ( .A0(n1071), .A1(n4170), .B0(n1086), .B1(n3991), .C0(n542), 
        .C1(readRequesterAddress[5]), .Y(n2194) );
  NAND4X1TS U3710 ( .A(n2188), .B(n2189), .C(n2190), .D(n2191), .Y(n2436) );
  AOI221X1TS U3711 ( .A0(n1025), .A1(n3187), .B0(n1009), .B1(n694), .C0(n2192), 
        .Y(n2191) );
  AOI222XLTS U3712 ( .A0(n938), .A1(n90), .B0(n768), .B1(n3126), .C0(n556), 
        .C1(n3125), .Y(n2190) );
  AOI222XLTS U3713 ( .A0(n1071), .A1(n4167), .B0(n1086), .B1(n3988), .C0(n542), 
        .C1(readRequesterAddress[4]), .Y(n2188) );
  NAND4X1TS U3714 ( .A(n2182), .B(n2183), .C(n2184), .D(n2185), .Y(n2437) );
  AOI221X1TS U3715 ( .A0(n1026), .A1(n3188), .B0(n1010), .B1(n693), .C0(n2186), 
        .Y(n2185) );
  AOI222XLTS U3716 ( .A0(n959), .A1(n37), .B0(n770), .B1(n3129), .C0(n557), 
        .C1(n3127), .Y(n2184) );
  AOI222XLTS U3717 ( .A0(n1072), .A1(n4164), .B0(n1089), .B1(n3985), .C0(n543), 
        .C1(readRequesterAddress[3]), .Y(n2182) );
  NAND4X1TS U3718 ( .A(n2176), .B(n2177), .C(n2178), .D(n2179), .Y(n2438) );
  AOI221X1TS U3719 ( .A0(n1026), .A1(n3189), .B0(n1010), .B1(n746), .C0(n2180), 
        .Y(n2179) );
  AOI222XLTS U3720 ( .A0(n959), .A1(n38), .B0(n770), .B1(n3131), .C0(n557), 
        .C1(n3130), .Y(n2178) );
  AOI222XLTS U3721 ( .A0(n1072), .A1(n4161), .B0(n1085), .B1(n3982), .C0(n543), 
        .C1(readRequesterAddress[2]), .Y(n2176) );
  NAND4X1TS U3722 ( .A(n2170), .B(n2171), .C(n2172), .D(n2173), .Y(n2439) );
  AOI221X1TS U3723 ( .A0(n1026), .A1(n3190), .B0(n1010), .B1(n692), .C0(n2174), 
        .Y(n2173) );
  AOI222XLTS U3724 ( .A0(n959), .A1(n39), .B0(n770), .B1(n3133), .C0(n557), 
        .C1(n3132), .Y(n2172) );
  AOI222XLTS U3725 ( .A0(n1072), .A1(n4158), .B0(n1085), .B1(n3979), .C0(n543), 
        .C1(readRequesterAddress[1]), .Y(n2170) );
  NAND4X1TS U3726 ( .A(n2156), .B(n2157), .C(n2158), .D(n2159), .Y(n2440) );
  AOI221X1TS U3727 ( .A0(n1026), .A1(n3192), .B0(n1010), .B1(n691), .C0(n2162), 
        .Y(n2159) );
  AOI222XLTS U3728 ( .A0(n959), .A1(n91), .B0(n770), .B1(n3135), .C0(n557), 
        .C1(n3134), .Y(n2158) );
  AOI222XLTS U3729 ( .A0(n1072), .A1(n4155), .B0(n1085), .B1(n3976), .C0(n543), 
        .C1(readRequesterAddress[0]), .Y(n2156) );
  NAND4X1TS U3730 ( .A(n2218), .B(n2219), .C(n2220), .D(n2221), .Y(n2431) );
  AOI221X1TS U3731 ( .A0(n1024), .A1(n3012), .B0(n1008), .B1(
        \requesterAddressbuffer[2][3] ), .C0(n2222), .Y(n2221) );
  AOI222XLTS U3732 ( .A0(n937), .A1(\requesterAddressbuffer[0][3] ), .B0(n765), 
        .B1(\requesterAddressbuffer[6][3] ), .C0(n555), .C1(n3034), .Y(n2220)
         );
  AOI222XLTS U3733 ( .A0(n1070), .A1(n4493), .B0(n1087), .B1(n4025), .C0(n541), 
        .C1(readRequesterAddress[3]), .Y(n2218) );
  NAND4X1TS U3734 ( .A(n2200), .B(n2201), .C(n2202), .D(n2203), .Y(n2434) );
  AOI221X1TS U3735 ( .A0(n1025), .A1(n3013), .B0(n1009), .B1(
        \requesterAddressbuffer[2][0] ), .C0(n2204), .Y(n2203) );
  AOI222XLTS U3736 ( .A0(n938), .A1(\requesterAddressbuffer[0][0] ), .B0(n768), 
        .B1(\requesterAddressbuffer[6][0] ), .C0(n556), .C1(n3035), .Y(n2202)
         );
  AOI222XLTS U3737 ( .A0(n1071), .A1(n4484), .B0(n1086), .B1(n4016), .C0(n542), 
        .C1(readRequesterAddress[0]), .Y(n2200) );
  INVX2TS U3738 ( .A(writeIn_NORTH), .Y(n982) );
  AO21X1TS U3739 ( .A0(n939), .A1(n2089), .B0(n2090), .Y(n2088) );
  OAI33XLTS U3740 ( .A0(n2288), .A1(n2064), .A2(n2065), .B0(n2091), .B1(n4504), 
        .B2(n936), .Y(n2090) );
  NOR4XLTS U3741 ( .A(n2092), .B(n2093), .C(n2094), .D(n2095), .Y(n2091) );
  INVX2TS U3742 ( .A(n2089), .Y(n936) );
  OAI32X1TS U3743 ( .A0(n2286), .A1(n2064), .A2(n2065), .B0(n2066), .B1(n2067), 
        .Y(n2450) );
  NOR4BX1TS U3744 ( .AN(n2075), .B(n2076), .C(n2077), .D(n2078), .Y(n2066) );
  OAI31X1TS U3745 ( .A0(n2068), .A1(n443), .A2(n2069), .B0(n4503), .Y(n2067)
         );
  OAI22X1TS U3746 ( .A0(n2082), .A1(n752), .B0(n2083), .B1(n649), .Y(n2076) );
  OAI211X1TS U3747 ( .A0(n3974), .A1(n1044), .B0(n2148), .C0(n2149), .Y(n2441)
         );
  AOI22X1TS U3748 ( .A0(n153), .A1(n2150), .B0(n1113), .B1(
        destinationAddressOut[13]), .Y(n2148) );
  AOI222XLTS U3749 ( .A0(n1073), .A1(n4194), .B0(n1050), .B1(
        destinationAddressIn_NORTH[13]), .C0(n1083), .C1(
        destinationAddressIn_WEST[13]), .Y(n2149) );
  NAND4X1TS U3750 ( .A(n2151), .B(n2152), .C(n2153), .D(n2154), .Y(n2150) );
  OAI211X1TS U3751 ( .A0(n3971), .A1(n1044), .B0(n2141), .C0(n2142), .Y(n2442)
         );
  AOI22X1TS U3752 ( .A0(n240), .A1(n2143), .B0(n1113), .B1(
        destinationAddressOut[12]), .Y(n2141) );
  AOI222XLTS U3753 ( .A0(n1073), .A1(n4191), .B0(n1050), .B1(
        destinationAddressIn_NORTH[12]), .C0(n1083), .C1(
        destinationAddressIn_WEST[12]), .Y(n2142) );
  NAND4X1TS U3754 ( .A(n2144), .B(n2145), .C(n2146), .D(n2147), .Y(n2143) );
  OAI211X1TS U3755 ( .A0(n3968), .A1(n1044), .B0(n2134), .C0(n2135), .Y(n2443)
         );
  AOI22X1TS U3756 ( .A0(n242), .A1(n2136), .B0(n1113), .B1(
        destinationAddressOut[11]), .Y(n2134) );
  AOI222XLTS U3757 ( .A0(n1073), .A1(n4188), .B0(n1050), .B1(
        destinationAddressIn_NORTH[11]), .C0(n1083), .C1(
        destinationAddressIn_WEST[11]), .Y(n2135) );
  NAND4X1TS U3758 ( .A(n2137), .B(n2138), .C(n2139), .D(n2140), .Y(n2136) );
  OAI211X1TS U3759 ( .A0(n3965), .A1(n1045), .B0(n2127), .C0(n2128), .Y(n2444)
         );
  AOI22X1TS U3760 ( .A0(n240), .A1(n2129), .B0(n1113), .B1(
        destinationAddressOut[10]), .Y(n2127) );
  AOI222XLTS U3761 ( .A0(n1073), .A1(n4185), .B0(n1050), .B1(
        destinationAddressIn_NORTH[10]), .C0(n1082), .C1(
        destinationAddressIn_WEST[10]), .Y(n2128) );
  NAND4X1TS U3762 ( .A(n2130), .B(n2131), .C(n2132), .D(n2133), .Y(n2129) );
  OAI211X1TS U3763 ( .A0(n3962), .A1(n1045), .B0(n2120), .C0(n2121), .Y(n2445)
         );
  AOI22X1TS U3764 ( .A0(n154), .A1(n2122), .B0(n1114), .B1(
        destinationAddressOut[9]), .Y(n2120) );
  AOI222XLTS U3765 ( .A0(n1081), .A1(n4182), .B0(n1049), .B1(
        destinationAddressIn_NORTH[9]), .C0(n1083), .C1(
        destinationAddressIn_WEST[9]), .Y(n2121) );
  NAND4X1TS U3766 ( .A(n2123), .B(n2124), .C(n2125), .D(n2126), .Y(n2122) );
  OAI211X1TS U3767 ( .A0(n3959), .A1(n1045), .B0(n2113), .C0(n2114), .Y(n2446)
         );
  AOI22X1TS U3768 ( .A0(n241), .A1(n2115), .B0(n1114), .B1(
        destinationAddressOut[8]), .Y(n2113) );
  AOI222XLTS U3769 ( .A0(n1081), .A1(n4179), .B0(n1049), .B1(
        destinationAddressIn_NORTH[8]), .C0(n1082), .C1(
        destinationAddressIn_WEST[8]), .Y(n2114) );
  NAND4X1TS U3770 ( .A(n2116), .B(n2117), .C(n2118), .D(n2119), .Y(n2115) );
  OAI211X1TS U3771 ( .A0(n3956), .A1(n1046), .B0(n2106), .C0(n2107), .Y(n2447)
         );
  AOI22X1TS U3772 ( .A0(n1131), .A1(n2108), .B0(n1114), .B1(
        destinationAddressOut[7]), .Y(n2106) );
  AOI222XLTS U3773 ( .A0(n1081), .A1(n4176), .B0(n1049), .B1(
        destinationAddressIn_NORTH[7]), .C0(n1082), .C1(
        destinationAddressIn_WEST[7]), .Y(n2107) );
  NAND4X1TS U3774 ( .A(n2109), .B(n2110), .C(n2111), .D(n2112), .Y(n2108) );
  OAI211X1TS U3775 ( .A0(n3953), .A1(n1046), .B0(n2098), .C0(n2099), .Y(n2448)
         );
  AOI22X1TS U3776 ( .A0(n241), .A1(n2101), .B0(n1114), .B1(
        destinationAddressOut[6]), .Y(n2098) );
  AOI222XLTS U3777 ( .A0(n1080), .A1(n4173), .B0(n1049), .B1(
        destinationAddressIn_NORTH[6]), .C0(n1082), .C1(
        destinationAddressIn_WEST[6]), .Y(n2099) );
  NAND4X1TS U3778 ( .A(n2102), .B(n2103), .C(n2104), .D(n2105), .Y(n2101) );
  INVX2TS U3779 ( .A(readIn_SOUTH), .Y(n996) );
  INVX2TS U3780 ( .A(readIn_NORTH), .Y(n981) );
  INVX2TS U3781 ( .A(destinationAddressIn_NORTH[7]), .Y(n979) );
  INVX2TS U3782 ( .A(destinationAddressIn_NORTH[6]), .Y(n980) );
  OAI21X1TS U3783 ( .A0(n126), .A1(n1141), .B0(n4502), .Y(n1143) );
  AO22X1TS U3784 ( .A0(n939), .A1(n11), .B0(n160), .B1(n154), .Y(n2889) );
  NOR2X1TS U3785 ( .A(n1145), .B(n1143), .Y(n2883) );
  AOI21X1TS U3786 ( .A0(n166), .A1(n153), .B0(n165), .Y(n1145) );
  XNOR2X1TS U3787 ( .A(n2990), .B(n1142), .Y(n2988) );
  OAI22X1TS U3788 ( .A0(n165), .A1(n2991), .B0(n2994), .B1(n9), .Y(n2990) );
  NOR2X1TS U3789 ( .A(n758), .B(n125), .Y(n2994) );
  NAND3X1TS U3790 ( .A(n125), .B(n11), .C(n8), .Y(n2079) );
  NAND2X1TS U3791 ( .A(n123), .B(n199), .Y(n1985) );
  AO22X1TS U3792 ( .A0(n3271), .A1(n234), .B0(n3270), .B1(n237), .Y(n2093) );
  AOI21X1TS U3793 ( .A0(n166), .A1(n439), .B0(n758), .Y(n1138) );
  AOI22X1TS U3794 ( .A0(n436), .A1(n3280), .B0(n448), .B1(n3326), .Y(n2151) );
  AOI22X1TS U3795 ( .A0(n436), .A1(n3281), .B0(n448), .B1(n3325), .Y(n2144) );
  AOI22X1TS U3796 ( .A0(n436), .A1(n3282), .B0(n448), .B1(n3324), .Y(n2137) );
  AOI22X1TS U3797 ( .A0(n436), .A1(n3283), .B0(n448), .B1(n3323), .Y(n2130) );
  AOI22X1TS U3798 ( .A0(n437), .A1(n3284), .B0(n449), .B1(n3322), .Y(n2123) );
  AOI22X1TS U3799 ( .A0(n437), .A1(n3285), .B0(n449), .B1(n3321), .Y(n2116) );
  AOI22X1TS U3800 ( .A0(n437), .A1(n3286), .B0(n449), .B1(n3320), .Y(n2109) );
  AOI22X1TS U3801 ( .A0(n437), .A1(n3287), .B0(n449), .B1(n3319), .Y(n2102) );
  AOI22X1TS U3802 ( .A0(n175), .A1(n3272), .B0(n201), .B1(n3334), .Y(n2154) );
  AOI22X1TS U3803 ( .A0(n176), .A1(n3273), .B0(n762), .B1(n3333), .Y(n2147) );
  AOI22X1TS U3804 ( .A0(n175), .A1(n3274), .B0(n202), .B1(n3332), .Y(n2140) );
  AOI22X1TS U3805 ( .A0(n176), .A1(n3275), .B0(n201), .B1(n3331), .Y(n2133) );
  AOI22X1TS U3806 ( .A0(n175), .A1(n3276), .B0(n762), .B1(n3330), .Y(n2126) );
  AOI22X1TS U3807 ( .A0(n176), .A1(n3277), .B0(n202), .B1(n3329), .Y(n2119) );
  AOI22X1TS U3808 ( .A0(n175), .A1(n3278), .B0(n201), .B1(n3328), .Y(n2112) );
  AOI22X1TS U3809 ( .A0(n176), .A1(n3279), .B0(n762), .B1(n3327), .Y(n2105) );
  AOI22X1TS U3810 ( .A0(n178), .A1(n3304), .B0(n3303), .B1(n223), .Y(n2152) );
  AOI22X1TS U3811 ( .A0(n179), .A1(n3306), .B0(n3305), .B1(n222), .Y(n2145) );
  AOI22X1TS U3812 ( .A0(n179), .A1(n3308), .B0(n3307), .B1(n2096), .Y(n2138)
         );
  AOI22X1TS U3813 ( .A0(n178), .A1(n3310), .B0(n3309), .B1(n223), .Y(n2131) );
  AOI22X1TS U3814 ( .A0(n178), .A1(n3312), .B0(n3311), .B1(n222), .Y(n2124) );
  AOI22X1TS U3815 ( .A0(n179), .A1(n3314), .B0(n3313), .B1(n2096), .Y(n2117)
         );
  AOI22X1TS U3816 ( .A0(n178), .A1(n3316), .B0(n3315), .B1(n223), .Y(n2110) );
  AOI22X1TS U3817 ( .A0(n179), .A1(n3318), .B0(n3317), .B1(n222), .Y(n2103) );
  AOI22X1TS U3818 ( .A0(n237), .A1(n3289), .B0(n235), .B1(n3288), .Y(n2153) );
  AOI22X1TS U3819 ( .A0(n2084), .A1(n3291), .B0(n234), .B1(n3290), .Y(n2146)
         );
  AOI22X1TS U3820 ( .A0(n238), .A1(n3293), .B0(n753), .B1(n3292), .Y(n2139) );
  AOI22X1TS U3821 ( .A0(n237), .A1(n593), .B0(n235), .B1(n3294), .Y(n2132) );
  AOI22X1TS U3822 ( .A0(n2084), .A1(n3296), .B0(n234), .B1(n3295), .Y(n2125)
         );
  AOI22X1TS U3823 ( .A0(n238), .A1(n3298), .B0(n753), .B1(n3297), .Y(n2118) );
  AOI22X1TS U3824 ( .A0(n237), .A1(n3300), .B0(n235), .B1(n3299), .Y(n2111) );
  AOI22X1TS U3825 ( .A0(n2084), .A1(n3302), .B0(n234), .B1(n3301), .Y(n2104)
         );
  AOI221X1TS U3826 ( .A0(n202), .A1(\readOutbuffer[2] ), .B0(n238), .B1(
        readOutbuffer_7), .C0(n13), .Y(n2075) );
  AOI21XLTS U3827 ( .A0(n4142), .A1(n946), .B0(n134), .Y(n1809) );
  AOI32XLTS U3828 ( .A0(n132), .A1(n1824), .A2(n1825), .B0(n3576), .B1(n650), 
        .Y(n2568) );
  AOI32XLTS U3829 ( .A0(n447), .A1(n1827), .A2(n4147), .B0(n1828), .B1(n1829), 
        .Y(n1825) );
  AOI32XLTS U3830 ( .A0(n25), .A1(n1839), .A2(n1840), .B0(n3858), .B1(n648), 
        .Y(n2566) );
  OAI221XLTS U3831 ( .A0(n217), .A1(n185), .B0(n518), .B1(n592), .C0(n1976), 
        .Y(n2500) );
  OAI221XLTS U3832 ( .A0(n216), .A1(n182), .B0(n517), .B1(n578), .C0(n1977), 
        .Y(n2499) );
  OAI221XLTS U3833 ( .A0(n217), .A1(n197), .B0(n518), .B1(n589), .C0(n1978), 
        .Y(n2498) );
  OAI221XLTS U3834 ( .A0(n216), .A1(n190), .B0(n517), .B1(n590), .C0(n1979), 
        .Y(n2497) );
  OAI221XLTS U3835 ( .A0(n217), .A1(n195), .B0(n518), .B1(n579), .C0(n1980), 
        .Y(n2496) );
  OAI221XLTS U3836 ( .A0(n216), .A1(n189), .B0(n517), .B1(n594), .C0(n1981), 
        .Y(n2495) );
  OAI221XLTS U3837 ( .A0(n217), .A1(n193), .B0(n518), .B1(n591), .C0(n1982), 
        .Y(n2494) );
  OAI221XLTS U3838 ( .A0(n216), .A1(n186), .B0(n517), .B1(n580), .C0(n1983), 
        .Y(n2493) );
  OAI221XLTS U3839 ( .A0(n215), .A1(n204), .B0(n516), .B1(n748), .C0(n1799), 
        .Y(n2574) );
  AOI32XLTS U3840 ( .A0(n1841), .A1(n1842), .A2(n4147), .B0(n1843), .B1(n1844), 
        .Y(n1840) );
  AND3X2TS U3841 ( .A(n1843), .B(n139), .C(n25), .Y(n1217) );
  AOI32XLTS U3842 ( .A0(n137), .A1(n1831), .A2(n1832), .B0(n3787), .B1(n752), 
        .Y(n2567) );
  AOI21XLTS U3843 ( .A0(readIn_NORTH), .A1(n1833), .B0(n1834), .Y(n1832) );
  OAI221XLTS U3844 ( .A0(n231), .A1(n184), .B0(n151), .B1(n605), .C0(n1953), 
        .Y(n2514) );
  OAI221XLTS U3845 ( .A0(n1794), .A1(n182), .B0(n150), .B1(n606), .C0(n1954), 
        .Y(n2513) );
  OAI221XLTS U3846 ( .A0(n231), .A1(n196), .B0(n151), .B1(n607), .C0(n1955), 
        .Y(n2512) );
  OAI221XLTS U3847 ( .A0(n1794), .A1(n190), .B0(n150), .B1(n599), .C0(n1956), 
        .Y(n2511) );
  OAI221XLTS U3848 ( .A0(n231), .A1(n195), .B0(n151), .B1(n608), .C0(n1957), 
        .Y(n2510) );
  OAI221XLTS U3849 ( .A0(n1794), .A1(n188), .B0(n1795), .B1(n609), .C0(n1958), 
        .Y(n2509) );
  OAI221XLTS U3850 ( .A0(n231), .A1(n193), .B0(n1795), .B1(n610), .C0(n1959), 
        .Y(n2508) );
  OAI221XLTS U3851 ( .A0(n230), .A1(n187), .B0(n150), .B1(n600), .C0(n1960), 
        .Y(n2507) );
  OAI221XLTS U3852 ( .A0(n230), .A1(n982), .B0(n1795), .B1(n750), .C0(n1796), 
        .Y(n2575) );
endmodule


module outputPortArbiter_3 ( clk, reset, selectBit_NORTH, 
        destinationAddressIn_NORTH, requesterAddressIn_NORTH, readIn_NORTH, 
        writeIn_NORTH, dataIn_NORTH, selectBit_SOUTH, 
        destinationAddressIn_SOUTH, requesterAddressIn_SOUTH, readIn_SOUTH, 
        writeIn_SOUTH, dataIn_SOUTH, selectBit_EAST, destinationAddressIn_EAST, 
        requesterAddressIn_EAST, readIn_EAST, writeIn_EAST, dataIn_EAST, 
        selectBit_WEST, destinationAddressIn_WEST, requesterAddressIn_WEST, 
        readIn_WEST, dataIn_WEST, readReady, readRequesterAddress, 
        cacheDataOut, destinationAddressOut, requesterAddressOut, readOut, 
        writeOut, dataOut, writeIn_WEST_BAR );
  input [13:0] destinationAddressIn_NORTH;
  input [5:0] requesterAddressIn_NORTH;
  input [31:0] dataIn_NORTH;
  input [13:0] destinationAddressIn_SOUTH;
  input [5:0] requesterAddressIn_SOUTH;
  input [31:0] dataIn_SOUTH;
  input [13:0] destinationAddressIn_EAST;
  input [5:0] requesterAddressIn_EAST;
  input [31:0] dataIn_EAST;
  input [13:0] destinationAddressIn_WEST;
  input [5:0] requesterAddressIn_WEST;
  input [31:0] dataIn_WEST;
  input [5:0] readRequesterAddress;
  input [31:0] cacheDataOut;
  output [13:0] destinationAddressOut;
  output [5:0] requesterAddressOut;
  output [31:0] dataOut;
  input clk, reset, selectBit_NORTH, readIn_NORTH, writeIn_NORTH,
         selectBit_SOUTH, readIn_SOUTH, writeIn_SOUTH, selectBit_EAST,
         readIn_EAST, writeIn_EAST, selectBit_WEST, readIn_WEST, readReady,
         writeIn_WEST_BAR;
  output readOut, writeOut;
  wire   writeIn_WEST, n2457, n2458, n2456, n2499, n2496, n2493, n2528, n2527,
         n2526, n2525, n2524, n2523, n2522, n2521, n2498, n2497, n2494, n2500,
         n2495, n2541, n2540, n2537, n2535, n2511, n2507, n2556, n2555, n2554,
         n2552, n4796, n2551, n2550, n2549, n2553, n2542, n2539, n2538, n2536,
         n2514, n2513, n2512, n2510, n2509, n2508, n2638, n2544, n2609, n2608,
         n2607, n2606, n2605, n2604, n2603, n2602, n2601, n2600, n2599, n2598,
         n2594, n2593, n2592, n2591, n2590, n2589, n2588, n2587, n2586, n2585,
         n2584, n2583, n2582, n2581, n2580, n2579, n2561, n2560, n2559, n2557,
         n2642, n2640, n2639, n2637, n2635, n2634, n2633, n2631, n2612, n2611,
         n2562, n2558, n2641, n2636, n2632, n2548, n2547, n2546, n2545, n2543,
         n2876, \requesterAddressbuffer[6][0] , n2875,
         \requesterAddressbuffer[6][1] , n2874, \requesterAddressbuffer[6][2] ,
         n2873, \requesterAddressbuffer[6][3] , n2872,
         \requesterAddressbuffer[6][4] , n2871, \requesterAddressbuffer[6][5] ,
         n2850, \requesterAddressbuffer[2][2] , n2849,
         \requesterAddressbuffer[2][3] , n2847, \requesterAddressbuffer[2][5] ,
         n2840, \requesterAddressbuffer[0][0] , n2839,
         \requesterAddressbuffer[0][1] , n2838, \requesterAddressbuffer[0][2] ,
         n2836, \requesterAddressbuffer[0][4] , n2852,
         \requesterAddressbuffer[2][0] , n2851, \requesterAddressbuffer[2][1] ,
         n2848, \requesterAddressbuffer[2][4] , n2837,
         \requesterAddressbuffer[0][3] , n2835, \requesterAddressbuffer[0][5] ,
         n2566, \readOutbuffer[2] , readOutbuffer_7, n2569, n2578, n2568,
         n2564, n2563, n2882, n2881, n2879, n2576, n2880, n2878, n2877, n2770,
         n2768, n2764, n2754, n99, n2748, n98, n2746, n97, n2739, n96, n2834,
         n64, n2833, n63, n2832, n62, n2829, n61, n2825, n60, n2814, n59,
         n2811, n58, n2807, n57, n2806, n56, n2769, n95, n2760, n94, n2743,
         n93, n2492, n92, n2491, n91, n2489, n90, n2488, n89, n2487, n88,
         n2464, n55, n2460, n54, n2767, n87, n2766, n86, n2765, n85, n2763,
         n84, n2762, n83, n2761, n82, n2759, n81, n2758, n80, n2757, n79,
         n2756, n78, n2755, n77, n2753, n76, n2752, n75, n2751, n74, n2750,
         n73, n2749, n72, n2747, n71, n2745, n70, n2744, n69, n2742, n68,
         n2741, n67, n2740, n66, n2490, n65, n2831, n53, n2830, n52, n2828,
         n51, n2827, n50, n2826, n49, n2824, n48, n2823, n47, n2822, n46,
         n2821, n4592, n2820, n4579, n2819, n4572, n2818, n4561, n2817, n4552,
         n2816, n4543, n2815, n4534, n2813, n4520, n2812, n4505, n2810, n4489,
         n2809, n4480, n2808, n4473, n2805, n4448, n2804, n4437, n2803, n4424,
         n2463, n4752, n2462, n4747, n2461, n4736, n2459, n4716, n2571, n2574,
         n2577, n2575, n2570, n2565, n2567, n2889, n8, n2887, n5323, n4833,
         n2434, n4837, n2431, n4838, n2450, n4835, n2440, n4760, n2439, n4751,
         n2438, n4742, n2437, n4733, n2436, n4724, n2435, n4715, n2433, n4714,
         n2432, n4713, n2430, n4712, n2429, n4711, n2428, n4702, n2427, n4693,
         n2426, n4684, n2425, n4675, n2424, n4666, n2423, n4657, n2422, n4648,
         n2421, n4639, n2420, n4630, n2419, n4621, n2418, n4612, n2417, n4603,
         n2416, n4594, n2415, n4585, n2414, n4576, n2413, n4567, n2412, n4558,
         n2411, n4549, n2410, n4540, n2409, n4531, n2408, n4522, n2407, n4513,
         n2406, n4504, n2405, n4495, n2404, n4486, n2403, n4477, n2402, n4468,
         n2401, n4459, n2400, n4450, n2399, n4441, n2398, n4432, n2397, n4423,
         n2448, n2447, n2446, n2445, n2444, n2443, n2442, n2441, n2486, n2484,
         n2485, n2472, n2471, n2470, n2469, n2468, n2467, n2466, n2465, n2530,
         n2674, n2672, n2671, n2670, n2669, n2668, n2667, n2666, n2665, n2664,
         n2662, n2661, n2660, n2657, n2656, n2655, n2654, n2653, n2652, n2651,
         n2650, n2649, n2648, n2647, n2646, n2645, n2644, n2534, n2533, n2532,
         n2531, n2529, n2673, n2663, n2659, n2658, n2643, n2516, n2703, n2692,
         n2691, n2689, n2802, n2706, n2705, n2700, n2698, n2696, n2695, n2694,
         n2690, n2687, n2686, n2685, n2684, n2677, n2675, n2801, n2799, n2798,
         n2796, n2795, n2793, n2791, n2790, n2789, n2788, n2787, n2786, n2785,
         n2784, n2781, n2779, n2778, n2777, n2776, n2774, n2773, n2772, n2771,
         n2478, n2477, n2476, n2475, n2473, n2704, n2702, n2701, n2699, n2697,
         n2693, n2688, n2683, n2682, n2681, n2680, n2679, n2678, n2676, n2520,
         n2519, n2518, n2517, n2515, n2800, n2797, n2794, n2792, n2783, n2782,
         n2780, n2775, n2474, n2731, n6312, n2736, n6302, n2734, n6301, n2733,
         n6300, n2725, n6299, n2723, n6298, n2720, n6297, n2718, n6296, n2715,
         n6295, n2713, n6294, n2504, n6293, n2738, n6281, n2737, n6280, n2735,
         n6279, n2732, n6278, n2730, n6277, n2729, n6276, n2728, n6275, n2727,
         n6274, n2726, n6273, n2724, n6272, n2722, n6271, n2721, n6270, n2719,
         n6269, n2717, n6268, n2716, n6267, n2714, n6266, n2712, n6265, n2711,
         n6264, n2710, n6263, n2709, n6262, n2708, n6261, n2707, n6260, n2506,
         n6259, n2505, n6258, n2503, n6257, n2502, n6256, n2501, n6255, n2858,
         \requesterAddressbuffer[3][0] , n2857, \requesterAddressbuffer[3][1] ,
         n2856, \requesterAddressbuffer[3][2] , n2855,
         \requesterAddressbuffer[3][3] , n2853, \requesterAddressbuffer[3][5] ,
         n2854, \requesterAddressbuffer[3][4] , n2870, n2869, n2868, n2867,
         n2866, n2865, n2860, n2859, n2864, n2863, n2862, n2861, n2846, n2845,
         n2844, n2843, n2842, n2841, n2455, n2453, n2454, n2452, n2573, n2572,
         n2883, n2884, N4718, n6347, n2479, n2451, n2480, n2481, n2482, n2483,
         n2885, n6253, n2888, n5327, n2886, n2610, n2595, n2596, n2597, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n719, n720, n722,
         n724, n728, n730, n732, n734, n735, n736, n739, n740, n741, n742,
         n745, n746, n747, n748, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n927,
         n929, n930, n931, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n957, n958, n959, n960, n966, n967, n968, n969,
         n970, n971, n972, n973, n1028, n1083, n1086, n1087, n1088, n1089,
         n1090, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2449, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
         n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
         n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
         n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
         n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
         n3007, n3008, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n1, n2, n3, n4, n5, n6, n7, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n718, n721, n723, n725,
         n726, n727, n729, n731, n733, n737, n738, n743, n744, n749, n762,
         n912, n913, n924, n925, n926, n928, n932, n933, n956, n961, n962,
         n963, n964, n965, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1084, n1085,
         n1091, n1107, n1134, n1151, n1167, n1198, n1215, n1751, n1798, n1939,
         n2109, n2905, n2906, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n3009, n3010, n3011, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3152, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4433, n4434, n4435, n4436,
         n4438, n4439, n4440, n4442, n4443, n4444, n4445, n4446, n4447, n4449,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4469, n4470, n4471, n4472,
         n4474, n4475, n4476, n4478, n4479, n4481, n4482, n4483, n4484, n4485,
         n4487, n4488, n4490, n4491, n4492, n4493, n4494, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4514, n4515, n4516, n4517, n4518, n4519, n4521, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4532, n4533, n4535,
         n4536, n4537, n4538, n4539, n4541, n4542;
  assign writeIn_WEST = writeIn_WEST_BAR;

  AOI2BB1X4TS U1146 ( .A0N(n109), .A1N(n1914), .B0(n1790), .Y(n1786) );
  AO21X4TS U1147 ( .A0(n1844), .A1(n746), .B0(n1788), .Y(n1790) );
  DFFNSRX2TS \writeOutbuffer_reg[5]  ( .D(n2576), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n660) );
  DFFNSRX2TS \writeOutbuffer_reg[1]  ( .D(n2572), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n911) );
  DFFNSRX2TS \destinationAddressbuffer_reg[5][6]  ( .D(n2528), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3159), .QN(n559) );
  DFFNSRX2TS \destinationAddressbuffer_reg[5][7]  ( .D(n2527), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3157), .QN(n560) );
  DFFNSRX2TS \destinationAddressbuffer_reg[5][8]  ( .D(n2526), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3155), .QN(n561) );
  DFFNSRX2TS \destinationAddressbuffer_reg[1][6]  ( .D(n2472), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3137), .QN(n766) );
  DFFNSRX2TS \destinationAddressbuffer_reg[1][7]  ( .D(n2471), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3136), .QN(n767) );
  DFFNSRX2TS \destinationAddressbuffer_reg[1][8]  ( .D(n2470), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3134), .QN(n768) );
  DFFNSRX2TS empty_reg_reg ( .D(n2885), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        n6253), .QN(n469) );
  DFFNSRX2TS \read_reg_reg[1]  ( .D(n2883), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n5), .QN(n2) );
  DFFNSRX2TS \read_reg_reg[0]  ( .D(n2889), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n442), .QN(n8) );
  DFFNSRX2TS \read_reg_reg[2]  ( .D(n2884), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n913), .QN(n6) );
  DFFNSRX2TS \write_reg_reg[2]  ( .D(n2886), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1), .QN(n471) );
  DFFNSRX2TS writeOut_reg ( .D(n651), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        writeOut), .QN(n4833) );
  DFFNSRX2TS \requesterAddressOut_reg[0]  ( .D(n2434), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[0]), .QN(n4837) );
  DFFNSRX2TS \requesterAddressOut_reg[3]  ( .D(n2431), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[3]), .QN(n4838) );
  DFFNSRX2TS readOut_reg ( .D(n2450), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        readOut), .QN(n4835) );
  DFFNSRX2TS \destinationAddressOut_reg[0]  ( .D(n2440), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[0]), .QN(n4760) );
  DFFNSRX2TS \destinationAddressOut_reg[1]  ( .D(n2439), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[1]), .QN(n4751) );
  DFFNSRX2TS \destinationAddressOut_reg[2]  ( .D(n2438), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[2]), .QN(n4742) );
  DFFNSRX2TS \destinationAddressOut_reg[3]  ( .D(n2437), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[3]), .QN(n4733) );
  DFFNSRX2TS \destinationAddressOut_reg[4]  ( .D(n2436), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[4]), .QN(n4724) );
  DFFNSRX2TS \destinationAddressOut_reg[5]  ( .D(n2435), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[5]), .QN(n4715) );
  DFFNSRX2TS \requesterAddressOut_reg[1]  ( .D(n2433), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[1]), .QN(n4714) );
  DFFNSRX2TS \requesterAddressOut_reg[2]  ( .D(n2432), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[2]), .QN(n4713) );
  DFFNSRX2TS \requesterAddressOut_reg[4]  ( .D(n2430), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[4]), .QN(n4712) );
  DFFNSRX2TS \requesterAddressOut_reg[5]  ( .D(n2429), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[5]), .QN(n4711) );
  DFFNSRX2TS \dataOut_reg[0]  ( .D(n2428), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[0]), .QN(n4702) );
  DFFNSRX2TS \dataOut_reg[1]  ( .D(n2427), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[1]), .QN(n4693) );
  DFFNSRX2TS \dataOut_reg[2]  ( .D(n2426), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[2]), .QN(n4684) );
  DFFNSRX2TS \dataOut_reg[3]  ( .D(n2425), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[3]), .QN(n4675) );
  DFFNSRX2TS \dataOut_reg[4]  ( .D(n2424), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[4]), .QN(n4666) );
  DFFNSRX2TS \dataOut_reg[5]  ( .D(n2423), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[5]), .QN(n4657) );
  DFFNSRX2TS \dataOut_reg[6]  ( .D(n2422), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[6]), .QN(n4648) );
  DFFNSRX2TS \dataOut_reg[7]  ( .D(n2421), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[7]), .QN(n4639) );
  DFFNSRX2TS \dataOut_reg[8]  ( .D(n2420), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[8]), .QN(n4630) );
  DFFNSRX2TS \dataOut_reg[9]  ( .D(n2419), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[9]), .QN(n4621) );
  DFFNSRX2TS \dataOut_reg[10]  ( .D(n2418), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[10]), .QN(n4612) );
  DFFNSRX2TS \dataOut_reg[11]  ( .D(n2417), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[11]), .QN(n4603) );
  DFFNSRX2TS \dataOut_reg[12]  ( .D(n2416), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[12]), .QN(n4594) );
  DFFNSRX2TS \dataOut_reg[13]  ( .D(n2415), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[13]), .QN(n4585) );
  DFFNSRX2TS \dataOut_reg[14]  ( .D(n2414), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[14]), .QN(n4576) );
  DFFNSRX2TS \dataOut_reg[15]  ( .D(n2413), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[15]), .QN(n4567) );
  DFFNSRX2TS \dataOut_reg[16]  ( .D(n2412), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[16]), .QN(n4558) );
  DFFNSRX2TS \dataOut_reg[17]  ( .D(n2411), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[17]), .QN(n4549) );
  DFFNSRX2TS \dataOut_reg[18]  ( .D(n2410), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[18]), .QN(n4540) );
  DFFNSRX2TS \dataOut_reg[19]  ( .D(n2409), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[19]), .QN(n4531) );
  DFFNSRX2TS \dataOut_reg[20]  ( .D(n2408), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[20]), .QN(n4522) );
  DFFNSRX2TS \dataOut_reg[21]  ( .D(n2407), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[21]), .QN(n4513) );
  DFFNSRX2TS \dataOut_reg[22]  ( .D(n2406), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[22]), .QN(n4504) );
  DFFNSRX2TS \dataOut_reg[23]  ( .D(n2405), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[23]), .QN(n4495) );
  DFFNSRX2TS \dataOut_reg[24]  ( .D(n2404), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[24]), .QN(n4486) );
  DFFNSRX2TS \dataOut_reg[25]  ( .D(n2403), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[25]), .QN(n4477) );
  DFFNSRX2TS \dataOut_reg[26]  ( .D(n2402), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[26]), .QN(n4468) );
  DFFNSRX2TS \dataOut_reg[27]  ( .D(n2401), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[27]), .QN(n4459) );
  DFFNSRX2TS \dataOut_reg[28]  ( .D(n2400), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[28]), .QN(n4450) );
  DFFNSRX2TS \dataOut_reg[29]  ( .D(n2399), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[29]), .QN(n4441) );
  DFFNSRX2TS \dataOut_reg[30]  ( .D(n2398), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[30]), .QN(n4432) );
  DFFNSRX2TS \dataOut_reg[31]  ( .D(n2397), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[31]), .QN(n4423) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][4]  ( .D(n2558), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n639) );
  DFFNSRXLTS \dataoutbuffer_reg[7][1]  ( .D(n2609), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n596) );
  DFFNSRXLTS \dataoutbuffer_reg[7][2]  ( .D(n2608), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n597) );
  DFFNSRXLTS \dataoutbuffer_reg[7][3]  ( .D(n2607), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n598) );
  DFFNSRXLTS \dataoutbuffer_reg[7][4]  ( .D(n2606), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n599) );
  DFFNSRXLTS \dataoutbuffer_reg[7][5]  ( .D(n2605), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n600) );
  DFFNSRXLTS \dataoutbuffer_reg[7][6]  ( .D(n2604), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n601) );
  DFFNSRXLTS \dataoutbuffer_reg[7][7]  ( .D(n2603), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n602) );
  DFFNSRXLTS \dataoutbuffer_reg[7][8]  ( .D(n2602), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n603) );
  DFFNSRXLTS \dataoutbuffer_reg[7][9]  ( .D(n2601), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n604) );
  DFFNSRXLTS \dataoutbuffer_reg[7][10]  ( .D(n2600), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n605) );
  DFFNSRXLTS \dataoutbuffer_reg[7][11]  ( .D(n2599), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n606) );
  DFFNSRXLTS \dataoutbuffer_reg[7][12]  ( .D(n2598), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n607) );
  DFFNSRXLTS \dataoutbuffer_reg[7][16]  ( .D(n2594), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n608) );
  DFFNSRXLTS \dataoutbuffer_reg[7][17]  ( .D(n2593), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n609) );
  DFFNSRXLTS \dataoutbuffer_reg[7][18]  ( .D(n2592), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n610) );
  DFFNSRXLTS \dataoutbuffer_reg[7][19]  ( .D(n2591), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n611) );
  DFFNSRXLTS \dataoutbuffer_reg[7][20]  ( .D(n2590), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n612) );
  DFFNSRXLTS \dataoutbuffer_reg[7][21]  ( .D(n2589), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n613) );
  DFFNSRXLTS \dataoutbuffer_reg[7][22]  ( .D(n2588), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n614) );
  DFFNSRXLTS \dataoutbuffer_reg[7][23]  ( .D(n2587), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n615) );
  DFFNSRXLTS \dataoutbuffer_reg[7][24]  ( .D(n2586), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n616) );
  DFFNSRXLTS \dataoutbuffer_reg[7][25]  ( .D(n2585), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n617) );
  DFFNSRXLTS \dataoutbuffer_reg[7][26]  ( .D(n2584), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n618) );
  DFFNSRXLTS \dataoutbuffer_reg[7][27]  ( .D(n2583), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n619) );
  DFFNSRXLTS \dataoutbuffer_reg[7][28]  ( .D(n2582), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n620) );
  DFFNSRXLTS \dataoutbuffer_reg[7][29]  ( .D(n2581), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n621) );
  DFFNSRXLTS \dataoutbuffer_reg[7][30]  ( .D(n2580), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n622) );
  DFFNSRXLTS \dataoutbuffer_reg[7][31]  ( .D(n2579), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n623) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][1]  ( .D(n2561), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n624) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][2]  ( .D(n2560), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n625) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][3]  ( .D(n2559), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n626) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][5]  ( .D(n2557), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n627) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][0]  ( .D(n2562), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n638) );
  DFFNSRXLTS \requesterAddressbuffer_reg[7][0]  ( .D(n2882), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n657) );
  DFFNSRXLTS \requesterAddressbuffer_reg[7][1]  ( .D(n2881), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n658) );
  DFFNSRXLTS \requesterAddressbuffer_reg[7][3]  ( .D(n2879), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n659) );
  DFFNSRXLTS \requesterAddressbuffer_reg[7][2]  ( .D(n2880), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n661) );
  DFFNSRXLTS \requesterAddressbuffer_reg[7][4]  ( .D(n2878), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n662) );
  DFFNSRXLTS \requesterAddressbuffer_reg[7][5]  ( .D(n2877), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n663) );
  DFFNSRXLTS \dataoutbuffer_reg[7][0]  ( .D(n2610), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n934) );
  DFFNSRXLTS \dataoutbuffer_reg[7][15]  ( .D(n2595), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n935) );
  DFFNSRXLTS \dataoutbuffer_reg[7][14]  ( .D(n2596), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n936) );
  DFFNSRXLTS \dataoutbuffer_reg[7][13]  ( .D(n2597), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n937) );
  DFFNSRXLTS \requesterAddressbuffer_reg[2][2]  ( .D(n2850), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][2] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[2][3]  ( .D(n2849), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][3] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[2][5]  ( .D(n2847), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][5] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[2][0]  ( .D(n2852), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][0] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[2][1]  ( .D(n2851), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][1] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[2][4]  ( .D(n2848), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][4] ) );
  DFFNSRXLTS \dataoutbuffer_reg[2][16]  ( .D(n2754), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n99) );
  DFFNSRXLTS \dataoutbuffer_reg[2][22]  ( .D(n2748), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n98) );
  DFFNSRXLTS \dataoutbuffer_reg[2][24]  ( .D(n2746), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n97) );
  DFFNSRXLTS \dataoutbuffer_reg[2][31]  ( .D(n2739), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n96) );
  DFFNSRXLTS \dataoutbuffer_reg[2][1]  ( .D(n2769), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n95) );
  DFFNSRXLTS \dataoutbuffer_reg[2][10]  ( .D(n2760), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n94) );
  DFFNSRXLTS \dataoutbuffer_reg[2][27]  ( .D(n2743), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n93) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][0]  ( .D(n2492), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n92) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][1]  ( .D(n2491), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n91) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][3]  ( .D(n2489), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n90) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][4]  ( .D(n2488), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n89) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][5]  ( .D(n2487), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n88) );
  DFFNSRXLTS \dataoutbuffer_reg[2][3]  ( .D(n2767), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n87) );
  DFFNSRXLTS \dataoutbuffer_reg[2][4]  ( .D(n2766), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n86) );
  DFFNSRXLTS \dataoutbuffer_reg[2][5]  ( .D(n2765), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n85) );
  DFFNSRXLTS \dataoutbuffer_reg[2][7]  ( .D(n2763), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n84) );
  DFFNSRXLTS \dataoutbuffer_reg[2][8]  ( .D(n2762), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n83) );
  DFFNSRXLTS \dataoutbuffer_reg[2][9]  ( .D(n2761), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n82) );
  DFFNSRXLTS \dataoutbuffer_reg[2][11]  ( .D(n2759), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n81) );
  DFFNSRXLTS \dataoutbuffer_reg[2][12]  ( .D(n2758), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n80) );
  DFFNSRXLTS \dataoutbuffer_reg[2][13]  ( .D(n2757), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n79) );
  DFFNSRXLTS \dataoutbuffer_reg[2][14]  ( .D(n2756), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n78) );
  DFFNSRXLTS \dataoutbuffer_reg[2][15]  ( .D(n2755), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n77) );
  DFFNSRXLTS \dataoutbuffer_reg[2][17]  ( .D(n2753), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n76) );
  DFFNSRXLTS \dataoutbuffer_reg[2][18]  ( .D(n2752), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n75) );
  DFFNSRXLTS \dataoutbuffer_reg[2][19]  ( .D(n2751), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n74) );
  DFFNSRXLTS \dataoutbuffer_reg[2][20]  ( .D(n2750), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n73) );
  DFFNSRXLTS \dataoutbuffer_reg[2][21]  ( .D(n2749), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n72) );
  DFFNSRXLTS \dataoutbuffer_reg[2][23]  ( .D(n2747), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n71) );
  DFFNSRXLTS \dataoutbuffer_reg[2][25]  ( .D(n2745), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n70) );
  DFFNSRXLTS \dataoutbuffer_reg[2][26]  ( .D(n2744), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n69) );
  DFFNSRXLTS \dataoutbuffer_reg[2][28]  ( .D(n2742), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n68) );
  DFFNSRXLTS \dataoutbuffer_reg[2][29]  ( .D(n2741), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n67) );
  DFFNSRXLTS \dataoutbuffer_reg[2][30]  ( .D(n2740), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n66) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][2]  ( .D(n2490), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n65) );
  DFFNSRXLTS \dataoutbuffer_reg[1][0]  ( .D(n2802), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3043), .QN(n812) );
  DFFNSRXLTS \dataoutbuffer_reg[1][1]  ( .D(n2801), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3042), .QN(n813) );
  DFFNSRXLTS \dataoutbuffer_reg[1][3]  ( .D(n2799), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3040), .QN(n814) );
  DFFNSRXLTS \dataoutbuffer_reg[1][4]  ( .D(n2798), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3039), .QN(n815) );
  DFFNSRXLTS \dataoutbuffer_reg[1][6]  ( .D(n2796), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3037), .QN(n816) );
  DFFNSRXLTS \dataoutbuffer_reg[1][7]  ( .D(n2795), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3036), .QN(n817) );
  DFFNSRXLTS \dataoutbuffer_reg[1][9]  ( .D(n2793), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3034), .QN(n818) );
  DFFNSRXLTS \dataoutbuffer_reg[1][11]  ( .D(n2791), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3032), .QN(n819) );
  DFFNSRXLTS \dataoutbuffer_reg[1][12]  ( .D(n2790), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3031), .QN(n820) );
  DFFNSRXLTS \dataoutbuffer_reg[1][13]  ( .D(n2789), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3030), .QN(n821) );
  DFFNSRXLTS \dataoutbuffer_reg[1][14]  ( .D(n2788), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3029), .QN(n822) );
  DFFNSRXLTS \dataoutbuffer_reg[1][15]  ( .D(n2787), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3028), .QN(n823) );
  DFFNSRXLTS \dataoutbuffer_reg[1][16]  ( .D(n2786), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3027), .QN(n824) );
  DFFNSRXLTS \dataoutbuffer_reg[1][17]  ( .D(n2785), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3026), .QN(n825) );
  DFFNSRXLTS \dataoutbuffer_reg[1][18]  ( .D(n2784), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3025), .QN(n826) );
  DFFNSRXLTS \dataoutbuffer_reg[1][21]  ( .D(n2781), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3022), .QN(n827) );
  DFFNSRXLTS \dataoutbuffer_reg[1][23]  ( .D(n2779), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3020), .QN(n828) );
  DFFNSRXLTS \dataoutbuffer_reg[1][24]  ( .D(n2778), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3019), .QN(n829) );
  DFFNSRXLTS \dataoutbuffer_reg[1][25]  ( .D(n2777), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3018), .QN(n830) );
  DFFNSRXLTS \dataoutbuffer_reg[1][26]  ( .D(n2776), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3017), .QN(n831) );
  DFFNSRXLTS \dataoutbuffer_reg[1][28]  ( .D(n2774), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3015), .QN(n832) );
  DFFNSRXLTS \dataoutbuffer_reg[1][29]  ( .D(n2773), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3014), .QN(n833) );
  DFFNSRXLTS \dataoutbuffer_reg[1][30]  ( .D(n2772), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3013), .QN(n834) );
  DFFNSRXLTS \dataoutbuffer_reg[1][31]  ( .D(n2771), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3012), .QN(n835) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][0]  ( .D(n2478), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3049), .QN(n836) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][1]  ( .D(n2477), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3048), .QN(n837) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][2]  ( .D(n2476), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3047), .QN(n838) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][3]  ( .D(n2475), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3046), .QN(n839) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][5]  ( .D(n2473), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3044), .QN(n840) );
  DFFNSRXLTS \dataoutbuffer_reg[1][2]  ( .D(n2800), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3041), .QN(n841) );
  DFFNSRXLTS \dataoutbuffer_reg[1][5]  ( .D(n2797), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3038), .QN(n842) );
  DFFNSRXLTS \dataoutbuffer_reg[1][8]  ( .D(n2794), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3035), .QN(n843) );
  DFFNSRXLTS \dataoutbuffer_reg[1][10]  ( .D(n2792), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3033), .QN(n844) );
  DFFNSRXLTS \dataoutbuffer_reg[1][19]  ( .D(n2783), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3024), .QN(n845) );
  DFFNSRXLTS \dataoutbuffer_reg[1][20]  ( .D(n2782), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3023), .QN(n846) );
  DFFNSRXLTS \dataoutbuffer_reg[1][22]  ( .D(n2780), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3021), .QN(n847) );
  DFFNSRXLTS \dataoutbuffer_reg[1][27]  ( .D(n2775), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3016), .QN(n848) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][0]  ( .D(n2846), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2914), .QN(n900) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][1]  ( .D(n2845), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2912), .QN(n901) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][2]  ( .D(n2844), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2911), .QN(n902) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][3]  ( .D(n2843), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2913), .QN(n903) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][4]  ( .D(n2842), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2910), .QN(n904) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][5]  ( .D(n2841), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2909), .QN(n905) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][4]  ( .D(n2474), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3045), .QN(n849) );
  DFFNSRXLTS \writeOutbuffer_reg[7]  ( .D(n2578), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n653) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][4]  ( .D(n2544), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3000) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][0]  ( .D(n2548), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3008) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][1]  ( .D(n2547), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3006) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][2]  ( .D(n2546), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3004) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][3]  ( .D(n2545), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3002) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][5]  ( .D(n2543), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2998) );
  DFFNSRXLTS \requesterAddressbuffer_reg[6][0]  ( .D(n2876), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][0] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[6][1]  ( .D(n2875), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][1] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[6][2]  ( .D(n2874), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][2] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[6][3]  ( .D(n2873), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][3] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[6][4]  ( .D(n2872), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][4] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[6][5]  ( .D(n2871), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][5] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[0][0]  ( .D(n2840), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][0] ), .QN(n643) );
  DFFNSRXLTS \requesterAddressbuffer_reg[0][1]  ( .D(n2839), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][1] ), .QN(n644) );
  DFFNSRXLTS \requesterAddressbuffer_reg[0][2]  ( .D(n2838), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][2] ), .QN(n645) );
  DFFNSRXLTS \requesterAddressbuffer_reg[0][4]  ( .D(n2836), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][4] ), .QN(n646) );
  DFFNSRXLTS \requesterAddressbuffer_reg[0][3]  ( .D(n2837), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][3] ), .QN(n647) );
  DFFNSRXLTS \requesterAddressbuffer_reg[0][5]  ( .D(n2835), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][5] ), .QN(n648) );
  DFFNSRXLTS \dataoutbuffer_reg[0][0]  ( .D(n2834), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n64), .QN(n667) );
  DFFNSRXLTS \dataoutbuffer_reg[0][1]  ( .D(n2833), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n63), .QN(n668) );
  DFFNSRXLTS \dataoutbuffer_reg[0][2]  ( .D(n2832), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n62), .QN(n669) );
  DFFNSRXLTS \dataoutbuffer_reg[0][5]  ( .D(n2829), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n61), .QN(n670) );
  DFFNSRXLTS \dataoutbuffer_reg[0][9]  ( .D(n2825), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n60), .QN(n671) );
  DFFNSRXLTS \dataoutbuffer_reg[0][20]  ( .D(n2814), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n59), .QN(n672) );
  DFFNSRXLTS \dataoutbuffer_reg[0][23]  ( .D(n2811), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n58), .QN(n673) );
  DFFNSRXLTS \dataoutbuffer_reg[0][27]  ( .D(n2807), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n57), .QN(n674) );
  DFFNSRXLTS \dataoutbuffer_reg[0][28]  ( .D(n2806), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n56), .QN(n675) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][0]  ( .D(n2464), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n55), .QN(n676) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][4]  ( .D(n2460), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n54), .QN(n677) );
  DFFNSRXLTS \dataoutbuffer_reg[0][3]  ( .D(n2831), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n53), .QN(n678) );
  DFFNSRXLTS \dataoutbuffer_reg[0][4]  ( .D(n2830), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n52), .QN(n679) );
  DFFNSRXLTS \dataoutbuffer_reg[0][6]  ( .D(n2828), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n51), .QN(n680) );
  DFFNSRXLTS \dataoutbuffer_reg[0][7]  ( .D(n2827), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n50), .QN(n681) );
  DFFNSRXLTS \dataoutbuffer_reg[0][8]  ( .D(n2826), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n49), .QN(n682) );
  DFFNSRXLTS \dataoutbuffer_reg[0][10]  ( .D(n2824), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n48), .QN(n683) );
  DFFNSRXLTS \dataoutbuffer_reg[0][11]  ( .D(n2823), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n47), .QN(n684) );
  DFFNSRXLTS \dataoutbuffer_reg[0][12]  ( .D(n2822), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n46), .QN(n685) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][6]  ( .D(n2556), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3160), .QN(n578) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][7]  ( .D(n2555), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3158), .QN(n579) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][8]  ( .D(n2554), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3156), .QN(n580) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][11]  ( .D(n2551), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3151), .QN(n581) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][12]  ( .D(n2550), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3149), .QN(n582) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][13]  ( .D(n2549), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3147), .QN(n583) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][9]  ( .D(n2553), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3154), .QN(n584) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][5]  ( .D(n2459), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n704), .QN(n4716) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][3]  ( .D(n2461), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n703), .QN(n4736) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][2]  ( .D(n2462), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n702), .QN(n4747) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][1]  ( .D(n2463), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n701), .QN(n4752) );
  DFFNSRXLTS \dataoutbuffer_reg[0][31]  ( .D(n2803), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n700), .QN(n4424) );
  DFFNSRXLTS \dataoutbuffer_reg[0][30]  ( .D(n2804), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n699), .QN(n4437) );
  DFFNSRXLTS \dataoutbuffer_reg[0][29]  ( .D(n2805), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n698), .QN(n4448) );
  DFFNSRXLTS \dataoutbuffer_reg[0][26]  ( .D(n2808), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n697), .QN(n4473) );
  DFFNSRXLTS \dataoutbuffer_reg[0][25]  ( .D(n2809), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n696), .QN(n4480) );
  DFFNSRXLTS \dataoutbuffer_reg[0][24]  ( .D(n2810), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n695), .QN(n4489) );
  DFFNSRXLTS \dataoutbuffer_reg[0][22]  ( .D(n2812), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n694), .QN(n4505) );
  DFFNSRXLTS \dataoutbuffer_reg[0][21]  ( .D(n2813), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n693), .QN(n4520) );
  DFFNSRXLTS \dataoutbuffer_reg[0][19]  ( .D(n2815), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n692), .QN(n4534) );
  DFFNSRXLTS \dataoutbuffer_reg[0][18]  ( .D(n2816), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n691), .QN(n4543) );
  DFFNSRXLTS \dataoutbuffer_reg[0][17]  ( .D(n2817), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n690), .QN(n4552) );
  DFFNSRXLTS \dataoutbuffer_reg[0][16]  ( .D(n2818), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n689), .QN(n4561) );
  DFFNSRXLTS \dataoutbuffer_reg[0][15]  ( .D(n2819), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n688), .QN(n4572) );
  DFFNSRXLTS \dataoutbuffer_reg[0][14]  ( .D(n2820), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n687), .QN(n4579) );
  DFFNSRXLTS \dataoutbuffer_reg[0][13]  ( .D(n2821), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n686), .QN(n4592) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][10]  ( .D(n2552), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n4796) );
  DFFNSRXLTS \dataoutbuffer_reg[2][6]  ( .D(n2764), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n666) );
  DFFNSRXLTS \dataoutbuffer_reg[2][2]  ( .D(n2768), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n665) );
  DFFNSRXLTS \dataoutbuffer_reg[2][0]  ( .D(n2770), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n664) );
  DFFNSRXLTS \write_reg_reg[0]  ( .D(n2888), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n4), .QN(n5327) );
  DFFNSRXLTS \write_reg_reg[1]  ( .D(n2887), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n3), .QN(n5323) );
  DFFNSRXLTS full_reg_reg ( .D(N4718), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(
        n6347) );
  DFFNSRXLTS \destinationAddressOut_reg[7]  ( .D(n2447), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[7]) );
  DFFNSRXLTS \destinationAddressOut_reg[6]  ( .D(n2448), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[6]) );
  DFFNSRXLTS \destinationAddressOut_reg[9]  ( .D(n2445), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[9]) );
  DFFNSRXLTS \destinationAddressOut_reg[8]  ( .D(n2446), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[8]) );
  DFFNSRXLTS \destinationAddressOut_reg[13]  ( .D(n2441), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[13]) );
  DFFNSRXLTS \destinationAddressOut_reg[12]  ( .D(n2442), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[12]) );
  DFFNSRXLTS \destinationAddressOut_reg[11]  ( .D(n2443), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[11]) );
  DFFNSRXLTS \destinationAddressOut_reg[10]  ( .D(n2444), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[10]) );
  DFFNSRXLTS \readOutbuffer_reg[1]  ( .D(n2564), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n655) );
  DFFNSRXLTS \readOutbuffer_reg[0]  ( .D(n2563), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n656) );
  DFFNSRXLTS \readOutbuffer_reg[7]  ( .D(n2570), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer_7) );
  DFFNSRXLTS \readOutbuffer_reg[5]  ( .D(n2568), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n654) );
  DFFNSRXLTS \readOutbuffer_reg[6]  ( .D(n2569), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n650) );
  DFFNSRXLTS \readOutbuffer_reg[4]  ( .D(n2567), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n710) );
  DFFNSRXLTS \readOutbuffer_reg[2]  ( .D(n2565), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\readOutbuffer[2] ), .QN(n709) );
  DFFNSRXLTS \readOutbuffer_reg[3]  ( .D(n2566), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n649) );
  DFFNSRXLTS \writeOutbuffer_reg[0]  ( .D(n2571), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n705) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][8]  ( .D(n2456), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3179), .QN(n555) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][7]  ( .D(n2457), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3178), .QN(n553) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][6]  ( .D(n2458), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3177), .QN(n554) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][12]  ( .D(n2452), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3183), .QN(n909) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][11]  ( .D(n2453), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3182), .QN(n907) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][10]  ( .D(n2454), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3181), .QN(n908) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][9]  ( .D(n2455), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3180), .QN(n906) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][13]  ( .D(n2451), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3184), .QN(n917) );
  DFFNSRXLTS \dataoutbuffer_reg[6][27]  ( .D(n2615), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2942), .QN(n940) );
  DFFNSRXLTS \dataoutbuffer_reg[6][26]  ( .D(n2616), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2944), .QN(n941) );
  DFFNSRXLTS \dataoutbuffer_reg[6][25]  ( .D(n2617), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2946), .QN(n942) );
  DFFNSRXLTS \dataoutbuffer_reg[6][24]  ( .D(n2618), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2948), .QN(n943) );
  DFFNSRXLTS \dataoutbuffer_reg[6][23]  ( .D(n2619), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2950), .QN(n944) );
  DFFNSRXLTS \dataoutbuffer_reg[6][22]  ( .D(n2620), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2952), .QN(n945) );
  DFFNSRXLTS \dataoutbuffer_reg[6][21]  ( .D(n2621), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2954), .QN(n946) );
  DFFNSRXLTS \dataoutbuffer_reg[6][20]  ( .D(n2622), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2956), .QN(n947) );
  DFFNSRXLTS \dataoutbuffer_reg[6][31]  ( .D(n2611), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2934), .QN(n637) );
  DFFNSRXLTS \dataoutbuffer_reg[6][30]  ( .D(n2612), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2936), .QN(n636) );
  DFFNSRXLTS \dataoutbuffer_reg[6][29]  ( .D(n2613), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2938), .QN(n938) );
  DFFNSRXLTS \dataoutbuffer_reg[6][28]  ( .D(n2614), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2940), .QN(n939) );
  DFFNSRXLTS \writeOutbuffer_reg[2]  ( .D(n2573), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n910) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][8]  ( .D(n2484), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3186), .QN(n764) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][7]  ( .D(n2485), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3135), .QN(n765) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][6]  ( .D(n2486), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3185), .QN(n763) );
  DFFNSRXLTS \dataoutbuffer_reg[6][3]  ( .D(n2639), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n2990), .QN(n630) );
  DFFNSRXLTS \dataoutbuffer_reg[6][2]  ( .D(n2640), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n2992), .QN(n629) );
  DFFNSRXLTS \dataoutbuffer_reg[6][1]  ( .D(n2641), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n2994), .QN(n640) );
  DFFNSRXLTS \dataoutbuffer_reg[6][0]  ( .D(n2642), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n2996), .QN(n628) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][12]  ( .D(n2480), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3190), .QN(n918) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][11]  ( .D(n2481), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3189), .QN(n919) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][10]  ( .D(n2482), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3188), .QN(n920) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][9]  ( .D(n2483), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3187), .QN(n921) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][5]  ( .D(n2853), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][5] ), .QN(n892) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][4]  ( .D(n2854), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][4] ), .QN(n893) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][3]  ( .D(n2855), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][3] ), .QN(n891) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][2]  ( .D(n2856), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][2] ), .QN(n890) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][1]  ( .D(n2857), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][1] ), .QN(n889) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][0]  ( .D(n2858), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][0] ), .QN(n888) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][13]  ( .D(n2479), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3191), .QN(n916) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][4]  ( .D(n2530), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n774) );
  DFFNSRXLTS \dataoutbuffer_reg[6][19]  ( .D(n2623), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2958), .QN(n948) );
  DFFNSRXLTS \dataoutbuffer_reg[6][18]  ( .D(n2624), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2960), .QN(n949) );
  DFFNSRXLTS \dataoutbuffer_reg[6][17]  ( .D(n2625), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2962), .QN(n950) );
  DFFNSRXLTS \dataoutbuffer_reg[6][16]  ( .D(n2626), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2964), .QN(n951) );
  DFFNSRXLTS \dataoutbuffer_reg[6][15]  ( .D(n2627), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2966), .QN(n952) );
  DFFNSRXLTS \dataoutbuffer_reg[6][14]  ( .D(n2628), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2968), .QN(n953) );
  DFFNSRXLTS \dataoutbuffer_reg[6][13]  ( .D(n2629), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2970), .QN(n954) );
  DFFNSRXLTS \dataoutbuffer_reg[6][12]  ( .D(n2630), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2972), .QN(n955) );
  DFFNSRXLTS \dataoutbuffer_reg[6][11]  ( .D(n2631), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2974), .QN(n635) );
  DFFNSRXLTS \dataoutbuffer_reg[6][10]  ( .D(n2632), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2976), .QN(n642) );
  DFFNSRXLTS \dataoutbuffer_reg[6][9]  ( .D(n2633), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n2978), .QN(n634) );
  DFFNSRXLTS \dataoutbuffer_reg[6][8]  ( .D(n2634), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n2980), .QN(n633) );
  DFFNSRXLTS \dataoutbuffer_reg[6][7]  ( .D(n2635), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n2982), .QN(n632) );
  DFFNSRXLTS \dataoutbuffer_reg[6][6]  ( .D(n2636), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n2984), .QN(n641) );
  DFFNSRXLTS \dataoutbuffer_reg[6][5]  ( .D(n2637), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n2986), .QN(n631) );
  DFFNSRXLTS \dataoutbuffer_reg[6][4]  ( .D(n2638), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n2988), .QN(n595) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][12]  ( .D(n2494), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3163), .QN(n569) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][11]  ( .D(n2495), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3165), .QN(n571) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][10]  ( .D(n2496), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3167), .QN(n557) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][9]  ( .D(n2497), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3169), .QN(n568) );
  DFFNSRXLTS \requesterAddressbuffer_reg[4][3]  ( .D(n2861), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2931) );
  DFFNSRXLTS \requesterAddressbuffer_reg[4][2]  ( .D(n2862), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2929) );
  DFFNSRXLTS \requesterAddressbuffer_reg[4][1]  ( .D(n2863), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2930) );
  DFFNSRXLTS \requesterAddressbuffer_reg[4][0]  ( .D(n2864), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2932) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][13]  ( .D(n2493), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3161), .QN(n558) );
  DFFNSRXLTS \dataoutbuffer_reg[3][1]  ( .D(n2737), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n6280), .QN(n862) );
  DFFNSRXLTS \dataoutbuffer_reg[3][0]  ( .D(n2738), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n6281), .QN(n861) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][13]  ( .D(n2521), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3146), .QN(n566) );
  DFFNSRXLTS \writeOutbuffer_reg[3]  ( .D(n2574), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n706) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][8]  ( .D(n2498), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3171), .QN(n567) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][7]  ( .D(n2499), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3173), .QN(n556) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][6]  ( .D(n2500), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3175), .QN(n570) );
  DFFNSRXLTS \requesterAddressbuffer_reg[4][5]  ( .D(n2859), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2927) );
  DFFNSRXLTS \requesterAddressbuffer_reg[4][4]  ( .D(n2860), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2928) );
  DFFNSRXLTS \writeOutbuffer_reg[4]  ( .D(n2575), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n708) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][8]  ( .D(n2512), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3143), .QN(n591) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][7]  ( .D(n2513), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3144), .QN(n590) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][6]  ( .D(n2514), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3145), .QN(n589) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][11]  ( .D(n2537), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3166), .QN(n574) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][9]  ( .D(n2539), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3170), .QN(n586) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][7]  ( .D(n2541), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3174), .QN(n572) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][6]  ( .D(n2542), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3176), .QN(n585) );
  DFFNSRXLTS \writeOutbuffer_reg[6]  ( .D(n2577), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n707) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][12]  ( .D(n2536), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3164), .QN(n588) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][10]  ( .D(n2538), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3168), .QN(n587) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][8]  ( .D(n2540), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3172), .QN(n573) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][13]  ( .D(n2465), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3129), .QN(n773) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][12]  ( .D(n2466), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3130), .QN(n772) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][11]  ( .D(n2467), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3131), .QN(n771) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][10]  ( .D(n2468), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3132), .QN(n770) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][9]  ( .D(n2469), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3133), .QN(n769) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][12]  ( .D(n2522), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3148), .QN(n565) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][11]  ( .D(n2523), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3150), .QN(n564) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][10]  ( .D(n2524), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .QN(n563) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][9]  ( .D(n2525), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3153), .QN(n562) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][5]  ( .D(n2501), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n6255), .QN(n887) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][4]  ( .D(n2502), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n6256), .QN(n886) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][3]  ( .D(n2503), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n6257), .QN(n885) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][2]  ( .D(n2504), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n6293), .QN(n860) );
  DFFNSRXLTS \dataoutbuffer_reg[5][31]  ( .D(n2643), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n811) );
  DFFNSRXLTS \dataoutbuffer_reg[5][30]  ( .D(n2644), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n801) );
  DFFNSRXLTS \dataoutbuffer_reg[5][29]  ( .D(n2645), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n800) );
  DFFNSRXLTS \dataoutbuffer_reg[5][28]  ( .D(n2646), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n799) );
  DFFNSRXLTS \dataoutbuffer_reg[5][27]  ( .D(n2647), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n798) );
  DFFNSRXLTS \dataoutbuffer_reg[5][26]  ( .D(n2648), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n797) );
  DFFNSRXLTS \dataoutbuffer_reg[5][25]  ( .D(n2649), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n796) );
  DFFNSRXLTS \dataoutbuffer_reg[5][24]  ( .D(n2650), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n795) );
  DFFNSRXLTS \dataoutbuffer_reg[5][23]  ( .D(n2651), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n794) );
  DFFNSRXLTS \dataoutbuffer_reg[5][22]  ( .D(n2652), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n793) );
  DFFNSRXLTS \dataoutbuffer_reg[5][21]  ( .D(n2653), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n792) );
  DFFNSRXLTS \dataoutbuffer_reg[5][20]  ( .D(n2654), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n791) );
  DFFNSRXLTS \dataoutbuffer_reg[5][19]  ( .D(n2655), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n790) );
  DFFNSRXLTS \dataoutbuffer_reg[5][18]  ( .D(n2656), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n789) );
  DFFNSRXLTS \dataoutbuffer_reg[5][17]  ( .D(n2657), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n788) );
  DFFNSRXLTS \dataoutbuffer_reg[5][16]  ( .D(n2658), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n810) );
  DFFNSRXLTS \dataoutbuffer_reg[5][15]  ( .D(n2659), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n809) );
  DFFNSRXLTS \dataoutbuffer_reg[5][14]  ( .D(n2660), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n787) );
  DFFNSRXLTS \dataoutbuffer_reg[5][13]  ( .D(n2661), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n786) );
  DFFNSRXLTS \dataoutbuffer_reg[5][12]  ( .D(n2662), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n785) );
  DFFNSRXLTS \dataoutbuffer_reg[5][11]  ( .D(n2663), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n808) );
  DFFNSRXLTS \dataoutbuffer_reg[5][10]  ( .D(n2664), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n784) );
  DFFNSRXLTS \dataoutbuffer_reg[5][9]  ( .D(n2665), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n783) );
  DFFNSRXLTS \dataoutbuffer_reg[5][8]  ( .D(n2666), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n782) );
  DFFNSRXLTS \dataoutbuffer_reg[5][7]  ( .D(n2667), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n781) );
  DFFNSRXLTS \dataoutbuffer_reg[5][6]  ( .D(n2668), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n780) );
  DFFNSRXLTS \dataoutbuffer_reg[5][5]  ( .D(n2669), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n779) );
  DFFNSRXLTS \dataoutbuffer_reg[5][4]  ( .D(n2670), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n778) );
  DFFNSRXLTS \dataoutbuffer_reg[5][3]  ( .D(n2671), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n777) );
  DFFNSRXLTS \dataoutbuffer_reg[5][2]  ( .D(n2672), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n776) );
  DFFNSRXLTS \dataoutbuffer_reg[5][1]  ( .D(n2673), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n807) );
  DFFNSRXLTS \dataoutbuffer_reg[5][0]  ( .D(n2674), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n775) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][5]  ( .D(n2529), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n806) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][3]  ( .D(n2531), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n805) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][2]  ( .D(n2532), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n804) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][1]  ( .D(n2533), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n803) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][0]  ( .D(n2534), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n802) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][13]  ( .D(n2535), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3162), .QN(n575) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][12]  ( .D(n2508), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3139), .QN(n594) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][11]  ( .D(n2509), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3140), .QN(n593) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][10]  ( .D(n2510), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3141), .QN(n592) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][9]  ( .D(n2511), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3142), .QN(n576) );
  DFFNSRXLTS \requesterAddressbuffer_reg[5][5]  ( .D(n2865), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n899) );
  DFFNSRXLTS \requesterAddressbuffer_reg[5][4]  ( .D(n2866), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n898) );
  DFFNSRXLTS \requesterAddressbuffer_reg[5][0]  ( .D(n2870), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n894) );
  DFFNSRXLTS \requesterAddressbuffer_reg[5][3]  ( .D(n2867), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n897) );
  DFFNSRXLTS \requesterAddressbuffer_reg[5][2]  ( .D(n2868), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n896) );
  DFFNSRXLTS \requesterAddressbuffer_reg[5][1]  ( .D(n2869), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n895) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][13]  ( .D(n2507), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3138), .QN(n577) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][1]  ( .D(n2519), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3005) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][0]  ( .D(n2520), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3007) );
  DFFNSRXLTS \dataoutbuffer_reg[4][31]  ( .D(n2675), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2933) );
  DFFNSRXLTS \dataoutbuffer_reg[4][30]  ( .D(n2676), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2935) );
  DFFNSRXLTS \dataoutbuffer_reg[4][29]  ( .D(n2677), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2937) );
  DFFNSRXLTS \dataoutbuffer_reg[4][28]  ( .D(n2678), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2939) );
  DFFNSRXLTS \dataoutbuffer_reg[4][27]  ( .D(n2679), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2941) );
  DFFNSRXLTS \dataoutbuffer_reg[4][26]  ( .D(n2680), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2943) );
  DFFNSRXLTS \dataoutbuffer_reg[4][25]  ( .D(n2681), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2945) );
  DFFNSRXLTS \dataoutbuffer_reg[4][24]  ( .D(n2682), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2947) );
  DFFNSRXLTS \dataoutbuffer_reg[4][23]  ( .D(n2683), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2949) );
  DFFNSRXLTS \dataoutbuffer_reg[4][22]  ( .D(n2684), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2951) );
  DFFNSRXLTS \dataoutbuffer_reg[4][21]  ( .D(n2685), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2953) );
  DFFNSRXLTS \dataoutbuffer_reg[4][20]  ( .D(n2686), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2955) );
  DFFNSRXLTS \dataoutbuffer_reg[4][19]  ( .D(n2687), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2957) );
  DFFNSRXLTS \dataoutbuffer_reg[4][18]  ( .D(n2688), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2959) );
  DFFNSRXLTS \dataoutbuffer_reg[4][17]  ( .D(n2689), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2961) );
  DFFNSRXLTS \dataoutbuffer_reg[4][16]  ( .D(n2690), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2963) );
  DFFNSRXLTS \dataoutbuffer_reg[4][15]  ( .D(n2691), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2965) );
  DFFNSRXLTS \dataoutbuffer_reg[4][14]  ( .D(n2692), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2967) );
  DFFNSRXLTS \dataoutbuffer_reg[4][13]  ( .D(n2693), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2969) );
  DFFNSRXLTS \dataoutbuffer_reg[4][12]  ( .D(n2694), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2971) );
  DFFNSRXLTS \dataoutbuffer_reg[4][11]  ( .D(n2695), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2973) );
  DFFNSRXLTS \dataoutbuffer_reg[4][10]  ( .D(n2696), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2975) );
  DFFNSRXLTS \dataoutbuffer_reg[4][9]  ( .D(n2697), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n2977) );
  DFFNSRXLTS \dataoutbuffer_reg[4][8]  ( .D(n2698), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n2979) );
  DFFNSRXLTS \dataoutbuffer_reg[4][7]  ( .D(n2699), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n2981) );
  DFFNSRXLTS \dataoutbuffer_reg[4][6]  ( .D(n2700), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n2983) );
  DFFNSRXLTS \dataoutbuffer_reg[4][5]  ( .D(n2701), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n2985) );
  DFFNSRXLTS \dataoutbuffer_reg[4][4]  ( .D(n2702), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n2987) );
  DFFNSRXLTS \dataoutbuffer_reg[4][3]  ( .D(n2703), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n2989) );
  DFFNSRXLTS \dataoutbuffer_reg[4][2]  ( .D(n2704), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n2991) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][1]  ( .D(n2505), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n6258), .QN(n884) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][0]  ( .D(n2506), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n6259), .QN(n883) );
  DFFNSRXLTS \dataoutbuffer_reg[3][31]  ( .D(n2707), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6260), .QN(n882) );
  DFFNSRXLTS \dataoutbuffer_reg[3][30]  ( .D(n2708), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6261), .QN(n881) );
  DFFNSRXLTS \dataoutbuffer_reg[3][29]  ( .D(n2709), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6262), .QN(n880) );
  DFFNSRXLTS \dataoutbuffer_reg[3][28]  ( .D(n2710), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6263), .QN(n879) );
  DFFNSRXLTS \dataoutbuffer_reg[3][27]  ( .D(n2711), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6264), .QN(n878) );
  DFFNSRXLTS \dataoutbuffer_reg[3][26]  ( .D(n2712), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6265), .QN(n877) );
  DFFNSRXLTS \dataoutbuffer_reg[3][25]  ( .D(n2713), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6294), .QN(n859) );
  DFFNSRXLTS \dataoutbuffer_reg[3][24]  ( .D(n2714), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6266), .QN(n876) );
  DFFNSRXLTS \dataoutbuffer_reg[3][23]  ( .D(n2715), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6295), .QN(n858) );
  DFFNSRXLTS \dataoutbuffer_reg[3][22]  ( .D(n2716), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6267), .QN(n875) );
  DFFNSRXLTS \dataoutbuffer_reg[3][21]  ( .D(n2717), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6268), .QN(n874) );
  DFFNSRXLTS \dataoutbuffer_reg[3][20]  ( .D(n2718), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6296), .QN(n857) );
  DFFNSRXLTS \dataoutbuffer_reg[3][19]  ( .D(n2719), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6269), .QN(n873) );
  DFFNSRXLTS \dataoutbuffer_reg[3][18]  ( .D(n2720), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6297), .QN(n856) );
  DFFNSRXLTS \dataoutbuffer_reg[3][17]  ( .D(n2721), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6270), .QN(n872) );
  DFFNSRXLTS \dataoutbuffer_reg[3][16]  ( .D(n2722), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6271), .QN(n871) );
  DFFNSRXLTS \dataoutbuffer_reg[3][15]  ( .D(n2723), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6298), .QN(n855) );
  DFFNSRXLTS \dataoutbuffer_reg[3][14]  ( .D(n2724), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6272), .QN(n870) );
  DFFNSRXLTS \dataoutbuffer_reg[3][13]  ( .D(n2725), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6299), .QN(n854) );
  DFFNSRXLTS \dataoutbuffer_reg[3][12]  ( .D(n2726), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6273), .QN(n869) );
  DFFNSRXLTS \dataoutbuffer_reg[3][11]  ( .D(n2727), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6274), .QN(n868) );
  DFFNSRXLTS \dataoutbuffer_reg[3][10]  ( .D(n2728), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6275), .QN(n867) );
  DFFNSRXLTS \dataoutbuffer_reg[3][9]  ( .D(n2729), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n6276), .QN(n866) );
  DFFNSRXLTS \dataoutbuffer_reg[3][8]  ( .D(n2730), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n6277), .QN(n865) );
  DFFNSRXLTS \dataoutbuffer_reg[3][7]  ( .D(n2731), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n6312), .QN(n850) );
  DFFNSRXLTS \dataoutbuffer_reg[3][6]  ( .D(n2732), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n6278), .QN(n864) );
  DFFNSRXLTS \dataoutbuffer_reg[3][5]  ( .D(n2733), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n6300), .QN(n853) );
  DFFNSRXLTS \dataoutbuffer_reg[3][4]  ( .D(n2734), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n6301), .QN(n852) );
  DFFNSRXLTS \dataoutbuffer_reg[3][3]  ( .D(n2735), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n6279), .QN(n863) );
  DFFNSRXLTS \dataoutbuffer_reg[3][2]  ( .D(n2736), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n6302), .QN(n851) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][5]  ( .D(n2515), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2997) );
  DFFNSRXLTS \dataoutbuffer_reg[4][1]  ( .D(n2705), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n2993) );
  DFFNSRXLTS \dataoutbuffer_reg[4][0]  ( .D(n2706), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n2995) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][4]  ( .D(n2516), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2999) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][3]  ( .D(n2517), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3001) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][2]  ( .D(n2518), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3003) );
  NOR3BX1TS U2 ( .AN(n444), .B(n1789), .C(n452), .Y(n1156) );
  BUFX3TS U3 ( .A(n756), .Y(n44) );
  CLKAND2X3TS U4 ( .A(n1962), .B(selectBit_WEST), .Y(n1893) );
  BUFX3TS U5 ( .A(n3505), .Y(n3496) );
  BUFX2TS U6 ( .A(n3505), .Y(n3497) );
  BUFX3TS U7 ( .A(n3933), .Y(n3923) );
  CLKBUFX4TS U8 ( .A(n1783), .Y(n444) );
  CLKINVX4TS U9 ( .A(n1845), .Y(n756) );
  XOR2X2TS U10 ( .A(n2015), .B(n112), .Y(n1845) );
  NAND2X1TS U11 ( .A(n1768), .B(n2008), .Y(n1915) );
  CLKBUFX2TS U12 ( .A(n3862), .Y(n3861) );
  OA21XLTS U13 ( .A0(n1938), .A1(n1915), .B0(n1796), .Y(n1937) );
  AOI21X1TS U14 ( .A0(n931), .A1(n761), .B0(n1754), .Y(n1791) );
  NAND2X1TS U15 ( .A(selectBit_EAST), .B(n1915), .Y(n1961) );
  AND2X2TS U16 ( .A(n1791), .B(n751), .Y(n1753) );
  CLKBUFX2TS U17 ( .A(n3437), .Y(n3436) );
  CLKBUFX2TS U18 ( .A(n3420), .Y(n3419) );
  AOI21X1TS U19 ( .A0(n1794), .A1(n735), .B0(n755), .Y(n1796) );
  OAI21X1TS U20 ( .A0(n1832), .A1(n1870), .B0(n3098), .Y(n1775) );
  AOI222XLTS U21 ( .A0(n538), .A1(n3777), .B0(n4078), .B1(n3861), .C0(n6280), 
        .C1(n3842), .Y(n1427) );
  OA22X1TS U22 ( .A0(n1811), .A1(n171), .B0(n1842), .B1(n1976), .Y(n744) );
  INVX2TS U23 ( .A(n466), .Y(n722) );
  AND2X2TS U24 ( .A(n1786), .B(n1783), .Y(n1750) );
  OA22X2TS U25 ( .A0(n1786), .A1(n172), .B0(n1871), .B1(n106), .Y(n10) );
  OAI32XLTS U26 ( .A0(n4198), .A1(n754), .A2(n1803), .B0(n1804), .B1(n969), 
        .Y(n1802) );
  BUFX4TS U27 ( .A(n3471), .Y(n3469) );
  AND3XLTS U28 ( .A(n1796), .B(n109), .C(n1791), .Y(n1171) );
  AND3XLTS U29 ( .A(n1794), .B(n1795), .C(n1791), .Y(n1170) );
  INVX3TS U30 ( .A(n2014), .Y(n958) );
  AOI2BB1X2TS U31 ( .A0N(n454), .A1N(n973), .B0(n2907), .Y(n2017) );
  NAND3XLTS U32 ( .A(n1845), .B(n1847), .C(n930), .Y(n1869) );
  OR2X4TS U33 ( .A(selectBit_NORTH), .B(selectBit_SOUTH), .Y(n2384) );
  INVX2TS U34 ( .A(n449), .Y(n732) );
  INVX2TS U35 ( .A(n1753), .Y(n449) );
  CLKBUFX2TS U36 ( .A(n1156), .Y(n3477) );
  INVX2TS U37 ( .A(n718), .Y(n741) );
  CLKBUFX2TS U38 ( .A(n1221), .Y(n3193) );
  CLKBUFX2TS U39 ( .A(n1121), .Y(n3657) );
  INVX2TS U40 ( .A(n1775), .Y(n742) );
  CLKBUFX2TS U41 ( .A(n1187), .Y(n3360) );
  CLKBUFX2TS U42 ( .A(n1100), .Y(n3755) );
  CLKBUFX2TS U43 ( .A(n3426), .Y(n3420) );
  CLKBUFX2TS U44 ( .A(n3908), .Y(n3907) );
  OA21XLTS U45 ( .A0(n1937), .A1(n170), .B0(n1928), .Y(n1754) );
  CLKBUFX2TS U46 ( .A(n1218), .Y(n3241) );
  AOI21X1TS U47 ( .A0(n929), .A1(n761), .B0(n161), .Y(n1799) );
  OAI32X1TS U48 ( .A0(n2016), .A1(n5327), .A2(n958), .B0(n151), .B1(n2017), 
        .Y(n2015) );
  NOR2X1TS U49 ( .A(n1028), .B(n1962), .Y(n1847) );
  OA22X1TS U50 ( .A0(n1816), .A1(n172), .B0(n1871), .B1(n119), .Y(n749) );
  CLKBUFX2TS U51 ( .A(n3193), .Y(n3124) );
  CLKBUFX2TS U52 ( .A(n3797), .Y(n3793) );
  CLKBUFX2TS U53 ( .A(n3624), .Y(n3614) );
  CLKBUFX2TS U54 ( .A(n3504), .Y(n3503) );
  OAI22X1TS U55 ( .A0(n739), .A1(n170), .B0(n1871), .B1(n1938), .Y(n1757) );
  CLKBUFX2TS U56 ( .A(n3623), .Y(n3619) );
  CLKBUFX2TS U57 ( .A(n3235), .Y(n3234) );
  INVX2TS U58 ( .A(n1795), .Y(n755) );
  CLKBUFX2TS U59 ( .A(n3194), .Y(n3123) );
  CLKBUFX2TS U60 ( .A(n3626), .Y(n3623) );
  CLKBUFX2TS U61 ( .A(n741), .Y(n3798) );
  CLKBUFX2TS U62 ( .A(n1171), .Y(n3426) );
  AND2X2TS U63 ( .A(n6347), .B(n2050), .Y(n7) );
  XNOR2X1TS U64 ( .A(n107), .B(n151), .Y(n9) );
  NAND2X1TS U65 ( .A(n739), .B(n1799), .Y(n1756) );
  AND2X2TS U66 ( .A(n2011), .B(n119), .Y(n11) );
  CLKINVX2TS U67 ( .A(n1757), .Y(n161) );
  AND2X2TS U68 ( .A(n6253), .B(n4541), .Y(n12) );
  AND2X2TS U69 ( .A(n469), .B(n4541), .Y(n13) );
  INVXLTS U70 ( .A(n40), .Y(n14) );
  INVXLTS U71 ( .A(readRequesterAddress[0]), .Y(n15) );
  INVXLTS U72 ( .A(n15), .Y(n16) );
  INVXLTS U73 ( .A(n15), .Y(n17) );
  INVXLTS U74 ( .A(n15), .Y(n18) );
  INVXLTS U75 ( .A(n15), .Y(n19) );
  INVXLTS U76 ( .A(readRequesterAddress[1]), .Y(n20) );
  INVXLTS U77 ( .A(n20), .Y(n21) );
  INVXLTS U78 ( .A(n20), .Y(n22) );
  INVXLTS U79 ( .A(n20), .Y(n23) );
  INVXLTS U80 ( .A(n20), .Y(n24) );
  INVXLTS U81 ( .A(readRequesterAddress[2]), .Y(n25) );
  INVXLTS U82 ( .A(n25), .Y(n26) );
  INVXLTS U83 ( .A(n25), .Y(n27) );
  INVXLTS U84 ( .A(n25), .Y(n28) );
  INVXLTS U85 ( .A(n25), .Y(n29) );
  INVXLTS U86 ( .A(readRequesterAddress[3]), .Y(n30) );
  INVXLTS U87 ( .A(n30), .Y(n31) );
  INVXLTS U88 ( .A(n30), .Y(n32) );
  INVXLTS U89 ( .A(n30), .Y(n33) );
  INVXLTS U90 ( .A(n30), .Y(n34) );
  INVXLTS U91 ( .A(readRequesterAddress[4]), .Y(n35) );
  INVXLTS U92 ( .A(n35), .Y(n36) );
  INVXLTS U93 ( .A(n35), .Y(n37) );
  INVXLTS U94 ( .A(n35), .Y(n38) );
  INVXLTS U95 ( .A(n35), .Y(n39) );
  INVXLTS U96 ( .A(readRequesterAddress[5]), .Y(n40) );
  INVXLTS U97 ( .A(n40), .Y(n41) );
  INVXLTS U98 ( .A(n40), .Y(n42) );
  INVXLTS U99 ( .A(n40), .Y(n43) );
  INVXLTS U100 ( .A(n442), .Y(n45) );
  INVXLTS U101 ( .A(n120), .Y(n100) );
  CLKBUFX2TS U102 ( .A(n1776), .Y(n101) );
  INVXLTS U103 ( .A(n1799), .Y(n102) );
  INVXLTS U104 ( .A(n102), .Y(n103) );
  CLKBUFX2TS U105 ( .A(n1807), .Y(n104) );
  INVXLTS U106 ( .A(n1884), .Y(n105) );
  INVXLTS U107 ( .A(n105), .Y(n106) );
  CLKBUFX2TS U108 ( .A(n1985), .Y(n107) );
  INVXLTS U109 ( .A(n11), .Y(n108) );
  INVX1TS U110 ( .A(n11), .Y(n109) );
  NAND3X1TS U111 ( .A(n756), .B(n1846), .C(n1847), .Y(n1795) );
  INVXLTS U112 ( .A(n2009), .Y(n110) );
  INVXLTS U113 ( .A(n2009), .Y(n111) );
  INVXLTS U114 ( .A(n471), .Y(n112) );
  INVXLTS U115 ( .A(n112), .Y(n113) );
  INVXLTS U116 ( .A(n913), .Y(n114) );
  INVXLTS U117 ( .A(n114), .Y(n115) );
  INVXLTS U118 ( .A(n9), .Y(n116) );
  INVXLTS U119 ( .A(n9), .Y(n117) );
  INVXLTS U120 ( .A(n1976), .Y(n118) );
  INVXLTS U121 ( .A(n118), .Y(n119) );
  INVXLTS U122 ( .A(n5), .Y(n120) );
  INVXLTS U123 ( .A(n968), .Y(n121) );
  INVXLTS U124 ( .A(n121), .Y(n122) );
  INVXLTS U125 ( .A(n967), .Y(n123) );
  INVXLTS U126 ( .A(n123), .Y(n124) );
  INVXLTS U127 ( .A(destinationAddressIn_NORTH[12]), .Y(n125) );
  INVXLTS U128 ( .A(destinationAddressIn_NORTH[12]), .Y(n126) );
  INVXLTS U129 ( .A(destinationAddressIn_NORTH[11]), .Y(n127) );
  INVXLTS U130 ( .A(destinationAddressIn_NORTH[11]), .Y(n128) );
  INVXLTS U131 ( .A(destinationAddressIn_NORTH[9]), .Y(n129) );
  INVXLTS U132 ( .A(destinationAddressIn_NORTH[9]), .Y(n130) );
  INVXLTS U133 ( .A(destinationAddressIn_NORTH[8]), .Y(n131) );
  INVXLTS U134 ( .A(destinationAddressIn_NORTH[13]), .Y(n132) );
  INVXLTS U135 ( .A(destinationAddressIn_NORTH[13]), .Y(n133) );
  INVXLTS U136 ( .A(destinationAddressIn_NORTH[10]), .Y(n134) );
  INVXLTS U137 ( .A(destinationAddressIn_NORTH[10]), .Y(n135) );
  INVXLTS U138 ( .A(n45), .Y(n136) );
  INVXLTS U139 ( .A(n8), .Y(n137) );
  INVXLTS U140 ( .A(n13), .Y(n138) );
  INVXLTS U141 ( .A(n13), .Y(n139) );
  INVXLTS U142 ( .A(n720), .Y(n140) );
  INVXLTS U143 ( .A(n140), .Y(n141) );
  INVXLTS U144 ( .A(n140), .Y(n142) );
  INVXLTS U145 ( .A(n151), .Y(n143) );
  INVXLTS U146 ( .A(n719), .Y(n144) );
  INVXLTS U147 ( .A(n144), .Y(n145) );
  INVXLTS U148 ( .A(n144), .Y(n146) );
  INVXLTS U149 ( .A(n970), .Y(n147) );
  INVXLTS U150 ( .A(n147), .Y(n148) );
  INVXLTS U151 ( .A(n147), .Y(n149) );
  INVXLTS U152 ( .A(n926), .Y(n150) );
  INVXLTS U153 ( .A(n150), .Y(n151) );
  INVXLTS U154 ( .A(n12), .Y(n152) );
  INVXLTS U155 ( .A(n12), .Y(n153) );
  INVXLTS U156 ( .A(n12), .Y(n154) );
  INVXLTS U157 ( .A(n711), .Y(n155) );
  INVXLTS U158 ( .A(n155), .Y(n156) );
  INVXLTS U159 ( .A(n155), .Y(n157) );
  INVX2TS U160 ( .A(n10), .Y(n158) );
  INVXLTS U161 ( .A(n10), .Y(n159) );
  INVXLTS U162 ( .A(n10), .Y(n160) );
  INVX2TS U163 ( .A(n161), .Y(n162) );
  INVXLTS U164 ( .A(n161), .Y(n163) );
  INVXLTS U165 ( .A(n3838), .Y(n164) );
  INVXLTS U166 ( .A(n3838), .Y(n165) );
  INVXLTS U167 ( .A(n4), .Y(n166) );
  INVXLTS U168 ( .A(n2037), .Y(n167) );
  INVXLTS U169 ( .A(n167), .Y(n168) );
  INVXLTS U170 ( .A(n167), .Y(n169) );
  INVXLTS U171 ( .A(n7), .Y(n170) );
  INVXLTS U172 ( .A(n7), .Y(n171) );
  INVXLTS U173 ( .A(n7), .Y(n172) );
  NOR2X1TS U435 ( .A(n971), .B(n2010), .Y(n2006) );
  CLKBUFX2TS U436 ( .A(n969), .Y(n434) );
  CLKINVX2TS U437 ( .A(n2006), .Y(n435) );
  CLKBUFX2TS U438 ( .A(selectBit_SOUTH), .Y(n436) );
  NAND2XLTS U439 ( .A(n2010), .B(n436), .Y(n2009) );
  CLKBUFX2TS U440 ( .A(n959), .Y(n437) );
  CLKINVX2TS U441 ( .A(selectBit_NORTH), .Y(n959) );
  INVX2TS U442 ( .A(readIn_SOUTH), .Y(n438) );
  CLKBUFX2TS U443 ( .A(n1791), .Y(n439) );
  CLKBUFX2TS U444 ( .A(n1769), .Y(n440) );
  NOR2XLTS U445 ( .A(n1768), .B(n1769), .Y(n1103) );
  CLKBUFX2TS U446 ( .A(n2383), .Y(n441) );
  INVX2TS U447 ( .A(n746), .Y(n443) );
  INVX2TS U448 ( .A(n1789), .Y(n746) );
  OAI21X1TS U449 ( .A0(n1789), .A1(n1961), .B0(n2007), .Y(n1818) );
  AOI21X1TS U450 ( .A0(n929), .A1(n105), .B0(n3894), .Y(n1783) );
  INVX2TS U451 ( .A(n930), .Y(n445) );
  NAND3XLTS U452 ( .A(n756), .B(n445), .C(n1893), .Y(n1810) );
  NAND3XLTS U453 ( .A(n1845), .B(n1846), .C(n1893), .Y(n1780) );
  NOR3BX1TS U454 ( .AN(n1893), .B(n44), .C(n1846), .Y(n1788) );
  XNOR2X1TS U455 ( .A(n2014), .B(n166), .Y(n1846) );
  INVX2TS U456 ( .A(n1083), .Y(n446) );
  CLKBUFX2TS U457 ( .A(n1779), .Y(n447) );
  AND3X2TS U458 ( .A(n1779), .B(n1780), .C(n1776), .Y(n1139) );
  AOI21XLTS U459 ( .A0(n1779), .A1(n735), .B0(n753), .Y(n1811) );
  OAI221XLTS U460 ( .A0(n112), .A1(n748), .B0(n1803), .B1(n1961), .C0(n1805), 
        .Y(n1804) );
  INVX2TS U461 ( .A(n747), .Y(n448) );
  NOR2BX1TS U462 ( .AN(n1776), .B(n1812), .Y(n1137) );
  NOR2BX1TS U463 ( .AN(n1807), .B(n1812), .Y(n1201) );
  INVXLTS U464 ( .A(n1753), .Y(n450) );
  INVXLTS U465 ( .A(n1753), .Y(n451) );
  CLKBUFX2TS U466 ( .A(n1788), .Y(n452) );
  CLKBUFX2TS U467 ( .A(n1813), .Y(n453) );
  NOR3BX1TS U468 ( .AN(n1813), .B(n1818), .C(n927), .Y(n1221) );
  NOR3BX1TS U469 ( .AN(n1813), .B(n1789), .C(n752), .Y(n1218) );
  AOI21X1TS U470 ( .A0(n929), .A1(n118), .B0(n749), .Y(n1813) );
  CLKINVX2TS U471 ( .A(n2384), .Y(n454) );
  INVXLTS U472 ( .A(n2384), .Y(n455) );
  NAND3XLTS U473 ( .A(n2383), .B(n973), .C(n455), .Y(n2050) );
  CLKBUFX2TS U474 ( .A(n1832), .Y(n456) );
  OAI21X1TS U475 ( .A0(n1841), .A1(n456), .B0(n3754), .Y(n1769) );
  CLKBUFX2TS U476 ( .A(n2035), .Y(n712) );
  INVX2TS U477 ( .A(n712), .Y(n457) );
  INVX2TS U478 ( .A(n712), .Y(n458) );
  AND3X2TS U479 ( .A(n101), .B(n448), .C(n1781), .Y(n1748) );
  INVX2TS U480 ( .A(n1748), .Y(n459) );
  INVX2TS U481 ( .A(n1748), .Y(n460) );
  INVX2TS U482 ( .A(n1748), .Y(n461) );
  CLKBUFX2TS U483 ( .A(n2048), .Y(n462) );
  CLKAND2X2TS U484 ( .A(n1773), .B(n742), .Y(n1746) );
  INVX2TS U485 ( .A(n1746), .Y(n463) );
  INVX2TS U486 ( .A(n1746), .Y(n464) );
  INVX2TS U487 ( .A(n1746), .Y(n465) );
  CLKINVX2TS U488 ( .A(n1750), .Y(n466) );
  INVXLTS U489 ( .A(n1750), .Y(n467) );
  INVXLTS U490 ( .A(n1750), .Y(n468) );
  INVX2TS U491 ( .A(n1028), .Y(n470) );
  INVX2TS U492 ( .A(n726), .Y(n472) );
  INVXLTS U493 ( .A(selectBit_EAST), .Y(n726) );
  INVX2TS U494 ( .A(selectBit_EAST), .Y(n973) );
  CLKBUFX2TS U495 ( .A(n2034), .Y(n714) );
  INVX2TS U496 ( .A(n714), .Y(n473) );
  INVX2TS U497 ( .A(n714), .Y(n474) );
  CLKBUFX2TS U498 ( .A(n2036), .Y(n713) );
  INVX2TS U499 ( .A(n713), .Y(n475) );
  INVX2TS U500 ( .A(n713), .Y(n476) );
  CLKBUFX2TS U501 ( .A(cacheDataOut[28]), .Y(n477) );
  CLKBUFX2TS U502 ( .A(cacheDataOut[28]), .Y(n478) );
  CLKBUFX2TS U503 ( .A(cacheDataOut[27]), .Y(n479) );
  CLKBUFX2TS U504 ( .A(cacheDataOut[27]), .Y(n480) );
  CLKBUFX2TS U505 ( .A(cacheDataOut[23]), .Y(n481) );
  CLKBUFX2TS U506 ( .A(cacheDataOut[23]), .Y(n482) );
  CLKBUFX2TS U507 ( .A(cacheDataOut[20]), .Y(n483) );
  CLKBUFX2TS U508 ( .A(cacheDataOut[20]), .Y(n484) );
  CLKBUFX2TS U509 ( .A(cacheDataOut[12]), .Y(n485) );
  CLKBUFX2TS U510 ( .A(cacheDataOut[12]), .Y(n486) );
  CLKBUFX2TS U511 ( .A(cacheDataOut[11]), .Y(n487) );
  CLKBUFX2TS U512 ( .A(cacheDataOut[11]), .Y(n488) );
  CLKBUFX2TS U513 ( .A(cacheDataOut[10]), .Y(n489) );
  CLKBUFX2TS U514 ( .A(cacheDataOut[10]), .Y(n490) );
  CLKBUFX2TS U515 ( .A(cacheDataOut[9]), .Y(n491) );
  CLKBUFX2TS U516 ( .A(cacheDataOut[9]), .Y(n492) );
  CLKBUFX2TS U517 ( .A(cacheDataOut[8]), .Y(n493) );
  CLKBUFX2TS U518 ( .A(cacheDataOut[8]), .Y(n494) );
  CLKBUFX2TS U519 ( .A(cacheDataOut[7]), .Y(n495) );
  CLKBUFX2TS U520 ( .A(cacheDataOut[7]), .Y(n496) );
  CLKBUFX2TS U521 ( .A(cacheDataOut[6]), .Y(n497) );
  CLKBUFX2TS U522 ( .A(cacheDataOut[6]), .Y(n498) );
  CLKBUFX2TS U523 ( .A(cacheDataOut[5]), .Y(n499) );
  CLKBUFX2TS U524 ( .A(cacheDataOut[5]), .Y(n500) );
  CLKBUFX2TS U525 ( .A(cacheDataOut[4]), .Y(n501) );
  CLKBUFX2TS U526 ( .A(cacheDataOut[4]), .Y(n502) );
  CLKBUFX2TS U527 ( .A(cacheDataOut[3]), .Y(n503) );
  CLKBUFX2TS U528 ( .A(cacheDataOut[3]), .Y(n504) );
  CLKBUFX2TS U529 ( .A(cacheDataOut[2]), .Y(n505) );
  CLKBUFX2TS U530 ( .A(cacheDataOut[2]), .Y(n506) );
  CLKBUFX2TS U531 ( .A(cacheDataOut[30]), .Y(n507) );
  CLKBUFX2TS U532 ( .A(cacheDataOut[30]), .Y(n508) );
  CLKBUFX2TS U533 ( .A(cacheDataOut[16]), .Y(n509) );
  CLKBUFX2TS U534 ( .A(cacheDataOut[16]), .Y(n510) );
  CLKBUFX2TS U535 ( .A(cacheDataOut[31]), .Y(n511) );
  CLKBUFX2TS U536 ( .A(cacheDataOut[31]), .Y(n512) );
  CLKBUFX2TS U537 ( .A(cacheDataOut[29]), .Y(n513) );
  CLKBUFX2TS U538 ( .A(cacheDataOut[29]), .Y(n514) );
  CLKBUFX2TS U539 ( .A(cacheDataOut[26]), .Y(n515) );
  CLKBUFX2TS U540 ( .A(cacheDataOut[26]), .Y(n516) );
  CLKBUFX2TS U541 ( .A(cacheDataOut[25]), .Y(n517) );
  CLKBUFX2TS U542 ( .A(cacheDataOut[25]), .Y(n518) );
  CLKBUFX2TS U543 ( .A(cacheDataOut[24]), .Y(n519) );
  CLKBUFX2TS U544 ( .A(cacheDataOut[24]), .Y(n520) );
  CLKBUFX2TS U545 ( .A(cacheDataOut[22]), .Y(n521) );
  CLKBUFX2TS U546 ( .A(cacheDataOut[22]), .Y(n522) );
  CLKBUFX2TS U547 ( .A(cacheDataOut[21]), .Y(n523) );
  CLKBUFX2TS U548 ( .A(cacheDataOut[21]), .Y(n524) );
  CLKBUFX2TS U549 ( .A(cacheDataOut[19]), .Y(n525) );
  CLKBUFX2TS U550 ( .A(cacheDataOut[19]), .Y(n526) );
  CLKBUFX2TS U551 ( .A(cacheDataOut[18]), .Y(n527) );
  CLKBUFX2TS U552 ( .A(cacheDataOut[18]), .Y(n528) );
  CLKBUFX2TS U553 ( .A(cacheDataOut[17]), .Y(n529) );
  CLKBUFX2TS U554 ( .A(cacheDataOut[17]), .Y(n530) );
  CLKBUFX2TS U555 ( .A(cacheDataOut[15]), .Y(n531) );
  CLKBUFX2TS U556 ( .A(cacheDataOut[15]), .Y(n532) );
  CLKBUFX2TS U557 ( .A(cacheDataOut[14]), .Y(n533) );
  CLKBUFX2TS U558 ( .A(cacheDataOut[14]), .Y(n534) );
  CLKBUFX2TS U559 ( .A(cacheDataOut[13]), .Y(n535) );
  CLKBUFX2TS U560 ( .A(cacheDataOut[13]), .Y(n536) );
  CLKBUFX2TS U561 ( .A(cacheDataOut[1]), .Y(n537) );
  CLKBUFX2TS U562 ( .A(cacheDataOut[1]), .Y(n538) );
  CLKBUFX2TS U563 ( .A(cacheDataOut[0]), .Y(n539) );
  CLKBUFX2TS U564 ( .A(cacheDataOut[0]), .Y(n540) );
  AND3X2TS U565 ( .A(n104), .B(n448), .C(n1811), .Y(n1759) );
  INVX2TS U566 ( .A(n1759), .Y(n541) );
  INVX2TS U567 ( .A(n1759), .Y(n542) );
  INVX2TS U568 ( .A(n1759), .Y(n543) );
  AND2X2TS U569 ( .A(n752), .B(n453), .Y(n1761) );
  INVX2TS U570 ( .A(n1761), .Y(n544) );
  INVX2TS U571 ( .A(n1761), .Y(n545) );
  INVX2TS U572 ( .A(n1761), .Y(n546) );
  INVX1TS U573 ( .A(n1754), .Y(n547) );
  INVXLTS U574 ( .A(n1754), .Y(n548) );
  INVXLTS U575 ( .A(n1754), .Y(n549) );
  CLKINVX2TS U576 ( .A(n547), .Y(n734) );
  CLKBUFX2TS U577 ( .A(n139), .Y(n923) );
  INVX2TS U578 ( .A(n923), .Y(n550) );
  INVX2TS U579 ( .A(n923), .Y(n551) );
  INVX2TS U580 ( .A(n923), .Y(n552) );
  AND2XLTS U581 ( .A(n1772), .B(n742), .Y(n1118) );
  CLKINVX2TS U582 ( .A(n1118), .Y(n718) );
  INVXLTS U583 ( .A(n1118), .Y(n721) );
  INVXLTS U584 ( .A(n1118), .Y(n723) );
  INVXLTS U585 ( .A(n1118), .Y(n725) );
  AO21X4TS U586 ( .A0(n726), .A1(n727), .B0(n729), .Y(n2014) );
  XNOR2XLTS U587 ( .A(n959), .B(selectBit_SOUTH), .Y(n727) );
  OA21XLTS U588 ( .A0(n2907), .A1(n454), .B0(selectBit_EAST), .Y(n729) );
  INVXLTS U589 ( .A(n472), .Y(n731) );
  NOR2XLTS U590 ( .A(n1765), .B(n1769), .Y(n1105) );
  NAND2XLTS U591 ( .A(n171), .B(n4541), .Y(n1088) );
  NAND2X1TS U592 ( .A(n5327), .B(n915), .Y(n1871) );
  INVXLTS U593 ( .A(n3610), .Y(n3605) );
  INVXLTS U594 ( .A(n3610), .Y(n3604) );
  NOR2BXLTS U595 ( .AN(n1799), .B(n748), .Y(n1185) );
  INVX1TS U596 ( .A(n541), .Y(n730) );
  INVXLTS U597 ( .A(n1928), .Y(n760) );
  INVX1TS U598 ( .A(n2017), .Y(n957) );
  NAND3XLTS U599 ( .A(n1847), .B(n756), .C(n930), .Y(n1805) );
  INVXLTS U600 ( .A(n2006), .Y(n927) );
  NAND2XLTS U601 ( .A(n2006), .B(n117), .Y(n1914) );
  NOR2BXLTS U602 ( .AN(n1831), .B(n1976), .Y(n1202) );
  NAND2XLTS U603 ( .A(n915), .B(n4541), .Y(n1087) );
  OA22X1TS U604 ( .A0(n1781), .A1(n171), .B0(n1842), .B1(n1884), .Y(n733) );
  NOR2BXLTS U605 ( .AN(n1831), .B(n456), .Y(n1104) );
  NOR2BXLTS U606 ( .AN(n1831), .B(n1884), .Y(n1138) );
  AOI22XLTS U607 ( .A0(n3362), .A1(n43), .B0(n3345), .B1(n4034), .Y(n1196) );
  AOI22XLTS U608 ( .A0(n3361), .A1(n21), .B0(n3344), .B1(n4022), .Y(n1188) );
  AOI22XLTS U609 ( .A0(n3362), .A1(n16), .B0(n3345), .B1(n4019), .Y(n1183) );
  AOI22XLTS U610 ( .A0(n3361), .A1(n31), .B0(n3344), .B1(n4028), .Y(n1192) );
  AOI22XLTS U611 ( .A0(n3361), .A1(n26), .B0(n3344), .B1(n4025), .Y(n1190) );
  INVXLTS U612 ( .A(n3610), .Y(n3606) );
  INVXLTS U613 ( .A(selectBit_WEST), .Y(n1028) );
  NAND2XLTS U614 ( .A(n446), .B(n5327), .Y(n1870) );
  NAND2XLTS U615 ( .A(readReady), .B(n4), .Y(n1841) );
  NAND2XLTS U616 ( .A(selectBit_WEST), .B(readReady), .Y(n2903) );
  INVXLTS U617 ( .A(readReady), .Y(n1083) );
  INVXLTS U618 ( .A(n3457), .Y(n3452) );
  INVXLTS U619 ( .A(n3405), .Y(n3400) );
  INVXLTS U620 ( .A(n3456), .Y(n3453) );
  INVXLTS U621 ( .A(n3404), .Y(n3401) );
  INVXLTS U622 ( .A(n3455), .Y(n3454) );
  INVXLTS U623 ( .A(n3403), .Y(n3402) );
  INVX1TS U624 ( .A(n463), .Y(n740) );
  INVX1TS U625 ( .A(n544), .Y(n728) );
  INVX1TS U626 ( .A(n1182), .Y(n3409) );
  CLKAND2X2TS U627 ( .A(n1816), .B(n1813), .Y(n1219) );
  AND2XLTS U628 ( .A(n755), .B(n439), .Y(n737) );
  CLKBUFX2TS U629 ( .A(n3114), .Y(n3109) );
  CLKBUFX2TS U630 ( .A(n3114), .Y(n3108) );
  CLKBUFX2TS U631 ( .A(n3343), .Y(n3340) );
  CLKBUFX2TS U632 ( .A(n3343), .Y(n3341) );
  CLKBUFX2TS U633 ( .A(n3609), .Y(n3607) );
  CLKBUFX2TS U634 ( .A(n3260), .Y(n3257) );
  CLKBUFX2TS U635 ( .A(n3260), .Y(n3258) );
  CLKBUFX2TS U636 ( .A(n3096), .Y(n3092) );
  INVXLTS U637 ( .A(n1768), .Y(n750) );
  OAI31XLTS U638 ( .A0(n111), .A1(n107), .A2(n931), .B0(n915), .Y(n1842) );
  AOI21XLTS U639 ( .A0(n1844), .A1(n1779), .B0(n757), .Y(n1781) );
  NOR2BXLTS U640 ( .AN(n1776), .B(n1780), .Y(n1140) );
  NOR2BXLTS U641 ( .AN(n1807), .B(n1810), .Y(n1203) );
  NAND2XLTS U642 ( .A(n1794), .B(n1844), .Y(n1765) );
  OR4XLTS U643 ( .A(n440), .B(n745), .C(n759), .D(n750), .Y(n743) );
  CLKINVX2TS U644 ( .A(n108), .Y(n751) );
  AND2XLTS U645 ( .A(n452), .B(n444), .Y(n738) );
  OAI21XLTS U646 ( .A0(n957), .A1(n2904), .B0(n2392), .Y(n2890) );
  NAND2XLTS U647 ( .A(n957), .B(n2904), .Y(n2392) );
  OAI22XLTS U648 ( .A0(n109), .A1(n969), .B0(n751), .B1(n972), .Y(n1797) );
  NAND2XLTS U649 ( .A(n4190), .B(n755), .Y(n1792) );
  NAND3XLTS U650 ( .A(n1845), .B(n445), .C(n1847), .Y(n1766) );
  NAND2X1TS U651 ( .A(n110), .B(n5323), .Y(n1812) );
  OAI21XLTS U652 ( .A0(n926), .A1(n2009), .B0(n109), .Y(n2008) );
  AOI21XLTS U653 ( .A0(n971), .A1(n2010), .B0(n2006), .Y(n1940) );
  NOR2X2TS U654 ( .A(n959), .B(n971), .Y(n2907) );
  NAND3XLTS U655 ( .A(n930), .B(n44), .C(n1893), .Y(n2007) );
  CLKINVX2TS U656 ( .A(n1804), .Y(n739) );
  CLKINVX2TS U657 ( .A(n1616), .Y(n3115) );
  OAI22XLTS U658 ( .A0(n1773), .A1(n172), .B0(n1832), .B1(n1871), .Y(n1616) );
  NAND2XLTS U659 ( .A(n4189), .B(n753), .Y(n1808) );
  OAI21XLTS U660 ( .A0(n2383), .A1(n958), .B0(n2903), .Y(n2904) );
  AOI32XLTS U661 ( .A0(n101), .A1(n1777), .A2(n1778), .B0(n3610), .B1(n654), 
        .Y(n2568) );
  NAND2XLTS U662 ( .A(n4189), .B(n757), .Y(n1777) );
  AOI32XLTS U663 ( .A0(n447), .A1(n1780), .A2(n4195), .B0(n1781), .B1(n1782), 
        .Y(n1778) );
  OA21XLTS U664 ( .A0(n2893), .A1(n2894), .B0(n2895), .Y(n2391) );
  AOI22XLTS U665 ( .A0(n1768), .A1(n434), .B0(n750), .B1(n972), .Y(n1767) );
  OAI22XLTS U666 ( .A0(n747), .A1(n969), .B0(n448), .B1(n972), .Y(n1782) );
  NAND2X1TS U667 ( .A(n926), .B(n113), .Y(n1976) );
  NOR2X1TS U668 ( .A(readReady), .B(selectBit_WEST), .Y(n2383) );
  NAND2XLTS U669 ( .A(n4189), .B(n452), .Y(n1784) );
  AOI21XLTS U670 ( .A0(readIn_NORTH), .A1(n1816), .B0(n1817), .Y(n1815) );
  OAI211XLTS U671 ( .A0(n3100), .A1(n637), .B0(n1679), .C0(n1680), .Y(n2611)
         );
  OAI211XLTS U672 ( .A0(n3100), .A1(n636), .B0(n1677), .C0(n1678), .Y(n2612)
         );
  OAI211XLTS U673 ( .A0(n3595), .A1(n806), .B0(n1882), .C0(n1883), .Y(n2529)
         );
  OAI211XLTS U674 ( .A0(n3245), .A1(n646), .B0(n1228), .C0(n1229), .Y(n2836)
         );
  OAI211XLTS U675 ( .A0(n3245), .A1(n645), .B0(n1224), .C0(n1225), .Y(n2838)
         );
  OAI211XLTS U676 ( .A0(n3245), .A1(n644), .B0(n1222), .C0(n1223), .Y(n2839)
         );
  OAI211XLTS U677 ( .A0(n3328), .A1(n840), .B0(n1974), .C0(n1975), .Y(n2473)
         );
  OAI211XLTS U678 ( .A0(n3520), .A1(n4246), .B0(n1490), .C0(n1491), .Y(n2705)
         );
  OAI211XLTS U679 ( .A0(n3520), .A1(n4243), .B0(n1488), .C0(n1489), .Y(n2706)
         );
  OAI211XLTS U680 ( .A0(n3453), .A1(n4246), .B0(n1426), .C0(n1427), .Y(n2737)
         );
  OAI211XLTS U681 ( .A0(n3453), .A1(n4243), .B0(n1424), .C0(n1425), .Y(n2738)
         );
  OAI211XLTS U682 ( .A0(n3328), .A1(n903), .B0(n1209), .C0(n1210), .Y(n2843)
         );
  OAI211XLTS U683 ( .A0(n3328), .A1(n901), .B0(n1205), .C0(n1206), .Y(n2845)
         );
  OAI211XLTS U684 ( .A0(n3401), .A1(n4342), .B0(n1362), .C0(n1363), .Y(n2769)
         );
  OAI211XLTS U685 ( .A0(n3401), .A1(n4339), .B0(n1360), .C0(n1361), .Y(n2770)
         );
  OAI211XLTS U686 ( .A0(n3251), .A1(n675), .B0(n1288), .C0(n1289), .Y(n2806)
         );
  OAI211XLTS U687 ( .A0(n3251), .A1(n677), .B0(n1994), .C0(n1995), .Y(n2460)
         );
  OAI211XLTS U688 ( .A0(n3105), .A1(n955), .B0(n1641), .C0(n1642), .Y(n2630)
         );
  OAI211XLTS U689 ( .A0(n3105), .A1(n954), .B0(n1643), .C0(n1644), .Y(n2629)
         );
  OAI211XLTS U690 ( .A0(n3104), .A1(n953), .B0(n1645), .C0(n1646), .Y(n2628)
         );
  OAI211XLTS U691 ( .A0(n3104), .A1(n952), .B0(n1647), .C0(n1648), .Y(n2627)
         );
  OAI211XLTS U692 ( .A0(n3104), .A1(n951), .B0(n1649), .C0(n1650), .Y(n2626)
         );
  OAI211XLTS U693 ( .A0(n3104), .A1(n950), .B0(n1651), .C0(n1652), .Y(n2625)
         );
  OAI211XLTS U694 ( .A0(n3103), .A1(n949), .B0(n1653), .C0(n1654), .Y(n2624)
         );
  OAI211XLTS U695 ( .A0(n3103), .A1(n948), .B0(n1655), .C0(n1656), .Y(n2623)
         );
  OAI211XLTS U696 ( .A0(n3103), .A1(n947), .B0(n1657), .C0(n1658), .Y(n2622)
         );
  OAI211XLTS U697 ( .A0(n3103), .A1(n946), .B0(n1659), .C0(n1660), .Y(n2621)
         );
  OAI211XLTS U698 ( .A0(n3102), .A1(n945), .B0(n1661), .C0(n1662), .Y(n2620)
         );
  OAI211XLTS U699 ( .A0(n3102), .A1(n944), .B0(n1663), .C0(n1664), .Y(n2619)
         );
  OAI211XLTS U700 ( .A0(n3102), .A1(n943), .B0(n1665), .C0(n1666), .Y(n2618)
         );
  OAI211XLTS U701 ( .A0(n3102), .A1(n942), .B0(n1667), .C0(n1668), .Y(n2617)
         );
  OAI211XLTS U702 ( .A0(n3101), .A1(n941), .B0(n1669), .C0(n1670), .Y(n2616)
         );
  OAI211XLTS U703 ( .A0(n3101), .A1(n940), .B0(n1671), .C0(n1672), .Y(n2615)
         );
  OAI211XLTS U704 ( .A0(n3101), .A1(n939), .B0(n1673), .C0(n1674), .Y(n2614)
         );
  OAI211XLTS U705 ( .A0(n3101), .A1(n938), .B0(n1675), .C0(n1676), .Y(n2613)
         );
  OAI211XLTS U706 ( .A0(n3105), .A1(n642), .B0(n1637), .C0(n1638), .Y(n2632)
         );
  OAI211XLTS U707 ( .A0(n3106), .A1(n641), .B0(n1629), .C0(n1630), .Y(n2636)
         );
  OAI211XLTS U708 ( .A0(n3105), .A1(n635), .B0(n1639), .C0(n1640), .Y(n2631)
         );
  OAI211XLTS U709 ( .A0(n3106), .A1(n634), .B0(n1635), .C0(n1636), .Y(n2633)
         );
  OAI211XLTS U710 ( .A0(n3106), .A1(n633), .B0(n1633), .C0(n1634), .Y(n2634)
         );
  OAI211XLTS U711 ( .A0(n3106), .A1(n632), .B0(n1631), .C0(n1632), .Y(n2635)
         );
  OAI211XLTS U712 ( .A0(n3107), .A1(n631), .B0(n1627), .C0(n1628), .Y(n2637)
         );
  OAI211XLTS U713 ( .A0(n3107), .A1(n595), .B0(n1625), .C0(n1626), .Y(n2638)
         );
  OAI211XLTS U714 ( .A0(n3107), .A1(n630), .B0(n1623), .C0(n1624), .Y(n2639)
         );
  OAI211XLTS U715 ( .A0(n3107), .A1(n629), .B0(n1621), .C0(n1622), .Y(n2640)
         );
  OAI211XLTS U716 ( .A0(n3511), .A1(n3994), .B0(n1904), .C0(n1905), .Y(n2515)
         );
  OAI211XLTS U717 ( .A0(n3511), .A1(n3988), .B0(n1900), .C0(n1901), .Y(n2517)
         );
  OAI211XLTS U718 ( .A0(n3511), .A1(n3985), .B0(n1898), .C0(n1899), .Y(n2518)
         );
  OAI211XLTS U719 ( .A0(n3512), .A1(n3982), .B0(n1896), .C0(n1897), .Y(n2519)
         );
  OAI211XLTS U720 ( .A0(n3512), .A1(n3979), .B0(n1894), .C0(n1895), .Y(n2520)
         );
  OAI211XLTS U721 ( .A0(n3512), .A1(n4333), .B0(n1548), .C0(n1549), .Y(n2676)
         );
  OAI211XLTS U722 ( .A0(n3513), .A1(n4327), .B0(n1544), .C0(n1545), .Y(n2678)
         );
  OAI211XLTS U723 ( .A0(n3513), .A1(n4324), .B0(n1542), .C0(n1543), .Y(n2679)
         );
  OAI211XLTS U724 ( .A0(n3513), .A1(n4321), .B0(n1540), .C0(n1541), .Y(n2680)
         );
  OAI211XLTS U725 ( .A0(n3514), .A1(n4318), .B0(n1538), .C0(n1539), .Y(n2681)
         );
  OAI211XLTS U726 ( .A0(n3514), .A1(n4315), .B0(n1536), .C0(n1537), .Y(n2682)
         );
  OAI211XLTS U727 ( .A0(n3514), .A1(n4312), .B0(n1534), .C0(n1535), .Y(n2683)
         );
  OAI211XLTS U728 ( .A0(n3515), .A1(n4297), .B0(n1524), .C0(n1525), .Y(n2688)
         );
  OAI211XLTS U729 ( .A0(n3517), .A1(n4282), .B0(n1514), .C0(n1515), .Y(n2693)
         );
  OAI211XLTS U730 ( .A0(n3518), .A1(n4270), .B0(n1506), .C0(n1507), .Y(n2697)
         );
  OAI211XLTS U731 ( .A0(n3518), .A1(n4264), .B0(n1502), .C0(n1503), .Y(n2699)
         );
  OAI211XLTS U732 ( .A0(n3519), .A1(n4258), .B0(n1498), .C0(n1499), .Y(n2701)
         );
  OAI211XLTS U733 ( .A0(n3519), .A1(n4255), .B0(n1496), .C0(n1497), .Y(n2702)
         );
  OAI211XLTS U734 ( .A0(n3519), .A1(n4249), .B0(n1492), .C0(n1493), .Y(n2704)
         );
  OAI211XLTS U735 ( .A0(n3512), .A1(n4336), .B0(n1550), .C0(n1551), .Y(n2675)
         );
  OAI211XLTS U736 ( .A0(n3513), .A1(n4330), .B0(n1546), .C0(n1547), .Y(n2677)
         );
  OAI211XLTS U737 ( .A0(n3514), .A1(n4309), .B0(n1532), .C0(n1533), .Y(n2684)
         );
  OAI211XLTS U738 ( .A0(n3515), .A1(n4306), .B0(n1530), .C0(n1531), .Y(n2685)
         );
  OAI211XLTS U739 ( .A0(n3515), .A1(n4303), .B0(n1528), .C0(n1529), .Y(n2686)
         );
  OAI211XLTS U740 ( .A0(n3515), .A1(n4300), .B0(n1526), .C0(n1527), .Y(n2687)
         );
  OAI211XLTS U741 ( .A0(n3516), .A1(n4291), .B0(n1520), .C0(n1521), .Y(n2690)
         );
  OAI211XLTS U742 ( .A0(n3517), .A1(n4279), .B0(n1512), .C0(n1513), .Y(n2694)
         );
  OAI211XLTS U743 ( .A0(n3517), .A1(n4276), .B0(n1510), .C0(n1511), .Y(n2695)
         );
  OAI211XLTS U744 ( .A0(n3517), .A1(n4273), .B0(n1508), .C0(n1509), .Y(n2696)
         );
  OAI211XLTS U745 ( .A0(n3518), .A1(n4267), .B0(n1504), .C0(n1505), .Y(n2698)
         );
  OAI211XLTS U746 ( .A0(n3518), .A1(n4261), .B0(n1500), .C0(n1501), .Y(n2700)
         );
  OAI211XLTS U747 ( .A0(n3516), .A1(n4294), .B0(n1522), .C0(n1523), .Y(n2689)
         );
  OAI211XLTS U748 ( .A0(n3516), .A1(n4288), .B0(n1518), .C0(n1519), .Y(n2691)
         );
  OAI211XLTS U749 ( .A0(n3516), .A1(n4285), .B0(n1516), .C0(n1517), .Y(n2692)
         );
  OAI211XLTS U750 ( .A0(n3519), .A1(n4252), .B0(n1494), .C0(n1495), .Y(n2703)
         );
  OAI211XLTS U751 ( .A0(n3511), .A1(n3991), .B0(n1902), .C0(n1903), .Y(n2516)
         );
  OAI211XLTS U752 ( .A0(n3445), .A1(n3982), .B0(n1918), .C0(n1919), .Y(n2505)
         );
  OAI211XLTS U753 ( .A0(n3445), .A1(n3979), .B0(n1916), .C0(n1917), .Y(n2506)
         );
  OAI211XLTS U754 ( .A0(n3445), .A1(n4336), .B0(n1486), .C0(n1487), .Y(n2707)
         );
  OAI211XLTS U755 ( .A0(n3445), .A1(n4333), .B0(n1484), .C0(n1485), .Y(n2708)
         );
  OAI211XLTS U756 ( .A0(n3446), .A1(n4330), .B0(n1482), .C0(n1483), .Y(n2709)
         );
  OAI211XLTS U757 ( .A0(n3446), .A1(n4327), .B0(n1480), .C0(n1481), .Y(n2710)
         );
  OAI211XLTS U758 ( .A0(n3446), .A1(n4324), .B0(n1478), .C0(n1479), .Y(n2711)
         );
  OAI211XLTS U759 ( .A0(n3446), .A1(n4321), .B0(n1476), .C0(n1477), .Y(n2712)
         );
  OAI211XLTS U760 ( .A0(n3447), .A1(n4315), .B0(n1472), .C0(n1473), .Y(n2714)
         );
  OAI211XLTS U761 ( .A0(n3447), .A1(n4309), .B0(n1468), .C0(n1469), .Y(n2716)
         );
  OAI211XLTS U762 ( .A0(n3448), .A1(n4306), .B0(n1466), .C0(n1467), .Y(n2717)
         );
  OAI211XLTS U763 ( .A0(n3448), .A1(n4300), .B0(n1462), .C0(n1463), .Y(n2719)
         );
  OAI211XLTS U764 ( .A0(n3449), .A1(n4294), .B0(n1458), .C0(n1459), .Y(n2721)
         );
  OAI211XLTS U765 ( .A0(n3449), .A1(n4291), .B0(n1456), .C0(n1457), .Y(n2722)
         );
  OAI211XLTS U766 ( .A0(n3449), .A1(n4285), .B0(n1452), .C0(n1453), .Y(n2724)
         );
  OAI211XLTS U767 ( .A0(n3450), .A1(n4279), .B0(n1448), .C0(n1449), .Y(n2726)
         );
  OAI211XLTS U768 ( .A0(n3450), .A1(n4276), .B0(n1446), .C0(n1447), .Y(n2727)
         );
  OAI211XLTS U769 ( .A0(n3450), .A1(n4273), .B0(n1444), .C0(n1445), .Y(n2728)
         );
  OAI211XLTS U770 ( .A0(n3451), .A1(n4270), .B0(n1442), .C0(n1443), .Y(n2729)
         );
  OAI211XLTS U771 ( .A0(n3451), .A1(n4267), .B0(n1440), .C0(n1441), .Y(n2730)
         );
  OAI211XLTS U772 ( .A0(n3451), .A1(n4261), .B0(n1436), .C0(n1437), .Y(n2732)
         );
  OAI211XLTS U773 ( .A0(n3452), .A1(n4252), .B0(n1430), .C0(n1431), .Y(n2735)
         );
  OAI211XLTS U774 ( .A0(n3447), .A1(n4318), .B0(n1474), .C0(n1475), .Y(n2713)
         );
  OAI211XLTS U775 ( .A0(n3447), .A1(n4312), .B0(n1470), .C0(n1471), .Y(n2715)
         );
  OAI211XLTS U776 ( .A0(n3448), .A1(n4303), .B0(n1464), .C0(n1465), .Y(n2718)
         );
  OAI211XLTS U777 ( .A0(n3448), .A1(n4297), .B0(n1460), .C0(n1461), .Y(n2720)
         );
  OAI211XLTS U778 ( .A0(n3449), .A1(n4288), .B0(n1454), .C0(n1455), .Y(n2723)
         );
  OAI211XLTS U779 ( .A0(n3450), .A1(n4282), .B0(n1450), .C0(n1451), .Y(n2725)
         );
  OAI211XLTS U780 ( .A0(n3452), .A1(n4258), .B0(n1434), .C0(n1435), .Y(n2733)
         );
  OAI211XLTS U781 ( .A0(n3452), .A1(n4255), .B0(n1432), .C0(n1433), .Y(n2734)
         );
  OAI211XLTS U782 ( .A0(n3452), .A1(n4249), .B0(n1428), .C0(n1429), .Y(n2736)
         );
  OAI211XLTS U783 ( .A0(n3451), .A1(n4264), .B0(n1438), .C0(n1439), .Y(n2731)
         );
  OAI211XLTS U784 ( .A0(n3444), .A1(n3988), .B0(n1922), .C0(n1923), .Y(n2503)
         );
  OAI211XLTS U785 ( .A0(n3444), .A1(n3985), .B0(n1920), .C0(n1921), .Y(n2504)
         );
  OAI211XLTS U786 ( .A0(n3444), .A1(n3994), .B0(n1926), .C0(n1927), .Y(n2501)
         );
  OAI211XLTS U787 ( .A0(n3444), .A1(n3991), .B0(n1924), .C0(n1925), .Y(n2502)
         );
  OAI211XLTS U788 ( .A0(n3604), .A1(n811), .B0(n1614), .C0(n1615), .Y(n2643)
         );
  OAI211XLTS U789 ( .A0(n3601), .A1(n810), .B0(n1584), .C0(n1585), .Y(n2658)
         );
  OAI211XLTS U790 ( .A0(n3600), .A1(n809), .B0(n1582), .C0(n1583), .Y(n2659)
         );
  OAI211XLTS U791 ( .A0(n3599), .A1(n808), .B0(n1574), .C0(n1575), .Y(n2663)
         );
  OAI211XLTS U792 ( .A0(n3597), .A1(n807), .B0(n1554), .C0(n1555), .Y(n2673)
         );
  OAI211XLTS U793 ( .A0(n3604), .A1(n801), .B0(n1612), .C0(n1613), .Y(n2644)
         );
  OAI211XLTS U794 ( .A0(n3604), .A1(n800), .B0(n1610), .C0(n1611), .Y(n2645)
         );
  OAI211XLTS U795 ( .A0(n3604), .A1(n799), .B0(n1608), .C0(n1609), .Y(n2646)
         );
  OAI211XLTS U796 ( .A0(n3603), .A1(n798), .B0(n1606), .C0(n1607), .Y(n2647)
         );
  OAI211XLTS U797 ( .A0(n3603), .A1(n797), .B0(n1604), .C0(n1605), .Y(n2648)
         );
  OAI211XLTS U798 ( .A0(n3603), .A1(n796), .B0(n1602), .C0(n1603), .Y(n2649)
         );
  OAI211XLTS U799 ( .A0(n3603), .A1(n795), .B0(n1600), .C0(n1601), .Y(n2650)
         );
  OAI211XLTS U800 ( .A0(n3602), .A1(n794), .B0(n1598), .C0(n1599), .Y(n2651)
         );
  OAI211XLTS U801 ( .A0(n3602), .A1(n793), .B0(n1596), .C0(n1597), .Y(n2652)
         );
  OAI211XLTS U802 ( .A0(n3602), .A1(n792), .B0(n1594), .C0(n1595), .Y(n2653)
         );
  OAI211XLTS U803 ( .A0(n3602), .A1(n791), .B0(n1592), .C0(n1593), .Y(n2654)
         );
  OAI211XLTS U804 ( .A0(n3601), .A1(n790), .B0(n1590), .C0(n1591), .Y(n2655)
         );
  OAI211XLTS U805 ( .A0(n3601), .A1(n789), .B0(n1588), .C0(n1589), .Y(n2656)
         );
  OAI211XLTS U806 ( .A0(n3601), .A1(n788), .B0(n1586), .C0(n1587), .Y(n2657)
         );
  OAI211XLTS U807 ( .A0(n3600), .A1(n787), .B0(n1580), .C0(n1581), .Y(n2660)
         );
  OAI211XLTS U808 ( .A0(n3600), .A1(n786), .B0(n1578), .C0(n1579), .Y(n2661)
         );
  OAI211XLTS U809 ( .A0(n3599), .A1(n785), .B0(n1576), .C0(n1577), .Y(n2662)
         );
  OAI211XLTS U810 ( .A0(n3599), .A1(n784), .B0(n1572), .C0(n1573), .Y(n2664)
         );
  OAI211XLTS U811 ( .A0(n3599), .A1(n783), .B0(n1570), .C0(n1571), .Y(n2665)
         );
  OAI211XLTS U812 ( .A0(n3598), .A1(n782), .B0(n1568), .C0(n1569), .Y(n2666)
         );
  OAI211XLTS U813 ( .A0(n3598), .A1(n781), .B0(n1566), .C0(n1567), .Y(n2667)
         );
  OAI211XLTS U814 ( .A0(n3598), .A1(n780), .B0(n1564), .C0(n1565), .Y(n2668)
         );
  OAI211XLTS U815 ( .A0(n3598), .A1(n779), .B0(n1562), .C0(n1563), .Y(n2669)
         );
  OAI211XLTS U816 ( .A0(n3597), .A1(n778), .B0(n1560), .C0(n1561), .Y(n2670)
         );
  OAI211XLTS U817 ( .A0(n3597), .A1(n777), .B0(n1558), .C0(n1559), .Y(n2671)
         );
  OAI211XLTS U818 ( .A0(n3597), .A1(n776), .B0(n1556), .C0(n1557), .Y(n2672)
         );
  OAI211XLTS U819 ( .A0(n3596), .A1(n775), .B0(n1552), .C0(n1553), .Y(n2674)
         );
  OAI211XLTS U820 ( .A0(n3392), .A1(n3943), .B0(n1945), .C0(n1946), .Y(n2490)
         );
  OAI211XLTS U821 ( .A0(n3393), .A1(n4431), .B0(n1420), .C0(n1421), .Y(n2740)
         );
  OAI211XLTS U822 ( .A0(n3394), .A1(n4428), .B0(n1418), .C0(n1419), .Y(n2741)
         );
  OAI211XLTS U823 ( .A0(n3394), .A1(n4425), .B0(n1416), .C0(n1417), .Y(n2742)
         );
  OAI211XLTS U824 ( .A0(n3394), .A1(n4417), .B0(n1412), .C0(n1413), .Y(n2744)
         );
  OAI211XLTS U825 ( .A0(n3395), .A1(n4414), .B0(n1410), .C0(n1411), .Y(n2745)
         );
  OAI211XLTS U826 ( .A0(n3395), .A1(n4408), .B0(n1406), .C0(n1407), .Y(n2747)
         );
  OAI211XLTS U827 ( .A0(n3396), .A1(n4402), .B0(n1402), .C0(n1403), .Y(n2749)
         );
  OAI211XLTS U828 ( .A0(n3396), .A1(n4399), .B0(n1400), .C0(n1401), .Y(n2750)
         );
  OAI211XLTS U829 ( .A0(n3396), .A1(n4396), .B0(n1398), .C0(n1399), .Y(n2751)
         );
  OAI211XLTS U830 ( .A0(n3396), .A1(n4393), .B0(n1396), .C0(n1397), .Y(n2752)
         );
  OAI211XLTS U831 ( .A0(n3397), .A1(n4390), .B0(n1394), .C0(n1395), .Y(n2753)
         );
  OAI211XLTS U832 ( .A0(n3397), .A1(n4384), .B0(n1390), .C0(n1391), .Y(n2755)
         );
  OAI211XLTS U833 ( .A0(n3397), .A1(n4381), .B0(n1388), .C0(n1389), .Y(n2756)
         );
  OAI211XLTS U834 ( .A0(n3398), .A1(n4378), .B0(n1386), .C0(n1387), .Y(n2757)
         );
  OAI211XLTS U835 ( .A0(n3398), .A1(n4375), .B0(n1384), .C0(n1385), .Y(n2758)
         );
  OAI211XLTS U836 ( .A0(n3398), .A1(n4372), .B0(n1382), .C0(n1383), .Y(n2759)
         );
  OAI211XLTS U837 ( .A0(n3399), .A1(n4366), .B0(n1378), .C0(n1379), .Y(n2761)
         );
  OAI211XLTS U838 ( .A0(n3399), .A1(n4363), .B0(n1376), .C0(n1377), .Y(n2762)
         );
  OAI211XLTS U839 ( .A0(n3399), .A1(n4360), .B0(n1374), .C0(n1375), .Y(n2763)
         );
  OAI211XLTS U840 ( .A0(n3400), .A1(n4354), .B0(n1370), .C0(n1371), .Y(n2765)
         );
  OAI211XLTS U841 ( .A0(n3400), .A1(n4351), .B0(n1368), .C0(n1369), .Y(n2766)
         );
  OAI211XLTS U842 ( .A0(n3400), .A1(n4348), .B0(n1366), .C0(n1367), .Y(n2767)
         );
  OAI211XLTS U843 ( .A0(n3392), .A1(n3952), .B0(n1951), .C0(n1952), .Y(n2487)
         );
  OAI211XLTS U844 ( .A0(n3392), .A1(n3949), .B0(n1949), .C0(n1950), .Y(n2488)
         );
  OAI211XLTS U845 ( .A0(n3392), .A1(n3946), .B0(n1947), .C0(n1948), .Y(n2489)
         );
  OAI211XLTS U846 ( .A0(n3393), .A1(n3940), .B0(n1943), .C0(n1944), .Y(n2491)
         );
  OAI211XLTS U847 ( .A0(n3393), .A1(n3937), .B0(n1941), .C0(n1942), .Y(n2492)
         );
  OAI211XLTS U848 ( .A0(n3394), .A1(n4420), .B0(n1414), .C0(n1415), .Y(n2743)
         );
  OAI211XLTS U849 ( .A0(n3398), .A1(n4369), .B0(n1380), .C0(n1381), .Y(n2760)
         );
  OAI211XLTS U850 ( .A0(n3393), .A1(n4435), .B0(n1422), .C0(n1423), .Y(n2739)
         );
  OAI211XLTS U851 ( .A0(n3395), .A1(n4411), .B0(n1408), .C0(n1409), .Y(n2746)
         );
  OAI211XLTS U852 ( .A0(n3395), .A1(n4405), .B0(n1404), .C0(n1405), .Y(n2748)
         );
  OAI211XLTS U853 ( .A0(n3397), .A1(n4387), .B0(n1392), .C0(n1393), .Y(n2754)
         );
  OAI211XLTS U854 ( .A0(n3399), .A1(n4357), .B0(n1372), .C0(n1373), .Y(n2764)
         );
  OAI211XLTS U855 ( .A0(n3400), .A1(n4345), .B0(n1364), .C0(n1365), .Y(n2768)
         );
  OAI211XLTS U856 ( .A0(n3247), .A1(n669), .B0(n1236), .C0(n1237), .Y(n2832)
         );
  OAI211XLTS U857 ( .A0(n3246), .A1(n668), .B0(n1234), .C0(n1235), .Y(n2833)
         );
  OAI211XLTS U858 ( .A0(n3246), .A1(n667), .B0(n1232), .C0(n1233), .Y(n2834)
         );
  OAI211XLTS U859 ( .A0(n3249), .A1(n685), .B0(n1256), .C0(n1257), .Y(n2822)
         );
  OAI211XLTS U860 ( .A0(n3249), .A1(n684), .B0(n1254), .C0(n1255), .Y(n2823)
         );
  OAI211XLTS U861 ( .A0(n3249), .A1(n683), .B0(n1252), .C0(n1253), .Y(n2824)
         );
  OAI211XLTS U862 ( .A0(n3248), .A1(n682), .B0(n1248), .C0(n1249), .Y(n2826)
         );
  OAI211XLTS U863 ( .A0(n3248), .A1(n681), .B0(n1246), .C0(n1247), .Y(n2827)
         );
  OAI211XLTS U864 ( .A0(n3248), .A1(n680), .B0(n1244), .C0(n1245), .Y(n2828)
         );
  OAI211XLTS U865 ( .A0(n3247), .A1(n679), .B0(n1240), .C0(n1241), .Y(n2830)
         );
  OAI211XLTS U866 ( .A0(n3247), .A1(n678), .B0(n1238), .C0(n1239), .Y(n2831)
         );
  OAI211XLTS U867 ( .A0(n3250), .A1(n674), .B0(n1286), .C0(n1287), .Y(n2807)
         );
  OAI211XLTS U868 ( .A0(n3250), .A1(n673), .B0(n1278), .C0(n1279), .Y(n2811)
         );
  OAI211XLTS U869 ( .A0(n3250), .A1(n672), .B0(n1272), .C0(n1273), .Y(n2814)
         );
  OAI211XLTS U870 ( .A0(n3248), .A1(n671), .B0(n1250), .C0(n1251), .Y(n2825)
         );
  OAI211XLTS U871 ( .A0(n3247), .A1(n670), .B0(n1242), .C0(n1243), .Y(n2829)
         );
  OAI211XLTS U872 ( .A0(n3250), .A1(n676), .B0(n1986), .C0(n1987), .Y(n2464)
         );
  OAI211XLTS U873 ( .A0(n3246), .A1(n648), .B0(n1230), .C0(n1231), .Y(n2835)
         );
  OAI211XLTS U874 ( .A0(n3246), .A1(n647), .B0(n1226), .C0(n1227), .Y(n2837)
         );
  OAI211XLTS U875 ( .A0(n3249), .A1(n643), .B0(n1216), .C0(n1217), .Y(n2840)
         );
  OAI211XLTS U876 ( .A0(n3336), .A1(n848), .B0(n1350), .C0(n1351), .Y(n2775)
         );
  OAI211XLTS U877 ( .A0(n3335), .A1(n847), .B0(n1340), .C0(n1341), .Y(n2780)
         );
  OAI211XLTS U878 ( .A0(n3335), .A1(n846), .B0(n1336), .C0(n1337), .Y(n2782)
         );
  OAI211XLTS U879 ( .A0(n3334), .A1(n845), .B0(n1334), .C0(n1335), .Y(n2783)
         );
  OAI211XLTS U880 ( .A0(n3332), .A1(n844), .B0(n1316), .C0(n1317), .Y(n2792)
         );
  OAI211XLTS U881 ( .A0(n3331), .A1(n843), .B0(n1312), .C0(n1313), .Y(n2794)
         );
  OAI211XLTS U882 ( .A0(n3331), .A1(n842), .B0(n1306), .C0(n1307), .Y(n2797)
         );
  OAI211XLTS U883 ( .A0(n3330), .A1(n841), .B0(n1300), .C0(n1301), .Y(n2800)
         );
  OAI211XLTS U884 ( .A0(n3330), .A1(n813), .B0(n1298), .C0(n1299), .Y(n2801)
         );
  OAI211XLTS U885 ( .A0(n3329), .A1(n812), .B0(n1296), .C0(n1297), .Y(n2802)
         );
  OAI211XLTS U886 ( .A0(n3337), .A1(n835), .B0(n1358), .C0(n1359), .Y(n2771)
         );
  OAI211XLTS U887 ( .A0(n3337), .A1(n834), .B0(n1356), .C0(n1357), .Y(n2772)
         );
  OAI211XLTS U888 ( .A0(n3337), .A1(n833), .B0(n1354), .C0(n1355), .Y(n2773)
         );
  OAI211XLTS U889 ( .A0(n3337), .A1(n832), .B0(n1352), .C0(n1353), .Y(n2774)
         );
  OAI211XLTS U890 ( .A0(n3336), .A1(n831), .B0(n1348), .C0(n1349), .Y(n2776)
         );
  OAI211XLTS U891 ( .A0(n3336), .A1(n830), .B0(n1346), .C0(n1347), .Y(n2777)
         );
  OAI211XLTS U892 ( .A0(n3336), .A1(n829), .B0(n1344), .C0(n1345), .Y(n2778)
         );
  OAI211XLTS U893 ( .A0(n3335), .A1(n828), .B0(n1342), .C0(n1343), .Y(n2779)
         );
  OAI211XLTS U894 ( .A0(n3335), .A1(n827), .B0(n1338), .C0(n1339), .Y(n2781)
         );
  OAI211XLTS U895 ( .A0(n3334), .A1(n826), .B0(n1332), .C0(n1333), .Y(n2784)
         );
  OAI211XLTS U896 ( .A0(n3334), .A1(n825), .B0(n1330), .C0(n1331), .Y(n2785)
         );
  OAI211XLTS U897 ( .A0(n3334), .A1(n824), .B0(n1328), .C0(n1329), .Y(n2786)
         );
  OAI211XLTS U898 ( .A0(n3333), .A1(n823), .B0(n1326), .C0(n1327), .Y(n2787)
         );
  OAI211XLTS U899 ( .A0(n3333), .A1(n822), .B0(n1324), .C0(n1325), .Y(n2788)
         );
  OAI211XLTS U900 ( .A0(n3333), .A1(n821), .B0(n1322), .C0(n1323), .Y(n2789)
         );
  OAI211XLTS U901 ( .A0(n3332), .A1(n820), .B0(n1320), .C0(n1321), .Y(n2790)
         );
  OAI211XLTS U902 ( .A0(n3332), .A1(n819), .B0(n1318), .C0(n1319), .Y(n2791)
         );
  OAI211XLTS U903 ( .A0(n3332), .A1(n818), .B0(n1314), .C0(n1315), .Y(n2793)
         );
  OAI211XLTS U904 ( .A0(n3331), .A1(n817), .B0(n1310), .C0(n1311), .Y(n2795)
         );
  OAI211XLTS U905 ( .A0(n3331), .A1(n816), .B0(n1308), .C0(n1309), .Y(n2796)
         );
  OAI211XLTS U906 ( .A0(n3330), .A1(n815), .B0(n1304), .C0(n1305), .Y(n2798)
         );
  OAI211XLTS U907 ( .A0(n3330), .A1(n814), .B0(n1302), .C0(n1303), .Y(n2799)
         );
  OAI211XLTS U908 ( .A0(n3329), .A1(n902), .B0(n1207), .C0(n1208), .Y(n2844)
         );
  OAI211XLTS U909 ( .A0(n3329), .A1(n905), .B0(n1213), .C0(n1214), .Y(n2841)
         );
  OAI211XLTS U910 ( .A0(n3329), .A1(n904), .B0(n1211), .C0(n1212), .Y(n2842)
         );
  OAI211XLTS U911 ( .A0(n3333), .A1(n900), .B0(n1199), .C0(n1200), .Y(n2846)
         );
  OAI211XLTS U912 ( .A0(n3338), .A1(n839), .B0(n1970), .C0(n1971), .Y(n2475)
         );
  OAI211XLTS U913 ( .A0(n3338), .A1(n838), .B0(n1968), .C0(n1969), .Y(n2476)
         );
  OAI211XLTS U914 ( .A0(n3338), .A1(n837), .B0(n1966), .C0(n1967), .Y(n2477)
         );
  OAI211XLTS U915 ( .A0(n3338), .A1(n836), .B0(n1964), .C0(n1965), .Y(n2478)
         );
  OAI211XLTS U916 ( .A0(n1616), .A1(n640), .B0(n1619), .C0(n1620), .Y(n2641)
         );
  OAI211XLTS U917 ( .A0(n1616), .A1(n628), .B0(n1617), .C0(n1618), .Y(n2642)
         );
  OAI211XLTS U918 ( .A0(n4183), .A1(n3401), .B0(n1194), .C0(n1195), .Y(n2848)
         );
  OAI211XLTS U919 ( .A0(n4186), .A1(n3401), .B0(n1196), .C0(n1197), .Y(n2847)
         );
  OAI211XLTS U920 ( .A0(n4174), .A1(n3402), .B0(n1188), .C0(n1189), .Y(n2851)
         );
  OAI211XLTS U921 ( .A0(n4171), .A1(n3402), .B0(n1183), .C0(n1184), .Y(n2852)
         );
  OAI211XLTS U922 ( .A0(n4180), .A1(n3402), .B0(n1192), .C0(n1193), .Y(n2849)
         );
  OAI211XLTS U923 ( .A0(n4177), .A1(n3402), .B0(n1190), .C0(n1191), .Y(n2850)
         );
  OAI211XLTS U924 ( .A0(n4036), .A1(n3520), .B0(n1165), .C0(n1166), .Y(n2859)
         );
  OAI211XLTS U925 ( .A0(n4033), .A1(n3520), .B0(n1163), .C0(n1164), .Y(n2860)
         );
  OAI211XLTS U926 ( .A0(n4030), .A1(n3454), .B0(n1176), .C0(n1177), .Y(n2855)
         );
  OAI211XLTS U927 ( .A0(n4021), .A1(n3454), .B0(n1168), .C0(n1169), .Y(n2858)
         );
  OAI211XLTS U928 ( .A0(n4027), .A1(n3454), .B0(n1174), .C0(n1175), .Y(n2856)
         );
  OAI211XLTS U929 ( .A0(n4024), .A1(n3454), .B0(n1172), .C0(n1173), .Y(n2857)
         );
  OAI211XLTS U930 ( .A0(n4033), .A1(n3453), .B0(n1178), .C0(n1179), .Y(n2854)
         );
  OAI211XLTS U931 ( .A0(n4036), .A1(n3453), .B0(n1180), .C0(n1181), .Y(n2853)
         );
  OAI211XLTS U932 ( .A0(n4030), .A1(n3521), .B0(n1161), .C0(n1162), .Y(n2861)
         );
  OAI211XLTS U933 ( .A0(n4027), .A1(n3521), .B0(n1159), .C0(n1160), .Y(n2862)
         );
  OAI211XLTS U934 ( .A0(n4024), .A1(n3521), .B0(n1157), .C0(n1158), .Y(n2863)
         );
  OAI211XLTS U935 ( .A0(n4021), .A1(n3521), .B0(n1152), .C0(n1153), .Y(n2864)
         );
  OAI211XLTS U936 ( .A0(n3339), .A1(n849), .B0(n1972), .C0(n1973), .Y(n2474)
         );
  INVXLTS U937 ( .A(n3341), .Y(n3339) );
  OAI211XLTS U938 ( .A0(n4716), .A1(n3256), .B0(n1996), .C0(n1997), .Y(n2459)
         );
  INVXLTS U939 ( .A(n3257), .Y(n3256) );
  OAI211XLTS U940 ( .A0(n3748), .A1(n659), .B0(n1112), .C0(n1113), .Y(n2879)
         );
  OAI211XLTS U941 ( .A0(n3749), .A1(n658), .B0(n1108), .C0(n1109), .Y(n2881)
         );
  OAI211XLTS U942 ( .A0(n3748), .A1(n627), .B0(n1829), .C0(n1830), .Y(n2557)
         );
  OAI211XLTS U943 ( .A0(n3742), .A1(n937), .B0(n1707), .C0(n1708), .Y(n2597)
         );
  OAI211XLTS U944 ( .A0(n3742), .A1(n936), .B0(n1709), .C0(n1710), .Y(n2596)
         );
  OAI211XLTS U945 ( .A0(n3742), .A1(n935), .B0(n1711), .C0(n1712), .Y(n2595)
         );
  OAI211XLTS U946 ( .A0(n3753), .A1(n934), .B0(n1681), .C0(n1682), .Y(n2610)
         );
  OAI211XLTS U947 ( .A0(n3756), .A1(n663), .B0(n1116), .C0(n1117), .Y(n2877)
         );
  OAI211XLTS U948 ( .A0(n3753), .A1(n662), .B0(n1114), .C0(n1115), .Y(n2878)
         );
  OAI211XLTS U949 ( .A0(n3753), .A1(n661), .B0(n1110), .C0(n1111), .Y(n2880)
         );
  OAI211XLTS U950 ( .A0(n3743), .A1(n657), .B0(n1101), .C0(n1102), .Y(n2882)
         );
  OAI211XLTS U951 ( .A0(n3746), .A1(n623), .B0(n1743), .C0(n1744), .Y(n2579)
         );
  OAI211XLTS U952 ( .A0(n3746), .A1(n622), .B0(n1741), .C0(n1742), .Y(n2580)
         );
  OAI211XLTS U953 ( .A0(n3746), .A1(n621), .B0(n1739), .C0(n1740), .Y(n2581)
         );
  OAI211XLTS U954 ( .A0(n3746), .A1(n620), .B0(n1737), .C0(n1738), .Y(n2582)
         );
  OAI211XLTS U955 ( .A0(n3745), .A1(n619), .B0(n1735), .C0(n1736), .Y(n2583)
         );
  OAI211XLTS U956 ( .A0(n3745), .A1(n618), .B0(n1733), .C0(n1734), .Y(n2584)
         );
  OAI211XLTS U957 ( .A0(n3745), .A1(n617), .B0(n1731), .C0(n1732), .Y(n2585)
         );
  OAI211XLTS U958 ( .A0(n3745), .A1(n616), .B0(n1729), .C0(n1730), .Y(n2586)
         );
  OAI211XLTS U959 ( .A0(n3744), .A1(n615), .B0(n1727), .C0(n1728), .Y(n2587)
         );
  OAI211XLTS U960 ( .A0(n3744), .A1(n614), .B0(n1725), .C0(n1726), .Y(n2588)
         );
  OAI211XLTS U961 ( .A0(n3744), .A1(n613), .B0(n1723), .C0(n1724), .Y(n2589)
         );
  OAI211XLTS U962 ( .A0(n3744), .A1(n612), .B0(n1721), .C0(n1722), .Y(n2590)
         );
  OAI211XLTS U963 ( .A0(n3743), .A1(n611), .B0(n1719), .C0(n1720), .Y(n2591)
         );
  OAI211XLTS U964 ( .A0(n3743), .A1(n610), .B0(n1717), .C0(n1718), .Y(n2592)
         );
  OAI211XLTS U965 ( .A0(n3743), .A1(n609), .B0(n1715), .C0(n1716), .Y(n2593)
         );
  OAI211XLTS U966 ( .A0(n3742), .A1(n608), .B0(n1713), .C0(n1714), .Y(n2594)
         );
  OAI211XLTS U967 ( .A0(n3741), .A1(n607), .B0(n1705), .C0(n1706), .Y(n2598)
         );
  OAI211XLTS U968 ( .A0(n3741), .A1(n606), .B0(n1703), .C0(n1704), .Y(n2599)
         );
  OAI211XLTS U969 ( .A0(n3741), .A1(n605), .B0(n1701), .C0(n1702), .Y(n2600)
         );
  OAI211XLTS U970 ( .A0(n3741), .A1(n604), .B0(n1699), .C0(n1700), .Y(n2601)
         );
  OAI211XLTS U971 ( .A0(n3753), .A1(n603), .B0(n1697), .C0(n1698), .Y(n2602)
         );
  OAI211XLTS U972 ( .A0(n3749), .A1(n602), .B0(n1695), .C0(n1696), .Y(n2603)
         );
  OAI211XLTS U973 ( .A0(n3757), .A1(n601), .B0(n1693), .C0(n1694), .Y(n2604)
         );
  OAI211XLTS U974 ( .A0(n3757), .A1(n600), .B0(n1691), .C0(n1692), .Y(n2605)
         );
  OAI211XLTS U975 ( .A0(n3750), .A1(n599), .B0(n1689), .C0(n1690), .Y(n2606)
         );
  OAI211XLTS U976 ( .A0(n3751), .A1(n598), .B0(n1687), .C0(n1688), .Y(n2607)
         );
  OAI211XLTS U977 ( .A0(n3752), .A1(n597), .B0(n1685), .C0(n1686), .Y(n2608)
         );
  OAI211XLTS U978 ( .A0(n3750), .A1(n596), .B0(n1683), .C0(n1684), .Y(n2609)
         );
  OAI211XLTS U979 ( .A0(n3747), .A1(n638), .B0(n1819), .C0(n1820), .Y(n2562)
         );
  OAI211XLTS U980 ( .A0(n3747), .A1(n626), .B0(n1825), .C0(n1826), .Y(n2559)
         );
  OAI211XLTS U981 ( .A0(n3747), .A1(n625), .B0(n1823), .C0(n1824), .Y(n2560)
         );
  OAI211XLTS U982 ( .A0(n3747), .A1(n624), .B0(n1821), .C0(n1822), .Y(n2561)
         );
  OAI211XLTS U983 ( .A0(n3748), .A1(n639), .B0(n1827), .C0(n1828), .Y(n2558)
         );
  OAI211XLTS U984 ( .A0(n4424), .A1(n3254), .B0(n1294), .C0(n1295), .Y(n2803)
         );
  OAI211XLTS U985 ( .A0(n4437), .A1(n3254), .B0(n1292), .C0(n1293), .Y(n2804)
         );
  OAI211XLTS U986 ( .A0(n4448), .A1(n3254), .B0(n1290), .C0(n1291), .Y(n2805)
         );
  OAI211XLTS U987 ( .A0(n4473), .A1(n3253), .B0(n1284), .C0(n1285), .Y(n2808)
         );
  OAI211XLTS U988 ( .A0(n4480), .A1(n3253), .B0(n1282), .C0(n1283), .Y(n2809)
         );
  OAI211XLTS U989 ( .A0(n4489), .A1(n3253), .B0(n1280), .C0(n1281), .Y(n2810)
         );
  OAI211XLTS U990 ( .A0(n4505), .A1(n3255), .B0(n1276), .C0(n1277), .Y(n2812)
         );
  OAI211XLTS U991 ( .A0(n4520), .A1(n3253), .B0(n1274), .C0(n1275), .Y(n2813)
         );
  OAI211XLTS U992 ( .A0(n4534), .A1(n3252), .B0(n1270), .C0(n1271), .Y(n2815)
         );
  OAI211XLTS U993 ( .A0(n4543), .A1(n3252), .B0(n1268), .C0(n1269), .Y(n2816)
         );
  OAI211XLTS U994 ( .A0(n4552), .A1(n3251), .B0(n1266), .C0(n1267), .Y(n2817)
         );
  OAI211XLTS U995 ( .A0(n4561), .A1(n3252), .B0(n1264), .C0(n1265), .Y(n2818)
         );
  OAI211XLTS U996 ( .A0(n4572), .A1(n3251), .B0(n1262), .C0(n1263), .Y(n2819)
         );
  OAI211XLTS U997 ( .A0(n4579), .A1(n3254), .B0(n1260), .C0(n1261), .Y(n2820)
         );
  OAI211XLTS U998 ( .A0(n4592), .A1(n3252), .B0(n1258), .C0(n1259), .Y(n2821)
         );
  OAI211XLTS U999 ( .A0(n4736), .A1(n3255), .B0(n1992), .C0(n1993), .Y(n2461)
         );
  OAI211XLTS U1000 ( .A0(n4747), .A1(n3255), .B0(n1990), .C0(n1991), .Y(n2462)
         );
  OAI211XLTS U1001 ( .A0(n4752), .A1(n3255), .B0(n1988), .C0(n1989), .Y(n2463)
         );
  AOI22XLTS U1002 ( .A0(n1770), .A1(n1771), .B0(n3113), .B1(n650), .Y(n2569)
         );
  AOI2BB2XLTS U1003 ( .B0(n1763), .B1(n1764), .A0N(n3754), .A1N(
        readOutbuffer_7), .Y(n2570) );
  NAND4XLTS U1004 ( .A(n436), .B(n441), .C(n731), .D(n437), .Y(n2024) );
  NAND4XLTS U1005 ( .A(n470), .B(n455), .C(n1083), .D(n731), .Y(n2026) );
  NAND4XLTS U1006 ( .A(n446), .B(n455), .C(n731), .D(n1028), .Y(n2027) );
  NAND3XLTS U1007 ( .A(n455), .B(n441), .C(n472), .Y(n2025) );
  NAND4XLTS U1008 ( .A(selectBit_NORTH), .B(n441), .C(n731), .D(n971), .Y(
        n2023) );
  NAND2X1TS U1009 ( .A(n1), .B(n143), .Y(n1832) );
  CLKBUFX2TS U1010 ( .A(n5327), .Y(n925) );
  NAND2X1TS U1011 ( .A(n1), .B(n151), .Y(n1884) );
  XNOR2X1TS U1012 ( .A(n2899), .B(n2908), .Y(n1094) );
  NAND3X1TS U1013 ( .A(n45), .B(n2), .C(n6), .Y(n2034) );
  NAND3X1TS U1014 ( .A(n8), .B(n913), .C(n100), .Y(n2036) );
  NAND3X1TS U1015 ( .A(n120), .B(n136), .C(n6), .Y(n2033) );
  NAND3X1TS U1016 ( .A(n115), .B(n120), .C(n45), .Y(n2035) );
  NAND3X1TS U1017 ( .A(n100), .B(n8), .C(n6), .Y(n2049) );
  CLKBUFX2TS U1018 ( .A(n3891), .Y(n3882) );
  CLKBUFX2TS U1019 ( .A(n3810), .Y(n3799) );
  CLKBUFX2TS U1020 ( .A(n3889), .Y(n3886) );
  CLKBUFX2TS U1021 ( .A(n3890), .Y(n3885) );
  CLKBUFX2TS U1022 ( .A(n728), .Y(n3888) );
  CLKBUFX2TS U1023 ( .A(n3889), .Y(n3887) );
  CLKBUFX2TS U1024 ( .A(n3890), .Y(n3884) );
  CLKBUFX2TS U1025 ( .A(n3891), .Y(n3883) );
  CLKBUFX2TS U1026 ( .A(n3810), .Y(n3800) );
  CLKBUFX2TS U1027 ( .A(n3809), .Y(n3801) );
  CLKBUFX2TS U1028 ( .A(n3808), .Y(n3803) );
  CLKBUFX2TS U1029 ( .A(n3809), .Y(n3802) );
  CLKBUFX2TS U1030 ( .A(n3794), .Y(n3789) );
  CLKBUFX2TS U1031 ( .A(n3794), .Y(n3790) );
  CLKBUFX2TS U1032 ( .A(n3796), .Y(n3791) );
  CLKBUFX2TS U1033 ( .A(n3794), .Y(n3792) );
  CLKBUFX2TS U1034 ( .A(n3795), .Y(n3788) );
  CLKBUFX2TS U1035 ( .A(n3795), .Y(n3787) );
  CLKBUFX2TS U1036 ( .A(n3867), .Y(n3855) );
  CLKBUFX2TS U1037 ( .A(n3867), .Y(n3856) );
  CLKBUFX2TS U1038 ( .A(n3864), .Y(n3857) );
  CLKBUFX2TS U1039 ( .A(n3864), .Y(n3858) );
  CLKBUFX2TS U1040 ( .A(n3863), .Y(n3860) );
  CLKBUFX2TS U1041 ( .A(n3863), .Y(n3859) );
  CLKBUFX2TS U1042 ( .A(n3808), .Y(n3804) );
  CLKBUFX2TS U1043 ( .A(n3807), .Y(n3805) );
  CLKBUFX2TS U1044 ( .A(n3931), .Y(n3928) );
  CLKBUFX2TS U1045 ( .A(n3930), .Y(n3927) );
  CLKBUFX2TS U1046 ( .A(n3931), .Y(n3926) );
  CLKBUFX2TS U1047 ( .A(n3932), .Y(n3925) );
  CLKBUFX2TS U1048 ( .A(n3932), .Y(n3924) );
  CLKBUFX2TS U1049 ( .A(n3930), .Y(n3929) );
  CLKBUFX2TS U1050 ( .A(n3807), .Y(n3806) );
  CLKBUFX2TS U1051 ( .A(n3867), .Y(n3865) );
  CLKBUFX2TS U1052 ( .A(n732), .Y(n3862) );
  CLKBUFX2TS U1053 ( .A(n732), .Y(n3864) );
  CLKBUFX2TS U1054 ( .A(n732), .Y(n3863) );
  CLKBUFX2TS U1055 ( .A(n722), .Y(n3930) );
  CLKBUFX2TS U1056 ( .A(n3934), .Y(n3932) );
  CLKBUFX2TS U1057 ( .A(n1750), .Y(n3931) );
  CLKBUFX2TS U1058 ( .A(n3934), .Y(n3933) );
  CLKBUFX2TS U1059 ( .A(n3797), .Y(n3794) );
  CLKBUFX2TS U1060 ( .A(n728), .Y(n3889) );
  CLKBUFX2TS U1061 ( .A(n3893), .Y(n3890) );
  CLKBUFX2TS U1062 ( .A(n3893), .Y(n3891) );
  CLKBUFX2TS U1063 ( .A(n3811), .Y(n3810) );
  CLKBUFX2TS U1064 ( .A(n1746), .Y(n3808) );
  CLKBUFX2TS U1065 ( .A(n740), .Y(n3807) );
  CLKBUFX2TS U1066 ( .A(n3797), .Y(n3795) );
  CLKBUFX2TS U1067 ( .A(n740), .Y(n3809) );
  CLKBUFX2TS U1068 ( .A(n3441), .Y(n3427) );
  CLKBUFX2TS U1069 ( .A(n3438), .Y(n3434) );
  CLKBUFX2TS U1070 ( .A(n3438), .Y(n3433) );
  CLKBUFX2TS U1071 ( .A(n3437), .Y(n3435) );
  CLKBUFX2TS U1072 ( .A(n3439), .Y(n3432) );
  CLKBUFX2TS U1073 ( .A(n3439), .Y(n3431) );
  CLKBUFX2TS U1074 ( .A(n3442), .Y(n3430) );
  CLKBUFX2TS U1075 ( .A(n3440), .Y(n3428) );
  CLKBUFX2TS U1076 ( .A(n3440), .Y(n3429) );
  CLKBUFX2TS U1077 ( .A(n3358), .Y(n3344) );
  CLKBUFX2TS U1078 ( .A(n3892), .Y(n3881) );
  CLKBUFX2TS U1079 ( .A(n3893), .Y(n3892) );
  CLKBUFX2TS U1080 ( .A(n3878), .Y(n3869) );
  CLKBUFX2TS U1081 ( .A(n3358), .Y(n3345) );
  CLKBUFX2TS U1082 ( .A(n730), .Y(n3875) );
  CLKBUFX2TS U1083 ( .A(n3876), .Y(n3874) );
  CLKBUFX2TS U1084 ( .A(n3877), .Y(n3873) );
  CLKBUFX2TS U1085 ( .A(n3877), .Y(n3872) );
  CLKBUFX2TS U1086 ( .A(n3878), .Y(n3871) );
  CLKBUFX2TS U1087 ( .A(n3878), .Y(n3870) );
  CLKBUFX2TS U1088 ( .A(n3917), .Y(n3915) );
  CLKBUFX2TS U1089 ( .A(n3918), .Y(n3914) );
  CLKBUFX2TS U1090 ( .A(n3918), .Y(n3913) );
  CLKBUFX2TS U1091 ( .A(n3919), .Y(n3912) );
  CLKBUFX2TS U1092 ( .A(n3919), .Y(n3911) );
  CLKBUFX2TS U1093 ( .A(n3919), .Y(n3910) );
  CLKBUFX2TS U1094 ( .A(n3917), .Y(n3916) );
  CLKBUFX2TS U1095 ( .A(n3356), .Y(n3348) );
  CLKBUFX2TS U1096 ( .A(n3355), .Y(n3350) );
  CLKBUFX2TS U1097 ( .A(n3354), .Y(n3352) );
  CLKBUFX2TS U1098 ( .A(n3354), .Y(n3353) );
  CLKBUFX2TS U1099 ( .A(n3355), .Y(n3351) );
  CLKBUFX2TS U1100 ( .A(n3356), .Y(n3349) );
  CLKBUFX2TS U1101 ( .A(n3357), .Y(n3347) );
  CLKBUFX2TS U1102 ( .A(n3357), .Y(n3346) );
  CLKBUFX2TS U1103 ( .A(n3507), .Y(n3492) );
  CLKBUFX2TS U1104 ( .A(n3507), .Y(n3493) );
  CLKBUFX2TS U1105 ( .A(n3239), .Y(n3226) );
  CLKBUFX2TS U1106 ( .A(n3239), .Y(n3227) );
  CLKBUFX2TS U1107 ( .A(n3237), .Y(n3231) );
  CLKBUFX2TS U1108 ( .A(n3237), .Y(n3230) );
  CLKBUFX2TS U1109 ( .A(n3238), .Y(n3229) );
  CLKBUFX2TS U1110 ( .A(n3236), .Y(n3233) );
  CLKBUFX2TS U1111 ( .A(n3236), .Y(n3232) );
  CLKBUFX2TS U1112 ( .A(n3238), .Y(n3228) );
  CLKBUFX2TS U1113 ( .A(n3796), .Y(n3786) );
  CLKBUFX2TS U1114 ( .A(n3797), .Y(n3796) );
  CLKBUFX2TS U1115 ( .A(n3506), .Y(n3494) );
  CLKBUFX2TS U1116 ( .A(n3388), .Y(n3375) );
  CLKBUFX2TS U1117 ( .A(n3509), .Y(n3501) );
  CLKBUFX2TS U1118 ( .A(n3509), .Y(n3500) );
  CLKBUFX2TS U1119 ( .A(n3509), .Y(n3499) );
  CLKBUFX2TS U1120 ( .A(n3509), .Y(n3498) );
  CLKBUFX2TS U1121 ( .A(n3506), .Y(n3495) );
  CLKBUFX2TS U1122 ( .A(n3224), .Y(n3211) );
  CLKBUFX2TS U1123 ( .A(n3224), .Y(n3209) );
  CLKBUFX2TS U1124 ( .A(n3222), .Y(n3215) );
  CLKBUFX2TS U1125 ( .A(n3221), .Y(n3216) );
  CLKBUFX2TS U1126 ( .A(n3387), .Y(n3377) );
  CLKBUFX2TS U1127 ( .A(n3224), .Y(n3210) );
  CLKBUFX2TS U1128 ( .A(n3385), .Y(n3381) );
  CLKBUFX2TS U1129 ( .A(n3387), .Y(n3376) );
  CLKBUFX2TS U1130 ( .A(n3223), .Y(n3212) );
  CLKBUFX2TS U1131 ( .A(n3223), .Y(n3213) );
  CLKBUFX2TS U1132 ( .A(n3222), .Y(n3214) );
  CLKBUFX2TS U1133 ( .A(n3221), .Y(n3217) );
  CLKBUFX2TS U1134 ( .A(n3220), .Y(n3218) );
  CLKBUFX2TS U1135 ( .A(n3384), .Y(n3382) );
  CLKBUFX2TS U1136 ( .A(n3385), .Y(n3380) );
  CLKBUFX2TS U1137 ( .A(n3386), .Y(n3378) );
  CLKBUFX2TS U1138 ( .A(n3386), .Y(n3379) );
  CLKBUFX2TS U1139 ( .A(n3510), .Y(n3502) );
  CLKBUFX2TS U1140 ( .A(n3220), .Y(n3219) );
  CLKBUFX2TS U1141 ( .A(n3384), .Y(n3383) );
  CLKBUFX2TS U1142 ( .A(n3837), .Y(n3828) );
  CLKBUFX2TS U1143 ( .A(n3867), .Y(n3866) );
  CLKBUFX2TS U1144 ( .A(n3835), .Y(n3833) );
  CLKBUFX2TS U1145 ( .A(n3836), .Y(n3831) );
  CLKBUFX2TS U1148 ( .A(n3835), .Y(n3832) );
  CLKBUFX2TS U1149 ( .A(n3836), .Y(n3830) );
  CLKBUFX2TS U1150 ( .A(n3837), .Y(n3829) );
  CLKBUFX2TS U1151 ( .A(n3933), .Y(n3922) );
  INVX2TS U1152 ( .A(n4539), .Y(n4541) );
  CLKBUFX2TS U1153 ( .A(n3783), .Y(n3772) );
  CLKBUFX2TS U1154 ( .A(n3779), .Y(n3778) );
  CLKBUFX2TS U1155 ( .A(n3781), .Y(n3773) );
  CLKBUFX2TS U1156 ( .A(n3780), .Y(n3775) );
  CLKBUFX2TS U1157 ( .A(n3781), .Y(n3774) );
  CLKBUFX2TS U1158 ( .A(n3779), .Y(n3777) );
  CLKBUFX2TS U1159 ( .A(n3780), .Y(n3776) );
  CLKBUFX2TS U1160 ( .A(n1048), .Y(n1036) );
  CLKBUFX2TS U1161 ( .A(n2117), .Y(n1037) );
  CLKBUFX2TS U1162 ( .A(n1047), .Y(n1038) );
  CLKBUFX2TS U1163 ( .A(n1047), .Y(n1039) );
  CLKBUFX2TS U1164 ( .A(n1049), .Y(n1040) );
  CLKBUFX2TS U1165 ( .A(n1046), .Y(n1041) );
  CLKBUFX2TS U1166 ( .A(n1045), .Y(n1044) );
  CLKBUFX2TS U1167 ( .A(n1046), .Y(n1042) );
  CLKBUFX2TS U1168 ( .A(n1045), .Y(n1043) );
  INVX2TS U1169 ( .A(n4539), .Y(n4542) );
  CLKBUFX2TS U1170 ( .A(n3460), .Y(n3455) );
  CLKBUFX2TS U1171 ( .A(n3460), .Y(n3456) );
  CLKBUFX2TS U1172 ( .A(n3460), .Y(n3457) );
  CLKBUFX2TS U1173 ( .A(n3408), .Y(n3404) );
  CLKBUFX2TS U1174 ( .A(n3408), .Y(n3403) );
  CLKBUFX2TS U1175 ( .A(n3360), .Y(n3354) );
  CLKBUFX2TS U1176 ( .A(n3360), .Y(n3355) );
  CLKBUFX2TS U1177 ( .A(n3359), .Y(n3356) );
  CLKBUFX2TS U1178 ( .A(n3359), .Y(n3357) );
  CLKBUFX2TS U1179 ( .A(n3359), .Y(n3358) );
  CLKBUFX2TS U1180 ( .A(n3508), .Y(n3505) );
  CLKBUFX2TS U1181 ( .A(n3508), .Y(n3506) );
  CLKBUFX2TS U1182 ( .A(n1219), .Y(n3224) );
  CLKBUFX2TS U1183 ( .A(n3443), .Y(n3438) );
  CLKBUFX2TS U1184 ( .A(n3442), .Y(n3441) );
  CLKBUFX2TS U1185 ( .A(n3443), .Y(n3439) );
  CLKBUFX2TS U1186 ( .A(n3442), .Y(n3440) );
  CLKBUFX2TS U1187 ( .A(n3880), .Y(n3876) );
  CLKBUFX2TS U1188 ( .A(n730), .Y(n3877) );
  CLKBUFX2TS U1189 ( .A(n3880), .Y(n3878) );
  CLKBUFX2TS U1190 ( .A(n3921), .Y(n3918) );
  CLKBUFX2TS U1191 ( .A(n3921), .Y(n3919) );
  CLKBUFX2TS U1192 ( .A(n3921), .Y(n3917) );
  CLKBUFX2TS U1193 ( .A(n3390), .Y(n3389) );
  CLKBUFX2TS U1194 ( .A(n3390), .Y(n3387) );
  CLKBUFX2TS U1195 ( .A(n1219), .Y(n3223) );
  CLKBUFX2TS U1196 ( .A(n3225), .Y(n3222) );
  CLKBUFX2TS U1197 ( .A(n3225), .Y(n3221) );
  CLKBUFX2TS U1198 ( .A(n3840), .Y(n3834) );
  CLKBUFX2TS U1199 ( .A(n3391), .Y(n3385) );
  CLKBUFX2TS U1200 ( .A(n3840), .Y(n3835) );
  CLKBUFX2TS U1201 ( .A(n3391), .Y(n3386) );
  CLKBUFX2TS U1202 ( .A(n3839), .Y(n3836) );
  CLKBUFX2TS U1203 ( .A(n3390), .Y(n3388) );
  CLKBUFX2TS U1204 ( .A(n3225), .Y(n3220) );
  CLKBUFX2TS U1205 ( .A(n3391), .Y(n3384) );
  CLKBUFX2TS U1206 ( .A(n3839), .Y(n3837) );
  CLKBUFX2TS U1207 ( .A(n3443), .Y(n3437) );
  CLKBUFX2TS U1208 ( .A(n3240), .Y(n3237) );
  CLKBUFX2TS U1209 ( .A(n3241), .Y(n3236) );
  CLKBUFX2TS U1210 ( .A(n3240), .Y(n3238) );
  CLKBUFX2TS U1211 ( .A(n3240), .Y(n3239) );
  CLKBUFX2TS U1212 ( .A(n728), .Y(n3893) );
  CLKBUFX2TS U1213 ( .A(n732), .Y(n3867) );
  CLKBUFX2TS U1214 ( .A(n722), .Y(n3934) );
  CLKBUFX2TS U1215 ( .A(n740), .Y(n3811) );
  CLKBUFX2TS U1216 ( .A(n741), .Y(n3797) );
  CLKBUFX2TS U1217 ( .A(n3275), .Y(n3261) );
  CLKBUFX2TS U1218 ( .A(n3542), .Y(n3528) );
  CLKBUFX2TS U1219 ( .A(n3152), .Y(n3116) );
  CLKBUFX2TS U1220 ( .A(n3275), .Y(n3262) );
  CLKBUFX2TS U1221 ( .A(n3542), .Y(n3529) );
  CLKBUFX2TS U1222 ( .A(n3152), .Y(n3117) );
  CLKBUFX2TS U1223 ( .A(n3654), .Y(n3645) );
  CLKBUFX2TS U1224 ( .A(n3653), .Y(n3646) );
  CLKBUFX2TS U1225 ( .A(n3653), .Y(n3647) );
  CLKBUFX2TS U1226 ( .A(n3658), .Y(n3648) );
  CLKBUFX2TS U1227 ( .A(n3271), .Y(n3269) );
  CLKBUFX2TS U1228 ( .A(n3272), .Y(n3268) );
  CLKBUFX2TS U1229 ( .A(n3273), .Y(n3266) );
  CLKBUFX2TS U1230 ( .A(n3273), .Y(n3265) );
  CLKBUFX2TS U1231 ( .A(n3272), .Y(n3267) );
  CLKBUFX2TS U1232 ( .A(n3274), .Y(n3264) );
  CLKBUFX2TS U1233 ( .A(n3274), .Y(n3263) );
  CLKBUFX2TS U1234 ( .A(n3538), .Y(n3537) );
  CLKBUFX2TS U1235 ( .A(n3538), .Y(n3536) );
  CLKBUFX2TS U1236 ( .A(n3539), .Y(n3535) );
  CLKBUFX2TS U1237 ( .A(n3540), .Y(n3533) );
  CLKBUFX2TS U1238 ( .A(n3540), .Y(n3532) );
  CLKBUFX2TS U1239 ( .A(n3539), .Y(n3534) );
  CLKBUFX2TS U1240 ( .A(n3541), .Y(n3531) );
  CLKBUFX2TS U1241 ( .A(n3541), .Y(n3530) );
  CLKBUFX2TS U1242 ( .A(n3127), .Y(n3121) );
  CLKBUFX2TS U1243 ( .A(n3127), .Y(n3120) );
  CLKBUFX2TS U1244 ( .A(n3128), .Y(n3119) );
  CLKBUFX2TS U1245 ( .A(n3128), .Y(n3118) );
  CLKBUFX2TS U1246 ( .A(n3691), .Y(n3676) );
  CLKBUFX2TS U1247 ( .A(n3651), .Y(n3649) );
  CLKBUFX2TS U1248 ( .A(n3654), .Y(n3644) );
  CLKBUFX2TS U1249 ( .A(n3655), .Y(n3642) );
  CLKBUFX2TS U1250 ( .A(n3688), .Y(n3686) );
  CLKBUFX2TS U1251 ( .A(n3691), .Y(n3685) );
  CLKBUFX2TS U1252 ( .A(n3692), .Y(n3684) );
  CLKBUFX2TS U1253 ( .A(n3689), .Y(n3683) );
  CLKBUFX2TS U1254 ( .A(n3689), .Y(n3682) );
  CLKBUFX2TS U1255 ( .A(n1106), .Y(n3681) );
  CLKBUFX2TS U1256 ( .A(n3691), .Y(n3680) );
  CLKBUFX2TS U1257 ( .A(n3690), .Y(n3679) );
  CLKBUFX2TS U1258 ( .A(n3690), .Y(n3678) );
  CLKBUFX2TS U1259 ( .A(n3691), .Y(n3677) );
  CLKBUFX2TS U1260 ( .A(n3655), .Y(n3643) );
  CLKBUFX2TS U1261 ( .A(n3475), .Y(n3461) );
  CLKBUFX2TS U1262 ( .A(n3424), .Y(n3410) );
  CLKBUFX2TS U1263 ( .A(n3625), .Y(n3611) );
  CLKBUFX2TS U1264 ( .A(n3879), .Y(n3868) );
  CLKBUFX2TS U1265 ( .A(n3880), .Y(n3879) );
  CLKBUFX2TS U1266 ( .A(n3920), .Y(n3909) );
  CLKBUFX2TS U1267 ( .A(n724), .Y(n3920) );
  CLKBUFX2TS U1268 ( .A(n3424), .Y(n3411) );
  CLKBUFX2TS U1269 ( .A(n3475), .Y(n3462) );
  CLKBUFX2TS U1270 ( .A(n3625), .Y(n3612) );
  CLKBUFX2TS U1271 ( .A(n3624), .Y(n3613) );
  CLKBUFX2TS U1272 ( .A(n3471), .Y(n3467) );
  CLKBUFX2TS U1273 ( .A(n3420), .Y(n3418) );
  CLKBUFX2TS U1274 ( .A(n3421), .Y(n3417) );
  CLKBUFX2TS U1275 ( .A(n3421), .Y(n3416) );
  CLKBUFX2TS U1276 ( .A(n3422), .Y(n3415) );
  CLKBUFX2TS U1277 ( .A(n3422), .Y(n3414) );
  CLKBUFX2TS U1278 ( .A(n3423), .Y(n3412) );
  CLKBUFX2TS U1279 ( .A(n3423), .Y(n3413) );
  CLKBUFX2TS U1280 ( .A(n3474), .Y(n3464) );
  CLKBUFX2TS U1281 ( .A(n3473), .Y(n3466) );
  CLKBUFX2TS U1282 ( .A(n3473), .Y(n3465) );
  CLKBUFX2TS U1283 ( .A(n3474), .Y(n3463) );
  CLKBUFX2TS U1284 ( .A(n3470), .Y(n3468) );
  CLKBUFX2TS U1285 ( .A(n3508), .Y(n3507) );
  INVX2TS U1286 ( .A(n3670), .Y(n3669) );
  INVX2TS U1287 ( .A(n3672), .Y(n3667) );
  INVX2TS U1288 ( .A(n3671), .Y(n3668) );
  CLKBUFX2TS U1289 ( .A(n3907), .Y(n3894) );
  CLKBUFX2TS U1290 ( .A(n3324), .Y(n3309) );
  CLKBUFX2TS U1291 ( .A(n3592), .Y(n3576) );
  CLKBUFX2TS U1292 ( .A(n3324), .Y(n3310) );
  CLKBUFX2TS U1293 ( .A(n3592), .Y(n3577) );
  CLKBUFX2TS U1294 ( .A(n3271), .Y(n3270) );
  CLKBUFX2TS U1295 ( .A(n3903), .Y(n3901) );
  CLKBUFX2TS U1296 ( .A(n3321), .Y(n3317) );
  CLKBUFX2TS U1297 ( .A(n3320), .Y(n3316) );
  CLKBUFX2TS U1298 ( .A(n3320), .Y(n3315) );
  CLKBUFX2TS U1299 ( .A(n3322), .Y(n3314) );
  CLKBUFX2TS U1300 ( .A(n3322), .Y(n3313) );
  CLKBUFX2TS U1301 ( .A(n3323), .Y(n3312) );
  CLKBUFX2TS U1302 ( .A(n3323), .Y(n3311) );
  CLKBUFX2TS U1303 ( .A(n3904), .Y(n3902) );
  CLKBUFX2TS U1304 ( .A(n3904), .Y(n3900) );
  CLKBUFX2TS U1305 ( .A(n3905), .Y(n3898) );
  CLKBUFX2TS U1306 ( .A(n3906), .Y(n3897) );
  CLKBUFX2TS U1307 ( .A(n3907), .Y(n3895) );
  CLKBUFX2TS U1308 ( .A(n3905), .Y(n3899) );
  CLKBUFX2TS U1309 ( .A(n3906), .Y(n3896) );
  CLKBUFX2TS U1310 ( .A(n3588), .Y(n3583) );
  CLKBUFX2TS U1311 ( .A(n3588), .Y(n3582) );
  CLKBUFX2TS U1312 ( .A(n3590), .Y(n3581) );
  CLKBUFX2TS U1313 ( .A(n3590), .Y(n3580) );
  CLKBUFX2TS U1314 ( .A(n3591), .Y(n3579) );
  CLKBUFX2TS U1315 ( .A(n3591), .Y(n3578) );
  CLKBUFX2TS U1316 ( .A(n3587), .Y(n3584) );
  CLKBUFX2TS U1317 ( .A(n3821), .Y(n3819) );
  CLKBUFX2TS U1318 ( .A(n3824), .Y(n3813) );
  CLKBUFX2TS U1319 ( .A(n3822), .Y(n3818) );
  CLKBUFX2TS U1320 ( .A(n3822), .Y(n3817) );
  CLKBUFX2TS U1321 ( .A(n3823), .Y(n3816) );
  CLKBUFX2TS U1322 ( .A(n3823), .Y(n3815) );
  CLKBUFX2TS U1323 ( .A(n3738), .Y(n3724) );
  CLKBUFX2TS U1324 ( .A(n3824), .Y(n3814) );
  CLKBUFX2TS U1325 ( .A(n3825), .Y(n3812) );
  CLKBUFX2TS U1326 ( .A(n3733), .Y(n3730) );
  CLKBUFX2TS U1327 ( .A(n3734), .Y(n3729) );
  CLKBUFX2TS U1328 ( .A(n3734), .Y(n3728) );
  CLKBUFX2TS U1329 ( .A(n3735), .Y(n3727) );
  CLKBUFX2TS U1330 ( .A(n3735), .Y(n3726) );
  CLKBUFX2TS U1331 ( .A(n3738), .Y(n3725) );
  CLKBUFX2TS U1332 ( .A(n3688), .Y(n3687) );
  CLKBUFX2TS U1333 ( .A(n3623), .Y(n3615) );
  CLKBUFX2TS U1334 ( .A(n3293), .Y(n3278) );
  CLKBUFX2TS U1335 ( .A(n3293), .Y(n3279) );
  CLKBUFX2TS U1336 ( .A(n3558), .Y(n3545) );
  CLKBUFX2TS U1337 ( .A(n3558), .Y(n3546) );
  CLKBUFX2TS U1338 ( .A(n3707), .Y(n3693) );
  CLKBUFX2TS U1339 ( .A(n3707), .Y(n3694) );
  CLKBUFX2TS U1340 ( .A(n3292), .Y(n3280) );
  CLKBUFX2TS U1341 ( .A(n3557), .Y(n3547) );
  CLKBUFX2TS U1342 ( .A(n3557), .Y(n3548) );
  CLKBUFX2TS U1343 ( .A(n3292), .Y(n3281) );
  CLKBUFX2TS U1344 ( .A(n3623), .Y(n3616) );
  CLKBUFX2TS U1345 ( .A(n3706), .Y(n3695) );
  CLKBUFX2TS U1346 ( .A(n3620), .Y(n3618) );
  CLKBUFX2TS U1347 ( .A(n3555), .Y(n3551) );
  CLKBUFX2TS U1348 ( .A(n3555), .Y(n3552) );
  CLKBUFX2TS U1349 ( .A(n3556), .Y(n3550) );
  CLKBUFX2TS U1350 ( .A(n3556), .Y(n3549) );
  CLKBUFX2TS U1351 ( .A(n1201), .Y(n3318) );
  CLKBUFX2TS U1352 ( .A(n3622), .Y(n3617) );
  CLKBUFX2TS U1353 ( .A(n3587), .Y(n3585) );
  CLKBUFX2TS U1354 ( .A(n3851), .Y(n3847) );
  CLKBUFX2TS U1355 ( .A(n3853), .Y(n3841) );
  CLKBUFX2TS U1356 ( .A(n3850), .Y(n3848) );
  CLKBUFX2TS U1357 ( .A(n3851), .Y(n3846) );
  CLKBUFX2TS U1358 ( .A(n3852), .Y(n3845) );
  CLKBUFX2TS U1359 ( .A(n3852), .Y(n3844) );
  CLKBUFX2TS U1360 ( .A(n3850), .Y(n3842) );
  CLKBUFX2TS U1361 ( .A(n3854), .Y(n3843) );
  CLKBUFX2TS U1362 ( .A(n3288), .Y(n3287) );
  CLKBUFX2TS U1363 ( .A(n3288), .Y(n3286) );
  CLKBUFX2TS U1364 ( .A(n3289), .Y(n3285) );
  CLKBUFX2TS U1365 ( .A(n3289), .Y(n3284) );
  CLKBUFX2TS U1366 ( .A(n3290), .Y(n3282) );
  CLKBUFX2TS U1367 ( .A(n3290), .Y(n3283) );
  CLKBUFX2TS U1368 ( .A(n3706), .Y(n3696) );
  CLKBUFX2TS U1369 ( .A(n3704), .Y(n3700) );
  CLKBUFX2TS U1370 ( .A(n3703), .Y(n3702) );
  CLKBUFX2TS U1371 ( .A(n3703), .Y(n3701) );
  CLKBUFX2TS U1372 ( .A(n3704), .Y(n3699) );
  CLKBUFX2TS U1373 ( .A(n3705), .Y(n3698) );
  CLKBUFX2TS U1374 ( .A(n3705), .Y(n3697) );
  CLKBUFX2TS U1375 ( .A(n3733), .Y(n3731) );
  CLKBUFX2TS U1376 ( .A(n3838), .Y(n3827) );
  CLKBUFX2TS U1377 ( .A(n3839), .Y(n3838) );
  CLKBUFX2TS U1378 ( .A(n3821), .Y(n3820) );
  CLKBUFX2TS U1379 ( .A(n3850), .Y(n3849) );
  INVX2TS U1380 ( .A(n3524), .Y(n3519) );
  INVX2TS U1381 ( .A(n3523), .Y(n3520) );
  INVX2TS U1382 ( .A(n3522), .Y(n3521) );
  INVX2TS U1383 ( .A(n3458), .Y(n3445) );
  CLKBUFX2TS U1384 ( .A(n3459), .Y(n3458) );
  INVX2TS U1385 ( .A(n3458), .Y(n3446) );
  INVX2TS U1386 ( .A(n3459), .Y(n3444) );
  INVX2TS U1387 ( .A(n3459), .Y(n3447) );
  INVX2TS U1388 ( .A(n3459), .Y(n3448) );
  INVX2TS U1389 ( .A(n3458), .Y(n3449) );
  INVX2TS U1390 ( .A(n3458), .Y(n3450) );
  INVX2TS U1391 ( .A(n3460), .Y(n3451) );
  INVX2TS U1392 ( .A(n3407), .Y(n3396) );
  INVX2TS U1393 ( .A(n3406), .Y(n3392) );
  INVX2TS U1394 ( .A(n3407), .Y(n3394) );
  INVX2TS U1395 ( .A(n3405), .Y(n3398) );
  INVX2TS U1396 ( .A(n3405), .Y(n3393) );
  CLKBUFX2TS U1397 ( .A(n3406), .Y(n3405) );
  INVX2TS U1398 ( .A(n3407), .Y(n3395) );
  INVX2TS U1399 ( .A(n3405), .Y(n3397) );
  INVX2TS U1400 ( .A(n3407), .Y(n3399) );
  CLKBUFX2TS U1401 ( .A(reset), .Y(n4539) );
  CLKBUFX2TS U1402 ( .A(n3784), .Y(n3783) );
  CLKBUFX2TS U1403 ( .A(n3784), .Y(n3782) );
  CLKBUFX2TS U1404 ( .A(n3785), .Y(n3781) );
  CLKBUFX2TS U1405 ( .A(n3785), .Y(n3779) );
  CLKBUFX2TS U1406 ( .A(n3785), .Y(n3780) );
  CLKBUFX2TS U1407 ( .A(n3372), .Y(n3363) );
  CLKBUFX2TS U1408 ( .A(n3372), .Y(n3362) );
  CLKBUFX2TS U1409 ( .A(n3371), .Y(n3364) );
  CLKBUFX2TS U1410 ( .A(n3370), .Y(n3366) );
  CLKBUFX2TS U1411 ( .A(n3369), .Y(n3367) );
  CLKBUFX2TS U1412 ( .A(n3369), .Y(n3368) );
  CLKBUFX2TS U1413 ( .A(n3371), .Y(n3365) );
  CLKBUFX2TS U1414 ( .A(n3305), .Y(n3296) );
  CLKBUFX2TS U1415 ( .A(n3304), .Y(n3298) );
  CLKBUFX2TS U1416 ( .A(n3305), .Y(n3297) );
  CLKBUFX2TS U1417 ( .A(n3304), .Y(n3299) );
  CLKBUFX2TS U1418 ( .A(n3205), .Y(n3197) );
  CLKBUFX2TS U1419 ( .A(n3205), .Y(n3196) );
  CLKBUFX2TS U1420 ( .A(n3301), .Y(n3300) );
  CLKBUFX2TS U1421 ( .A(n3203), .Y(n3201) );
  CLKBUFX2TS U1422 ( .A(n3204), .Y(n3198) );
  CLKBUFX2TS U1423 ( .A(n3204), .Y(n3199) );
  CLKBUFX2TS U1424 ( .A(n3203), .Y(n3200) );
  CLKBUFX2TS U1425 ( .A(n1049), .Y(n1047) );
  CLKBUFX2TS U1426 ( .A(n1049), .Y(n1046) );
  CLKBUFX2TS U1427 ( .A(n1049), .Y(n1045) );
  CLKBUFX2TS U1428 ( .A(n2117), .Y(n1048) );
  CLKBUFX2TS U1429 ( .A(n1098), .Y(n3758) );
  CLKBUFX2TS U1430 ( .A(n1098), .Y(n3759) );
  CLKBUFX2TS U1431 ( .A(n3769), .Y(n3760) );
  CLKBUFX2TS U1432 ( .A(n3769), .Y(n3761) );
  CLKBUFX2TS U1433 ( .A(n3769), .Y(n3762) );
  CLKBUFX2TS U1434 ( .A(n3769), .Y(n3763) );
  CLKBUFX2TS U1435 ( .A(n3767), .Y(n3766) );
  CLKBUFX2TS U1436 ( .A(n3768), .Y(n3764) );
  CLKBUFX2TS U1437 ( .A(n3768), .Y(n3765) );
  CLKBUFX2TS U1438 ( .A(n1154), .Y(n3509) );
  CLKBUFX2TS U1439 ( .A(n3675), .Y(n3670) );
  CLKBUFX2TS U1440 ( .A(n3675), .Y(n3671) );
  CLKBUFX2TS U1441 ( .A(n3675), .Y(n3672) );
  CLKBUFX2TS U1442 ( .A(n3527), .Y(n3524) );
  CLKBUFX2TS U1443 ( .A(n3527), .Y(n3522) );
  CLKBUFX2TS U1444 ( .A(n3527), .Y(n3523) );
  CLKBUFX2TS U1445 ( .A(n3626), .Y(n3624) );
  CLKBUFX2TS U1446 ( .A(n1154), .Y(n3508) );
  CLKBUFX2TS U1447 ( .A(n1187), .Y(n3359) );
  CLKBUFX2TS U1448 ( .A(n3477), .Y(n3471) );
  CLKBUFX2TS U1449 ( .A(n3477), .Y(n3472) );
  CLKBUFX2TS U1450 ( .A(n3627), .Y(n3620) );
  CLKBUFX2TS U1451 ( .A(n3627), .Y(n3621) );
  CLKBUFX2TS U1452 ( .A(n3627), .Y(n3622) );
  CLKBUFX2TS U1453 ( .A(n3510), .Y(n3504) );
  CLKBUFX2TS U1454 ( .A(n1154), .Y(n3510) );
  CLKBUFX2TS U1455 ( .A(n3626), .Y(n3625) );
  CLKBUFX2TS U1456 ( .A(n3657), .Y(n3652) );
  CLKBUFX2TS U1457 ( .A(n3425), .Y(n3424) );
  CLKBUFX2TS U1458 ( .A(n3425), .Y(n3422) );
  CLKBUFX2TS U1459 ( .A(n3425), .Y(n3423) );
  CLKBUFX2TS U1460 ( .A(n3906), .Y(n3904) );
  CLKBUFX2TS U1461 ( .A(n3905), .Y(n3903) );
  CLKBUFX2TS U1462 ( .A(n3826), .Y(n3821) );
  CLKBUFX2TS U1463 ( .A(n3826), .Y(n3822) );
  CLKBUFX2TS U1464 ( .A(n3826), .Y(n3823) );
  CLKBUFX2TS U1465 ( .A(n3739), .Y(n3736) );
  CLKBUFX2TS U1466 ( .A(n3739), .Y(n3737) );
  CLKBUFX2TS U1467 ( .A(n3739), .Y(n3738) );
  CLKBUFX2TS U1468 ( .A(n3560), .Y(n3554) );
  CLKBUFX2TS U1469 ( .A(n3560), .Y(n3555) );
  CLKBUFX2TS U1470 ( .A(n3559), .Y(n3556) );
  CLKBUFX2TS U1471 ( .A(n1203), .Y(n3293) );
  CLKBUFX2TS U1472 ( .A(n3559), .Y(n3557) );
  CLKBUFX2TS U1473 ( .A(n3559), .Y(n3558) );
  CLKBUFX2TS U1474 ( .A(n1203), .Y(n3292) );
  CLKBUFX2TS U1475 ( .A(n3277), .Y(n3271) );
  CLKBUFX2TS U1476 ( .A(n1137), .Y(n3587) );
  CLKBUFX2TS U1477 ( .A(n3656), .Y(n3653) );
  CLKBUFX2TS U1478 ( .A(n3854), .Y(n3850) );
  CLKBUFX2TS U1479 ( .A(n3854), .Y(n3851) );
  CLKBUFX2TS U1480 ( .A(n3854), .Y(n3852) );
  CLKBUFX2TS U1481 ( .A(n3294), .Y(n3288) );
  CLKBUFX2TS U1482 ( .A(n3294), .Y(n3289) );
  CLKBUFX2TS U1483 ( .A(n3276), .Y(n3273) );
  CLKBUFX2TS U1484 ( .A(n3277), .Y(n3272) );
  CLKBUFX2TS U1485 ( .A(n3294), .Y(n3290) );
  CLKBUFX2TS U1486 ( .A(n3276), .Y(n3274) );
  CLKBUFX2TS U1487 ( .A(n3476), .Y(n3475) );
  CLKBUFX2TS U1488 ( .A(n3294), .Y(n3291) );
  CLKBUFX2TS U1489 ( .A(n3276), .Y(n3275) );
  CLKBUFX2TS U1490 ( .A(n3476), .Y(n3473) );
  CLKBUFX2TS U1491 ( .A(n3476), .Y(n3474) );
  CLKBUFX2TS U1492 ( .A(n1137), .Y(n3588) );
  CLKBUFX2TS U1493 ( .A(n3544), .Y(n3538) );
  CLKBUFX2TS U1494 ( .A(n3588), .Y(n3590) );
  CLKBUFX2TS U1495 ( .A(n3543), .Y(n3540) );
  CLKBUFX2TS U1496 ( .A(n1137), .Y(n3589) );
  CLKBUFX2TS U1497 ( .A(n3544), .Y(n3539) );
  CLKBUFX2TS U1498 ( .A(n3588), .Y(n3591) );
  CLKBUFX2TS U1499 ( .A(n3543), .Y(n3541) );
  CLKBUFX2TS U1500 ( .A(n1137), .Y(n3592) );
  CLKBUFX2TS U1501 ( .A(n3543), .Y(n3542) );
  CLKBUFX2TS U1502 ( .A(n3192), .Y(n3127) );
  CLKBUFX2TS U1503 ( .A(n3193), .Y(n3125) );
  CLKBUFX2TS U1504 ( .A(n3193), .Y(n3126) );
  CLKBUFX2TS U1505 ( .A(n3192), .Y(n3128) );
  CLKBUFX2TS U1506 ( .A(n3192), .Y(n3152) );
  CLKBUFX2TS U1507 ( .A(n3656), .Y(n3654) );
  CLKBUFX2TS U1508 ( .A(n3708), .Y(n3706) );
  CLKBUFX2TS U1509 ( .A(n3692), .Y(n3689) );
  CLKBUFX2TS U1510 ( .A(n3708), .Y(n3703) );
  CLKBUFX2TS U1511 ( .A(n1105), .Y(n3704) );
  CLKBUFX2TS U1512 ( .A(n1106), .Y(n3690) );
  CLKBUFX2TS U1513 ( .A(n3708), .Y(n3705) );
  CLKBUFX2TS U1514 ( .A(n3692), .Y(n3691) );
  CLKBUFX2TS U1515 ( .A(n3656), .Y(n3655) );
  CLKBUFX2TS U1516 ( .A(n3708), .Y(n3707) );
  CLKBUFX2TS U1517 ( .A(n3692), .Y(n3688) );
  CLKBUFX2TS U1518 ( .A(n3426), .Y(n3421) );
  CLKBUFX2TS U1519 ( .A(n1201), .Y(n3320) );
  CLKBUFX2TS U1520 ( .A(n3325), .Y(n3322) );
  CLKBUFX2TS U1521 ( .A(n1201), .Y(n3321) );
  CLKBUFX2TS U1522 ( .A(n3325), .Y(n3323) );
  CLKBUFX2TS U1523 ( .A(n3325), .Y(n3324) );
  CLKBUFX2TS U1524 ( .A(n3822), .Y(n3824) );
  CLKBUFX2TS U1525 ( .A(n3821), .Y(n3825) );
  CLKBUFX2TS U1526 ( .A(n3740), .Y(n3734) );
  CLKBUFX2TS U1527 ( .A(n3740), .Y(n3735) );
  CLKBUFX2TS U1528 ( .A(n3740), .Y(n3733) );
  CLKBUFX2TS U1529 ( .A(n3242), .Y(n3235) );
  CLKBUFX2TS U1530 ( .A(n1218), .Y(n3242) );
  CLKBUFX2TS U1531 ( .A(n3908), .Y(n3905) );
  CLKBUFX2TS U1532 ( .A(n3908), .Y(n3906) );
  CLKBUFX2TS U1533 ( .A(n1185), .Y(n3390) );
  CLKBUFX2TS U1534 ( .A(n1185), .Y(n3391) );
  CLKBUFX2TS U1535 ( .A(n730), .Y(n3880) );
  CLKBUFX2TS U1536 ( .A(n1219), .Y(n3225) );
  CLKBUFX2TS U1537 ( .A(n1170), .Y(n3442) );
  CLKBUFX2TS U1538 ( .A(n1170), .Y(n3443) );
  CLKBUFX2TS U1539 ( .A(n736), .Y(n3840) );
  CLKBUFX2TS U1540 ( .A(n736), .Y(n3839) );
  CLKBUFX2TS U1541 ( .A(n724), .Y(n3921) );
  CLKBUFX2TS U1542 ( .A(n1218), .Y(n3240) );
  INVX2TS U1543 ( .A(n3673), .Y(n3659) );
  CLKBUFX2TS U1544 ( .A(n3674), .Y(n3673) );
  INVX2TS U1545 ( .A(n3673), .Y(n3660) );
  INVX2TS U1546 ( .A(n3674), .Y(n3661) );
  INVX2TS U1547 ( .A(n3674), .Y(n3662) );
  INVX2TS U1548 ( .A(n3674), .Y(n3663) );
  INVX2TS U1549 ( .A(n3675), .Y(n3664) );
  INVX2TS U1550 ( .A(n3673), .Y(n3665) );
  INVX2TS U1551 ( .A(n743), .Y(n3666) );
  CLKBUFX2TS U1552 ( .A(n3477), .Y(n3470) );
  CLKBUFX2TS U1553 ( .A(n3409), .Y(n3406) );
  CLKBUFX2TS U1554 ( .A(n3409), .Y(n3407) );
  CLKBUFX2TS U1555 ( .A(n737), .Y(n3459) );
  CLKBUFX2TS U1556 ( .A(n3409), .Y(n3408) );
  CLKBUFX2TS U1557 ( .A(n737), .Y(n3460) );
  CLKBUFX2TS U1558 ( .A(n3123), .Y(n3122) );
  CLKBUFX2TS U1559 ( .A(n3651), .Y(n3650) );
  CLKBUFX2TS U1560 ( .A(n3561), .Y(n3553) );
  CLKBUFX2TS U1561 ( .A(n3325), .Y(n3319) );
  CLKBUFX2TS U1562 ( .A(n3589), .Y(n3586) );
  CLKBUFX2TS U1563 ( .A(n3735), .Y(n3732) );
  INVX2TS U1564 ( .A(n3115), .Y(n3098) );
  INVX2TS U1565 ( .A(n3525), .Y(n3512) );
  INVX2TS U1566 ( .A(n3525), .Y(n3513) );
  INVX2TS U1567 ( .A(n3526), .Y(n3514) );
  INVX2TS U1568 ( .A(n3526), .Y(n3515) );
  INVX2TS U1569 ( .A(n3525), .Y(n3517) );
  INVX2TS U1570 ( .A(n3526), .Y(n3518) );
  INVX2TS U1571 ( .A(n3526), .Y(n3516) );
  INVX2TS U1572 ( .A(n3525), .Y(n3511) );
  CLKBUFX2TS U1573 ( .A(n3750), .Y(n3746) );
  CLKBUFX2TS U1574 ( .A(n3750), .Y(n3745) );
  CLKBUFX2TS U1575 ( .A(n3751), .Y(n3744) );
  CLKBUFX2TS U1576 ( .A(n3751), .Y(n3743) );
  CLKBUFX2TS U1577 ( .A(n3752), .Y(n3742) );
  CLKBUFX2TS U1578 ( .A(n3752), .Y(n3741) );
  INVX2TS U1579 ( .A(n3112), .Y(n3100) );
  INVX2TS U1580 ( .A(n3109), .Y(n3104) );
  INVX2TS U1581 ( .A(n3109), .Y(n3103) );
  INVX2TS U1582 ( .A(n3108), .Y(n3102) );
  INVX2TS U1583 ( .A(n3114), .Y(n3101) );
  INVX2TS U1584 ( .A(n3109), .Y(n3105) );
  INVX2TS U1585 ( .A(n3108), .Y(n3106) );
  INVX2TS U1586 ( .A(n3108), .Y(n3107) );
  INVX2TS U1587 ( .A(n3608), .Y(n3603) );
  INVX2TS U1588 ( .A(n3609), .Y(n3602) );
  INVX2TS U1589 ( .A(n3607), .Y(n3601) );
  INVX2TS U1590 ( .A(n3340), .Y(n3336) );
  INVX2TS U1591 ( .A(n3340), .Y(n3335) );
  INVX2TS U1592 ( .A(n3340), .Y(n3334) );
  INVX2TS U1593 ( .A(n3343), .Y(n3328) );
  INVX2TS U1594 ( .A(n3608), .Y(n3595) );
  INVX2TS U1595 ( .A(n3258), .Y(n3245) );
  INVX2TS U1596 ( .A(n3341), .Y(n3333) );
  INVX2TS U1597 ( .A(n3341), .Y(n3332) );
  INVX2TS U1598 ( .A(n3341), .Y(n3331) );
  INVX2TS U1599 ( .A(n744), .Y(n3330) );
  INVX2TS U1600 ( .A(n744), .Y(n3329) );
  INVX2TS U1601 ( .A(n3607), .Y(n3600) );
  INVX2TS U1602 ( .A(n3607), .Y(n3599) );
  INVX2TS U1603 ( .A(n3607), .Y(n3598) );
  INVX2TS U1604 ( .A(n3608), .Y(n3597) );
  INVX2TS U1605 ( .A(n3608), .Y(n3596) );
  INVX2TS U1606 ( .A(n3257), .Y(n3250) );
  INVX2TS U1607 ( .A(n3257), .Y(n3248) );
  INVX2TS U1608 ( .A(n3258), .Y(n3247) );
  INVX2TS U1609 ( .A(n3258), .Y(n3246) );
  INVX2TS U1610 ( .A(n3257), .Y(n3249) );
  INVX2TS U1611 ( .A(n3258), .Y(n3251) );
  INVX2TS U1612 ( .A(n3259), .Y(n3253) );
  INVX2TS U1613 ( .A(n3260), .Y(n3252) );
  INVX2TS U1614 ( .A(n3113), .Y(n3099) );
  INVX2TS U1615 ( .A(n3259), .Y(n3243) );
  INVX2TS U1616 ( .A(n3342), .Y(n3326) );
  INVX2TS U1617 ( .A(n3342), .Y(n3327) );
  INVX2TS U1618 ( .A(n3609), .Y(n3593) );
  INVX2TS U1619 ( .A(n3609), .Y(n3594) );
  INVX2TS U1620 ( .A(n3259), .Y(n3244) );
  CLKBUFX2TS U1621 ( .A(n3308), .Y(n3301) );
  CLKBUFX2TS U1622 ( .A(n3307), .Y(n3305) );
  CLKBUFX2TS U1623 ( .A(n3308), .Y(n3303) );
  CLKBUFX2TS U1624 ( .A(n3308), .Y(n3302) );
  CLKBUFX2TS U1625 ( .A(n3307), .Y(n3304) );
  CLKBUFX2TS U1626 ( .A(n1186), .Y(n3369) );
  CLKBUFX2TS U1627 ( .A(n3207), .Y(n3204) );
  CLKBUFX2TS U1628 ( .A(n3208), .Y(n3203) );
  CLKBUFX2TS U1629 ( .A(n3208), .Y(n3202) );
  CLKBUFX2TS U1630 ( .A(n3374), .Y(n3371) );
  CLKBUFX2TS U1631 ( .A(n1186), .Y(n3370) );
  CLKBUFX2TS U1632 ( .A(n3207), .Y(n3205) );
  CLKBUFX2TS U1633 ( .A(n3374), .Y(n3372) );
  CLKBUFX2TS U1634 ( .A(n760), .Y(n3784) );
  CLKBUFX2TS U1635 ( .A(n760), .Y(n3785) );
  CLKBUFX2TS U1636 ( .A(n3488), .Y(n3479) );
  CLKBUFX2TS U1637 ( .A(n3488), .Y(n3480) );
  CLKBUFX2TS U1638 ( .A(n3373), .Y(n3361) );
  CLKBUFX2TS U1639 ( .A(n3374), .Y(n3373) );
  CLKBUFX2TS U1640 ( .A(n3487), .Y(n3481) );
  CLKBUFX2TS U1641 ( .A(n3487), .Y(n3482) );
  CLKBUFX2TS U1642 ( .A(n3485), .Y(n3483) );
  INVX2TS U1643 ( .A(n3096), .Y(n3081) );
  INVX2TS U1644 ( .A(n3096), .Y(n3082) );
  INVX2TS U1645 ( .A(n3097), .Y(n3091) );
  INVX2TS U1646 ( .A(n3097), .Y(n3090) );
  INVX2TS U1647 ( .A(n3095), .Y(n3089) );
  INVX2TS U1648 ( .A(n3095), .Y(n3088) );
  INVX2TS U1649 ( .A(n3092), .Y(n3087) );
  INVX2TS U1650 ( .A(n3092), .Y(n3085) );
  INVX2TS U1651 ( .A(n3092), .Y(n3084) );
  INVX2TS U1652 ( .A(n3092), .Y(n3086) );
  INVX2TS U1653 ( .A(n3096), .Y(n3083) );
  CLKBUFX2TS U1654 ( .A(n3306), .Y(n3295) );
  CLKBUFX2TS U1655 ( .A(n3307), .Y(n3306) );
  CLKBUFX2TS U1656 ( .A(n3057), .Y(n3055) );
  CLKBUFX2TS U1657 ( .A(n3061), .Y(n3009) );
  CLKBUFX2TS U1658 ( .A(n3060), .Y(n3010) );
  CLKBUFX2TS U1659 ( .A(n3060), .Y(n3011) );
  CLKBUFX2TS U1660 ( .A(n3059), .Y(n3050) );
  CLKBUFX2TS U1661 ( .A(n3059), .Y(n3051) );
  CLKBUFX2TS U1662 ( .A(n3057), .Y(n3054) );
  CLKBUFX2TS U1663 ( .A(n3058), .Y(n3052) );
  CLKBUFX2TS U1664 ( .A(n3058), .Y(n3053) );
  CLKBUFX2TS U1665 ( .A(n3637), .Y(n3630) );
  CLKBUFX2TS U1666 ( .A(n3637), .Y(n3629) );
  CLKBUFX2TS U1667 ( .A(n3638), .Y(n3628) );
  CLKBUFX2TS U1668 ( .A(n3574), .Y(n3562) );
  CLKBUFX2TS U1669 ( .A(n3573), .Y(n3564) );
  CLKBUFX2TS U1670 ( .A(n3574), .Y(n3563) );
  CLKBUFX2TS U1671 ( .A(n3575), .Y(n3565) );
  CLKBUFX2TS U1672 ( .A(n3573), .Y(n3566) );
  CLKBUFX2TS U1673 ( .A(n3572), .Y(n3567) );
  CLKBUFX2TS U1674 ( .A(n3719), .Y(n3718) );
  CLKBUFX2TS U1675 ( .A(n3636), .Y(n3631) );
  CLKBUFX2TS U1676 ( .A(n3636), .Y(n3632) );
  CLKBUFX2TS U1677 ( .A(n3635), .Y(n3634) );
  CLKBUFX2TS U1678 ( .A(n3722), .Y(n3710) );
  CLKBUFX2TS U1679 ( .A(n1104), .Y(n3711) );
  CLKBUFX2TS U1680 ( .A(n3721), .Y(n3712) );
  CLKBUFX2TS U1681 ( .A(n3721), .Y(n3713) );
  CLKBUFX2TS U1682 ( .A(n3723), .Y(n3714) );
  CLKBUFX2TS U1683 ( .A(n3720), .Y(n3715) );
  CLKBUFX2TS U1684 ( .A(n3720), .Y(n3716) );
  CLKBUFX2TS U1685 ( .A(n3719), .Y(n3717) );
  CLKBUFX2TS U1686 ( .A(n3635), .Y(n3633) );
  CLKBUFX2TS U1687 ( .A(n3078), .Y(n3065) );
  CLKBUFX2TS U1688 ( .A(n3078), .Y(n3064) );
  CLKBUFX2TS U1689 ( .A(n3572), .Y(n3568) );
  CLKBUFX2TS U1690 ( .A(n3571), .Y(n3569) );
  CLKBUFX2TS U1691 ( .A(n3571), .Y(n3570) );
  CLKBUFX2TS U1692 ( .A(n2924), .Y(n2109) );
  CLKBUFX2TS U1693 ( .A(n3074), .Y(n3072) );
  CLKBUFX2TS U1694 ( .A(n3074), .Y(n3071) );
  CLKBUFX2TS U1695 ( .A(n3076), .Y(n3069) );
  CLKBUFX2TS U1696 ( .A(n3080), .Y(n3070) );
  CLKBUFX2TS U1697 ( .A(n3077), .Y(n3066) );
  CLKBUFX2TS U1698 ( .A(n3076), .Y(n3068) );
  CLKBUFX2TS U1699 ( .A(n3077), .Y(n3067) );
  CLKBUFX2TS U1700 ( .A(n3206), .Y(n3195) );
  CLKBUFX2TS U1701 ( .A(n3207), .Y(n3206) );
  CLKBUFX2TS U1702 ( .A(n2920), .Y(n2919) );
  CLKBUFX2TS U1703 ( .A(n2920), .Y(n2918) );
  CLKBUFX2TS U1704 ( .A(n2921), .Y(n2917) );
  CLKBUFX2TS U1705 ( .A(n2921), .Y(n2916) );
  CLKBUFX2TS U1706 ( .A(n2924), .Y(n2905) );
  CLKBUFX2TS U1707 ( .A(n2923), .Y(n2915) );
  CLKBUFX2TS U1708 ( .A(n2923), .Y(n2906) );
  INVX2TS U1709 ( .A(n1167), .Y(n1151) );
  INVX2TS U1710 ( .A(n1198), .Y(n1134) );
  INVX2TS U1711 ( .A(n1215), .Y(n1107) );
  CLKBUFX2TS U1712 ( .A(n3771), .Y(n3770) );
  CLKBUFX2TS U1713 ( .A(n1098), .Y(n3769) );
  CLKBUFX2TS U1714 ( .A(n3771), .Y(n3767) );
  CLKBUFX2TS U1715 ( .A(n3771), .Y(n3768) );
  CLKBUFX2TS U1716 ( .A(n2117), .Y(n1049) );
  CLKBUFX2TS U1717 ( .A(n1034), .Y(n1021) );
  CLKBUFX2TS U1718 ( .A(n1034), .Y(n1022) );
  CLKBUFX2TS U1719 ( .A(n1033), .Y(n1023) );
  CLKBUFX2TS U1720 ( .A(n1035), .Y(n1024) );
  CLKBUFX2TS U1721 ( .A(n2118), .Y(n1025) );
  CLKBUFX2TS U1722 ( .A(n1032), .Y(n1026) );
  CLKBUFX2TS U1723 ( .A(n1031), .Y(n1030) );
  CLKBUFX2TS U1724 ( .A(n1032), .Y(n1027) );
  CLKBUFX2TS U1725 ( .A(n1031), .Y(n1029) );
  CLKBUFX2TS U1726 ( .A(n1018), .Y(n1008) );
  CLKBUFX2TS U1727 ( .A(n1017), .Y(n1009) );
  CLKBUFX2TS U1728 ( .A(n1017), .Y(n1010) );
  CLKBUFX2TS U1729 ( .A(n1016), .Y(n1011) );
  CLKBUFX2TS U1730 ( .A(n1015), .Y(n1014) );
  CLKBUFX2TS U1731 ( .A(n1016), .Y(n1012) );
  CLKBUFX2TS U1732 ( .A(n1015), .Y(n1013) );
  CLKBUFX2TS U1733 ( .A(n977), .Y(n928) );
  CLKBUFX2TS U1734 ( .A(n991), .Y(n979) );
  CLKBUFX2TS U1735 ( .A(n977), .Y(n932) );
  CLKBUFX2TS U1736 ( .A(n2121), .Y(n980) );
  CLKBUFX2TS U1737 ( .A(n976), .Y(n933) );
  CLKBUFX2TS U1738 ( .A(n990), .Y(n981) );
  CLKBUFX2TS U1739 ( .A(n990), .Y(n982) );
  CLKBUFX2TS U1740 ( .A(n978), .Y(n956) );
  CLKBUFX2TS U1741 ( .A(n976), .Y(n961) );
  CLKBUFX2TS U1742 ( .A(n992), .Y(n983) );
  CLKBUFX2TS U1743 ( .A(n975), .Y(n962) );
  CLKBUFX2TS U1744 ( .A(n989), .Y(n984) );
  CLKBUFX2TS U1745 ( .A(n974), .Y(n965) );
  CLKBUFX2TS U1746 ( .A(n988), .Y(n987) );
  CLKBUFX2TS U1747 ( .A(n975), .Y(n963) );
  CLKBUFX2TS U1748 ( .A(n989), .Y(n985) );
  CLKBUFX2TS U1749 ( .A(n974), .Y(n964) );
  CLKBUFX2TS U1750 ( .A(n988), .Y(n986) );
  CLKBUFX2TS U1751 ( .A(n1075), .Y(n1065) );
  CLKBUFX2TS U1752 ( .A(n1004), .Y(n994) );
  CLKBUFX2TS U1753 ( .A(n1075), .Y(n1066) );
  CLKBUFX2TS U1754 ( .A(n1004), .Y(n995) );
  CLKBUFX2TS U1755 ( .A(n1074), .Y(n1067) );
  CLKBUFX2TS U1756 ( .A(n1003), .Y(n996) );
  CLKBUFX2TS U1757 ( .A(n1074), .Y(n1068) );
  CLKBUFX2TS U1758 ( .A(n1003), .Y(n997) );
  CLKBUFX2TS U1759 ( .A(n1075), .Y(n1069) );
  CLKBUFX2TS U1760 ( .A(n1002), .Y(n998) );
  CLKBUFX2TS U1761 ( .A(n1073), .Y(n1072) );
  CLKBUFX2TS U1762 ( .A(n1002), .Y(n1001) );
  CLKBUFX2TS U1763 ( .A(n1076), .Y(n1070) );
  CLKBUFX2TS U1764 ( .A(n1002), .Y(n999) );
  CLKBUFX2TS U1765 ( .A(n1073), .Y(n1071) );
  CLKBUFX2TS U1766 ( .A(n1002), .Y(n1000) );
  CLKBUFX2TS U1767 ( .A(n1059), .Y(n1051) );
  CLKBUFX2TS U1768 ( .A(n1059), .Y(n1052) );
  CLKBUFX2TS U1769 ( .A(n1058), .Y(n1053) );
  CLKBUFX2TS U1770 ( .A(n1057), .Y(n1056) );
  CLKBUFX2TS U1771 ( .A(n1058), .Y(n1054) );
  CLKBUFX2TS U1772 ( .A(n1057), .Y(n1055) );
  NOR3BX1TS U1773 ( .AN(n444), .B(n1790), .C(n927), .Y(n1154) );
  CLKBUFX2TS U1774 ( .A(n1123), .Y(n3627) );
  CLKBUFX2TS U1775 ( .A(n1123), .Y(n3626) );
  CLKBUFX2TS U1776 ( .A(n1121), .Y(n3656) );
  CLKBUFX2TS U1777 ( .A(n1171), .Y(n3425) );
  CLKBUFX2TS U1778 ( .A(n1103), .Y(n3739) );
  CLKBUFX2TS U1779 ( .A(n161), .Y(n3826) );
  CLKBUFX2TS U1780 ( .A(n1221), .Y(n3194) );
  CLKBUFX2TS U1781 ( .A(n1139), .Y(n3561) );
  CLKBUFX2TS U1782 ( .A(n3658), .Y(n3651) );
  CLKBUFX2TS U1783 ( .A(n1121), .Y(n3658) );
  CLKBUFX2TS U1784 ( .A(n1105), .Y(n3709) );
  CLKBUFX2TS U1785 ( .A(n3755), .Y(n3754) );
  CLKBUFX2TS U1786 ( .A(n1221), .Y(n3192) );
  CLKBUFX2TS U1787 ( .A(n1204), .Y(n3277) );
  CLKBUFX2TS U1788 ( .A(n1204), .Y(n3276) );
  CLKBUFX2TS U1789 ( .A(n1203), .Y(n3294) );
  CLKBUFX2TS U1790 ( .A(n1105), .Y(n3708) );
  CLKBUFX2TS U1791 ( .A(n1106), .Y(n3692) );
  CLKBUFX2TS U1792 ( .A(n1156), .Y(n3476) );
  CLKBUFX2TS U1793 ( .A(n1140), .Y(n3544) );
  CLKBUFX2TS U1794 ( .A(n1140), .Y(n3543) );
  CLKBUFX2TS U1795 ( .A(n734), .Y(n3853) );
  CLKBUFX2TS U1796 ( .A(n734), .Y(n3854) );
  CLKBUFX2TS U1797 ( .A(n1139), .Y(n3560) );
  CLKBUFX2TS U1798 ( .A(n1139), .Y(n3559) );
  CLKBUFX2TS U1799 ( .A(n1201), .Y(n3325) );
  CLKBUFX2TS U1800 ( .A(n1103), .Y(n3740) );
  INVX2TS U1801 ( .A(n1806), .Y(n748) );
  INVX2TS U1802 ( .A(n1756), .Y(n736) );
  INVX2TS U1803 ( .A(n459), .Y(n724) );
  CLKBUFX2TS U1804 ( .A(n10), .Y(n3908) );
  CLKBUFX2TS U1805 ( .A(n743), .Y(n3674) );
  CLKBUFX2TS U1806 ( .A(n738), .Y(n3526) );
  CLKBUFX2TS U1807 ( .A(n738), .Y(n3525) );
  INVX2TS U1808 ( .A(n1765), .Y(n745) );
  CLKBUFX2TS U1809 ( .A(n743), .Y(n3675) );
  CLKBUFX2TS U1810 ( .A(n738), .Y(n3527) );
  CLKBUFX2TS U1811 ( .A(n3343), .Y(n3342) );
  CLKBUFX2TS U1812 ( .A(n3260), .Y(n3259) );
  CLKBUFX2TS U1813 ( .A(n3756), .Y(n3750) );
  CLKBUFX2TS U1814 ( .A(n3756), .Y(n3751) );
  CLKBUFX2TS U1815 ( .A(n3756), .Y(n3752) );
  CLKBUFX2TS U1816 ( .A(n3755), .Y(n3753) );
  CLKBUFX2TS U1817 ( .A(n3112), .Y(n3110) );
  CLKBUFX2TS U1818 ( .A(n3112), .Y(n3111) );
  CLKBUFX2TS U1819 ( .A(n3749), .Y(n3747) );
  CLKBUFX2TS U1820 ( .A(n3749), .Y(n3748) );
  INVX2TS U1821 ( .A(n3342), .Y(n3338) );
  INVX2TS U1822 ( .A(n3342), .Y(n3337) );
  INVX2TS U1823 ( .A(n749), .Y(n3255) );
  INVX2TS U1824 ( .A(n749), .Y(n3254) );
  CLKBUFX2TS U1825 ( .A(n762), .Y(n1167) );
  CLKBUFX2TS U1826 ( .A(n1751), .Y(n1198) );
  CLKBUFX2TS U1827 ( .A(n762), .Y(n1215) );
  CLKBUFX2TS U1828 ( .A(n3641), .Y(n3637) );
  CLKBUFX2TS U1829 ( .A(n3490), .Y(n3487) );
  CLKBUFX2TS U1830 ( .A(n3491), .Y(n3485) );
  CLKBUFX2TS U1831 ( .A(n3491), .Y(n3486) );
  CLKBUFX2TS U1832 ( .A(n3491), .Y(n3484) );
  CLKBUFX2TS U1833 ( .A(n3490), .Y(n3488) );
  CLKBUFX2TS U1834 ( .A(n3575), .Y(n3574) );
  CLKBUFX2TS U1835 ( .A(n3575), .Y(n3572) );
  CLKBUFX2TS U1836 ( .A(n1138), .Y(n3573) );
  CLKBUFX2TS U1837 ( .A(n3575), .Y(n3571) );
  CLKBUFX2TS U1838 ( .A(n3079), .Y(n3078) );
  CLKBUFX2TS U1839 ( .A(n3080), .Y(n3074) );
  CLKBUFX2TS U1840 ( .A(n2926), .Y(n2920) );
  CLKBUFX2TS U1841 ( .A(n3080), .Y(n3075) );
  CLKBUFX2TS U1842 ( .A(n2054), .Y(n2921) );
  CLKBUFX2TS U1843 ( .A(n3061), .Y(n3060) );
  CLKBUFX2TS U1844 ( .A(n2054), .Y(n2922) );
  CLKBUFX2TS U1845 ( .A(n3062), .Y(n3059) );
  CLKBUFX2TS U1846 ( .A(n2926), .Y(n2924) );
  CLKBUFX2TS U1847 ( .A(n3062), .Y(n3057) );
  CLKBUFX2TS U1848 ( .A(n3079), .Y(n3076) );
  CLKBUFX2TS U1849 ( .A(n2926), .Y(n2923) );
  CLKBUFX2TS U1850 ( .A(n3062), .Y(n3058) );
  CLKBUFX2TS U1851 ( .A(n3079), .Y(n3077) );
  CLKBUFX2TS U1852 ( .A(n3640), .Y(n3638) );
  CLKBUFX2TS U1853 ( .A(n3641), .Y(n3636) );
  CLKBUFX2TS U1854 ( .A(n3723), .Y(n3721) );
  CLKBUFX2TS U1855 ( .A(n3723), .Y(n3720) );
  CLKBUFX2TS U1856 ( .A(n3723), .Y(n3719) );
  CLKBUFX2TS U1857 ( .A(n3640), .Y(n3639) );
  CLKBUFX2TS U1858 ( .A(n3641), .Y(n3635) );
  CLKBUFX2TS U1859 ( .A(n1202), .Y(n3308) );
  CLKBUFX2TS U1860 ( .A(n1202), .Y(n3307) );
  CLKBUFX2TS U1861 ( .A(n1220), .Y(n3208) );
  CLKBUFX2TS U1862 ( .A(n1220), .Y(n3207) );
  CLKBUFX2TS U1863 ( .A(n1186), .Y(n3374) );
  CLKBUFX2TS U1864 ( .A(n3489), .Y(n3478) );
  CLKBUFX2TS U1865 ( .A(n3490), .Y(n3489) );
  CLKBUFX2TS U1866 ( .A(n3095), .Y(n3093) );
  CLKBUFX2TS U1867 ( .A(n3095), .Y(n3094) );
  CLKBUFX2TS U1868 ( .A(n1104), .Y(n3722) );
  INVX2TS U1869 ( .A(n1805), .Y(n754) );
  CLKBUFX2TS U1870 ( .A(n3063), .Y(n3056) );
  CLKBUFX2TS U1871 ( .A(n4217), .Y(n4219) );
  CLKBUFX2TS U1872 ( .A(n4220), .Y(n4222) );
  CLKBUFX2TS U1873 ( .A(n3079), .Y(n3073) );
  CLKBUFX2TS U1874 ( .A(n2925), .Y(n1939) );
  CLKBUFX2TS U1875 ( .A(n2926), .Y(n2925) );
  INVX2TS U1876 ( .A(n1215), .Y(n1078) );
  INVX2TS U1877 ( .A(n1751), .Y(n1079) );
  CLKBUFX2TS U1878 ( .A(n762), .Y(n1751) );
  INVX2TS U1879 ( .A(n1751), .Y(n1080) );
  INVX2TS U1880 ( .A(n1798), .Y(n1081) );
  INVX2TS U1881 ( .A(n1798), .Y(n1082) );
  INVX2TS U1882 ( .A(n1751), .Y(n1084) );
  INVX2TS U1883 ( .A(n1798), .Y(n1085) );
  INVX2TS U1884 ( .A(n1798), .Y(n1091) );
  NAND2X1TS U1885 ( .A(n141), .B(n550), .Y(n2117) );
  INVX2TS U1886 ( .A(n1087), .Y(n914) );
  CLKBUFX2TS U1887 ( .A(n1035), .Y(n1034) );
  CLKBUFX2TS U1888 ( .A(n2118), .Y(n1033) );
  CLKBUFX2TS U1889 ( .A(n1035), .Y(n1032) );
  CLKBUFX2TS U1890 ( .A(n1035), .Y(n1031) );
  CLKBUFX2TS U1891 ( .A(n978), .Y(n977) );
  CLKBUFX2TS U1892 ( .A(n1062), .Y(n1060) );
  CLKBUFX2TS U1893 ( .A(n2123), .Y(n976) );
  CLKBUFX2TS U1894 ( .A(n2114), .Y(n1075) );
  CLKBUFX2TS U1895 ( .A(n992), .Y(n990) );
  CLKBUFX2TS U1896 ( .A(n2120), .Y(n1004) );
  CLKBUFX2TS U1897 ( .A(n1063), .Y(n1059) );
  CLKBUFX2TS U1898 ( .A(n1077), .Y(n1074) );
  CLKBUFX2TS U1899 ( .A(n1006), .Y(n1003) );
  CLKBUFX2TS U1900 ( .A(n1020), .Y(n1017) );
  CLKBUFX2TS U1901 ( .A(n978), .Y(n975) );
  CLKBUFX2TS U1902 ( .A(n1063), .Y(n1058) );
  CLKBUFX2TS U1903 ( .A(n992), .Y(n989) );
  CLKBUFX2TS U1904 ( .A(n1020), .Y(n1016) );
  CLKBUFX2TS U1905 ( .A(n978), .Y(n974) );
  CLKBUFX2TS U1906 ( .A(n1063), .Y(n1057) );
  CLKBUFX2TS U1907 ( .A(n1077), .Y(n1073) );
  CLKBUFX2TS U1908 ( .A(n992), .Y(n988) );
  CLKBUFX2TS U1909 ( .A(n1006), .Y(n1002) );
  CLKBUFX2TS U1910 ( .A(n1020), .Y(n1015) );
  CLKBUFX2TS U1911 ( .A(n1098), .Y(n3771) );
  CLKBUFX2TS U1912 ( .A(n4217), .Y(n4218) );
  CLKBUFX2TS U1913 ( .A(n4220), .Y(n4221) );
  CLKBUFX2TS U1914 ( .A(n1018), .Y(n1007) );
  CLKBUFX2TS U1915 ( .A(n1019), .Y(n1018) );
  CLKBUFX2TS U1916 ( .A(n2121), .Y(n991) );
  CLKBUFX2TS U1917 ( .A(n1076), .Y(n1064) );
  CLKBUFX2TS U1918 ( .A(n2114), .Y(n1076) );
  CLKBUFX2TS U1919 ( .A(n1005), .Y(n993) );
  CLKBUFX2TS U1920 ( .A(n2120), .Y(n1005) );
  CLKBUFX2TS U1921 ( .A(n1061), .Y(n1050) );
  CLKBUFX2TS U1922 ( .A(n1062), .Y(n1061) );
  INVX2TS U1923 ( .A(n4197), .Y(n4195) );
  NOR2X1TS U1924 ( .A(n1766), .B(n1769), .Y(n1106) );
  NOR2BX1TS U1925 ( .AN(n1844), .B(n1803), .Y(n1772) );
  AOI21X1TS U1926 ( .A0(n931), .A1(n105), .B0(n733), .Y(n1776) );
  NOR2BX1TS U1927 ( .AN(n117), .B(n1940), .Y(n1779) );
  XNOR2X1TS U1928 ( .A(n2396), .B(n2394), .Y(n1089) );
  XOR2X1TS U1929 ( .A(n3), .B(n2393), .Y(n2396) );
  OAI211X1TS U1930 ( .A0(n111), .A1(n116), .B0(n1812), .C0(n1940), .Y(n1789)
         );
  AOI2BB1X1TS U1931 ( .A0N(n751), .A1N(n1914), .B0(n1818), .Y(n1816) );
  NOR3X1TS U1932 ( .A(n1772), .B(n1774), .C(n758), .Y(n1773) );
  NAND3X1TS U1933 ( .A(n110), .B(n3), .C(n751), .Y(n1768) );
  NOR2X1TS U1934 ( .A(n435), .B(n116), .Y(n1806) );
  NOR2X1TS U1935 ( .A(n116), .B(n1940), .Y(n1794) );
  INVX2TS U1936 ( .A(n1846), .Y(n930) );
  AOI21X1TS U1937 ( .A0(n931), .A1(n118), .B0(n744), .Y(n1807) );
  NOR2X1TS U1938 ( .A(n2890), .B(n2391), .Y(n2393) );
  INVX2TS U1939 ( .A(n1780), .Y(n757) );
  CLKBUFX2TS U1940 ( .A(n733), .Y(n3610) );
  INVX2TS U1941 ( .A(n1810), .Y(n753) );
  INVX2TS U1942 ( .A(n1766), .Y(n759) );
  OAI21X1TS U1943 ( .A0(n747), .A1(n1963), .B0(n1940), .Y(n1803) );
  NOR2X1TS U1944 ( .A(n111), .B(n117), .Y(n1963) );
  AO21X1TS U1945 ( .A0(n2393), .A1(n2394), .B0(n143), .Y(n2395) );
  INVX2TS U1946 ( .A(n1869), .Y(n758) );
  CLKBUFX2TS U1947 ( .A(n3115), .Y(n3113) );
  INVX2TS U1948 ( .A(n1812), .Y(n747) );
  NAND2X1TS U1949 ( .A(n761), .B(n1831), .Y(n1928) );
  INVX2TS U1950 ( .A(n2007), .Y(n752) );
  CLKBUFX2TS U1951 ( .A(n1100), .Y(n3756) );
  CLKBUFX2TS U1952 ( .A(n733), .Y(n3609) );
  CLKBUFX2TS U1953 ( .A(n3115), .Y(n3112) );
  CLKBUFX2TS U1954 ( .A(n3115), .Y(n3114) );
  CLKBUFX2TS U1955 ( .A(n733), .Y(n3608) );
  CLKBUFX2TS U1956 ( .A(n744), .Y(n3343) );
  CLKBUFX2TS U1957 ( .A(n749), .Y(n3260) );
  CLKBUFX2TS U1958 ( .A(n3757), .Y(n3749) );
  CLKBUFX2TS U1959 ( .A(n1100), .Y(n3757) );
  NOR2BX1TS U1960 ( .AN(n1860), .B(n119), .Y(n1220) );
  NOR2BX1TS U1961 ( .AN(n1860), .B(n1938), .Y(n1186) );
  CLKBUFX2TS U1962 ( .A(n3097), .Y(n3096) );
  CLKBUFX2TS U1963 ( .A(n3097), .Y(n3095) );
  CLKBUFX2TS U1964 ( .A(destinationAddressIn_SOUTH[6]), .Y(n4217) );
  CLKBUFX2TS U1965 ( .A(destinationAddressIn_SOUTH[7]), .Y(n4220) );
  CLKBUFX2TS U1966 ( .A(n2040), .Y(n3063) );
  CLKBUFX2TS U1967 ( .A(n1155), .Y(n3491) );
  CLKBUFX2TS U1968 ( .A(n1155), .Y(n3490) );
  CLKBUFX2TS U1969 ( .A(n1138), .Y(n3575) );
  CLKBUFX2TS U1970 ( .A(n1104), .Y(n3723) );
  CLKBUFX2TS U1971 ( .A(n1122), .Y(n3640) );
  CLKBUFX2TS U1972 ( .A(n1122), .Y(n3641) );
  CLKBUFX2TS U1973 ( .A(n2040), .Y(n3061) );
  CLKBUFX2TS U1974 ( .A(n2039), .Y(n3080) );
  CLKBUFX2TS U1975 ( .A(n2054), .Y(n2926) );
  CLKBUFX2TS U1976 ( .A(n2040), .Y(n3062) );
  CLKBUFX2TS U1977 ( .A(n2039), .Y(n3079) );
  CLKBUFX2TS U1978 ( .A(n762), .Y(n1798) );
  INVX2TS U1979 ( .A(n2050), .Y(n960) );
  CLKBUFX2TS U1980 ( .A(n4198), .Y(n4197) );
  NAND2X1TS U1981 ( .A(n462), .B(n550), .Y(n1098) );
  INVX2TS U1982 ( .A(n4191), .Y(n4189) );
  CLKBUFX2TS U1983 ( .A(n2115), .Y(n1062) );
  CLKBUFX2TS U1984 ( .A(n2119), .Y(n1019) );
  CLKBUFX2TS U1985 ( .A(n2115), .Y(n1063) );
  CLKBUFX2TS U1986 ( .A(n2114), .Y(n1077) );
  CLKBUFX2TS U1987 ( .A(n2121), .Y(n992) );
  CLKBUFX2TS U1988 ( .A(n2120), .Y(n1006) );
  CLKBUFX2TS U1989 ( .A(n2119), .Y(n1020) );
  CLKBUFX2TS U1990 ( .A(n2123), .Y(n978) );
  CLKBUFX2TS U1991 ( .A(n2118), .Y(n1035) );
  CLKBUFX2TS U1992 ( .A(n4118), .Y(n4119) );
  CLKBUFX2TS U1993 ( .A(n4115), .Y(n4116) );
  CLKBUFX2TS U1994 ( .A(n4112), .Y(n4113) );
  CLKBUFX2TS U1995 ( .A(n4073), .Y(n4074) );
  CLKBUFX2TS U1996 ( .A(n4166), .Y(n4167) );
  CLKBUFX2TS U1997 ( .A(n4163), .Y(n4164) );
  CLKBUFX2TS U1998 ( .A(n4160), .Y(n4161) );
  CLKBUFX2TS U1999 ( .A(n4157), .Y(n4158) );
  CLKBUFX2TS U2000 ( .A(n4154), .Y(n4155) );
  CLKBUFX2TS U2001 ( .A(n4151), .Y(n4152) );
  CLKBUFX2TS U2002 ( .A(n4148), .Y(n4149) );
  CLKBUFX2TS U2003 ( .A(n4145), .Y(n4146) );
  CLKBUFX2TS U2004 ( .A(n4142), .Y(n4143) );
  CLKBUFX2TS U2005 ( .A(n4139), .Y(n4140) );
  CLKBUFX2TS U2006 ( .A(n4136), .Y(n4137) );
  CLKBUFX2TS U2007 ( .A(n4133), .Y(n4134) );
  CLKBUFX2TS U2008 ( .A(n4130), .Y(n4131) );
  CLKBUFX2TS U2009 ( .A(n4127), .Y(n4128) );
  CLKBUFX2TS U2010 ( .A(n4124), .Y(n4125) );
  CLKBUFX2TS U2011 ( .A(n4121), .Y(n4122) );
  CLKBUFX2TS U2012 ( .A(n4109), .Y(n4110) );
  CLKBUFX2TS U2013 ( .A(n4106), .Y(n4107) );
  CLKBUFX2TS U2014 ( .A(n4103), .Y(n4104) );
  CLKBUFX2TS U2015 ( .A(n4100), .Y(n4101) );
  CLKBUFX2TS U2016 ( .A(n4097), .Y(n4098) );
  CLKBUFX2TS U2017 ( .A(n4094), .Y(n4095) );
  CLKBUFX2TS U2018 ( .A(n4091), .Y(n4092) );
  CLKBUFX2TS U2019 ( .A(n4088), .Y(n4089) );
  CLKBUFX2TS U2020 ( .A(n4082), .Y(n4083) );
  CLKBUFX2TS U2021 ( .A(n4079), .Y(n4080) );
  CLKBUFX2TS U2022 ( .A(n4076), .Y(n4077) );
  CLKBUFX2TS U2023 ( .A(n4085), .Y(n4086) );
  INVX2TS U2024 ( .A(n4288), .Y(n4286) );
  INVX2TS U2025 ( .A(n4285), .Y(n4283) );
  INVX2TS U2026 ( .A(n4282), .Y(n4280) );
  INVX2TS U2027 ( .A(n4243), .Y(n4241) );
  INVX2TS U2028 ( .A(n3979), .Y(n3977) );
  INVX2TS U2029 ( .A(n3994), .Y(n3992) );
  INVX2TS U2030 ( .A(n3988), .Y(n3986) );
  INVX2TS U2031 ( .A(n3985), .Y(n3983) );
  INVX2TS U2032 ( .A(n3982), .Y(n3980) );
  INVX2TS U2033 ( .A(n4336), .Y(n4334) );
  INVX2TS U2034 ( .A(n4333), .Y(n4331) );
  INVX2TS U2035 ( .A(n4330), .Y(n4328) );
  INVX2TS U2036 ( .A(n4327), .Y(n4325) );
  INVX2TS U2037 ( .A(n4324), .Y(n4322) );
  INVX2TS U2038 ( .A(n4321), .Y(n4319) );
  INVX2TS U2039 ( .A(n4318), .Y(n4316) );
  INVX2TS U2040 ( .A(n4315), .Y(n4313) );
  INVX2TS U2041 ( .A(n4312), .Y(n4310) );
  INVX2TS U2042 ( .A(n4309), .Y(n4307) );
  INVX2TS U2043 ( .A(n4306), .Y(n4304) );
  INVX2TS U2044 ( .A(n4303), .Y(n4301) );
  INVX2TS U2045 ( .A(n4300), .Y(n4298) );
  INVX2TS U2046 ( .A(n4297), .Y(n4295) );
  INVX2TS U2047 ( .A(n4294), .Y(n4292) );
  INVX2TS U2048 ( .A(n4291), .Y(n4289) );
  INVX2TS U2049 ( .A(n4279), .Y(n4277) );
  INVX2TS U2050 ( .A(n4276), .Y(n4274) );
  INVX2TS U2051 ( .A(n4273), .Y(n4271) );
  INVX2TS U2052 ( .A(n4270), .Y(n4268) );
  INVX2TS U2053 ( .A(n4267), .Y(n4265) );
  INVX2TS U2054 ( .A(n4264), .Y(n4262) );
  INVX2TS U2055 ( .A(n4261), .Y(n4259) );
  INVX2TS U2056 ( .A(n4258), .Y(n4256) );
  INVX2TS U2057 ( .A(n4255), .Y(n4253) );
  INVX2TS U2058 ( .A(n4252), .Y(n4250) );
  INVX2TS U2059 ( .A(n4249), .Y(n4247) );
  INVX2TS U2060 ( .A(n4246), .Y(n4244) );
  INVX2TS U2061 ( .A(n3991), .Y(n3989) );
  CLKBUFX2TS U2062 ( .A(n4516), .Y(n4517) );
  CLKBUFX2TS U2063 ( .A(n4508), .Y(n4509) );
  CLKBUFX2TS U2064 ( .A(n4506), .Y(n4507) );
  CLKBUFX2TS U2065 ( .A(n4497), .Y(n4498) );
  CLKBUFX2TS U2066 ( .A(n4494), .Y(n4496) );
  CLKBUFX2TS U2067 ( .A(n4488), .Y(n4490) );
  CLKBUFX2TS U2068 ( .A(n4485), .Y(n4487) );
  CLKBUFX2TS U2069 ( .A(n4483), .Y(n4484) );
  CLKBUFX2TS U2070 ( .A(n4479), .Y(n4481) );
  CLKBUFX2TS U2071 ( .A(n4476), .Y(n4478) );
  CLKBUFX2TS U2072 ( .A(n4472), .Y(n4474) );
  CLKBUFX2TS U2073 ( .A(n4467), .Y(n4469) );
  CLKBUFX2TS U2074 ( .A(n4511), .Y(n4512) );
  CLKBUFX2TS U2075 ( .A(n4499), .Y(n4500) );
  CLKBUFX2TS U2076 ( .A(n4491), .Y(n4492) );
  CLKBUFX2TS U2077 ( .A(n4453), .Y(n4454) );
  CLKBUFX2TS U2078 ( .A(n4439), .Y(n4440) );
  CLKBUFX2TS U2079 ( .A(n4521), .Y(n4523) );
  CLKBUFX2TS U2080 ( .A(n4465), .Y(n4466) );
  CLKBUFX2TS U2081 ( .A(n4460), .Y(n4461) );
  CLKBUFX2TS U2082 ( .A(n4457), .Y(n4458) );
  CLKBUFX2TS U2083 ( .A(n4451), .Y(n4452) );
  CLKBUFX2TS U2084 ( .A(n4442), .Y(n4443) );
  CLKBUFX2TS U2085 ( .A(n4446), .Y(n4447) );
  INVX2TS U2086 ( .A(n4036), .Y(n4034) );
  INVX2TS U2087 ( .A(n4033), .Y(n4031) );
  INVX2TS U2088 ( .A(n4030), .Y(n4028) );
  INVX2TS U2089 ( .A(n4027), .Y(n4025) );
  INVX2TS U2090 ( .A(n4024), .Y(n4022) );
  INVX2TS U2091 ( .A(n4021), .Y(n4019) );
  CLKBUFX2TS U2092 ( .A(n4037), .Y(n4038) );
  CLKBUFX2TS U2093 ( .A(n4052), .Y(n4053) );
  CLKBUFX2TS U2094 ( .A(n4046), .Y(n4047) );
  CLKBUFX2TS U2095 ( .A(n4043), .Y(n4044) );
  CLKBUFX2TS U2096 ( .A(n4040), .Y(n4041) );
  CLKBUFX2TS U2097 ( .A(n4049), .Y(n4050) );
  CLKBUFX2TS U2098 ( .A(n4070), .Y(n4071) );
  CLKBUFX2TS U2099 ( .A(n4067), .Y(n4068) );
  CLKBUFX2TS U2100 ( .A(n4061), .Y(n4062) );
  CLKBUFX2TS U2101 ( .A(n4064), .Y(n4065) );
  CLKBUFX2TS U2102 ( .A(n4058), .Y(n4059) );
  CLKBUFX2TS U2103 ( .A(n4055), .Y(n4056) );
  INVX2TS U2104 ( .A(n3952), .Y(n3950) );
  INVX2TS U2105 ( .A(n3946), .Y(n3944) );
  INVX2TS U2106 ( .A(n3943), .Y(n3941) );
  INVX2TS U2107 ( .A(n3940), .Y(n3938) );
  INVX2TS U2108 ( .A(n3949), .Y(n3947) );
  INVX2TS U2109 ( .A(n3937), .Y(n3935) );
  INVX2TS U2110 ( .A(n4420), .Y(n4418) );
  INVX2TS U2111 ( .A(n4425), .Y(n4421) );
  INVX2TS U2112 ( .A(n4417), .Y(n4415) );
  INVX2TS U2113 ( .A(n4414), .Y(n4412) );
  INVX2TS U2114 ( .A(n4411), .Y(n4409) );
  INVX2TS U2115 ( .A(n4408), .Y(n4406) );
  INVX2TS U2116 ( .A(n4393), .Y(n4391) );
  INVX2TS U2117 ( .A(n4378), .Y(n4376) );
  INVX2TS U2118 ( .A(n4428), .Y(n4426) );
  INVX2TS U2119 ( .A(n4405), .Y(n4403) );
  INVX2TS U2120 ( .A(n4402), .Y(n4400) );
  INVX2TS U2121 ( .A(n4399), .Y(n4397) );
  INVX2TS U2122 ( .A(n4396), .Y(n4394) );
  INVX2TS U2123 ( .A(n4387), .Y(n4385) );
  INVX2TS U2124 ( .A(n4375), .Y(n4373) );
  INVX2TS U2125 ( .A(n4390), .Y(n4388) );
  INVX2TS U2126 ( .A(n4384), .Y(n4382) );
  INVX2TS U2127 ( .A(n4381), .Y(n4379) );
  INVX2TS U2128 ( .A(n4369), .Y(n4367) );
  INVX2TS U2129 ( .A(n4357), .Y(n4355) );
  INVX2TS U2130 ( .A(n4342), .Y(n4340) );
  INVX2TS U2131 ( .A(n4435), .Y(n4433) );
  INVX2TS U2132 ( .A(n4431), .Y(n4429) );
  INVX2TS U2133 ( .A(n4372), .Y(n4370) );
  INVX2TS U2134 ( .A(n4366), .Y(n4364) );
  INVX2TS U2135 ( .A(n4363), .Y(n4361) );
  INVX2TS U2136 ( .A(n4360), .Y(n4358) );
  INVX2TS U2137 ( .A(n4354), .Y(n4352) );
  INVX2TS U2138 ( .A(n4348), .Y(n4346) );
  INVX2TS U2139 ( .A(n4345), .Y(n4343) );
  INVX2TS U2140 ( .A(n4339), .Y(n4337) );
  INVX2TS U2141 ( .A(n4351), .Y(n4349) );
  CLKBUFX2TS U2142 ( .A(n4212), .Y(n4213) );
  CLKBUFX2TS U2143 ( .A(n4202), .Y(n4203) );
  CLKBUFX2TS U2144 ( .A(n4214), .Y(n4215) );
  CLKBUFX2TS U2145 ( .A(n4207), .Y(n4208) );
  CLKBUFX2TS U2146 ( .A(n4204), .Y(n4205) );
  CLKBUFX2TS U2147 ( .A(n4537), .Y(n4538) );
  CLKBUFX2TS U2148 ( .A(n4532), .Y(n4533) );
  CLKBUFX2TS U2149 ( .A(n4535), .Y(n4536) );
  CLKBUFX2TS U2150 ( .A(n4527), .Y(n4528) );
  CLKBUFX2TS U2151 ( .A(n4524), .Y(n4525) );
  INVX2TS U2152 ( .A(n4186), .Y(n4184) );
  INVX2TS U2153 ( .A(n4180), .Y(n4178) );
  INVX2TS U2154 ( .A(n4183), .Y(n4181) );
  INVX2TS U2155 ( .A(n4177), .Y(n4175) );
  INVX2TS U2156 ( .A(n4174), .Y(n4172) );
  INVX2TS U2157 ( .A(n4171), .Y(n4169) );
  INVX2TS U2158 ( .A(n4191), .Y(n4190) );
  CLKBUFX2TS U2159 ( .A(n4199), .Y(n4200) );
  CLKBUFX2TS U2160 ( .A(n4235), .Y(n4236) );
  CLKBUFX2TS U2161 ( .A(n4229), .Y(n4230) );
  CLKBUFX2TS U2162 ( .A(n4226), .Y(n4227) );
  CLKBUFX2TS U2163 ( .A(n4238), .Y(n4239) );
  CLKBUFX2TS U2164 ( .A(n4232), .Y(n4233) );
  CLKBUFX2TS U2165 ( .A(n4223), .Y(n4224) );
  CLKBUFX2TS U2166 ( .A(n4472), .Y(n4475) );
  CLKBUFX2TS U2167 ( .A(n4470), .Y(n4471) );
  CLKBUFX2TS U2168 ( .A(n4436), .Y(n4438) );
  CLKBUFX2TS U2169 ( .A(n4518), .Y(n4519) );
  CLKBUFX2TS U2170 ( .A(n4514), .Y(n4515) );
  CLKBUFX2TS U2171 ( .A(n4508), .Y(n4510) );
  CLKBUFX2TS U2172 ( .A(n4502), .Y(n4503) );
  CLKBUFX2TS U2173 ( .A(n4499), .Y(n4501) );
  CLKBUFX2TS U2174 ( .A(n4491), .Y(n4493) );
  CLKBUFX2TS U2175 ( .A(n4479), .Y(n4482) );
  CLKBUFX2TS U2176 ( .A(n4463), .Y(n4464) );
  CLKBUFX2TS U2177 ( .A(n4460), .Y(n4462) );
  CLKBUFX2TS U2178 ( .A(n4455), .Y(n4456) );
  CLKBUFX2TS U2179 ( .A(n4446), .Y(n4449) );
  CLKBUFX2TS U2180 ( .A(n4444), .Y(n4445) );
  CLKBUFX2TS U2181 ( .A(n4214), .Y(n4216) );
  CLKBUFX2TS U2182 ( .A(n4210), .Y(n4211) );
  CLKBUFX2TS U2183 ( .A(n4207), .Y(n4209) );
  CLKBUFX2TS U2184 ( .A(n4204), .Y(n4206) );
  CLKBUFX2TS U2185 ( .A(n4524), .Y(n4526) );
  CLKBUFX2TS U2186 ( .A(n4529), .Y(n4530) );
  CLKBUFX2TS U2187 ( .A(n4235), .Y(n4237) );
  CLKBUFX2TS U2188 ( .A(n4232), .Y(n4234) );
  CLKBUFX2TS U2189 ( .A(n4226), .Y(n4228) );
  CLKBUFX2TS U2190 ( .A(n4223), .Y(n4225) );
  CLKBUFX2TS U2191 ( .A(n4238), .Y(n4240) );
  CLKBUFX2TS U2192 ( .A(n4229), .Y(n4231) );
  CLKBUFX2TS U2193 ( .A(n4199), .Y(n4201) );
  CLKBUFX2TS U2194 ( .A(n4043), .Y(n4045) );
  CLKBUFX2TS U2195 ( .A(n4163), .Y(n4165) );
  CLKBUFX2TS U2196 ( .A(n4160), .Y(n4162) );
  CLKBUFX2TS U2197 ( .A(n4151), .Y(n4153) );
  CLKBUFX2TS U2198 ( .A(n4148), .Y(n4150) );
  CLKBUFX2TS U2199 ( .A(n4136), .Y(n4138) );
  CLKBUFX2TS U2200 ( .A(n4130), .Y(n4132) );
  CLKBUFX2TS U2201 ( .A(n4127), .Y(n4129) );
  CLKBUFX2TS U2202 ( .A(n4124), .Y(n4126) );
  CLKBUFX2TS U2203 ( .A(n4118), .Y(n4120) );
  CLKBUFX2TS U2204 ( .A(n4115), .Y(n4117) );
  CLKBUFX2TS U2205 ( .A(n4112), .Y(n4114) );
  CLKBUFX2TS U2206 ( .A(n4109), .Y(n4111) );
  CLKBUFX2TS U2207 ( .A(n4106), .Y(n4108) );
  CLKBUFX2TS U2208 ( .A(n4097), .Y(n4099) );
  CLKBUFX2TS U2209 ( .A(n4094), .Y(n4096) );
  CLKBUFX2TS U2210 ( .A(n4085), .Y(n4087) );
  CLKBUFX2TS U2211 ( .A(n4082), .Y(n4084) );
  CLKBUFX2TS U2212 ( .A(n4052), .Y(n4054) );
  CLKBUFX2TS U2213 ( .A(n4049), .Y(n4051) );
  CLKBUFX2TS U2214 ( .A(n4046), .Y(n4048) );
  CLKBUFX2TS U2215 ( .A(n4040), .Y(n4042) );
  CLKBUFX2TS U2216 ( .A(n4037), .Y(n4039) );
  CLKBUFX2TS U2217 ( .A(n4103), .Y(n4105) );
  CLKBUFX2TS U2218 ( .A(n4157), .Y(n4159) );
  CLKBUFX2TS U2219 ( .A(n4154), .Y(n4156) );
  CLKBUFX2TS U2220 ( .A(n4142), .Y(n4144) );
  CLKBUFX2TS U2221 ( .A(n4133), .Y(n4135) );
  CLKBUFX2TS U2222 ( .A(n4100), .Y(n4102) );
  CLKBUFX2TS U2223 ( .A(n4088), .Y(n4090) );
  CLKBUFX2TS U2224 ( .A(n4076), .Y(n4078) );
  CLKBUFX2TS U2225 ( .A(n4166), .Y(n4168) );
  CLKBUFX2TS U2226 ( .A(n4145), .Y(n4147) );
  CLKBUFX2TS U2227 ( .A(n4139), .Y(n4141) );
  CLKBUFX2TS U2228 ( .A(n4121), .Y(n4123) );
  CLKBUFX2TS U2229 ( .A(n4091), .Y(n4093) );
  CLKBUFX2TS U2230 ( .A(n4079), .Y(n4081) );
  CLKBUFX2TS U2231 ( .A(n4073), .Y(n4075) );
  CLKBUFX2TS U2232 ( .A(n4070), .Y(n4072) );
  CLKBUFX2TS U2233 ( .A(n4067), .Y(n4069) );
  CLKBUFX2TS U2234 ( .A(n4064), .Y(n4066) );
  CLKBUFX2TS U2235 ( .A(n4061), .Y(n4063) );
  CLKBUFX2TS U2236 ( .A(n4058), .Y(n4060) );
  CLKBUFX2TS U2237 ( .A(n4055), .Y(n4057) );
  INVX2TS U2238 ( .A(n3994), .Y(n3993) );
  INVX2TS U2239 ( .A(n3988), .Y(n3987) );
  INVX2TS U2240 ( .A(n3985), .Y(n3984) );
  INVX2TS U2241 ( .A(n3982), .Y(n3981) );
  INVX2TS U2242 ( .A(n3991), .Y(n3990) );
  INVX2TS U2243 ( .A(n3979), .Y(n3978) );
  INVX2TS U2244 ( .A(n4036), .Y(n4035) );
  INVX2TS U2245 ( .A(n4030), .Y(n4029) );
  INVX2TS U2246 ( .A(n4033), .Y(n4032) );
  INVX2TS U2247 ( .A(n4027), .Y(n4026) );
  INVX2TS U2248 ( .A(n4024), .Y(n4023) );
  INVX2TS U2249 ( .A(n4021), .Y(n4020) );
  INVX2TS U2250 ( .A(n3997), .Y(n3995) );
  INVX2TS U2251 ( .A(n4000), .Y(n3998) );
  INVX2TS U2252 ( .A(n4015), .Y(n4013) );
  INVX2TS U2253 ( .A(n4012), .Y(n4010) );
  INVX2TS U2254 ( .A(n4006), .Y(n4004) );
  INVX2TS U2255 ( .A(n4003), .Y(n4001) );
  INVX2TS U2256 ( .A(n4018), .Y(n4016) );
  INVX2TS U2257 ( .A(n4009), .Y(n4007) );
  INVX2TS U2258 ( .A(n4194), .Y(n4192) );
  INVX2TS U2259 ( .A(n3973), .Y(n3971) );
  INVX2TS U2260 ( .A(n3967), .Y(n3965) );
  INVX2TS U2261 ( .A(n3964), .Y(n3962) );
  INVX2TS U2262 ( .A(n3976), .Y(n3974) );
  INVX2TS U2263 ( .A(n3970), .Y(n3968) );
  INVX2TS U2264 ( .A(n3961), .Y(n3959) );
  INVX2TS U2265 ( .A(n3955), .Y(n3953) );
  INVX2TS U2266 ( .A(n3958), .Y(n3956) );
  INVX2TS U2267 ( .A(n4384), .Y(n4383) );
  INVX2TS U2268 ( .A(n4381), .Y(n4380) );
  INVX2TS U2269 ( .A(n4378), .Y(n4377) );
  INVX2TS U2270 ( .A(n4339), .Y(n4338) );
  INVX2TS U2271 ( .A(n4435), .Y(n4434) );
  INVX2TS U2272 ( .A(n4431), .Y(n4430) );
  INVX2TS U2273 ( .A(n4428), .Y(n4427) );
  INVX2TS U2274 ( .A(n4425), .Y(n4422) );
  INVX2TS U2275 ( .A(n4420), .Y(n4419) );
  INVX2TS U2276 ( .A(n4417), .Y(n4416) );
  INVX2TS U2277 ( .A(n4414), .Y(n4413) );
  INVX2TS U2278 ( .A(n4411), .Y(n4410) );
  INVX2TS U2279 ( .A(n4408), .Y(n4407) );
  INVX2TS U2280 ( .A(n4405), .Y(n4404) );
  INVX2TS U2281 ( .A(n4402), .Y(n4401) );
  INVX2TS U2282 ( .A(n4399), .Y(n4398) );
  INVX2TS U2283 ( .A(n4396), .Y(n4395) );
  INVX2TS U2284 ( .A(n4393), .Y(n4392) );
  INVX2TS U2285 ( .A(n4390), .Y(n4389) );
  INVX2TS U2286 ( .A(n4387), .Y(n4386) );
  INVX2TS U2287 ( .A(n4375), .Y(n4374) );
  INVX2TS U2288 ( .A(n4372), .Y(n4371) );
  INVX2TS U2289 ( .A(n4369), .Y(n4368) );
  INVX2TS U2290 ( .A(n4366), .Y(n4365) );
  INVX2TS U2291 ( .A(n4363), .Y(n4362) );
  INVX2TS U2292 ( .A(n4360), .Y(n4359) );
  INVX2TS U2293 ( .A(n4357), .Y(n4356) );
  INVX2TS U2294 ( .A(n4354), .Y(n4353) );
  INVX2TS U2295 ( .A(n4351), .Y(n4350) );
  INVX2TS U2296 ( .A(n4348), .Y(n4347) );
  INVX2TS U2297 ( .A(n4345), .Y(n4344) );
  INVX2TS U2298 ( .A(n4342), .Y(n4341) );
  INVX2TS U2299 ( .A(n4194), .Y(n4193) );
  INVX2TS U2300 ( .A(n3973), .Y(n3972) );
  INVX2TS U2301 ( .A(n3970), .Y(n3969) );
  INVX2TS U2302 ( .A(n3964), .Y(n3963) );
  INVX2TS U2303 ( .A(n3961), .Y(n3960) );
  INVX2TS U2304 ( .A(n3955), .Y(n3954) );
  INVX2TS U2305 ( .A(n3976), .Y(n3975) );
  INVX2TS U2306 ( .A(n3967), .Y(n3966) );
  INVX2TS U2307 ( .A(n3958), .Y(n3957) );
  INVX2TS U2308 ( .A(n3997), .Y(n3996) );
  INVX2TS U2309 ( .A(n4000), .Y(n3999) );
  INVX2TS U2310 ( .A(n4015), .Y(n4014) );
  INVX2TS U2311 ( .A(n4009), .Y(n4008) );
  INVX2TS U2312 ( .A(n4006), .Y(n4005) );
  INVX2TS U2313 ( .A(n4018), .Y(n4017) );
  INVX2TS U2314 ( .A(n4012), .Y(n4011) );
  INVX2TS U2315 ( .A(n4003), .Y(n4002) );
  INVX2TS U2316 ( .A(n4330), .Y(n4329) );
  INVX2TS U2317 ( .A(n4327), .Y(n4326) );
  INVX2TS U2318 ( .A(n4324), .Y(n4323) );
  INVX2TS U2319 ( .A(n4321), .Y(n4320) );
  INVX2TS U2320 ( .A(n4318), .Y(n4317) );
  INVX2TS U2321 ( .A(n4315), .Y(n4314) );
  INVX2TS U2322 ( .A(n4312), .Y(n4311) );
  INVX2TS U2323 ( .A(n4309), .Y(n4308) );
  INVX2TS U2324 ( .A(n4306), .Y(n4305) );
  INVX2TS U2325 ( .A(n4303), .Y(n4302) );
  INVX2TS U2326 ( .A(n4300), .Y(n4299) );
  INVX2TS U2327 ( .A(n4297), .Y(n4296) );
  INVX2TS U2328 ( .A(n4294), .Y(n4293) );
  INVX2TS U2329 ( .A(n4291), .Y(n4290) );
  INVX2TS U2330 ( .A(n4288), .Y(n4287) );
  INVX2TS U2331 ( .A(n4285), .Y(n4284) );
  INVX2TS U2332 ( .A(n4282), .Y(n4281) );
  INVX2TS U2333 ( .A(n4279), .Y(n4278) );
  INVX2TS U2334 ( .A(n4273), .Y(n4272) );
  INVX2TS U2335 ( .A(n4261), .Y(n4260) );
  INVX2TS U2336 ( .A(n4246), .Y(n4245) );
  INVX2TS U2337 ( .A(n4336), .Y(n4335) );
  INVX2TS U2338 ( .A(n4333), .Y(n4332) );
  INVX2TS U2339 ( .A(n4276), .Y(n4275) );
  INVX2TS U2340 ( .A(n4270), .Y(n4269) );
  INVX2TS U2341 ( .A(n4267), .Y(n4266) );
  INVX2TS U2342 ( .A(n4264), .Y(n4263) );
  INVX2TS U2343 ( .A(n4258), .Y(n4257) );
  INVX2TS U2344 ( .A(n4252), .Y(n4251) );
  INVX2TS U2345 ( .A(n4249), .Y(n4248) );
  INVX2TS U2346 ( .A(n4243), .Y(n4242) );
  INVX2TS U2347 ( .A(n4255), .Y(n4254) );
  INVX2TS U2348 ( .A(n3949), .Y(n3948) );
  INVX2TS U2349 ( .A(n3937), .Y(n3936) );
  INVX2TS U2350 ( .A(n3952), .Y(n3951) );
  INVX2TS U2351 ( .A(n3946), .Y(n3945) );
  INVX2TS U2352 ( .A(n3943), .Y(n3942) );
  INVX2TS U2353 ( .A(n3940), .Y(n3939) );
  INVX2TS U2354 ( .A(n4186), .Y(n4185) );
  INVX2TS U2355 ( .A(n4183), .Y(n4182) );
  INVX2TS U2356 ( .A(n4177), .Y(n4176) );
  INVX2TS U2357 ( .A(n4180), .Y(n4179) );
  INVX2TS U2358 ( .A(n4174), .Y(n4173) );
  INVX2TS U2359 ( .A(n4171), .Y(n4170) );
  INVX2TS U2360 ( .A(n1938), .Y(n761) );
  INVX2TS U2361 ( .A(n924), .Y(n717) );
  INVX2TS U2362 ( .A(n2896), .Y(n716) );
  INVX2TS U2363 ( .A(n2032), .Y(n720) );
  AOI21X1TS U2364 ( .A0(n437), .A1(n925), .B0(n1985), .Y(n2010) );
  AOI222XLTS U2365 ( .A0(n4200), .A1(n3375), .B0(n4188), .B1(n3360), .C0(n4192), .C1(n3409), .Y(n1758) );
  AOI222XLTS U2366 ( .A0(n4187), .A1(n3457), .B0(n4193), .B1(n3436), .C0(n4201), .C1(n3419), .Y(n1755) );
  NOR3X1TS U2367 ( .A(n2449), .B(n166), .C(n2391), .Y(n2394) );
  OAI21X1TS U2368 ( .A0(n456), .A1(n1842), .B0(n1843), .Y(n1100) );
  OAI21X1TS U2369 ( .A0(n759), .A1(n745), .B0(n915), .Y(n1843) );
  XNOR2X1TS U2370 ( .A(n4), .B(n2892), .Y(n1086) );
  NOR2X1TS U2371 ( .A(n2391), .B(n2449), .Y(n2892) );
  NOR2X1TS U2372 ( .A(n959), .B(n166), .Y(n1985) );
  NOR2X1TS U2373 ( .A(n1915), .B(n973), .Y(n1844) );
  OAI2BB2XLTS U2374 ( .B0(n1985), .B1(n471), .A0N(n1832), .A1N(n1985), .Y(
        n2011) );
  OAI22X1TS U2375 ( .A0(n1090), .A1(n1087), .B0(n1088), .B1(n113), .Y(n2886)
         );
  INVX2TS U2376 ( .A(n170), .Y(n915) );
  XOR2X1TS U2377 ( .A(n1086), .B(n137), .Y(n2891) );
  XOR2X1TS U2378 ( .A(n2012), .B(n2013), .Y(n1962) );
  NAND2X1TS U2379 ( .A(n4), .B(n2014), .Y(n2012) );
  XOR2X1TS U2380 ( .A(n3), .B(n957), .Y(n2013) );
  OAI22X1TS U2381 ( .A0(n1094), .A1(n2890), .B0(n2897), .B1(n2392), .Y(n2894)
         );
  AOI32X1TS U2382 ( .A0(n1096), .A1(n715), .A2(n2896), .B0(n2897), .B1(n2392), 
        .Y(n2895) );
  AOI211XLTS U2383 ( .A0(n1094), .A1(n2890), .B0(n716), .C0(n2449), .Y(n2893)
         );
  OAI221XLTS U2384 ( .A0(n541), .A1(n149), .B0(n3328), .B1(n911), .C0(n1760), 
        .Y(n2572) );
  AOI222XLTS U2385 ( .A0(n4192), .A1(n3270), .B0(n4188), .B1(n3280), .C0(n4201), .C1(n3318), .Y(n1760) );
  OAI221XLTS U2386 ( .A0(n466), .A1(n148), .B0(n158), .B1(n708), .C0(n1752), 
        .Y(n2575) );
  AOI222XLTS U2387 ( .A0(n4200), .A1(n3494), .B0(n4193), .B1(n3472), .C0(n4187), .C1(n3524), .Y(n1752) );
  OAI221XLTS U2388 ( .A0(n459), .A1(n134), .B0(n3593), .B1(n563), .C0(n1889), 
        .Y(n2524) );
  AOI222XLTS U2389 ( .A0(n4007), .A1(n3538), .B0(n3966), .B1(n3545), .C0(n4231), .C1(n3586), .Y(n1889) );
  OAI221XLTS U2390 ( .A0(n463), .A1(n149), .B0(n3100), .B1(n707), .C0(n1747), 
        .Y(n2577) );
  AOI222XLTS U2391 ( .A0(n4200), .A1(n3652), .B0(n4188), .B1(n3615), .C0(n4192), .C1(n3798), .Y(n1747) );
  OAI221XLTS U2392 ( .A0(n461), .A1(n148), .B0(n3595), .B1(n660), .C0(n1749), 
        .Y(n2576) );
  AOI222XLTS U2393 ( .A0(n4187), .A1(n3544), .B0(n4193), .B1(n3547), .C0(n4201), .C1(n3585), .Y(n1749) );
  OAI221XLTS U2394 ( .A0(n3672), .A1(n148), .B0(n3751), .B1(n653), .C0(n1745), 
        .Y(n2578) );
  AOI222XLTS U2395 ( .A0(n4187), .A1(n3687), .B0(n4193), .B1(n3695), .C0(n4201), .C1(n3731), .Y(n1745) );
  INVX2TS U2396 ( .A(n1961), .Y(n735) );
  NOR2X1TS U2397 ( .A(n1841), .B(n171), .Y(n1831) );
  NOR2X1TS U2398 ( .A(n748), .B(n471), .Y(n1774) );
  INVX2TS U2399 ( .A(n1841), .Y(n931) );
  INVX2TS U2400 ( .A(n2018), .Y(n3097) );
  NAND4BX1TS U2401 ( .AN(n152), .B(n2382), .C(n2025), .D(n2023), .Y(n2018) );
  AND3X2TS U2402 ( .A(n2026), .B(n2024), .C(n2027), .Y(n2382) );
  NOR2BX1TS U2403 ( .AN(n1860), .B(n456), .Y(n1122) );
  NOR2BX1TS U2404 ( .AN(n1860), .B(n106), .Y(n1155) );
  NOR2X1TS U2405 ( .A(n2023), .B(n152), .Y(n2054) );
  NOR2X1TS U2406 ( .A(n2024), .B(n153), .Y(n2040) );
  NOR2X1TS U2407 ( .A(n2026), .B(n154), .Y(n2039) );
  INVX2TS U2408 ( .A(n2038), .Y(n651) );
  AOI221X1TS U2409 ( .A0(n4188), .A1(n3080), .B0(writeIn_SOUTH), .B1(n3063), 
        .C0(n2041), .Y(n2038) );
  NOR2X1TS U2410 ( .A(n1870), .B(n170), .Y(n1860) );
  INVX2TS U2411 ( .A(writeIn_EAST), .Y(n4194) );
  INVX2TS U2412 ( .A(n1870), .Y(n929) );
  OR2X2TS U2413 ( .A(n2025), .B(n154), .Y(n762) );
  OAI221XLTS U2414 ( .A0(n4198), .A1(n2025), .B0(n4191), .B1(n2026), .C0(n2027), .Y(n2021) );
  OAI22X1TS U2415 ( .A0(n811), .A1(n1048), .B0(n623), .B1(n2118), .Y(n2380) );
  OAI22X1TS U2416 ( .A0(n801), .A1(n1048), .B0(n622), .B1(n1033), .Y(n2374) );
  OAI22X1TS U2417 ( .A0(n800), .A1(n1048), .B0(n621), .B1(n1034), .Y(n2368) );
  OAI22X1TS U2418 ( .A0(n799), .A1(n1047), .B0(n620), .B1(n1033), .Y(n2362) );
  OAI22X1TS U2419 ( .A0(n798), .A1(n1036), .B0(n619), .B1(n1021), .Y(n2356) );
  OAI22X1TS U2420 ( .A0(n797), .A1(n1036), .B0(n618), .B1(n1021), .Y(n2350) );
  OAI22X1TS U2421 ( .A0(n796), .A1(n1036), .B0(n617), .B1(n1021), .Y(n2344) );
  OAI22X1TS U2422 ( .A0(n795), .A1(n1036), .B0(n616), .B1(n1021), .Y(n2338) );
  OAI22X1TS U2423 ( .A0(n794), .A1(n1037), .B0(n615), .B1(n1022), .Y(n2332) );
  OAI22X1TS U2424 ( .A0(n793), .A1(n1037), .B0(n614), .B1(n1022), .Y(n2326) );
  OAI22X1TS U2425 ( .A0(n792), .A1(n1037), .B0(n613), .B1(n1022), .Y(n2320) );
  OAI22X1TS U2426 ( .A0(n791), .A1(n1037), .B0(n612), .B1(n1022), .Y(n2314) );
  OAI22X1TS U2427 ( .A0(n790), .A1(n1038), .B0(n611), .B1(n1023), .Y(n2308) );
  OAI22X1TS U2428 ( .A0(n789), .A1(n1038), .B0(n610), .B1(n1023), .Y(n2302) );
  OAI22X1TS U2429 ( .A0(n788), .A1(n1038), .B0(n609), .B1(n1023), .Y(n2296) );
  OAI22X1TS U2430 ( .A0(n810), .A1(n1038), .B0(n608), .B1(n1023), .Y(n2290) );
  OAI22X1TS U2431 ( .A0(n809), .A1(n1039), .B0(n935), .B1(n1033), .Y(n2284) );
  OAI22X1TS U2432 ( .A0(n787), .A1(n1039), .B0(n936), .B1(n1032), .Y(n2278) );
  OAI22X1TS U2433 ( .A0(n786), .A1(n1039), .B0(n937), .B1(n1031), .Y(n2272) );
  OAI22X1TS U2434 ( .A0(n785), .A1(n1039), .B0(n607), .B1(n1032), .Y(n2266) );
  OAI22X1TS U2435 ( .A0(n808), .A1(n1047), .B0(n606), .B1(n1024), .Y(n2260) );
  OAI22X1TS U2436 ( .A0(n784), .A1(n1046), .B0(n605), .B1(n1024), .Y(n2254) );
  OAI22X1TS U2437 ( .A0(n783), .A1(n1045), .B0(n604), .B1(n1024), .Y(n2248) );
  OAI22X1TS U2438 ( .A0(n782), .A1(n1046), .B0(n603), .B1(n1024), .Y(n2242) );
  OAI22X1TS U2439 ( .A0(n781), .A1(n1040), .B0(n602), .B1(n1025), .Y(n2236) );
  OAI22X1TS U2440 ( .A0(n780), .A1(n1040), .B0(n601), .B1(n1025), .Y(n2230) );
  OAI22X1TS U2441 ( .A0(n779), .A1(n1040), .B0(n600), .B1(n1025), .Y(n2224) );
  OAI22X1TS U2442 ( .A0(n778), .A1(n1040), .B0(n599), .B1(n1025), .Y(n2218) );
  OAI22X1TS U2443 ( .A0(n777), .A1(n1041), .B0(n598), .B1(n1026), .Y(n2212) );
  OAI22X1TS U2444 ( .A0(n776), .A1(n1041), .B0(n597), .B1(n1026), .Y(n2206) );
  OAI22X1TS U2445 ( .A0(n807), .A1(n1041), .B0(n596), .B1(n1026), .Y(n2200) );
  OAI22X1TS U2446 ( .A0(n775), .A1(n1041), .B0(n934), .B1(n1026), .Y(n2194) );
  OAI22X1TS U2447 ( .A0(n899), .A1(n1042), .B0(n663), .B1(n1027), .Y(n2188) );
  OAI22X1TS U2448 ( .A0(n898), .A1(n1042), .B0(n662), .B1(n1027), .Y(n2182) );
  OAI22X1TS U2449 ( .A0(n896), .A1(n1042), .B0(n661), .B1(n1027), .Y(n2170) );
  OAI22X1TS U2450 ( .A0(n895), .A1(n1043), .B0(n658), .B1(n1029), .Y(n2164) );
  OAI22X1TS U2451 ( .A0(n806), .A1(n1043), .B0(n627), .B1(n1029), .Y(n2152) );
  OAI22X1TS U2452 ( .A0(n774), .A1(n1043), .B0(n639), .B1(n1029), .Y(n2146) );
  OAI22X1TS U2453 ( .A0(n805), .A1(n1044), .B0(n626), .B1(n1030), .Y(n2140) );
  OAI22X1TS U2454 ( .A0(n804), .A1(n1044), .B0(n625), .B1(n1030), .Y(n2134) );
  OAI22X1TS U2455 ( .A0(n803), .A1(n1044), .B0(n624), .B1(n1030), .Y(n2128) );
  OAI22X1TS U2456 ( .A0(n802), .A1(n1044), .B0(n638), .B1(n1030), .Y(n2116) );
  OAI22X1TS U2457 ( .A0(n897), .A1(n1042), .B0(n659), .B1(n1027), .Y(n2176) );
  OAI22X1TS U2458 ( .A0(n894), .A1(n1043), .B0(n657), .B1(n1029), .Y(n2158) );
  OAI22X1TS U2459 ( .A0(n434), .A1(n2023), .B0(n438), .B1(n2024), .Y(n2022) );
  NOR2X1TS U2460 ( .A(n2034), .B(n139), .Y(n2119) );
  NOR2X1TS U2461 ( .A(n2036), .B(n138), .Y(n2120) );
  NOR2X1TS U2462 ( .A(n2049), .B(n138), .Y(n2115) );
  NOR2X1TS U2463 ( .A(n2033), .B(n139), .Y(n2114) );
  NOR2X1TS U2464 ( .A(n2035), .B(n138), .Y(n2121) );
  NOR2X1TS U2465 ( .A(n2027), .B(n153), .Y(n2123) );
  INVX2TS U2466 ( .A(requesterAddressIn_WEST[4]), .Y(n4033) );
  INVX2TS U2467 ( .A(requesterAddressIn_WEST[5]), .Y(n4036) );
  INVX2TS U2468 ( .A(requesterAddressIn_WEST[3]), .Y(n4030) );
  INVX2TS U2469 ( .A(requesterAddressIn_WEST[2]), .Y(n4027) );
  INVX2TS U2470 ( .A(requesterAddressIn_WEST[1]), .Y(n4024) );
  INVX2TS U2471 ( .A(requesterAddressIn_WEST[0]), .Y(n4021) );
  INVX2TS U2472 ( .A(requesterAddressIn_EAST[5]), .Y(n4186) );
  INVX2TS U2473 ( .A(requesterAddressIn_EAST[4]), .Y(n4183) );
  INVX2TS U2474 ( .A(requesterAddressIn_EAST[3]), .Y(n4180) );
  INVX2TS U2475 ( .A(requesterAddressIn_EAST[2]), .Y(n4177) );
  INVX2TS U2476 ( .A(requesterAddressIn_EAST[1]), .Y(n4174) );
  INVX2TS U2477 ( .A(requesterAddressIn_EAST[0]), .Y(n4171) );
  INVX2TS U2478 ( .A(destinationAddressIn_WEST[5]), .Y(n3994) );
  INVX2TS U2479 ( .A(destinationAddressIn_WEST[3]), .Y(n3988) );
  INVX2TS U2480 ( .A(destinationAddressIn_WEST[2]), .Y(n3985) );
  INVX2TS U2481 ( .A(destinationAddressIn_WEST[1]), .Y(n3982) );
  INVX2TS U2482 ( .A(destinationAddressIn_WEST[0]), .Y(n3979) );
  INVX2TS U2483 ( .A(dataIn_WEST[30]), .Y(n4333) );
  INVX2TS U2484 ( .A(dataIn_WEST[28]), .Y(n4327) );
  INVX2TS U2485 ( .A(dataIn_WEST[27]), .Y(n4324) );
  INVX2TS U2486 ( .A(dataIn_WEST[26]), .Y(n4321) );
  INVX2TS U2487 ( .A(dataIn_WEST[25]), .Y(n4318) );
  INVX2TS U2488 ( .A(dataIn_WEST[24]), .Y(n4315) );
  INVX2TS U2489 ( .A(dataIn_WEST[23]), .Y(n4312) );
  INVX2TS U2490 ( .A(dataIn_WEST[18]), .Y(n4297) );
  INVX2TS U2491 ( .A(dataIn_WEST[13]), .Y(n4282) );
  INVX2TS U2492 ( .A(dataIn_WEST[9]), .Y(n4270) );
  INVX2TS U2493 ( .A(dataIn_WEST[7]), .Y(n4264) );
  INVX2TS U2494 ( .A(dataIn_WEST[5]), .Y(n4258) );
  INVX2TS U2495 ( .A(dataIn_WEST[4]), .Y(n4255) );
  INVX2TS U2496 ( .A(dataIn_WEST[2]), .Y(n4249) );
  INVX2TS U2497 ( .A(dataIn_WEST[31]), .Y(n4336) );
  INVX2TS U2498 ( .A(dataIn_WEST[29]), .Y(n4330) );
  INVX2TS U2499 ( .A(dataIn_WEST[22]), .Y(n4309) );
  INVX2TS U2500 ( .A(dataIn_WEST[21]), .Y(n4306) );
  INVX2TS U2501 ( .A(dataIn_WEST[20]), .Y(n4303) );
  INVX2TS U2502 ( .A(dataIn_WEST[19]), .Y(n4300) );
  INVX2TS U2503 ( .A(dataIn_WEST[16]), .Y(n4291) );
  INVX2TS U2504 ( .A(dataIn_WEST[12]), .Y(n4279) );
  INVX2TS U2505 ( .A(dataIn_WEST[11]), .Y(n4276) );
  INVX2TS U2506 ( .A(dataIn_WEST[10]), .Y(n4273) );
  INVX2TS U2507 ( .A(dataIn_WEST[8]), .Y(n4267) );
  INVX2TS U2508 ( .A(dataIn_WEST[6]), .Y(n4261) );
  INVX2TS U2509 ( .A(dataIn_WEST[1]), .Y(n4246) );
  INVX2TS U2510 ( .A(dataIn_WEST[0]), .Y(n4243) );
  INVX2TS U2511 ( .A(dataIn_WEST[17]), .Y(n4294) );
  INVX2TS U2512 ( .A(dataIn_WEST[15]), .Y(n4288) );
  INVX2TS U2513 ( .A(dataIn_WEST[14]), .Y(n4285) );
  INVX2TS U2514 ( .A(dataIn_WEST[3]), .Y(n4252) );
  INVX2TS U2515 ( .A(destinationAddressIn_WEST[4]), .Y(n3991) );
  INVX2TS U2516 ( .A(destinationAddressIn_EAST[5]), .Y(n3952) );
  INVX2TS U2517 ( .A(destinationAddressIn_EAST[3]), .Y(n3946) );
  INVX2TS U2518 ( .A(destinationAddressIn_EAST[2]), .Y(n3943) );
  INVX2TS U2519 ( .A(destinationAddressIn_EAST[1]), .Y(n3940) );
  INVX2TS U2520 ( .A(destinationAddressIn_EAST[0]), .Y(n3937) );
  INVX2TS U2521 ( .A(destinationAddressIn_EAST[4]), .Y(n3949) );
  NAND2X1TS U2522 ( .A(n169), .B(n550), .Y(n2118) );
  INVX2TS U2523 ( .A(readIn_WEST), .Y(n4191) );
  INVX2TS U2524 ( .A(destinationAddressIn_EAST[12]), .Y(n3973) );
  INVX2TS U2525 ( .A(destinationAddressIn_EAST[11]), .Y(n3970) );
  INVX2TS U2526 ( .A(destinationAddressIn_EAST[9]), .Y(n3964) );
  INVX2TS U2527 ( .A(destinationAddressIn_EAST[13]), .Y(n3976) );
  INVX2TS U2528 ( .A(destinationAddressIn_EAST[10]), .Y(n3967) );
  INVX2TS U2529 ( .A(destinationAddressIn_EAST[8]), .Y(n3961) );
  INVX2TS U2530 ( .A(destinationAddressIn_EAST[6]), .Y(n3955) );
  INVX2TS U2531 ( .A(destinationAddressIn_EAST[7]), .Y(n3958) );
  INVX2TS U2532 ( .A(dataIn_EAST[15]), .Y(n4384) );
  INVX2TS U2533 ( .A(dataIn_EAST[14]), .Y(n4381) );
  INVX2TS U2534 ( .A(dataIn_EAST[13]), .Y(n4378) );
  INVX2TS U2535 ( .A(dataIn_EAST[0]), .Y(n4339) );
  INVX2TS U2536 ( .A(dataIn_EAST[31]), .Y(n4435) );
  INVX2TS U2537 ( .A(dataIn_EAST[30]), .Y(n4431) );
  INVX2TS U2538 ( .A(dataIn_EAST[29]), .Y(n4428) );
  INVX2TS U2539 ( .A(dataIn_EAST[28]), .Y(n4425) );
  INVX2TS U2540 ( .A(dataIn_EAST[27]), .Y(n4420) );
  INVX2TS U2541 ( .A(dataIn_EAST[26]), .Y(n4417) );
  INVX2TS U2542 ( .A(dataIn_EAST[25]), .Y(n4414) );
  INVX2TS U2543 ( .A(dataIn_EAST[24]), .Y(n4411) );
  INVX2TS U2544 ( .A(dataIn_EAST[23]), .Y(n4408) );
  INVX2TS U2545 ( .A(dataIn_EAST[22]), .Y(n4405) );
  INVX2TS U2546 ( .A(dataIn_EAST[21]), .Y(n4402) );
  INVX2TS U2547 ( .A(dataIn_EAST[20]), .Y(n4399) );
  INVX2TS U2548 ( .A(dataIn_EAST[19]), .Y(n4396) );
  INVX2TS U2549 ( .A(dataIn_EAST[18]), .Y(n4393) );
  INVX2TS U2550 ( .A(dataIn_EAST[17]), .Y(n4390) );
  INVX2TS U2551 ( .A(dataIn_EAST[16]), .Y(n4387) );
  INVX2TS U2552 ( .A(dataIn_EAST[12]), .Y(n4375) );
  INVX2TS U2553 ( .A(dataIn_EAST[11]), .Y(n4372) );
  INVX2TS U2554 ( .A(dataIn_EAST[10]), .Y(n4369) );
  INVX2TS U2555 ( .A(dataIn_EAST[9]), .Y(n4366) );
  INVX2TS U2556 ( .A(dataIn_EAST[8]), .Y(n4363) );
  INVX2TS U2557 ( .A(dataIn_EAST[7]), .Y(n4360) );
  INVX2TS U2558 ( .A(dataIn_EAST[6]), .Y(n4357) );
  INVX2TS U2559 ( .A(dataIn_EAST[5]), .Y(n4354) );
  INVX2TS U2560 ( .A(dataIn_EAST[3]), .Y(n4348) );
  INVX2TS U2561 ( .A(dataIn_EAST[2]), .Y(n4345) );
  INVX2TS U2562 ( .A(dataIn_EAST[1]), .Y(n4342) );
  INVX2TS U2563 ( .A(dataIn_EAST[4]), .Y(n4351) );
  INVX2TS U2564 ( .A(destinationAddressIn_WEST[6]), .Y(n3997) );
  INVX2TS U2565 ( .A(destinationAddressIn_WEST[7]), .Y(n4000) );
  INVX2TS U2566 ( .A(destinationAddressIn_WEST[12]), .Y(n4015) );
  INVX2TS U2567 ( .A(destinationAddressIn_WEST[11]), .Y(n4012) );
  INVX2TS U2568 ( .A(destinationAddressIn_WEST[9]), .Y(n4006) );
  INVX2TS U2569 ( .A(destinationAddressIn_WEST[8]), .Y(n4003) );
  INVX2TS U2570 ( .A(destinationAddressIn_WEST[13]), .Y(n4018) );
  INVX2TS U2571 ( .A(destinationAddressIn_WEST[10]), .Y(n4009) );
  CLKBUFX2TS U2572 ( .A(dataIn_SOUTH[15]), .Y(n4476) );
  CLKBUFX2TS U2573 ( .A(dataIn_SOUTH[14]), .Y(n4472) );
  CLKBUFX2TS U2574 ( .A(dataIn_SOUTH[13]), .Y(n4470) );
  CLKBUFX2TS U2575 ( .A(requesterAddressIn_SOUTH[4]), .Y(n4535) );
  CLKBUFX2TS U2576 ( .A(requesterAddressIn_SOUTH[1]), .Y(n4527) );
  CLKBUFX2TS U2577 ( .A(requesterAddressIn_SOUTH[0]), .Y(n4524) );
  CLKBUFX2TS U2578 ( .A(requesterAddressIn_SOUTH[5]), .Y(n4537) );
  CLKBUFX2TS U2579 ( .A(requesterAddressIn_SOUTH[3]), .Y(n4532) );
  CLKBUFX2TS U2580 ( .A(requesterAddressIn_SOUTH[2]), .Y(n4529) );
  CLKBUFX2TS U2581 ( .A(destinationAddressIn_SOUTH[0]), .Y(n4202) );
  CLKBUFX2TS U2582 ( .A(dataIn_SOUTH[0]), .Y(n4436) );
  CLKBUFX2TS U2583 ( .A(destinationAddressIn_SOUTH[5]), .Y(n4214) );
  CLKBUFX2TS U2584 ( .A(destinationAddressIn_SOUTH[3]), .Y(n4210) );
  CLKBUFX2TS U2585 ( .A(destinationAddressIn_SOUTH[2]), .Y(n4207) );
  CLKBUFX2TS U2586 ( .A(destinationAddressIn_SOUTH[1]), .Y(n4204) );
  CLKBUFX2TS U2587 ( .A(dataIn_SOUTH[31]), .Y(n4521) );
  CLKBUFX2TS U2588 ( .A(dataIn_SOUTH[30]), .Y(n4518) );
  CLKBUFX2TS U2589 ( .A(dataIn_SOUTH[29]), .Y(n4516) );
  CLKBUFX2TS U2590 ( .A(dataIn_SOUTH[28]), .Y(n4514) );
  CLKBUFX2TS U2591 ( .A(dataIn_SOUTH[27]), .Y(n4511) );
  CLKBUFX2TS U2592 ( .A(dataIn_SOUTH[26]), .Y(n4508) );
  CLKBUFX2TS U2593 ( .A(dataIn_SOUTH[25]), .Y(n4506) );
  CLKBUFX2TS U2594 ( .A(dataIn_SOUTH[24]), .Y(n4502) );
  CLKBUFX2TS U2595 ( .A(dataIn_SOUTH[23]), .Y(n4499) );
  CLKBUFX2TS U2596 ( .A(dataIn_SOUTH[22]), .Y(n4497) );
  CLKBUFX2TS U2597 ( .A(dataIn_SOUTH[21]), .Y(n4494) );
  CLKBUFX2TS U2598 ( .A(dataIn_SOUTH[20]), .Y(n4491) );
  CLKBUFX2TS U2599 ( .A(dataIn_SOUTH[19]), .Y(n4488) );
  CLKBUFX2TS U2600 ( .A(dataIn_SOUTH[18]), .Y(n4485) );
  CLKBUFX2TS U2601 ( .A(dataIn_SOUTH[17]), .Y(n4483) );
  CLKBUFX2TS U2602 ( .A(dataIn_SOUTH[16]), .Y(n4479) );
  CLKBUFX2TS U2603 ( .A(dataIn_SOUTH[12]), .Y(n4467) );
  CLKBUFX2TS U2604 ( .A(dataIn_SOUTH[11]), .Y(n4465) );
  CLKBUFX2TS U2605 ( .A(dataIn_SOUTH[10]), .Y(n4463) );
  CLKBUFX2TS U2606 ( .A(dataIn_SOUTH[9]), .Y(n4460) );
  CLKBUFX2TS U2607 ( .A(dataIn_SOUTH[8]), .Y(n4457) );
  CLKBUFX2TS U2608 ( .A(dataIn_SOUTH[7]), .Y(n4455) );
  CLKBUFX2TS U2609 ( .A(dataIn_SOUTH[6]), .Y(n4453) );
  CLKBUFX2TS U2610 ( .A(dataIn_SOUTH[5]), .Y(n4451) );
  CLKBUFX2TS U2611 ( .A(dataIn_SOUTH[3]), .Y(n4444) );
  CLKBUFX2TS U2612 ( .A(dataIn_SOUTH[2]), .Y(n4442) );
  CLKBUFX2TS U2613 ( .A(dataIn_SOUTH[1]), .Y(n4439) );
  CLKBUFX2TS U2614 ( .A(destinationAddressIn_SOUTH[4]), .Y(n4212) );
  CLKBUFX2TS U2615 ( .A(dataIn_SOUTH[4]), .Y(n4446) );
  CLKBUFX2TS U2616 ( .A(writeIn_SOUTH), .Y(n4199) );
  CLKBUFX2TS U2617 ( .A(destinationAddressIn_SOUTH[12]), .Y(n4235) );
  CLKBUFX2TS U2618 ( .A(destinationAddressIn_SOUTH[11]), .Y(n4232) );
  CLKBUFX2TS U2619 ( .A(destinationAddressIn_SOUTH[9]), .Y(n4226) );
  CLKBUFX2TS U2620 ( .A(destinationAddressIn_SOUTH[13]), .Y(n4238) );
  CLKBUFX2TS U2621 ( .A(destinationAddressIn_SOUTH[10]), .Y(n4229) );
  CLKBUFX2TS U2622 ( .A(destinationAddressIn_SOUTH[8]), .Y(n4223) );
  CLKBUFX2TS U2623 ( .A(dataIn_NORTH[15]), .Y(n4118) );
  CLKBUFX2TS U2624 ( .A(dataIn_NORTH[14]), .Y(n4115) );
  CLKBUFX2TS U2625 ( .A(dataIn_NORTH[13]), .Y(n4112) );
  CLKBUFX2TS U2626 ( .A(requesterAddressIn_NORTH[5]), .Y(n4070) );
  CLKBUFX2TS U2627 ( .A(requesterAddressIn_NORTH[4]), .Y(n4067) );
  CLKBUFX2TS U2628 ( .A(requesterAddressIn_NORTH[3]), .Y(n4064) );
  CLKBUFX2TS U2629 ( .A(requesterAddressIn_NORTH[2]), .Y(n4061) );
  CLKBUFX2TS U2630 ( .A(requesterAddressIn_NORTH[1]), .Y(n4058) );
  CLKBUFX2TS U2631 ( .A(requesterAddressIn_NORTH[0]), .Y(n4055) );
  CLKBUFX2TS U2632 ( .A(destinationAddressIn_NORTH[0]), .Y(n4037) );
  CLKBUFX2TS U2633 ( .A(dataIn_NORTH[0]), .Y(n4073) );
  CLKBUFX2TS U2634 ( .A(destinationAddressIn_NORTH[5]), .Y(n4052) );
  CLKBUFX2TS U2635 ( .A(destinationAddressIn_NORTH[3]), .Y(n4046) );
  CLKBUFX2TS U2636 ( .A(destinationAddressIn_NORTH[2]), .Y(n4043) );
  CLKBUFX2TS U2637 ( .A(destinationAddressIn_NORTH[1]), .Y(n4040) );
  CLKBUFX2TS U2638 ( .A(dataIn_NORTH[31]), .Y(n4166) );
  CLKBUFX2TS U2639 ( .A(dataIn_NORTH[30]), .Y(n4163) );
  CLKBUFX2TS U2640 ( .A(dataIn_NORTH[29]), .Y(n4160) );
  CLKBUFX2TS U2641 ( .A(dataIn_NORTH[28]), .Y(n4157) );
  CLKBUFX2TS U2642 ( .A(dataIn_NORTH[27]), .Y(n4154) );
  CLKBUFX2TS U2643 ( .A(dataIn_NORTH[26]), .Y(n4151) );
  CLKBUFX2TS U2644 ( .A(dataIn_NORTH[25]), .Y(n4148) );
  CLKBUFX2TS U2645 ( .A(dataIn_NORTH[24]), .Y(n4145) );
  CLKBUFX2TS U2646 ( .A(dataIn_NORTH[23]), .Y(n4142) );
  CLKBUFX2TS U2647 ( .A(dataIn_NORTH[22]), .Y(n4139) );
  CLKBUFX2TS U2648 ( .A(dataIn_NORTH[21]), .Y(n4136) );
  CLKBUFX2TS U2649 ( .A(dataIn_NORTH[20]), .Y(n4133) );
  CLKBUFX2TS U2650 ( .A(dataIn_NORTH[19]), .Y(n4130) );
  CLKBUFX2TS U2651 ( .A(dataIn_NORTH[18]), .Y(n4127) );
  CLKBUFX2TS U2652 ( .A(dataIn_NORTH[17]), .Y(n4124) );
  CLKBUFX2TS U2653 ( .A(dataIn_NORTH[16]), .Y(n4121) );
  CLKBUFX2TS U2654 ( .A(dataIn_NORTH[12]), .Y(n4109) );
  CLKBUFX2TS U2655 ( .A(dataIn_NORTH[11]), .Y(n4106) );
  CLKBUFX2TS U2656 ( .A(dataIn_NORTH[10]), .Y(n4103) );
  CLKBUFX2TS U2657 ( .A(dataIn_NORTH[9]), .Y(n4100) );
  CLKBUFX2TS U2658 ( .A(dataIn_NORTH[8]), .Y(n4097) );
  CLKBUFX2TS U2659 ( .A(dataIn_NORTH[7]), .Y(n4094) );
  CLKBUFX2TS U2660 ( .A(dataIn_NORTH[6]), .Y(n4091) );
  CLKBUFX2TS U2661 ( .A(dataIn_NORTH[5]), .Y(n4088) );
  CLKBUFX2TS U2662 ( .A(dataIn_NORTH[3]), .Y(n4082) );
  CLKBUFX2TS U2663 ( .A(dataIn_NORTH[2]), .Y(n4079) );
  CLKBUFX2TS U2664 ( .A(dataIn_NORTH[1]), .Y(n4076) );
  CLKBUFX2TS U2665 ( .A(destinationAddressIn_NORTH[4]), .Y(n4049) );
  CLKBUFX2TS U2666 ( .A(dataIn_NORTH[4]), .Y(n4085) );
  NOR2X1TS U2667 ( .A(n914), .B(n1092), .Y(n2885) );
  AOI31X1TS U2668 ( .A0(n1093), .A1(n716), .A2(n1094), .B0(n139), .Y(n1092) );
  XNOR2X1TS U2669 ( .A(n1095), .B(n1096), .Y(n1093) );
  INVX2TS U2670 ( .A(readIn_EAST), .Y(n4198) );
  INVX2TS U2671 ( .A(writeIn_WEST), .Y(n4187) );
  INVX2TS U2672 ( .A(writeIn_WEST), .Y(n4188) );
  XNOR2X1TS U2673 ( .A(n2898), .B(n1096), .Y(n2897) );
  OAI2BB1X1TS U2674 ( .A0N(n120), .A1N(n2899), .B0(n2900), .Y(n2898) );
  OAI21X1TS U2675 ( .A0(n2899), .A1(n2), .B0(n3), .Y(n2900) );
  NOR2X1TS U2676 ( .A(n136), .B(n166), .Y(n2899) );
  XOR2X1TS U2677 ( .A(n115), .B(n113), .Y(n1096) );
  INVX2TS U2678 ( .A(n1094), .Y(n715) );
  OAI22X1TS U2679 ( .A0(n717), .A1(n706), .B0(n707), .B1(n2036), .Y(n2046) );
  OAI22X1TS U2680 ( .A0(n660), .A1(n2032), .B0(n653), .B1(n167), .Y(n2045) );
  AOI21X1TS U2681 ( .A0(n137), .A1(n925), .B0(n2899), .Y(n2896) );
  NAND2X1TS U2682 ( .A(n143), .B(n113), .Y(n1938) );
  CLKBUFX2TS U2683 ( .A(n2048), .Y(n924) );
  NOR2X1TS U2684 ( .A(n1095), .B(n913), .Y(n2048) );
  OAI22X1TS U2685 ( .A0(n910), .A1(n2049), .B0(n911), .B1(n2033), .Y(n2044) );
  OAI22X1TS U2686 ( .A0(n705), .A1(n2034), .B0(n708), .B1(n2035), .Y(n2047) );
  OAI22X1TS U2687 ( .A0(n717), .A1(n649), .B0(n2032), .B1(n654), .Y(n2031) );
  OAI22X1TS U2688 ( .A0(n2033), .A1(n655), .B0(n2034), .B1(n656), .Y(n2030) );
  NAND3X1TS U2689 ( .A(n2), .B(n137), .C(n115), .Y(n2032) );
  INVX2TS U2690 ( .A(n2033), .Y(n719) );
  INVX2TS U2691 ( .A(n2049), .Y(n711) );
  AOI222XLTS U2692 ( .A0(n4227), .A1(n3389), .B0(n4005), .B1(n3354), .C0(n3962), .C1(n3404), .Y(n1956) );
  AOI222XLTS U2693 ( .A0(n4230), .A1(n3389), .B0(n4008), .B1(n3355), .C0(n3965), .C1(n3404), .Y(n1957) );
  AOI222XLTS U2694 ( .A0(n4233), .A1(n3388), .B0(n4011), .B1(n3354), .C0(n3968), .C1(n3403), .Y(n1958) );
  AOI222XLTS U2695 ( .A0(n4236), .A1(n3384), .B0(n4014), .B1(n3355), .C0(n3971), .C1(n3403), .Y(n1959) );
  AOI222XLTS U2696 ( .A0(n4239), .A1(n3388), .B0(n4017), .B1(n3359), .C0(n3974), .C1(n3403), .Y(n1960) );
  AOI222XLTS U2697 ( .A0(n4221), .A1(n3387), .B0(n3999), .B1(n1187), .C0(n3956), .C1(n3406), .Y(n1954) );
  AOI222XLTS U2698 ( .A0(n4224), .A1(n3385), .B0(n4002), .B1(n3360), .C0(n3959), .C1(n3404), .Y(n1955) );
  AOI222XLTS U2699 ( .A0(n4218), .A1(n3386), .B0(n3996), .B1(n1187), .C0(n3953), .C1(n3406), .Y(n1953) );
  AOI222XLTS U2700 ( .A0(n4010), .A1(n3455), .B0(n3969), .B1(n3438), .C0(n4234), .C1(n3420), .Y(n1934) );
  AOI222XLTS U2701 ( .A0(n3995), .A1(n3457), .B0(n3954), .B1(n3436), .C0(n4219), .C1(n3419), .Y(n1929) );
  AOI222XLTS U2702 ( .A0(n4013), .A1(n3455), .B0(n3972), .B1(n3439), .C0(n4237), .C1(n3426), .Y(n1935) );
  AOI222XLTS U2703 ( .A0(n4004), .A1(n3456), .B0(n3963), .B1(n3438), .C0(n4228), .C1(n1171), .Y(n1932) );
  AOI222XLTS U2704 ( .A0(n4001), .A1(n3456), .B0(n3960), .B1(n3436), .C0(n4225), .C1(n3419), .Y(n1931) );
  AOI222XLTS U2705 ( .A0(n4016), .A1(n3455), .B0(n3975), .B1(n3442), .C0(n4240), .C1(n3425), .Y(n1936) );
  AOI222XLTS U2706 ( .A0(n4007), .A1(n3456), .B0(n3966), .B1(n3439), .C0(n4231), .C1(n1171), .Y(n1933) );
  AOI222XLTS U2707 ( .A0(n3998), .A1(n3457), .B0(n3957), .B1(n3436), .C0(n4222), .C1(n3419), .Y(n1930) );
  AOI22X1TS U2708 ( .A0(n3639), .A1(n43), .B0(n3992), .B1(n3612), .Y(n1858) );
  AOI222XLTS U2709 ( .A0(n2998), .A1(n3112), .B0(n4216), .B1(n3655), .C0(n4053), .C1(n3806), .Y(n1859) );
  AOI22X1TS U2710 ( .A0(n3639), .A1(n32), .B0(n3986), .B1(n3613), .Y(n1854) );
  AOI222XLTS U2711 ( .A0(n3002), .A1(n3111), .B0(n4211), .B1(n3657), .C0(n4047), .C1(n3806), .Y(n1855) );
  AOI22X1TS U2712 ( .A0(n3636), .A1(n29), .B0(n3983), .B1(n3612), .Y(n1852) );
  AOI222XLTS U2713 ( .A0(n3004), .A1(n3111), .B0(n4209), .B1(n3658), .C0(n4044), .C1(n3806), .Y(n1853) );
  AOI22X1TS U2714 ( .A0(n3639), .A1(n22), .B0(n3980), .B1(n3613), .Y(n1850) );
  AOI222XLTS U2715 ( .A0(n3006), .A1(n3111), .B0(n4206), .B1(n3655), .C0(n4041), .C1(n3805), .Y(n1851) );
  AOI22X1TS U2716 ( .A0(n3640), .A1(n17), .B0(n3977), .B1(n3613), .Y(n1848) );
  AOI222XLTS U2717 ( .A0(n3008), .A1(n3110), .B0(n4202), .B1(n3653), .C0(n4038), .C1(n3805), .Y(n1849) );
  AOI22X1TS U2718 ( .A0(n3637), .A1(n36), .B0(n3989), .B1(n3613), .Y(n1856) );
  AOI222XLTS U2719 ( .A0(n3000), .A1(n3111), .B0(n4212), .B1(n3653), .C0(n4050), .C1(n3806), .Y(n1857) );
  AOI22X1TS U2720 ( .A0(n3635), .A1(n14), .B0(n3612), .B1(n4034), .Y(n1132) );
  AOI222XLTS U2721 ( .A0(\requesterAddressbuffer[6][5] ), .A1(n3110), .B0(
        n3654), .B1(requesterAddressIn_SOUTH[5]), .C0(n3805), .C1(n4072), .Y(
        n1133) );
  AOI22X1TS U2722 ( .A0(n3635), .A1(n37), .B0(n3611), .B1(n4031), .Y(n1130) );
  AOI222XLTS U2723 ( .A0(\requesterAddressbuffer[6][4] ), .A1(n3113), .B0(
        n3650), .B1(requesterAddressIn_SOUTH[4]), .C0(n3804), .C1(n4069), .Y(
        n1131) );
  AOI22X1TS U2724 ( .A0(n3639), .A1(n32), .B0(n3611), .B1(n4028), .Y(n1128) );
  AOI222XLTS U2725 ( .A0(\requesterAddressbuffer[6][3] ), .A1(n3110), .B0(
        n3650), .B1(requesterAddressIn_SOUTH[3]), .C0(n3804), .C1(n4066), .Y(
        n1129) );
  AOI22X1TS U2726 ( .A0(n3640), .A1(n27), .B0(n3611), .B1(n4025), .Y(n1126) );
  AOI222XLTS U2727 ( .A0(\requesterAddressbuffer[6][2] ), .A1(n3109), .B0(
        n3650), .B1(requesterAddressIn_SOUTH[2]), .C0(n3804), .C1(n4063), .Y(
        n1127) );
  AOI22X1TS U2728 ( .A0(n3641), .A1(n22), .B0(n3612), .B1(n4022), .Y(n1124) );
  AOI222XLTS U2729 ( .A0(\requesterAddressbuffer[6][1] ), .A1(n3108), .B0(
        n3650), .B1(requesterAddressIn_SOUTH[1]), .C0(n3804), .C1(n4060), .Y(
        n1125) );
  AOI22X1TS U2730 ( .A0(n3638), .A1(n17), .B0(n3611), .B1(n4019), .Y(n1119) );
  AOI222XLTS U2731 ( .A0(\requesterAddressbuffer[6][0] ), .A1(n3110), .B0(
        n3656), .B1(requesterAddressIn_SOUTH[0]), .C0(n3805), .C1(n4057), .Y(
        n1120) );
  AOI222XLTS U2732 ( .A0(n4195), .A1(n1772), .B0(readIn_NORTH), .B1(n1773), 
        .C0(n4190), .C1(n758), .Y(n1771) );
  INVX2TS U2733 ( .A(n4197), .Y(n4196) );
  XOR2X1TS U2734 ( .A(n2388), .B(n2389), .Y(n1090) );
  XOR2X1TS U2735 ( .A(n1), .B(n2390), .Y(n2389) );
  OAI21X1TS U2736 ( .A0(n2393), .A1(n2394), .B0(n2395), .Y(n2388) );
  NOR2X1TS U2737 ( .A(n2391), .B(n2392), .Y(n2390) );
  INVX2TS U2738 ( .A(selectBit_SOUTH), .Y(n971) );
  OAI32X1TS U2739 ( .A0(n2385), .A1(n2386), .A2(n2387), .B0(n6347), .B1(n154), 
        .Y(N4718) );
  NAND2X1TS U2740 ( .A(n2891), .B(n914), .Y(n2385) );
  XOR2X1TS U2741 ( .A(n1089), .B(n2), .Y(n2386) );
  XOR2X1TS U2742 ( .A(n1090), .B(n6), .Y(n2387) );
  NOR2BX1TS U2743 ( .AN(n2903), .B(n2383), .Y(n2901) );
  XOR2X1TS U2744 ( .A(n1083), .B(n470), .Y(n2902) );
  OAI221XLTS U2745 ( .A0(n543), .A1(n132), .B0(n3326), .B1(n773), .C0(n1984), 
        .Y(n2465) );
  AOI222XLTS U2746 ( .A0(n3974), .A1(n3276), .B0(n4017), .B1(n3278), .C0(n4240), .C1(n3320), .Y(n1984) );
  OAI221XLTS U2747 ( .A0(n542), .A1(n125), .B0(n3326), .B1(n772), .C0(n1983), 
        .Y(n2466) );
  AOI222XLTS U2748 ( .A0(n3971), .A1(n1204), .B0(n4014), .B1(n3278), .C0(n4237), .C1(n3319), .Y(n1983) );
  OAI221XLTS U2749 ( .A0(n543), .A1(n127), .B0(n3326), .B1(n771), .C0(n1982), 
        .Y(n2467) );
  AOI222XLTS U2750 ( .A0(n3968), .A1(n3272), .B0(n4011), .B1(n3278), .C0(n4234), .C1(n3319), .Y(n1982) );
  OAI221XLTS U2751 ( .A0(n542), .A1(n135), .B0(n3326), .B1(n770), .C0(n1981), 
        .Y(n2468) );
  AOI222XLTS U2752 ( .A0(n3965), .A1(n1204), .B0(n4008), .B1(n3278), .C0(n4231), .C1(n3319), .Y(n1981) );
  OAI221XLTS U2753 ( .A0(n543), .A1(n129), .B0(n3327), .B1(n769), .C0(n1980), 
        .Y(n2469) );
  AOI222XLTS U2754 ( .A0(n3962), .A1(n3272), .B0(n4005), .B1(n3279), .C0(n4228), .C1(n3319), .Y(n1980) );
  OAI221XLTS U2755 ( .A0(n542), .A1(n131), .B0(n3327), .B1(n768), .C0(n1979), 
        .Y(n2470) );
  AOI222XLTS U2756 ( .A0(n3959), .A1(n3270), .B0(n4002), .B1(n3279), .C0(n4225), .C1(n3318), .Y(n1979) );
  OAI221XLTS U2757 ( .A0(n543), .A1(n124), .B0(n3327), .B1(n767), .C0(n1978), 
        .Y(n2471) );
  AOI222XLTS U2758 ( .A0(n3956), .A1(n3270), .B0(n3999), .B1(n3279), .C0(n4222), .C1(n3318), .Y(n1978) );
  OAI221XLTS U2759 ( .A0(n542), .A1(n122), .B0(n3327), .B1(n766), .C0(n1977), 
        .Y(n2472) );
  AOI222XLTS U2760 ( .A0(n3953), .A1(n3270), .B0(n3996), .B1(n3279), .C0(n4219), .C1(n3318), .Y(n1977) );
  OAI221XLTS U2761 ( .A0(n468), .A1(n126), .B0(n160), .B1(n594), .C0(n1912), 
        .Y(n2508) );
  AOI222XLTS U2762 ( .A0(n4236), .A1(n3492), .B0(n3972), .B1(n3469), .C0(n4013), .C1(n3522), .Y(n1912) );
  OAI221XLTS U2763 ( .A0(n467), .A1(n127), .B0(n159), .B1(n593), .C0(n1911), 
        .Y(n2509) );
  AOI222XLTS U2764 ( .A0(n4233), .A1(n3492), .B0(n3969), .B1(n3469), .C0(n4010), .C1(n3522), .Y(n1911) );
  OAI221XLTS U2765 ( .A0(n468), .A1(n135), .B0(n160), .B1(n592), .C0(n1910), 
        .Y(n2510) );
  AOI222XLTS U2766 ( .A0(n4230), .A1(n3492), .B0(n3966), .B1(n3469), .C0(n4007), .C1(n3523), .Y(n1910) );
  OAI221XLTS U2767 ( .A0(n467), .A1(n966), .B0(n159), .B1(n591), .C0(n1908), 
        .Y(n2512) );
  AOI222XLTS U2768 ( .A0(n4224), .A1(n3493), .B0(n3960), .B1(n3470), .C0(n4001), .C1(n3523), .Y(n1908) );
  OAI221XLTS U2769 ( .A0(n468), .A1(n124), .B0(n160), .B1(n590), .C0(n1907), 
        .Y(n2513) );
  AOI222XLTS U2770 ( .A0(n4221), .A1(n3493), .B0(n3957), .B1(n3472), .C0(n3998), .C1(n3524), .Y(n1907) );
  OAI221XLTS U2771 ( .A0(n467), .A1(n968), .B0(n159), .B1(n589), .C0(n1906), 
        .Y(n2514) );
  AOI222XLTS U2772 ( .A0(n4218), .A1(n3493), .B0(n3954), .B1(n3470), .C0(n3995), .C1(n3524), .Y(n1906) );
  OAI221XLTS U2773 ( .A0(n468), .A1(n129), .B0(n160), .B1(n576), .C0(n1909), 
        .Y(n2511) );
  AOI222XLTS U2774 ( .A0(n4227), .A1(n3493), .B0(n3963), .B1(n3469), .C0(n4004), .C1(n3523), .Y(n1909) );
  OAI221XLTS U2775 ( .A0(n544), .A1(n4018), .B0(n3243), .B1(n917), .C0(n2005), 
        .Y(n2451) );
  AOI222XLTS U2776 ( .A0(n4239), .A1(n3192), .B0(
        destinationAddressIn_NORTH[13]), .B1(n3220), .C0(n3974), .C1(n3241), 
        .Y(n2005) );
  OAI221XLTS U2777 ( .A0(n546), .A1(n4015), .B0(n3243), .B1(n909), .C0(n2004), 
        .Y(n2452) );
  AOI222XLTS U2778 ( .A0(n4236), .A1(n3122), .B0(
        destinationAddressIn_NORTH[12]), .B1(n3220), .C0(n3971), .C1(n3234), 
        .Y(n2004) );
  OAI221XLTS U2779 ( .A0(n545), .A1(n4009), .B0(n3243), .B1(n908), .C0(n2002), 
        .Y(n2454) );
  AOI222XLTS U2780 ( .A0(n4230), .A1(n3122), .B0(
        destinationAddressIn_NORTH[10]), .B1(n3223), .C0(n3965), .C1(n3234), 
        .Y(n2002) );
  OAI221XLTS U2781 ( .A0(n546), .A1(n4012), .B0(n3243), .B1(n907), .C0(n2003), 
        .Y(n2453) );
  AOI222XLTS U2782 ( .A0(n4233), .A1(n3122), .B0(
        destinationAddressIn_NORTH[11]), .B1(n3223), .C0(n3968), .C1(n3234), 
        .Y(n2003) );
  OAI221XLTS U2783 ( .A0(n545), .A1(n4006), .B0(n3244), .B1(n906), .C0(n2001), 
        .Y(n2455) );
  AOI222XLTS U2784 ( .A0(n4227), .A1(n3122), .B0(destinationAddressIn_NORTH[9]), .B1(n3209), .C0(n3962), .C1(n3234), .Y(n2001) );
  OAI221XLTS U2785 ( .A0(n465), .A1(n134), .B0(n3099), .B1(n587), .C0(n1865), 
        .Y(n2538) );
  AOI222XLTS U2786 ( .A0(n4230), .A1(n3652), .B0(n4008), .B1(n3615), .C0(n3965), .C1(n3793), .Y(n1865) );
  OAI221XLTS U2787 ( .A0(n465), .A1(n130), .B0(n3099), .B1(n586), .C0(n1864), 
        .Y(n2539) );
  AOI222XLTS U2788 ( .A0(n4227), .A1(n3652), .B0(n4005), .B1(n3614), .C0(n3962), .C1(n3793), .Y(n1864) );
  OAI221XLTS U2789 ( .A0(n464), .A1(n131), .B0(n3099), .B1(n573), .C0(n1863), 
        .Y(n2540) );
  AOI222XLTS U2790 ( .A0(n4224), .A1(n3657), .B0(n4002), .B1(n3615), .C0(n3959), .C1(n3798), .Y(n1863) );
  OAI221XLTS U2791 ( .A0(n464), .A1(n967), .B0(n3099), .B1(n572), .C0(n1862), 
        .Y(n2541) );
  AOI222XLTS U2792 ( .A0(n4221), .A1(n3652), .B0(n3999), .B1(n3614), .C0(n3956), .C1(n3798), .Y(n1862) );
  OAI221XLTS U2793 ( .A0(n460), .A1(n133), .B0(n3593), .B1(n566), .C0(n1892), 
        .Y(n2521) );
  AOI222XLTS U2794 ( .A0(n4016), .A1(n3543), .B0(n3975), .B1(n3545), .C0(n4240), .C1(n3589), .Y(n1892) );
  OAI221XLTS U2795 ( .A0(n461), .A1(n126), .B0(n3593), .B1(n565), .C0(n1891), 
        .Y(n2522) );
  AOI222XLTS U2796 ( .A0(n4013), .A1(n3539), .B0(n3972), .B1(n3545), .C0(n4237), .C1(n3586), .Y(n1891) );
  OAI221XLTS U2797 ( .A0(n460), .A1(n128), .B0(n3593), .B1(n564), .C0(n1890), 
        .Y(n2523) );
  AOI222XLTS U2798 ( .A0(n4010), .A1(n3538), .B0(n3969), .B1(n3545), .C0(n4234), .C1(n3586), .Y(n1890) );
  OAI221XLTS U2799 ( .A0(n461), .A1(n130), .B0(n3594), .B1(n562), .C0(n1888), 
        .Y(n2525) );
  AOI222XLTS U2800 ( .A0(n4004), .A1(n3539), .B0(n3963), .B1(n3546), .C0(n4228), .C1(n3586), .Y(n1888) );
  OAI221XLTS U2801 ( .A0(n460), .A1(n966), .B0(n3594), .B1(n561), .C0(n1887), 
        .Y(n2526) );
  AOI222XLTS U2802 ( .A0(n4001), .A1(n3544), .B0(n3960), .B1(n3546), .C0(n4225), .C1(n3585), .Y(n1887) );
  OAI221XLTS U2803 ( .A0(n461), .A1(n967), .B0(n3594), .B1(n560), .C0(n1886), 
        .Y(n2527) );
  AOI222XLTS U2804 ( .A0(n3998), .A1(n1140), .B0(n3957), .B1(n3546), .C0(n4222), .C1(n3585), .Y(n1886) );
  OAI221XLTS U2805 ( .A0(n460), .A1(n968), .B0(n3594), .B1(n559), .C0(n1885), 
        .Y(n2528) );
  AOI222XLTS U2806 ( .A0(n3995), .A1(n1140), .B0(n3954), .B1(n3546), .C0(n4219), .C1(n3585), .Y(n1885) );
  OAI221XLTS U2807 ( .A0(n546), .A1(n4003), .B0(n3244), .B1(n555), .C0(n2000), 
        .Y(n2456) );
  AOI222XLTS U2808 ( .A0(n4224), .A1(n3193), .B0(destinationAddressIn_NORTH[8]), .B1(n3209), .C0(n3959), .C1(n3241), .Y(n2000) );
  OAI221XLTS U2809 ( .A0(n545), .A1(n3997), .B0(n3244), .B1(n554), .C0(n1998), 
        .Y(n2458) );
  AOI222XLTS U2810 ( .A0(n4218), .A1(n3124), .B0(destinationAddressIn_NORTH[6]), .B1(n3209), .C0(n3953), .C1(n3241), .Y(n1998) );
  OAI221XLTS U2811 ( .A0(n546), .A1(n4000), .B0(n3244), .B1(n553), .C0(n1999), 
        .Y(n2457) );
  AOI222XLTS U2812 ( .A0(n4221), .A1(n3124), .B0(destinationAddressIn_NORTH[7]), .B1(n3209), .C0(n3956), .C1(n1218), .Y(n1999) );
  OAI221XLTS U2813 ( .A0(n545), .A1(writeIn_WEST), .B0(n3245), .B1(n705), .C0(
        n1762), .Y(n2571) );
  AOI222XLTS U2814 ( .A0(n4200), .A1(n3124), .B0(writeIn_NORTH), .B1(n3211), 
        .C0(n4192), .C1(n3242), .Y(n1762) );
  OAI221XLTS U2815 ( .A0(n465), .A1(n122), .B0(n3100), .B1(n585), .C0(n1861), 
        .Y(n2542) );
  AOI222XLTS U2816 ( .A0(n4218), .A1(n1121), .B0(n3996), .B1(n3616), .C0(n3953), .C1(n3798), .Y(n1861) );
  OAI221XLTS U2817 ( .A0(n464), .A1(n125), .B0(n3098), .B1(n588), .C0(n1867), 
        .Y(n2536) );
  AOI222XLTS U2818 ( .A0(n4236), .A1(n3657), .B0(n4014), .B1(n3615), .C0(n3971), .C1(n3793), .Y(n1867) );
  OAI221XLTS U2819 ( .A0(n465), .A1(n133), .B0(n3098), .B1(n575), .C0(n1868), 
        .Y(n2535) );
  AOI222XLTS U2820 ( .A0(n4239), .A1(n3658), .B0(n4017), .B1(n3614), .C0(n3974), .C1(n3795), .Y(n1868) );
  OAI221XLTS U2821 ( .A0(n464), .A1(n128), .B0(n3098), .B1(n574), .C0(n1866), 
        .Y(n2537) );
  AOI222XLTS U2822 ( .A0(n4233), .A1(n3654), .B0(n4011), .B1(n3614), .C0(n3968), .C1(n3793), .Y(n1866) );
  OAI221XLTS U2823 ( .A0(n3671), .A1(n135), .B0(n4796), .B1(n3748), .C0(n1837), 
        .Y(n2552) );
  AOI222XLTS U2824 ( .A0(n4007), .A1(n3690), .B0(n3966), .B1(n3693), .C0(
        destinationAddressIn_SOUTH[10]), .C1(n3732), .Y(n1837) );
  OAI221XLTS U2825 ( .A0(n3671), .A1(n129), .B0(n3757), .B1(n584), .C0(n1836), 
        .Y(n2553) );
  AOI222XLTS U2826 ( .A0(n4004), .A1(n3689), .B0(n3963), .B1(n3694), .C0(
        destinationAddressIn_SOUTH[9]), .C1(n3732), .Y(n1836) );
  OAI221XLTS U2827 ( .A0(n3670), .A1(n127), .B0(n3755), .B1(n581), .C0(n1838), 
        .Y(n2551) );
  AOI222XLTS U2828 ( .A0(n4010), .A1(n3690), .B0(n3969), .B1(n3693), .C0(
        destinationAddressIn_SOUTH[11]), .C1(n3732), .Y(n1838) );
  OAI221XLTS U2829 ( .A0(n3671), .A1(n966), .B0(n1100), .B1(n580), .C0(n1835), 
        .Y(n2554) );
  AOI222XLTS U2830 ( .A0(n4001), .A1(n3687), .B0(n3960), .B1(n3694), .C0(
        destinationAddressIn_SOUTH[8]), .C1(n3731), .Y(n1835) );
  OAI221XLTS U2831 ( .A0(n3672), .A1(n124), .B0(n3752), .B1(n579), .C0(n1834), 
        .Y(n2555) );
  AOI222XLTS U2832 ( .A0(n3998), .A1(n3687), .B0(n3957), .B1(n3694), .C0(n4220), .C1(n3731), .Y(n1834) );
  OAI221XLTS U2833 ( .A0(n3672), .A1(n968), .B0(n3755), .B1(n578), .C0(n1833), 
        .Y(n2556) );
  AOI222XLTS U2834 ( .A0(n3995), .A1(n3687), .B0(n3954), .B1(n3694), .C0(n4217), .C1(n3731), .Y(n1833) );
  OAI221XLTS U2835 ( .A0(n3670), .A1(n132), .B0(n3754), .B1(n583), .C0(n1840), 
        .Y(n2549) );
  AOI222XLTS U2836 ( .A0(n4016), .A1(n1106), .B0(n3975), .B1(n3693), .C0(
        destinationAddressIn_SOUTH[13]), .C1(n3739), .Y(n1840) );
  OAI221XLTS U2837 ( .A0(n3670), .A1(n126), .B0(n3754), .B1(n582), .C0(n1839), 
        .Y(n2550) );
  AOI222XLTS U2838 ( .A0(n4013), .A1(n3689), .B0(n3972), .B1(n3693), .C0(
        destinationAddressIn_SOUTH[12]), .C1(n3732), .Y(n1839) );
  OAI211X1TS U2839 ( .A0(n3596), .A1(n899), .B0(n1149), .C0(n1150), .Y(n2865)
         );
  AOI22X1TS U2840 ( .A0(n3529), .A1(n4034), .B0(n3918), .B1(n4071), .Y(n1149)
         );
  AOI222XLTS U2841 ( .A0(n3577), .A1(n4537), .B0(n3569), .B1(n42), .C0(n3548), 
        .C1(n4185), .Y(n1150) );
  OAI211X1TS U2842 ( .A0(n3596), .A1(n898), .B0(n1147), .C0(n1148), .Y(n2866)
         );
  AOI22X1TS U2843 ( .A0(n3528), .A1(n4031), .B0(n3920), .B1(n4068), .Y(n1147)
         );
  AOI222XLTS U2844 ( .A0(n3576), .A1(n4535), .B0(n3569), .B1(n38), .C0(n3548), 
        .C1(n4182), .Y(n1148) );
  OAI211X1TS U2845 ( .A0(n3595), .A1(n897), .B0(n1145), .C0(n1146), .Y(n2867)
         );
  AOI22X1TS U2846 ( .A0(n3528), .A1(n4028), .B0(n3909), .B1(n4065), .Y(n1145)
         );
  AOI222XLTS U2847 ( .A0(n3576), .A1(n4532), .B0(n3568), .B1(n34), .C0(n3547), 
        .C1(n4179), .Y(n1146) );
  OAI211X1TS U2848 ( .A0(n3596), .A1(n896), .B0(n1143), .C0(n1144), .Y(n2868)
         );
  AOI22X1TS U2849 ( .A0(n3528), .A1(n4025), .B0(n3909), .B1(n4062), .Y(n1143)
         );
  AOI222XLTS U2850 ( .A0(n3576), .A1(n4530), .B0(n3568), .B1(n29), .C0(n3547), 
        .C1(n4176), .Y(n1144) );
  OAI211X1TS U2851 ( .A0(n3595), .A1(n895), .B0(n1141), .C0(n1142), .Y(n2869)
         );
  AOI22X1TS U2852 ( .A0(n3528), .A1(n4022), .B0(n3909), .B1(n4059), .Y(n1141)
         );
  AOI222XLTS U2853 ( .A0(n3576), .A1(n4527), .B0(n3568), .B1(n24), .C0(n3547), 
        .C1(n4173), .Y(n1142) );
  OAI211X1TS U2854 ( .A0(n3600), .A1(n894), .B0(n1135), .C0(n1136), .Y(n2870)
         );
  AOI22X1TS U2855 ( .A0(n3529), .A1(n4019), .B0(n3909), .B1(n4056), .Y(n1135)
         );
  AOI222XLTS U2856 ( .A0(n3577), .A1(n4526), .B0(n3569), .B1(n19), .C0(n3548), 
        .C1(n4170), .Y(n1136) );
  AOI222XLTS U2857 ( .A0(n4212), .A1(n3317), .B0(n3300), .B1(n38), .C0(n3990), 
        .C1(n1203), .Y(n1973) );
  AOI22X1TS U2858 ( .A0(n3262), .A1(n4184), .B0(n3869), .B1(n4071), .Y(n1213)
         );
  AOI222XLTS U2859 ( .A0(n3310), .A1(n4537), .B0(n3301), .B1(n42), .C0(n3281), 
        .C1(n4035), .Y(n1214) );
  AOI22X1TS U2860 ( .A0(n3261), .A1(n4181), .B0(n3869), .B1(n4068), .Y(n1211)
         );
  AOI222XLTS U2861 ( .A0(n3309), .A1(n4535), .B0(n3307), .B1(n39), .C0(n3281), 
        .C1(n4032), .Y(n1212) );
  AOI22X1TS U2862 ( .A0(n3261), .A1(n4178), .B0(n3868), .B1(n4065), .Y(n1209)
         );
  AOI222XLTS U2863 ( .A0(n3309), .A1(n4532), .B0(n3301), .B1(n33), .C0(n3280), 
        .C1(n4029), .Y(n1210) );
  AOI22X1TS U2864 ( .A0(n3261), .A1(n4175), .B0(n3868), .B1(n4062), .Y(n1207)
         );
  AOI222XLTS U2865 ( .A0(n3309), .A1(n4530), .B0(n3301), .B1(n28), .C0(n3280), 
        .C1(n4026), .Y(n1208) );
  AOI22X1TS U2866 ( .A0(n3261), .A1(n4172), .B0(n3868), .B1(n4059), .Y(n1205)
         );
  AOI222XLTS U2867 ( .A0(n3309), .A1(n4527), .B0(n3302), .B1(n23), .C0(n3280), 
        .C1(n4023), .Y(n1206) );
  AOI22X1TS U2868 ( .A0(n3262), .A1(n4169), .B0(n3868), .B1(n4056), .Y(n1199)
         );
  AOI222XLTS U2869 ( .A0(n3310), .A1(n4526), .B0(n3304), .B1(n18), .C0(n3281), 
        .C1(n4020), .Y(n1200) );
  AOI22X1TS U2870 ( .A0(n3950), .A1(n3435), .B0(n4215), .B1(n3418), .Y(n1926)
         );
  AOI222XLTS U2871 ( .A0(n3780), .A1(n41), .B0(n4054), .B1(n3866), .C0(n6255), 
        .C1(n3853), .Y(n1927) );
  AOI22X1TS U2872 ( .A0(n3947), .A1(n3435), .B0(n4213), .B1(n3418), .Y(n1924)
         );
  AOI222XLTS U2873 ( .A0(n3779), .A1(n39), .B0(n4051), .B1(n3866), .C0(n6256), 
        .C1(n3849), .Y(n1925) );
  AOI22X1TS U2874 ( .A0(n3944), .A1(n3435), .B0(n4210), .B1(n3418), .Y(n1922)
         );
  AOI222XLTS U2875 ( .A0(n3783), .A1(n34), .B0(n4048), .B1(n3866), .C0(n6257), 
        .C1(n3848), .Y(n1923) );
  AOI22X1TS U2876 ( .A0(n3938), .A1(n3434), .B0(n4205), .B1(n3424), .Y(n1918)
         );
  AOI222XLTS U2877 ( .A0(n3772), .A1(n24), .B0(n4042), .B1(n3865), .C0(n6258), 
        .C1(n3848), .Y(n1919) );
  AOI22X1TS U2878 ( .A0(n3935), .A1(n3434), .B0(n4203), .B1(n3424), .Y(n1916)
         );
  AOI222XLTS U2879 ( .A0(n3785), .A1(n19), .B0(n4039), .B1(n3865), .C0(n6259), 
        .C1(n3848), .Y(n1917) );
  AOI22X1TS U2880 ( .A0(n3941), .A1(n3435), .B0(n4208), .B1(n3418), .Y(n1920)
         );
  AOI222XLTS U2881 ( .A0(n3783), .A1(n29), .B0(n4045), .B1(n1753), .C0(n6293), 
        .C1(n3848), .Y(n1921) );
  AOI22X1TS U2882 ( .A0(n4215), .A1(n3124), .B0(n3993), .B1(n3892), .Y(n1996)
         );
  AOI222XLTS U2883 ( .A0(n3950), .A1(n3236), .B0(n4054), .B1(n3210), .C0(n3195), .C1(n14), .Y(n1997) );
  AOI22X1TS U2884 ( .A0(n4210), .A1(n1221), .B0(n3987), .B1(n3891), .Y(n1992)
         );
  AOI222XLTS U2885 ( .A0(n3944), .A1(n3237), .B0(n4048), .B1(n3210), .C0(n3197), .C1(n31), .Y(n1993) );
  AOI22X1TS U2886 ( .A0(n4208), .A1(n3194), .B0(n3984), .B1(n3889), .Y(n1990)
         );
  AOI222XLTS U2887 ( .A0(n3941), .A1(n3238), .B0(n4045), .B1(n3210), .C0(n3197), .C1(n26), .Y(n1991) );
  AOI22X1TS U2888 ( .A0(n4205), .A1(n3125), .B0(n3981), .B1(n3890), .Y(n1988)
         );
  AOI222XLTS U2889 ( .A0(n3938), .A1(n3242), .B0(n4042), .B1(n3211), .C0(n3196), .C1(n21), .Y(n1989) );
  AOI22X1TS U2890 ( .A0(n4523), .A1(n3128), .B0(n4334), .B1(n3891), .Y(n1294)
         );
  AOI222XLTS U2891 ( .A0(n4434), .A1(n3242), .B0(n4168), .B1(n3211), .C0(n512), 
        .C1(n3206), .Y(n1295) );
  AOI22X1TS U2892 ( .A0(n4518), .A1(n3194), .B0(n4331), .B1(n728), .Y(n1292)
         );
  AOI222XLTS U2893 ( .A0(n4430), .A1(n3239), .B0(n4165), .B1(n3212), .C0(n508), 
        .C1(n3198), .Y(n1293) );
  AOI22X1TS U2894 ( .A0(n4517), .A1(n3152), .B0(n4328), .B1(n3892), .Y(n1290)
         );
  AOI222XLTS U2895 ( .A0(n4427), .A1(n3236), .B0(n4162), .B1(n3212), .C0(n514), 
        .C1(n3198), .Y(n1291) );
  AOI22X1TS U2896 ( .A0(n4509), .A1(n3152), .B0(n4319), .B1(n3893), .Y(n1284)
         );
  AOI222XLTS U2897 ( .A0(n4416), .A1(n3237), .B0(n4153), .B1(n3213), .C0(n516), 
        .C1(n3202), .Y(n1285) );
  AOI22X1TS U2898 ( .A0(n4507), .A1(n3126), .B0(n4316), .B1(n3888), .Y(n1282)
         );
  AOI222XLTS U2899 ( .A0(n4413), .A1(n3233), .B0(n4150), .B1(n3213), .C0(n518), 
        .C1(n3198), .Y(n1283) );
  AOI22X1TS U2900 ( .A0(n4502), .A1(n3126), .B0(n4313), .B1(n3888), .Y(n1280)
         );
  AOI222XLTS U2901 ( .A0(n4410), .A1(n3233), .B0(n4147), .B1(n3213), .C0(n520), 
        .C1(n3199), .Y(n1281) );
  AOI22X1TS U2902 ( .A0(n4498), .A1(n3127), .B0(n4307), .B1(n3888), .Y(n1276)
         );
  AOI222XLTS U2903 ( .A0(n4404), .A1(n3233), .B0(n4141), .B1(n3214), .C0(n522), 
        .C1(n3199), .Y(n1277) );
  AOI22X1TS U2904 ( .A0(n4496), .A1(n3126), .B0(n4304), .B1(n3887), .Y(n1274)
         );
  AOI222XLTS U2905 ( .A0(n4401), .A1(n3232), .B0(n4138), .B1(n3214), .C0(n524), 
        .C1(n3200), .Y(n1275) );
  AOI22X1TS U2906 ( .A0(n4490), .A1(n3125), .B0(n4298), .B1(n3887), .Y(n1270)
         );
  AOI222XLTS U2907 ( .A0(n4395), .A1(n3232), .B0(n4132), .B1(n3214), .C0(n526), 
        .C1(n3200), .Y(n1271) );
  AOI22X1TS U2908 ( .A0(n4487), .A1(n3121), .B0(n4295), .B1(n3887), .Y(n1268)
         );
  AOI222XLTS U2909 ( .A0(n4392), .A1(n3231), .B0(n4129), .B1(n3215), .C0(n528), 
        .C1(n3201), .Y(n1269) );
  AOI22X1TS U2910 ( .A0(n4484), .A1(n3121), .B0(n4292), .B1(n3886), .Y(n1266)
         );
  AOI222XLTS U2911 ( .A0(n4389), .A1(n3231), .B0(n4126), .B1(n3215), .C0(n530), 
        .C1(n3200), .Y(n1267) );
  AOI22X1TS U2912 ( .A0(n4481), .A1(n3121), .B0(n4289), .B1(n3886), .Y(n1264)
         );
  AOI222XLTS U2913 ( .A0(n4386), .A1(n3231), .B0(n4123), .B1(n3215), .C0(n510), 
        .C1(n3201), .Y(n1265) );
  AOI22X1TS U2914 ( .A0(n4478), .A1(n3121), .B0(n4286), .B1(n3886), .Y(n1262)
         );
  AOI222XLTS U2915 ( .A0(n4383), .A1(n3231), .B0(n4120), .B1(n3215), .C0(n532), 
        .C1(n3202), .Y(n1263) );
  AOI22X1TS U2916 ( .A0(n4474), .A1(n3120), .B0(n4283), .B1(n3886), .Y(n1260)
         );
  AOI222XLTS U2917 ( .A0(n4380), .A1(n3230), .B0(n4117), .B1(n3216), .C0(n534), 
        .C1(n3201), .Y(n1261) );
  AOI22X1TS U2918 ( .A0(n4470), .A1(n3120), .B0(n4280), .B1(n3885), .Y(n1258)
         );
  AOI222XLTS U2919 ( .A0(n4377), .A1(n3230), .B0(n4114), .B1(n3216), .C0(n536), 
        .C1(n3201), .Y(n1259) );
  AOI22X1TS U2920 ( .A0(n3478), .A1(n31), .B0(n3461), .B1(n4178), .Y(n1161) );
  AOI222XLTS U2921 ( .A0(n2931), .A1(n3895), .B0(n3503), .B1(
        requesterAddressIn_SOUTH[3]), .C0(n3922), .C1(n4066), .Y(n1162) );
  AOI22X1TS U2922 ( .A0(n3478), .A1(n26), .B0(n3461), .B1(n4175), .Y(n1159) );
  AOI222XLTS U2923 ( .A0(n2929), .A1(n3894), .B0(n3503), .B1(n4530), .C0(n3922), .C1(n4063), .Y(n1160) );
  AOI22X1TS U2924 ( .A0(n3478), .A1(n21), .B0(n3461), .B1(n4172), .Y(n1157) );
  AOI222XLTS U2925 ( .A0(n2930), .A1(n3894), .B0(n3503), .B1(
        requesterAddressIn_SOUTH[1]), .C0(n3922), .C1(n4060), .Y(n1158) );
  AOI22X1TS U2926 ( .A0(n3479), .A1(n16), .B0(n3462), .B1(n4169), .Y(n1152) );
  AOI222XLTS U2927 ( .A0(n2932), .A1(n3899), .B0(n3503), .B1(n4526), .C0(n3922), .C1(n4057), .Y(n1153) );
  AOI22X1TS U2928 ( .A0(n3427), .A1(n4178), .B0(n3410), .B1(n4533), .Y(n1176)
         );
  AOI222XLTS U2929 ( .A0(n3783), .A1(n33), .B0(n3862), .B1(n4065), .C0(
        \requesterAddressbuffer[3][3] ), .C1(n3841), .Y(n1177) );
  AOI22X1TS U2930 ( .A0(n3427), .A1(n4175), .B0(n3410), .B1(n4529), .Y(n1174)
         );
  AOI222XLTS U2931 ( .A0(n3784), .A1(n28), .B0(n3862), .B1(n4062), .C0(
        \requesterAddressbuffer[3][2] ), .C1(n3853), .Y(n1175) );
  AOI22X1TS U2932 ( .A0(n3427), .A1(n4172), .B0(n3410), .B1(n4528), .Y(n1172)
         );
  AOI222XLTS U2933 ( .A0(n3784), .A1(n23), .B0(n3862), .B1(n4059), .C0(
        \requesterAddressbuffer[3][1] ), .C1(n3853), .Y(n1173) );
  AOI22X1TS U2934 ( .A0(n1170), .A1(n4169), .B0(n3411), .B1(n4525), .Y(n1168)
         );
  AOI222XLTS U2935 ( .A0(n3772), .A1(n18), .B0(n3866), .B1(n4056), .C0(
        \requesterAddressbuffer[3][0] ), .C1(n3849), .Y(n1169) );
  AOI222XLTS U2936 ( .A0(\requesterAddressbuffer[2][1] ), .A1(n3812), .B0(
        n3389), .B1(n4527), .C0(n3827), .C1(n4060), .Y(n1189) );
  AOI222XLTS U2937 ( .A0(\requesterAddressbuffer[2][0] ), .A1(n3814), .B0(
        n3387), .B1(n4526), .C0(n3827), .C1(n4057), .Y(n1184) );
  AOI222XLTS U2938 ( .A0(\requesterAddressbuffer[2][3] ), .A1(n3812), .B0(
        n3385), .B1(n4532), .C0(n3827), .C1(n4066), .Y(n1193) );
  AOI222XLTS U2939 ( .A0(\requesterAddressbuffer[2][2] ), .A1(n3812), .B0(
        n3386), .B1(n4530), .C0(n3827), .C1(n4063), .Y(n1191) );
  AOI22X1TS U2940 ( .A0(n3479), .A1(readRequesterAddress[5]), .B0(n3462), .B1(
        n4184), .Y(n1165) );
  AOI222XLTS U2941 ( .A0(n2927), .A1(n3895), .B0(n3502), .B1(
        requesterAddressIn_SOUTH[5]), .C0(n3923), .C1(n4072), .Y(n1166) );
  AOI22X1TS U2942 ( .A0(n3479), .A1(n39), .B0(n3461), .B1(n4181), .Y(n1163) );
  AOI222XLTS U2943 ( .A0(n2928), .A1(n3895), .B0(n3504), .B1(
        requesterAddressIn_SOUTH[4]), .C0(n3923), .C1(n4069), .Y(n1164) );
  AOI22X1TS U2944 ( .A0(n3427), .A1(n4181), .B0(n3410), .B1(n4536), .Y(n1178)
         );
  AOI222XLTS U2945 ( .A0(n3772), .A1(n38), .B0(n3861), .B1(n4068), .C0(
        \requesterAddressbuffer[3][4] ), .C1(n3841), .Y(n1179) );
  AOI22X1TS U2946 ( .A0(n1170), .A1(n4184), .B0(n3411), .B1(n4538), .Y(n1180)
         );
  AOI222XLTS U2947 ( .A0(n3772), .A1(readRequesterAddress[5]), .B0(n3861), 
        .B1(n4071), .C0(\requesterAddressbuffer[3][5] ), .C1(n3841), .Y(n1181)
         );
  AOI222XLTS U2948 ( .A0(\requesterAddressbuffer[2][4] ), .A1(n3823), .B0(
        n3389), .B1(n4535), .C0(n3828), .C1(n4069), .Y(n1195) );
  AOI22X1TS U2949 ( .A0(n3362), .A1(n36), .B0(n3344), .B1(n4031), .Y(n1194) );
  AOI222XLTS U2950 ( .A0(\requesterAddressbuffer[2][5] ), .A1(n3823), .B0(
        n3383), .B1(n4537), .C0(n3828), .C1(n4072), .Y(n1197) );
  AOI22X1TS U2951 ( .A0(n4280), .A1(n3680), .B0(n4113), .B1(n3665), .Y(n1707)
         );
  AOI222XLTS U2952 ( .A0(n4471), .A1(n3736), .B0(n535), .B1(n3714), .C0(n4377), 
        .C1(n3700), .Y(n1708) );
  AOI22X1TS U2953 ( .A0(n4283), .A1(n3680), .B0(n4116), .B1(n3664), .Y(n1709)
         );
  AOI222XLTS U2954 ( .A0(n4475), .A1(n3736), .B0(n533), .B1(n1104), .C0(n4380), 
        .C1(n3700), .Y(n1710) );
  AOI22X1TS U2955 ( .A0(n4286), .A1(n3681), .B0(n4119), .B1(n3664), .Y(n1711)
         );
  AOI222XLTS U2956 ( .A0(n4476), .A1(n3736), .B0(n531), .B1(n3719), .C0(n4383), 
        .C1(n3700), .Y(n1712) );
  AOI22X1TS U2957 ( .A0(n4241), .A1(n3677), .B0(n4074), .B1(n3668), .Y(n1681)
         );
  AOI222XLTS U2958 ( .A0(n4438), .A1(n3725), .B0(n539), .B1(n3717), .C0(n4338), 
        .C1(n3696), .Y(n1682) );
  AOI22X1TS U2959 ( .A0(n4034), .A1(n3677), .B0(n4071), .B1(n3668), .Y(n1116)
         );
  AOI222XLTS U2960 ( .A0(n4538), .A1(n3725), .B0(n14), .B1(n3717), .C0(n4185), 
        .C1(n3696), .Y(n1117) );
  AOI22X1TS U2961 ( .A0(n4031), .A1(n3676), .B0(n4068), .B1(n3668), .Y(n1114)
         );
  AOI222XLTS U2962 ( .A0(n4536), .A1(n3724), .B0(n36), .B1(n3717), .C0(n4182), 
        .C1(n3696), .Y(n1115) );
  AOI22X1TS U2963 ( .A0(n4025), .A1(n3676), .B0(n4062), .B1(n3669), .Y(n1110)
         );
  AOI222XLTS U2964 ( .A0(n4529), .A1(n3724), .B0(n26), .B1(n3718), .C0(n4176), 
        .C1(n3696), .Y(n1111) );
  AOI22X1TS U2965 ( .A0(n4028), .A1(n3676), .B0(n4065), .B1(n3669), .Y(n1112)
         );
  AOI222XLTS U2966 ( .A0(n4533), .A1(n3724), .B0(n31), .B1(n3718), .C0(n4179), 
        .C1(n3695), .Y(n1113) );
  AOI22X1TS U2967 ( .A0(n4022), .A1(n3676), .B0(n4059), .B1(n3669), .Y(n1108)
         );
  AOI222XLTS U2968 ( .A0(n4528), .A1(n3724), .B0(n21), .B1(n3718), .C0(n4173), 
        .C1(n3695), .Y(n1109) );
  AOI22X1TS U2969 ( .A0(n4019), .A1(n3682), .B0(n4056), .B1(n3669), .Y(n1101)
         );
  AOI222XLTS U2970 ( .A0(n4525), .A1(n3726), .B0(n16), .B1(n3718), .C0(n4170), 
        .C1(n3700), .Y(n1102) );
  AOI22X1TS U2971 ( .A0(n3989), .A1(n3686), .B0(n4050), .B1(n3659), .Y(n1827)
         );
  AOI222XLTS U2972 ( .A0(n4213), .A1(n3730), .B0(n37), .B1(n3722), .C0(n3948), 
        .C1(n3709), .Y(n1828) );
  AOI22X1TS U2973 ( .A0(n3977), .A1(n3685), .B0(n4038), .B1(n3660), .Y(n1819)
         );
  AOI222XLTS U2974 ( .A0(n4203), .A1(n3729), .B0(n17), .B1(n3710), .C0(n3936), 
        .C1(n3709), .Y(n1820) );
  AOI22X1TS U2975 ( .A0(n3992), .A1(n3686), .B0(n4053), .B1(n3659), .Y(n1829)
         );
  AOI222XLTS U2976 ( .A0(n4215), .A1(n3730), .B0(n42), .B1(n3722), .C0(n3951), 
        .C1(n3695), .Y(n1830) );
  AOI22X1TS U2977 ( .A0(n3986), .A1(n3686), .B0(n4047), .B1(n3659), .Y(n1825)
         );
  AOI222XLTS U2978 ( .A0(n4210), .A1(n3730), .B0(n32), .B1(n3722), .C0(n3945), 
        .C1(n3704), .Y(n1826) );
  AOI22X1TS U2979 ( .A0(n3983), .A1(n3686), .B0(n4044), .B1(n3659), .Y(n1823)
         );
  AOI222XLTS U2980 ( .A0(n4208), .A1(n3730), .B0(n27), .B1(n3719), .C0(n3942), 
        .C1(n3704), .Y(n1824) );
  AOI22X1TS U2981 ( .A0(n3980), .A1(n3685), .B0(n4041), .B1(n3660), .Y(n1821)
         );
  AOI222XLTS U2982 ( .A0(n4205), .A1(n3729), .B0(n22), .B1(n3710), .C0(n3939), 
        .C1(n3703), .Y(n1822) );
  AOI22X1TS U2983 ( .A0(n4334), .A1(n3685), .B0(n4167), .B1(n3660), .Y(n1743)
         );
  AOI222XLTS U2984 ( .A0(n4521), .A1(n3729), .B0(n511), .B1(n3710), .C0(n4434), 
        .C1(n1105), .Y(n1744) );
  AOI22X1TS U2985 ( .A0(n4331), .A1(n3685), .B0(n4164), .B1(n3660), .Y(n1741)
         );
  AOI222XLTS U2986 ( .A0(n4519), .A1(n3729), .B0(n507), .B1(n3710), .C0(n4430), 
        .C1(n3705), .Y(n1742) );
  AOI22X1TS U2987 ( .A0(n4328), .A1(n3684), .B0(n4161), .B1(n3661), .Y(n1739)
         );
  AOI222XLTS U2988 ( .A0(n4516), .A1(n3728), .B0(n513), .B1(n3711), .C0(n4427), 
        .C1(n3705), .Y(n1740) );
  AOI22X1TS U2989 ( .A0(n4325), .A1(n3684), .B0(n4158), .B1(n3661), .Y(n1737)
         );
  AOI222XLTS U2990 ( .A0(n4515), .A1(n3728), .B0(n477), .B1(n3711), .C0(n4422), 
        .C1(n3707), .Y(n1738) );
  AOI22X1TS U2991 ( .A0(n4322), .A1(n3684), .B0(n4155), .B1(n3661), .Y(n1735)
         );
  AOI222XLTS U2992 ( .A0(n4511), .A1(n3728), .B0(n479), .B1(n3711), .C0(n4419), 
        .C1(n3709), .Y(n1736) );
  AOI22X1TS U2993 ( .A0(n4319), .A1(n3684), .B0(n4152), .B1(n3661), .Y(n1733)
         );
  AOI222XLTS U2994 ( .A0(n4510), .A1(n3728), .B0(n515), .B1(n3711), .C0(n4416), 
        .C1(n3709), .Y(n1734) );
  AOI22X1TS U2995 ( .A0(n4316), .A1(n3683), .B0(n4149), .B1(n3662), .Y(n1731)
         );
  AOI222XLTS U2996 ( .A0(n4506), .A1(n3727), .B0(n517), .B1(n3712), .C0(n4413), 
        .C1(n3707), .Y(n1732) );
  AOI22X1TS U2997 ( .A0(n4313), .A1(n3683), .B0(n4146), .B1(n3662), .Y(n1729)
         );
  AOI222XLTS U2998 ( .A0(n4503), .A1(n3727), .B0(n519), .B1(n3712), .C0(n4410), 
        .C1(n3706), .Y(n1730) );
  AOI22X1TS U2999 ( .A0(n4310), .A1(n3683), .B0(n4143), .B1(n3662), .Y(n1727)
         );
  AOI222XLTS U3000 ( .A0(n4501), .A1(n3727), .B0(n481), .B1(n3712), .C0(n4407), 
        .C1(n3702), .Y(n1728) );
  AOI22X1TS U3001 ( .A0(n4307), .A1(n3683), .B0(n4140), .B1(n3662), .Y(n1725)
         );
  AOI222XLTS U3002 ( .A0(n4497), .A1(n3727), .B0(n521), .B1(n3712), .C0(n4404), 
        .C1(n3702), .Y(n1726) );
  AOI22X1TS U3003 ( .A0(n4304), .A1(n3682), .B0(n4137), .B1(n3663), .Y(n1723)
         );
  AOI222XLTS U3004 ( .A0(n4494), .A1(n3726), .B0(n523), .B1(n3713), .C0(n4401), 
        .C1(n3702), .Y(n1724) );
  AOI22X1TS U3005 ( .A0(n4301), .A1(n3682), .B0(n4134), .B1(n3663), .Y(n1721)
         );
  AOI222XLTS U3006 ( .A0(n4493), .A1(n3726), .B0(n483), .B1(n3713), .C0(n4398), 
        .C1(n3702), .Y(n1722) );
  AOI22X1TS U3007 ( .A0(n4298), .A1(n3682), .B0(n4131), .B1(n3663), .Y(n1719)
         );
  AOI222XLTS U3008 ( .A0(n4488), .A1(n3726), .B0(n525), .B1(n3713), .C0(n4395), 
        .C1(n3701), .Y(n1720) );
  AOI22X1TS U3009 ( .A0(n4295), .A1(n3681), .B0(n4128), .B1(n3663), .Y(n1717)
         );
  AOI222XLTS U3010 ( .A0(n4485), .A1(n3735), .B0(n527), .B1(n3713), .C0(n4392), 
        .C1(n3701), .Y(n1718) );
  AOI22X1TS U3011 ( .A0(n4292), .A1(n3681), .B0(n4125), .B1(n3664), .Y(n1715)
         );
  AOI222XLTS U3012 ( .A0(n4483), .A1(n3740), .B0(n529), .B1(n3721), .C0(n4389), 
        .C1(n3701), .Y(n1716) );
  AOI22X1TS U3013 ( .A0(n4289), .A1(n3681), .B0(n4122), .B1(n3664), .Y(n1713)
         );
  AOI222XLTS U3014 ( .A0(n4482), .A1(n1103), .B0(n509), .B1(n3720), .C0(n4386), 
        .C1(n3701), .Y(n1714) );
  AOI22X1TS U3015 ( .A0(n4277), .A1(n3680), .B0(n4110), .B1(n3665), .Y(n1705)
         );
  AOI222XLTS U3016 ( .A0(n4467), .A1(n3738), .B0(n485), .B1(n3714), .C0(n4374), 
        .C1(n3699), .Y(n1706) );
  AOI22X1TS U3017 ( .A0(n4274), .A1(n3680), .B0(n4107), .B1(n3665), .Y(n1703)
         );
  AOI222XLTS U3018 ( .A0(n4465), .A1(n3733), .B0(n487), .B1(n3714), .C0(n4371), 
        .C1(n3699), .Y(n1704) );
  AOI22X1TS U3019 ( .A0(n4271), .A1(n3679), .B0(n4104), .B1(n3665), .Y(n1701)
         );
  AOI222XLTS U3020 ( .A0(n4464), .A1(n3737), .B0(n489), .B1(n3714), .C0(n4368), 
        .C1(n3699), .Y(n1702) );
  AOI22X1TS U3021 ( .A0(n4268), .A1(n3679), .B0(n4101), .B1(n3666), .Y(n1699)
         );
  AOI222XLTS U3022 ( .A0(n4462), .A1(n3737), .B0(n491), .B1(n3715), .C0(n4365), 
        .C1(n3699), .Y(n1700) );
  AOI22X1TS U3023 ( .A0(n4265), .A1(n3679), .B0(n4098), .B1(n3666), .Y(n1697)
         );
  AOI222XLTS U3024 ( .A0(n4457), .A1(n3738), .B0(n493), .B1(n3715), .C0(n4362), 
        .C1(n3698), .Y(n1698) );
  AOI22X1TS U3025 ( .A0(n4262), .A1(n3679), .B0(n4095), .B1(n3666), .Y(n1695)
         );
  AOI222XLTS U3026 ( .A0(n4456), .A1(n3736), .B0(n495), .B1(n3715), .C0(n4359), 
        .C1(n3698), .Y(n1696) );
  AOI22X1TS U3027 ( .A0(n4259), .A1(n3678), .B0(n4092), .B1(n3666), .Y(n1693)
         );
  AOI222XLTS U3028 ( .A0(n4453), .A1(n3734), .B0(n497), .B1(n3715), .C0(n4356), 
        .C1(n3698), .Y(n1694) );
  AOI22X1TS U3029 ( .A0(n4256), .A1(n3678), .B0(n4089), .B1(n3667), .Y(n1691)
         );
  AOI222XLTS U3030 ( .A0(n4451), .A1(n3737), .B0(n499), .B1(n3716), .C0(n4353), 
        .C1(n3698), .Y(n1692) );
  AOI22X1TS U3031 ( .A0(n4253), .A1(n3678), .B0(n4086), .B1(n3667), .Y(n1689)
         );
  AOI222XLTS U3032 ( .A0(n4449), .A1(n3734), .B0(n501), .B1(n3716), .C0(n4350), 
        .C1(n3697), .Y(n1690) );
  AOI22X1TS U3033 ( .A0(n4250), .A1(n3678), .B0(n4083), .B1(n3667), .Y(n1687)
         );
  AOI222XLTS U3034 ( .A0(n4445), .A1(n3737), .B0(n503), .B1(n3716), .C0(n4347), 
        .C1(n3697), .Y(n1688) );
  AOI22X1TS U3035 ( .A0(n4247), .A1(n3677), .B0(n4080), .B1(n3667), .Y(n1685)
         );
  AOI222XLTS U3036 ( .A0(n4442), .A1(n3725), .B0(n505), .B1(n3716), .C0(n4344), 
        .C1(n3697), .Y(n1686) );
  AOI22X1TS U3037 ( .A0(n4244), .A1(n3677), .B0(n4077), .B1(n3668), .Y(n1683)
         );
  AOI222XLTS U3038 ( .A0(n4439), .A1(n3725), .B0(n537), .B1(n3717), .C0(n4341), 
        .C1(n3697), .Y(n1684) );
  AOI22X1TS U3039 ( .A0(n4469), .A1(n3645), .B0(n4110), .B1(n3802), .Y(n1641)
         );
  AOI222XLTS U3040 ( .A0(n4373), .A1(n3789), .B0(n486), .B1(n3631), .C0(n4278), 
        .C1(n3621), .Y(n1642) );
  AOI22X1TS U3041 ( .A0(n4470), .A1(n3645), .B0(n4113), .B1(n3800), .Y(n1643)
         );
  AOI222XLTS U3042 ( .A0(n4376), .A1(n3789), .B0(n536), .B1(n3630), .C0(n4281), 
        .C1(n3621), .Y(n1644) );
  AOI22X1TS U3043 ( .A0(n4474), .A1(n3645), .B0(n4116), .B1(n3801), .Y(n1645)
         );
  AOI222XLTS U3044 ( .A0(n4379), .A1(n3789), .B0(n534), .B1(n3630), .C0(n4284), 
        .C1(n3621), .Y(n1646) );
  AOI22X1TS U3045 ( .A0(n4478), .A1(n3645), .B0(n4119), .B1(n3811), .Y(n1647)
         );
  AOI222XLTS U3046 ( .A0(n4382), .A1(n3789), .B0(n532), .B1(n3631), .C0(n4287), 
        .C1(n3621), .Y(n1648) );
  AOI22X1TS U3047 ( .A0(n4481), .A1(n3646), .B0(n4122), .B1(n3799), .Y(n1649)
         );
  AOI222XLTS U3048 ( .A0(n4385), .A1(n3790), .B0(n510), .B1(n3630), .C0(n4290), 
        .C1(n3620), .Y(n1650) );
  AOI22X1TS U3049 ( .A0(n4484), .A1(n3646), .B0(n4125), .B1(n3810), .Y(n1651)
         );
  AOI222XLTS U3050 ( .A0(n4388), .A1(n3790), .B0(n530), .B1(n3629), .C0(n4293), 
        .C1(n3622), .Y(n1652) );
  AOI22X1TS U3051 ( .A0(n4487), .A1(n3646), .B0(n4128), .B1(n3800), .Y(n1653)
         );
  AOI222XLTS U3052 ( .A0(n4391), .A1(n3790), .B0(n528), .B1(n3630), .C0(n4296), 
        .C1(n3618), .Y(n1654) );
  AOI22X1TS U3053 ( .A0(n4490), .A1(n3646), .B0(n4131), .B1(n3810), .Y(n1655)
         );
  AOI222XLTS U3054 ( .A0(n4394), .A1(n3790), .B0(n526), .B1(n3629), .C0(n4299), 
        .C1(n3618), .Y(n1656) );
  AOI22X1TS U3055 ( .A0(n4492), .A1(n3647), .B0(n4134), .B1(n3800), .Y(n1657)
         );
  AOI222XLTS U3056 ( .A0(n4397), .A1(n3791), .B0(n484), .B1(n3629), .C0(n4302), 
        .C1(n3618), .Y(n1658) );
  AOI22X1TS U3057 ( .A0(n4496), .A1(n3647), .B0(n4137), .B1(n3799), .Y(n1659)
         );
  AOI222XLTS U3058 ( .A0(n4400), .A1(n3791), .B0(n524), .B1(n3629), .C0(n4305), 
        .C1(n3618), .Y(n1660) );
  AOI22X1TS U3059 ( .A0(n4498), .A1(n3647), .B0(n4140), .B1(n3809), .Y(n1661)
         );
  AOI222XLTS U3060 ( .A0(n4403), .A1(n3791), .B0(n522), .B1(n3628), .C0(n4308), 
        .C1(n3620), .Y(n1662) );
  AOI22X1TS U3061 ( .A0(n4500), .A1(n3647), .B0(n4143), .B1(n3799), .Y(n1663)
         );
  AOI222XLTS U3062 ( .A0(n4406), .A1(n3791), .B0(n482), .B1(n3628), .C0(n4311), 
        .C1(n3620), .Y(n1664) );
  AOI22X1TS U3063 ( .A0(n4502), .A1(n3648), .B0(n4146), .B1(n3799), .Y(n1665)
         );
  AOI222XLTS U3064 ( .A0(n4409), .A1(n3792), .B0(n520), .B1(n3628), .C0(n4314), 
        .C1(n3626), .Y(n1666) );
  AOI22X1TS U3065 ( .A0(n4507), .A1(n3648), .B0(n4149), .B1(n3809), .Y(n1667)
         );
  AOI222XLTS U3066 ( .A0(n4412), .A1(n3792), .B0(n518), .B1(n3638), .C0(n4317), 
        .C1(n3622), .Y(n1668) );
  AOI22X1TS U3067 ( .A0(n4509), .A1(n3648), .B0(n4152), .B1(n3808), .Y(n1669)
         );
  AOI222XLTS U3068 ( .A0(n4415), .A1(n3792), .B0(n516), .B1(n3631), .C0(n4320), 
        .C1(n3619), .Y(n1670) );
  AOI22X1TS U3069 ( .A0(n4512), .A1(n3648), .B0(n4155), .B1(n3808), .Y(n1671)
         );
  AOI222XLTS U3070 ( .A0(n4418), .A1(n3792), .B0(n480), .B1(n3628), .C0(n4323), 
        .C1(n3619), .Y(n1672) );
  AOI22X1TS U3071 ( .A0(n4514), .A1(n3649), .B0(n4158), .B1(n3807), .Y(n1673)
         );
  AOI222XLTS U3072 ( .A0(n4421), .A1(n3796), .B0(n478), .B1(n3637), .C0(n4326), 
        .C1(n3619), .Y(n1674) );
  AOI22X1TS U3073 ( .A0(n4517), .A1(n3649), .B0(n4161), .B1(n3811), .Y(n1675)
         );
  AOI222XLTS U3074 ( .A0(n4426), .A1(n3796), .B0(n514), .B1(n3636), .C0(n4329), 
        .C1(n3619), .Y(n1676) );
  AOI22X1TS U3075 ( .A0(n4334), .A1(n3537), .B0(n4167), .B1(n3915), .Y(n1614)
         );
  AOI222XLTS U3076 ( .A0(n4521), .A1(n3583), .B0(n512), .B1(n3562), .C0(n4434), 
        .C1(n3554), .Y(n1615) );
  AOI22X1TS U3077 ( .A0(n4289), .A1(n3533), .B0(n4122), .B1(n3911), .Y(n1584)
         );
  AOI222XLTS U3078 ( .A0(n4482), .A1(n3581), .B0(n509), .B1(n1138), .C0(n4386), 
        .C1(n3561), .Y(n1585) );
  AOI22X1TS U3079 ( .A0(n4286), .A1(n3533), .B0(n4119), .B1(n3911), .Y(n1582)
         );
  AOI222XLTS U3080 ( .A0(n4476), .A1(n3581), .B0(n531), .B1(n3564), .C0(n4383), 
        .C1(n3552), .Y(n1583) );
  AOI22X1TS U3081 ( .A0(n4274), .A1(n3532), .B0(n4107), .B1(n3920), .Y(n1574)
         );
  AOI222XLTS U3082 ( .A0(n4465), .A1(n3580), .B0(n488), .B1(n3566), .C0(n4371), 
        .C1(n3551), .Y(n1575) );
  AOI22X1TS U3083 ( .A0(n4244), .A1(n3529), .B0(n4077), .B1(n3921), .Y(n1554)
         );
  AOI222XLTS U3084 ( .A0(n4439), .A1(n3577), .B0(n538), .B1(n3567), .C0(n4341), 
        .C1(n3549), .Y(n1555) );
  AOI22X1TS U3085 ( .A0(n3992), .A1(n3540), .B0(n4053), .B1(n3916), .Y(n1882)
         );
  AOI222XLTS U3086 ( .A0(n4215), .A1(n3584), .B0(n3568), .B1(n41), .C0(n3951), 
        .C1(n3548), .Y(n1883) );
  OAI211X1TS U3087 ( .A0(n3605), .A1(n805), .B0(n1878), .C0(n1879), .Y(n2531)
         );
  AOI22X1TS U3088 ( .A0(n3986), .A1(n3540), .B0(n4047), .B1(n3916), .Y(n1878)
         );
  AOI222XLTS U3089 ( .A0(destinationAddressIn_SOUTH[3]), .A1(n3584), .B0(n3570), .B1(n33), .C0(n3945), .C1(n3553), .Y(n1879) );
  OAI211X1TS U3090 ( .A0(n3605), .A1(n804), .B0(n1876), .C0(n1877), .Y(n2532)
         );
  AOI22X1TS U3091 ( .A0(n3983), .A1(n3541), .B0(n4044), .B1(n3916), .Y(n1876)
         );
  AOI222XLTS U3092 ( .A0(n4208), .A1(n3584), .B0(n3570), .B1(n28), .C0(n3942), 
        .C1(n3553), .Y(n1877) );
  OAI211X1TS U3093 ( .A0(n3605), .A1(n803), .B0(n1874), .C0(n1875), .Y(n2533)
         );
  AOI22X1TS U3094 ( .A0(n3980), .A1(n3537), .B0(n4041), .B1(n3915), .Y(n1874)
         );
  AOI222XLTS U3095 ( .A0(n4205), .A1(n3583), .B0(n3570), .B1(n23), .C0(n3939), 
        .C1(n3553), .Y(n1875) );
  OAI211X1TS U3096 ( .A0(n3605), .A1(n802), .B0(n1872), .C0(n1873), .Y(n2534)
         );
  AOI22X1TS U3097 ( .A0(n3977), .A1(n3537), .B0(n4038), .B1(n3915), .Y(n1872)
         );
  AOI222XLTS U3098 ( .A0(n4203), .A1(n3583), .B0(n3569), .B1(n18), .C0(n3936), 
        .C1(n3553), .Y(n1873) );
  AOI22X1TS U3099 ( .A0(n4331), .A1(n3537), .B0(n4164), .B1(n3915), .Y(n1612)
         );
  AOI222XLTS U3100 ( .A0(n4519), .A1(n3583), .B0(n508), .B1(n1138), .C0(n4430), 
        .C1(n3557), .Y(n1613) );
  AOI22X1TS U3101 ( .A0(n4328), .A1(n3536), .B0(n4161), .B1(n3914), .Y(n1610)
         );
  AOI222XLTS U3102 ( .A0(n4516), .A1(n3582), .B0(n513), .B1(n3562), .C0(n4427), 
        .C1(n3555), .Y(n1611) );
  AOI22X1TS U3103 ( .A0(n4325), .A1(n3536), .B0(n4158), .B1(n3914), .Y(n1608)
         );
  AOI222XLTS U3104 ( .A0(n4515), .A1(n3582), .B0(n477), .B1(n3574), .C0(n4422), 
        .C1(n3557), .Y(n1609) );
  AOI22X1TS U3105 ( .A0(n4322), .A1(n3536), .B0(n4155), .B1(n3914), .Y(n1606)
         );
  AOI222XLTS U3106 ( .A0(n4511), .A1(n3582), .B0(n479), .B1(n3573), .C0(n4419), 
        .C1(n3554), .Y(n1607) );
  AOI22X1TS U3107 ( .A0(n4319), .A1(n3536), .B0(n4152), .B1(n3914), .Y(n1604)
         );
  AOI222XLTS U3108 ( .A0(n4510), .A1(n3582), .B0(n515), .B1(n3563), .C0(n4416), 
        .C1(n3554), .Y(n1605) );
  AOI22X1TS U3109 ( .A0(n4316), .A1(n3535), .B0(n4149), .B1(n3913), .Y(n1602)
         );
  AOI222XLTS U3110 ( .A0(n4506), .A1(n3589), .B0(n517), .B1(n3563), .C0(n4413), 
        .C1(n1139), .Y(n1603) );
  AOI22X1TS U3111 ( .A0(n4313), .A1(n3535), .B0(n4146), .B1(n3913), .Y(n1600)
         );
  AOI222XLTS U3112 ( .A0(n4503), .A1(n3590), .B0(n519), .B1(n3562), .C0(n4410), 
        .C1(n3558), .Y(n1601) );
  AOI22X1TS U3113 ( .A0(n4310), .A1(n3535), .B0(n4143), .B1(n3913), .Y(n1598)
         );
  AOI222XLTS U3114 ( .A0(n4501), .A1(n3591), .B0(n481), .B1(n3564), .C0(n4407), 
        .C1(n3560), .Y(n1599) );
  AOI22X1TS U3115 ( .A0(n4307), .A1(n3535), .B0(n4140), .B1(n3913), .Y(n1596)
         );
  AOI222XLTS U3116 ( .A0(n4497), .A1(n3590), .B0(n521), .B1(n3564), .C0(n4404), 
        .C1(n3556), .Y(n1597) );
  AOI22X1TS U3117 ( .A0(n4304), .A1(n3534), .B0(n4137), .B1(n3912), .Y(n1594)
         );
  AOI222XLTS U3118 ( .A0(n4494), .A1(n3592), .B0(n523), .B1(n3562), .C0(n4401), 
        .C1(n3560), .Y(n1595) );
  AOI22X1TS U3119 ( .A0(n4301), .A1(n3534), .B0(n4134), .B1(n3912), .Y(n1592)
         );
  AOI222XLTS U3120 ( .A0(n4493), .A1(n3592), .B0(n483), .B1(n3564), .C0(n4398), 
        .C1(n3556), .Y(n1593) );
  AOI22X1TS U3121 ( .A0(n4298), .A1(n3534), .B0(n4131), .B1(n3912), .Y(n1590)
         );
  AOI222XLTS U3122 ( .A0(n4488), .A1(n3589), .B0(n525), .B1(n3573), .C0(n4395), 
        .C1(n3561), .Y(n1591) );
  AOI22X1TS U3123 ( .A0(n4295), .A1(n3533), .B0(n4128), .B1(n3912), .Y(n1588)
         );
  AOI222XLTS U3124 ( .A0(n4485), .A1(n3581), .B0(n527), .B1(n3563), .C0(n4392), 
        .C1(n3554), .Y(n1589) );
  AOI22X1TS U3125 ( .A0(n4292), .A1(n3533), .B0(n4125), .B1(n3911), .Y(n1586)
         );
  AOI222XLTS U3126 ( .A0(n4483), .A1(n3581), .B0(n529), .B1(n3572), .C0(n4389), 
        .C1(n3555), .Y(n1587) );
  AOI22X1TS U3127 ( .A0(n4283), .A1(n3532), .B0(n4116), .B1(n3911), .Y(n1580)
         );
  AOI222XLTS U3128 ( .A0(n4475), .A1(n3580), .B0(n533), .B1(n3563), .C0(n4380), 
        .C1(n3552), .Y(n1581) );
  AOI22X1TS U3129 ( .A0(n4280), .A1(n3532), .B0(n4113), .B1(n3917), .Y(n1578)
         );
  AOI222XLTS U3130 ( .A0(n4471), .A1(n3580), .B0(n535), .B1(n3565), .C0(n4377), 
        .C1(n3552), .Y(n1579) );
  AOI22X1TS U3131 ( .A0(n4277), .A1(n3532), .B0(n4110), .B1(n724), .Y(n1576)
         );
  AOI222XLTS U3132 ( .A0(n4467), .A1(n3580), .B0(n485), .B1(n3571), .C0(n4374), 
        .C1(n3551), .Y(n1577) );
  AOI22X1TS U3133 ( .A0(n4271), .A1(n3531), .B0(n4104), .B1(n3920), .Y(n1572)
         );
  AOI222XLTS U3134 ( .A0(n4464), .A1(n3579), .B0(n490), .B1(n3566), .C0(n4368), 
        .C1(n3551), .Y(n1573) );
  AOI22X1TS U3135 ( .A0(n4268), .A1(n3534), .B0(n4101), .B1(n3917), .Y(n1570)
         );
  AOI222XLTS U3136 ( .A0(n4462), .A1(n3587), .B0(n492), .B1(n3565), .C0(n4365), 
        .C1(n3551), .Y(n1571) );
  AOI22X1TS U3137 ( .A0(n4265), .A1(n3531), .B0(n4098), .B1(n3919), .Y(n1568)
         );
  AOI222XLTS U3138 ( .A0(n4457), .A1(n3579), .B0(n494), .B1(n3566), .C0(n4362), 
        .C1(n3550), .Y(n1569) );
  AOI22X1TS U3139 ( .A0(n4262), .A1(n3531), .B0(n4095), .B1(n724), .Y(n1566)
         );
  AOI222XLTS U3140 ( .A0(n4456), .A1(n3579), .B0(n496), .B1(n3565), .C0(n4359), 
        .C1(n3550), .Y(n1567) );
  AOI22X1TS U3141 ( .A0(n4259), .A1(n3531), .B0(n4092), .B1(n1748), .Y(n1564)
         );
  AOI222XLTS U3142 ( .A0(n4453), .A1(n3579), .B0(n498), .B1(n3565), .C0(n4356), 
        .C1(n3552), .Y(n1565) );
  AOI22X1TS U3143 ( .A0(n4256), .A1(n3530), .B0(n4089), .B1(n3910), .Y(n1562)
         );
  AOI222XLTS U3144 ( .A0(n4451), .A1(n3578), .B0(n500), .B1(n3567), .C0(n4353), 
        .C1(n3550), .Y(n1563) );
  AOI22X1TS U3145 ( .A0(n4253), .A1(n3530), .B0(n4086), .B1(n3910), .Y(n1560)
         );
  AOI222XLTS U3146 ( .A0(n4449), .A1(n3578), .B0(n502), .B1(n3567), .C0(n4350), 
        .C1(n3550), .Y(n1561) );
  AOI22X1TS U3147 ( .A0(n4250), .A1(n3530), .B0(n4083), .B1(n3910), .Y(n1558)
         );
  AOI222XLTS U3148 ( .A0(n4445), .A1(n3578), .B0(n504), .B1(n3566), .C0(n4347), 
        .C1(n3549), .Y(n1559) );
  AOI22X1TS U3149 ( .A0(n4247), .A1(n3530), .B0(n4080), .B1(n3910), .Y(n1556)
         );
  AOI222XLTS U3150 ( .A0(n4442), .A1(n3578), .B0(n506), .B1(n3567), .C0(n4344), 
        .C1(n3549), .Y(n1557) );
  AOI22X1TS U3151 ( .A0(n4241), .A1(n3529), .B0(n4074), .B1(n3918), .Y(n1552)
         );
  AOI222XLTS U3152 ( .A0(n4438), .A1(n3577), .B0(n540), .B1(n3572), .C0(n4338), 
        .C1(n3549), .Y(n1553) );
  AOI22X1TS U3153 ( .A0(n4463), .A1(n3644), .B0(n4104), .B1(n3801), .Y(n1637)
         );
  AOI222XLTS U3154 ( .A0(n4367), .A1(n3788), .B0(n489), .B1(n3634), .C0(n4272), 
        .C1(n3625), .Y(n1638) );
  AOI22X1TS U3155 ( .A0(n4454), .A1(n3643), .B0(n4092), .B1(n3803), .Y(n1629)
         );
  AOI222XLTS U3156 ( .A0(n4355), .A1(n3787), .B0(n497), .B1(n3633), .C0(n4260), 
        .C1(n3627), .Y(n1630) );
  AOI22X1TS U3157 ( .A0(n4523), .A1(n3649), .B0(n4167), .B1(n3811), .Y(n1679)
         );
  AOI222XLTS U3158 ( .A0(n4433), .A1(n3794), .B0(n511), .B1(n3634), .C0(n4335), 
        .C1(n3616), .Y(n1680) );
  AOI22X1TS U3159 ( .A0(n4518), .A1(n3649), .B0(n4164), .B1(n740), .Y(n1677)
         );
  AOI222XLTS U3160 ( .A0(n4429), .A1(n3795), .B0(n507), .B1(n3638), .C0(n4332), 
        .C1(n3625), .Y(n1678) );
  AOI22X1TS U3161 ( .A0(n4466), .A1(n3644), .B0(n4107), .B1(n3802), .Y(n1639)
         );
  AOI222XLTS U3162 ( .A0(n4370), .A1(n3788), .B0(n487), .B1(n3631), .C0(n4275), 
        .C1(n3623), .Y(n1640) );
  AOI22X1TS U3163 ( .A0(n4461), .A1(n3644), .B0(n4101), .B1(n3802), .Y(n1635)
         );
  AOI222XLTS U3164 ( .A0(n4364), .A1(n3788), .B0(n491), .B1(n3632), .C0(n4269), 
        .C1(n3624), .Y(n1636) );
  AOI22X1TS U3165 ( .A0(n4458), .A1(n3644), .B0(n4098), .B1(n3801), .Y(n1633)
         );
  AOI222XLTS U3166 ( .A0(n4361), .A1(n3788), .B0(n493), .B1(n3632), .C0(n4266), 
        .C1(n3622), .Y(n1634) );
  AOI22X1TS U3167 ( .A0(n4455), .A1(n3643), .B0(n4095), .B1(n3801), .Y(n1631)
         );
  AOI222XLTS U3168 ( .A0(n4358), .A1(n3787), .B0(n495), .B1(n3632), .C0(n4263), 
        .C1(n3624), .Y(n1632) );
  AOI22X1TS U3169 ( .A0(n4452), .A1(n3643), .B0(n4089), .B1(n3803), .Y(n1627)
         );
  AOI222XLTS U3170 ( .A0(n4352), .A1(n3787), .B0(n499), .B1(n3632), .C0(n4257), 
        .C1(n3617), .Y(n1628) );
  AOI22X1TS U3171 ( .A0(n4444), .A1(n3642), .B0(n4083), .B1(n3803), .Y(n1623)
         );
  AOI222XLTS U3172 ( .A0(n4346), .A1(n3786), .B0(n503), .B1(n3634), .C0(n4251), 
        .C1(n3617), .Y(n1624) );
  AOI22X1TS U3173 ( .A0(n4443), .A1(n3642), .B0(n4080), .B1(n3803), .Y(n1621)
         );
  AOI222XLTS U3174 ( .A0(n4343), .A1(n3786), .B0(n505), .B1(n3633), .C0(n4248), 
        .C1(n3616), .Y(n1622) );
  AOI22X1TS U3175 ( .A0(n4447), .A1(n3643), .B0(n4086), .B1(n3802), .Y(n1625)
         );
  AOI222XLTS U3176 ( .A0(n4349), .A1(n3787), .B0(n501), .B1(n3633), .C0(n4254), 
        .C1(n3617), .Y(n1626) );
  AOI22X1TS U3177 ( .A0(n4418), .A1(n3273), .B0(n4155), .B1(n3874), .Y(n1350)
         );
  AOI222XLTS U3178 ( .A0(n4512), .A1(n3315), .B0(n479), .B1(n3295), .C0(n4323), 
        .C1(n3286), .Y(n1351) );
  AOI22X1TS U3179 ( .A0(n4403), .A1(n3268), .B0(n4140), .B1(n3878), .Y(n1340)
         );
  AOI222XLTS U3180 ( .A0(n4498), .A1(n3321), .B0(n521), .B1(n3298), .C0(n4308), 
        .C1(n3285), .Y(n1341) );
  AOI22X1TS U3181 ( .A0(n4397), .A1(n3267), .B0(n4134), .B1(n3873), .Y(n1336)
         );
  AOI222XLTS U3182 ( .A0(n4492), .A1(n3321), .B0(n483), .B1(n3298), .C0(n4302), 
        .C1(n3285), .Y(n1337) );
  AOI22X1TS U3183 ( .A0(n4394), .A1(n3267), .B0(n4131), .B1(n3873), .Y(n1334)
         );
  AOI222XLTS U3184 ( .A0(n4490), .A1(n3321), .B0(n525), .B1(n3299), .C0(n4299), 
        .C1(n3284), .Y(n1335) );
  AOI22X1TS U3185 ( .A0(n4367), .A1(n3264), .B0(n4104), .B1(n3877), .Y(n1316)
         );
  AOI222XLTS U3186 ( .A0(dataIn_SOUTH[10]), .A1(n3312), .B0(n489), .B1(n3303), 
        .C0(n4272), .C1(n3282), .Y(n1317) );
  AOI22X1TS U3187 ( .A0(n4361), .A1(n3264), .B0(n4098), .B1(n3871), .Y(n1312)
         );
  AOI222XLTS U3188 ( .A0(n4458), .A1(n3312), .B0(n493), .B1(n3303), .C0(n4266), 
        .C1(n3291), .Y(n1313) );
  AOI22X1TS U3189 ( .A0(n4352), .A1(n3263), .B0(n4089), .B1(n3870), .Y(n1306)
         );
  AOI222XLTS U3190 ( .A0(n4452), .A1(n3311), .B0(n499), .B1(n3302), .C0(n4257), 
        .C1(n3291), .Y(n1307) );
  AOI22X1TS U3191 ( .A0(n4343), .A1(n3263), .B0(n4080), .B1(n3870), .Y(n1300)
         );
  AOI222XLTS U3192 ( .A0(n4443), .A1(n3311), .B0(n505), .B1(n3302), .C0(n4248), 
        .C1(n3291), .Y(n1301) );
  AOI22X1TS U3193 ( .A0(n3950), .A1(n3269), .B0(n4053), .B1(n3879), .Y(n1974)
         );
  AOI222XLTS U3194 ( .A0(n4216), .A1(n3317), .B0(n3306), .B1(n43), .C0(n3993), 
        .C1(n3281), .Y(n1975) );
  AOI22X1TS U3195 ( .A0(n3944), .A1(n3269), .B0(n4047), .B1(n730), .Y(n1970)
         );
  AOI222XLTS U3196 ( .A0(n4211), .A1(n3317), .B0(n3300), .B1(n34), .C0(n3987), 
        .C1(n3293), .Y(n1971) );
  AOI22X1TS U3197 ( .A0(n3941), .A1(n3269), .B0(n4044), .B1(n3879), .Y(n1968)
         );
  AOI222XLTS U3198 ( .A0(n4209), .A1(n3317), .B0(n3300), .B1(n29), .C0(n3984), 
        .C1(n3292), .Y(n1969) );
  AOI22X1TS U3199 ( .A0(n3938), .A1(n3277), .B0(n4041), .B1(n3875), .Y(n1966)
         );
  AOI222XLTS U3200 ( .A0(n4206), .A1(n3316), .B0(n3300), .B1(n24), .C0(n3981), 
        .C1(n3293), .Y(n1967) );
  AOI22X1TS U3201 ( .A0(n3935), .A1(n3277), .B0(n4038), .B1(n3875), .Y(n1964)
         );
  AOI222XLTS U3202 ( .A0(n4202), .A1(n3316), .B0(n3306), .B1(n19), .C0(n3978), 
        .C1(n3292), .Y(n1965) );
  AOI22X1TS U3203 ( .A0(n4433), .A1(n3274), .B0(n4167), .B1(n3875), .Y(n1358)
         );
  AOI222XLTS U3204 ( .A0(n4523), .A1(n3316), .B0(n511), .B1(n3296), .C0(n4335), 
        .C1(n3287), .Y(n1359) );
  AOI22X1TS U3205 ( .A0(n4429), .A1(n3275), .B0(n4164), .B1(n3875), .Y(n1356)
         );
  AOI222XLTS U3206 ( .A0(dataIn_SOUTH[30]), .A1(n3316), .B0(n507), .B1(n3295), 
        .C0(n4332), .C1(n3287), .Y(n1357) );
  AOI22X1TS U3207 ( .A0(n4426), .A1(n3274), .B0(n4161), .B1(n3874), .Y(n1354)
         );
  AOI222XLTS U3208 ( .A0(n4517), .A1(n3315), .B0(n513), .B1(n3296), .C0(n4329), 
        .C1(n3287), .Y(n1355) );
  AOI22X1TS U3209 ( .A0(n4421), .A1(n3275), .B0(n4158), .B1(n3874), .Y(n1352)
         );
  AOI222XLTS U3210 ( .A0(dataIn_SOUTH[28]), .A1(n3315), .B0(n477), .B1(n3295), 
        .C0(n4326), .C1(n3287), .Y(n1353) );
  AOI22X1TS U3211 ( .A0(n4415), .A1(n3273), .B0(n4152), .B1(n3874), .Y(n1348)
         );
  AOI222XLTS U3212 ( .A0(n4509), .A1(n3315), .B0(n515), .B1(n3297), .C0(n4320), 
        .C1(n3286), .Y(n1349) );
  AOI22X1TS U3213 ( .A0(n4412), .A1(n3268), .B0(n4149), .B1(n3879), .Y(n1346)
         );
  AOI222XLTS U3214 ( .A0(n4507), .A1(n3323), .B0(n517), .B1(n3297), .C0(n4317), 
        .C1(n3286), .Y(n1347) );
  AOI22X1TS U3215 ( .A0(n4409), .A1(n3268), .B0(n4146), .B1(n3880), .Y(n1344)
         );
  AOI222XLTS U3216 ( .A0(dataIn_SOUTH[24]), .A1(n3324), .B0(n519), .B1(n3296), 
        .C0(n4314), .C1(n3286), .Y(n1345) );
  AOI22X1TS U3217 ( .A0(n4406), .A1(n3268), .B0(n4143), .B1(n3876), .Y(n1342)
         );
  AOI222XLTS U3218 ( .A0(n4500), .A1(n3323), .B0(n481), .B1(n3298), .C0(n4311), 
        .C1(n3285), .Y(n1343) );
  AOI22X1TS U3219 ( .A0(n4400), .A1(n3267), .B0(n4137), .B1(n3873), .Y(n1338)
         );
  AOI222XLTS U3220 ( .A0(n4496), .A1(n3320), .B0(n523), .B1(n3296), .C0(n4305), 
        .C1(n3285), .Y(n1339) );
  AOI22X1TS U3221 ( .A0(n4391), .A1(n3266), .B0(n4128), .B1(n3873), .Y(n1332)
         );
  AOI222XLTS U3222 ( .A0(n4487), .A1(n3314), .B0(n527), .B1(n3297), .C0(n4296), 
        .C1(n3284), .Y(n1333) );
  AOI22X1TS U3223 ( .A0(n4388), .A1(n3266), .B0(n4125), .B1(n3872), .Y(n1330)
         );
  AOI222XLTS U3224 ( .A0(n4484), .A1(n3314), .B0(n529), .B1(n3299), .C0(n4293), 
        .C1(n3284), .Y(n1331) );
  AOI22X1TS U3225 ( .A0(n4385), .A1(n3266), .B0(n4122), .B1(n3872), .Y(n1328)
         );
  AOI222XLTS U3226 ( .A0(n4481), .A1(n3314), .B0(n509), .B1(n3295), .C0(n4290), 
        .C1(n3284), .Y(n1329) );
  AOI22X1TS U3227 ( .A0(n4382), .A1(n3266), .B0(n4119), .B1(n3872), .Y(n1326)
         );
  AOI222XLTS U3228 ( .A0(n4478), .A1(n3314), .B0(n531), .B1(n3298), .C0(n4287), 
        .C1(n3283), .Y(n1327) );
  AOI22X1TS U3229 ( .A0(n4379), .A1(n3265), .B0(n4116), .B1(n3872), .Y(n1324)
         );
  AOI222XLTS U3230 ( .A0(n4474), .A1(n3313), .B0(n533), .B1(n3297), .C0(n4284), 
        .C1(n3283), .Y(n1325) );
  AOI22X1TS U3231 ( .A0(n4376), .A1(n3265), .B0(n4113), .B1(n3877), .Y(n1322)
         );
  AOI222XLTS U3232 ( .A0(dataIn_SOUTH[13]), .A1(n3313), .B0(n535), .B1(n3303), 
        .C0(n4281), .C1(n3283), .Y(n1323) );
  AOI22X1TS U3233 ( .A0(n4373), .A1(n3265), .B0(n4110), .B1(n3876), .Y(n1320)
         );
  AOI222XLTS U3234 ( .A0(n4469), .A1(n3313), .B0(n485), .B1(n3299), .C0(n4278), 
        .C1(n3282), .Y(n1321) );
  AOI22X1TS U3235 ( .A0(n4370), .A1(n3265), .B0(n4107), .B1(n3876), .Y(n1318)
         );
  AOI222XLTS U3236 ( .A0(n4466), .A1(n3313), .B0(n487), .B1(n3304), .C0(n4275), 
        .C1(n3282), .Y(n1319) );
  AOI22X1TS U3237 ( .A0(n4364), .A1(n3267), .B0(n4101), .B1(n3871), .Y(n1314)
         );
  AOI222XLTS U3238 ( .A0(n4461), .A1(n3322), .B0(n491), .B1(n3303), .C0(n4269), 
        .C1(n3282), .Y(n1315) );
  AOI22X1TS U3239 ( .A0(n4358), .A1(n3264), .B0(n4095), .B1(n3871), .Y(n1310)
         );
  AOI222XLTS U3240 ( .A0(dataIn_SOUTH[7]), .A1(n3312), .B0(n495), .B1(n3308), 
        .C0(n4263), .C1(n3290), .Y(n1311) );
  AOI22X1TS U3241 ( .A0(n4355), .A1(n3264), .B0(n4092), .B1(n3871), .Y(n1308)
         );
  AOI222XLTS U3242 ( .A0(n4454), .A1(n3312), .B0(n497), .B1(n3305), .C0(n4260), 
        .C1(n3283), .Y(n1309) );
  AOI22X1TS U3243 ( .A0(n4349), .A1(n3263), .B0(n4086), .B1(n3870), .Y(n1304)
         );
  AOI222XLTS U3244 ( .A0(n4447), .A1(n3311), .B0(n501), .B1(n3302), .C0(n4254), 
        .C1(n3290), .Y(n1305) );
  AOI22X1TS U3245 ( .A0(n4346), .A1(n3263), .B0(n4083), .B1(n3870), .Y(n1302)
         );
  AOI222XLTS U3246 ( .A0(dataIn_SOUTH[3]), .A1(n3311), .B0(n503), .B1(n3306), 
        .C0(n4251), .C1(n3291), .Y(n1303) );
  AOI22X1TS U3247 ( .A0(n4340), .A1(n3262), .B0(n4077), .B1(n3869), .Y(n1298)
         );
  AOI222XLTS U3248 ( .A0(n4440), .A1(n3310), .B0(n537), .B1(n3305), .C0(n4245), 
        .C1(n3288), .Y(n1299) );
  AOI22X1TS U3249 ( .A0(n4337), .A1(n3262), .B0(n4074), .B1(n3869), .Y(n1296)
         );
  AOI222XLTS U3250 ( .A0(dataIn_SOUTH[0]), .A1(n3310), .B0(n539), .B1(n3299), 
        .C0(n4242), .C1(n3289), .Y(n1297) );
  AOI22X1TS U3251 ( .A0(n4469), .A1(n3120), .B0(n4277), .B1(n3885), .Y(n1256)
         );
  AOI222XLTS U3252 ( .A0(n4374), .A1(n3230), .B0(n4111), .B1(n3216), .C0(n486), 
        .C1(n3204), .Y(n1257) );
  AOI22X1TS U3253 ( .A0(n4466), .A1(n3120), .B0(n4274), .B1(n3885), .Y(n1254)
         );
  AOI222XLTS U3254 ( .A0(n4371), .A1(n3230), .B0(n4108), .B1(n3216), .C0(n488), 
        .C1(n3203), .Y(n1255) );
  AOI22X1TS U3255 ( .A0(n4463), .A1(n3119), .B0(n4271), .B1(n3885), .Y(n1252)
         );
  AOI222XLTS U3256 ( .A0(n4368), .A1(n3229), .B0(n4105), .B1(n3217), .C0(n490), 
        .C1(n3205), .Y(n1253) );
  AOI22X1TS U3257 ( .A0(n4458), .A1(n3119), .B0(n4265), .B1(n3884), .Y(n1248)
         );
  AOI222XLTS U3258 ( .A0(n4362), .A1(n3229), .B0(n4099), .B1(n3217), .C0(n494), 
        .C1(n3202), .Y(n1249) );
  AOI22X1TS U3259 ( .A0(n4455), .A1(n3119), .B0(n4262), .B1(n3884), .Y(n1246)
         );
  AOI222XLTS U3260 ( .A0(n4359), .A1(n3229), .B0(n4096), .B1(n3217), .C0(n496), 
        .C1(n3202), .Y(n1247) );
  AOI22X1TS U3261 ( .A0(n4454), .A1(n3119), .B0(n4259), .B1(n3884), .Y(n1244)
         );
  AOI222XLTS U3262 ( .A0(n4356), .A1(n3229), .B0(n4093), .B1(n3218), .C0(n498), 
        .C1(n3208), .Y(n1245) );
  AOI22X1TS U3263 ( .A0(n4447), .A1(n3118), .B0(n4253), .B1(n3883), .Y(n1240)
         );
  AOI222XLTS U3264 ( .A0(n4350), .A1(n3228), .B0(n4087), .B1(n3218), .C0(n502), 
        .C1(n3204), .Y(n1241) );
  AOI22X1TS U3265 ( .A0(n4444), .A1(n3118), .B0(n4250), .B1(n3883), .Y(n1238)
         );
  AOI222XLTS U3266 ( .A0(n4347), .A1(n3228), .B0(n4084), .B1(n3218), .C0(n504), 
        .C1(n3206), .Y(n1239) );
  AOI22X1TS U3267 ( .A0(n4213), .A1(n3123), .B0(n3990), .B1(n3889), .Y(n1994)
         );
  AOI222XLTS U3268 ( .A0(n3947), .A1(n3239), .B0(n4051), .B1(n3210), .C0(n3197), .C1(n36), .Y(n1995) );
  AOI22X1TS U3269 ( .A0(n4203), .A1(n3194), .B0(n3978), .B1(n3890), .Y(n1986)
         );
  AOI222XLTS U3270 ( .A0(n3935), .A1(n3240), .B0(n4039), .B1(n3211), .C0(n3197), .C1(n16), .Y(n1987) );
  AOI22X1TS U3271 ( .A0(n4514), .A1(n3125), .B0(n4325), .B1(n3892), .Y(n1288)
         );
  AOI222XLTS U3272 ( .A0(n4422), .A1(n3238), .B0(n4159), .B1(n3212), .C0(n478), 
        .C1(n3198), .Y(n1289) );
  AOI22X1TS U3273 ( .A0(n4512), .A1(n3127), .B0(n4322), .B1(n1761), .Y(n1286)
         );
  AOI222XLTS U3274 ( .A0(n4419), .A1(n3235), .B0(n4156), .B1(n3212), .C0(n480), 
        .C1(n3199), .Y(n1287) );
  AOI22X1TS U3275 ( .A0(n4500), .A1(n3128), .B0(n4310), .B1(n3888), .Y(n1278)
         );
  AOI222XLTS U3276 ( .A0(n4407), .A1(n3233), .B0(n4144), .B1(n3213), .C0(n482), 
        .C1(n3199), .Y(n1279) );
  AOI22X1TS U3277 ( .A0(n4492), .A1(n3126), .B0(n4301), .B1(n3887), .Y(n1272)
         );
  AOI222XLTS U3278 ( .A0(n4398), .A1(n3232), .B0(n4135), .B1(n3214), .C0(n484), 
        .C1(n3200), .Y(n1273) );
  AOI22X1TS U3279 ( .A0(n4461), .A1(n3125), .B0(n4268), .B1(n3884), .Y(n1250)
         );
  AOI222XLTS U3280 ( .A0(n4365), .A1(n3232), .B0(n4102), .B1(n3217), .C0(n492), 
        .C1(n3207), .Y(n1251) );
  AOI22X1TS U3281 ( .A0(n4452), .A1(n3118), .B0(n4256), .B1(n3883), .Y(n1242)
         );
  AOI222XLTS U3282 ( .A0(n4353), .A1(n3228), .B0(n4090), .B1(n3218), .C0(n500), 
        .C1(n3203), .Y(n1243) );
  AOI22X1TS U3283 ( .A0(n4443), .A1(n3118), .B0(n4247), .B1(n3883), .Y(n1236)
         );
  AOI222XLTS U3284 ( .A0(n4344), .A1(n3228), .B0(n4081), .B1(n3219), .C0(n506), 
        .C1(n3208), .Y(n1237) );
  AOI22X1TS U3285 ( .A0(n4440), .A1(n3117), .B0(n4244), .B1(n3882), .Y(n1234)
         );
  AOI222XLTS U3286 ( .A0(n4341), .A1(n3227), .B0(n4078), .B1(n3219), .C0(n538), 
        .C1(n3205), .Y(n1235) );
  AOI22X1TS U3287 ( .A0(n4436), .A1(n3117), .B0(n4241), .B1(n3882), .Y(n1232)
         );
  AOI222XLTS U3288 ( .A0(n4338), .A1(n3227), .B0(n4075), .B1(n3219), .C0(n540), 
        .C1(n3206), .Y(n1233) );
  AOI22X1TS U3289 ( .A0(n3117), .A1(n4538), .B0(n3882), .B1(n4035), .Y(n1230)
         );
  AOI222XLTS U3290 ( .A0(n3227), .A1(n4184), .B0(n3219), .B1(n4072), .C0(n3196), .C1(n43), .Y(n1231) );
  AOI22X1TS U3291 ( .A0(n3116), .A1(n4533), .B0(n3881), .B1(n4029), .Y(n1226)
         );
  AOI222XLTS U3292 ( .A0(n3226), .A1(n4178), .B0(n1219), .B1(n4066), .C0(n3195), .C1(n32), .Y(n1227) );
  AOI22X1TS U3293 ( .A0(n3116), .A1(n4536), .B0(n3882), .B1(n4032), .Y(n1228)
         );
  AOI222XLTS U3294 ( .A0(n3226), .A1(n4181), .B0(n3224), .B1(n4069), .C0(n3196), .C1(n37), .Y(n1229) );
  AOI22X1TS U3295 ( .A0(n3116), .A1(n4529), .B0(n3881), .B1(n4026), .Y(n1224)
         );
  AOI222XLTS U3296 ( .A0(n3226), .A1(n4175), .B0(n3222), .B1(n4063), .C0(n3195), .C1(n27), .Y(n1225) );
  AOI22X1TS U3297 ( .A0(n3116), .A1(n4528), .B0(n3881), .B1(n4023), .Y(n1222)
         );
  AOI222XLTS U3298 ( .A0(n3226), .A1(n4172), .B0(n3221), .B1(n4060), .C0(n3195), .C1(n22), .Y(n1223) );
  AOI22X1TS U3299 ( .A0(n3117), .A1(n4525), .B0(n3881), .B1(n4020), .Y(n1216)
         );
  AOI222XLTS U3300 ( .A0(n3227), .A1(n4169), .B0(n3225), .B1(n4057), .C0(n3196), .C1(n17), .Y(n1217) );
  AOI22X1TS U3301 ( .A0(n4433), .A1(n3434), .B0(n4523), .B1(n3423), .Y(n1486)
         );
  AOI222XLTS U3302 ( .A0(n512), .A1(n3778), .B0(n4168), .B1(n3865), .C0(n6260), 
        .C1(n3847), .Y(n1487) );
  AOI22X1TS U3303 ( .A0(n4429), .A1(n3434), .B0(n4518), .B1(n3422), .Y(n1484)
         );
  AOI222XLTS U3304 ( .A0(n508), .A1(n3782), .B0(n4165), .B1(n3865), .C0(n6261), 
        .C1(n3847), .Y(n1485) );
  AOI22X1TS U3305 ( .A0(n4426), .A1(n3433), .B0(n4517), .B1(n3421), .Y(n1482)
         );
  AOI222XLTS U3306 ( .A0(n514), .A1(n3782), .B0(n4162), .B1(n3863), .C0(n6262), 
        .C1(n3847), .Y(n1483) );
  AOI22X1TS U3307 ( .A0(n4421), .A1(n3433), .B0(n4514), .B1(n3421), .Y(n1480)
         );
  AOI222XLTS U3308 ( .A0(n478), .A1(n3782), .B0(n4159), .B1(n3864), .C0(n6263), 
        .C1(n3847), .Y(n1481) );
  AOI22X1TS U3309 ( .A0(n4418), .A1(n3433), .B0(n4512), .B1(n3423), .Y(n1478)
         );
  AOI222XLTS U3310 ( .A0(n480), .A1(n3781), .B0(n4156), .B1(n3863), .C0(n6264), 
        .C1(n3846), .Y(n1479) );
  AOI22X1TS U3311 ( .A0(n4415), .A1(n3433), .B0(n4509), .B1(n3422), .Y(n1476)
         );
  AOI222XLTS U3312 ( .A0(n516), .A1(n3775), .B0(n4153), .B1(n3864), .C0(n6265), 
        .C1(n3846), .Y(n1477) );
  AOI22X1TS U3313 ( .A0(n4409), .A1(n3432), .B0(n4502), .B1(n3417), .Y(n1472)
         );
  AOI222XLTS U3314 ( .A0(n520), .A1(n3779), .B0(n4147), .B1(n3855), .C0(n6266), 
        .C1(n3846), .Y(n1473) );
  AOI22X1TS U3315 ( .A0(n4403), .A1(n3432), .B0(n4498), .B1(n3417), .Y(n1468)
         );
  AOI222XLTS U3316 ( .A0(n522), .A1(n3781), .B0(n4141), .B1(n3855), .C0(n6267), 
        .C1(n3845), .Y(n1469) );
  AOI22X1TS U3317 ( .A0(n4400), .A1(n3431), .B0(n4496), .B1(n3416), .Y(n1466)
         );
  AOI222XLTS U3318 ( .A0(n524), .A1(n3773), .B0(n4138), .B1(n3856), .C0(n6268), 
        .C1(n3845), .Y(n1467) );
  AOI22X1TS U3319 ( .A0(n4394), .A1(n3431), .B0(n4490), .B1(n3416), .Y(n1462)
         );
  AOI222XLTS U3320 ( .A0(n526), .A1(n3773), .B0(n4132), .B1(n3856), .C0(n6269), 
        .C1(n3844), .Y(n1463) );
  AOI22X1TS U3321 ( .A0(n4388), .A1(n3440), .B0(n4484), .B1(n3415), .Y(n1458)
         );
  AOI222XLTS U3322 ( .A0(n530), .A1(n3773), .B0(n4126), .B1(n3857), .C0(n6270), 
        .C1(n3844), .Y(n1459) );
  AOI22X1TS U3323 ( .A0(n4385), .A1(n3440), .B0(n4481), .B1(n3415), .Y(n1456)
         );
  AOI222XLTS U3324 ( .A0(n510), .A1(n3774), .B0(n4123), .B1(n3857), .C0(n6271), 
        .C1(n3844), .Y(n1457) );
  AOI22X1TS U3325 ( .A0(n4379), .A1(n3430), .B0(n4474), .B1(n3414), .Y(n1452)
         );
  AOI222XLTS U3326 ( .A0(n534), .A1(n3774), .B0(n4117), .B1(n3857), .C0(n6272), 
        .C1(n3852), .Y(n1453) );
  AOI22X1TS U3327 ( .A0(n4373), .A1(n3430), .B0(n4469), .B1(n3414), .Y(n1448)
         );
  AOI222XLTS U3328 ( .A0(n486), .A1(n3775), .B0(n4111), .B1(n3858), .C0(n6273), 
        .C1(n3851), .Y(n1449) );
  AOI22X1TS U3329 ( .A0(n4370), .A1(n3430), .B0(n4466), .B1(n3414), .Y(n1446)
         );
  AOI222XLTS U3330 ( .A0(n488), .A1(n3775), .B0(n4108), .B1(n3858), .C0(n6274), 
        .C1(n3851), .Y(n1447) );
  AOI22X1TS U3331 ( .A0(n4367), .A1(n3429), .B0(n4463), .B1(n3413), .Y(n1444)
         );
  AOI222XLTS U3332 ( .A0(n490), .A1(n3778), .B0(n4105), .B1(n3858), .C0(n6275), 
        .C1(n3852), .Y(n1445) );
  AOI22X1TS U3333 ( .A0(n4364), .A1(n3431), .B0(n4461), .B1(n3416), .Y(n1442)
         );
  AOI222XLTS U3334 ( .A0(n492), .A1(n3776), .B0(n4102), .B1(n3859), .C0(n6276), 
        .C1(n3850), .Y(n1443) );
  AOI22X1TS U3335 ( .A0(n4361), .A1(n3429), .B0(n4458), .B1(n3413), .Y(n1440)
         );
  AOI222XLTS U3336 ( .A0(n494), .A1(n3776), .B0(n4099), .B1(n3859), .C0(n6277), 
        .C1(n3843), .Y(n1441) );
  AOI22X1TS U3337 ( .A0(n4355), .A1(n3429), .B0(n4454), .B1(n3413), .Y(n1436)
         );
  AOI222XLTS U3338 ( .A0(n498), .A1(n3777), .B0(n4093), .B1(n3859), .C0(n6278), 
        .C1(n3843), .Y(n1437) );
  AOI22X1TS U3339 ( .A0(n4346), .A1(n3428), .B0(n4444), .B1(n3412), .Y(n1430)
         );
  AOI222XLTS U3340 ( .A0(n504), .A1(n3778), .B0(n4084), .B1(n3860), .C0(n6279), 
        .C1(n3842), .Y(n1431) );
  AOI22X1TS U3341 ( .A0(n4340), .A1(n3443), .B0(n4440), .B1(n3411), .Y(n1426)
         );
  AOI22X1TS U3342 ( .A0(n4337), .A1(n3441), .B0(n4436), .B1(n3411), .Y(n1424)
         );
  AOI222XLTS U3343 ( .A0(n540), .A1(n3778), .B0(n4075), .B1(n3861), .C0(n6281), 
        .C1(n3841), .Y(n1425) );
  AOI22X1TS U3344 ( .A0(n4412), .A1(n3432), .B0(n4507), .B1(n3417), .Y(n1474)
         );
  AOI222XLTS U3345 ( .A0(n518), .A1(n3780), .B0(n4150), .B1(n3855), .C0(n6294), 
        .C1(n3846), .Y(n1475) );
  AOI22X1TS U3346 ( .A0(n4406), .A1(n3432), .B0(n4500), .B1(n3417), .Y(n1470)
         );
  AOI222XLTS U3347 ( .A0(n482), .A1(n3782), .B0(n4144), .B1(n3855), .C0(n6295), 
        .C1(n3845), .Y(n1471) );
  AOI22X1TS U3348 ( .A0(n4397), .A1(n3431), .B0(n4492), .B1(n3416), .Y(n1464)
         );
  AOI222XLTS U3349 ( .A0(n484), .A1(n3773), .B0(n4135), .B1(n3856), .C0(n6296), 
        .C1(n3845), .Y(n1465) );
  AOI22X1TS U3350 ( .A0(n4391), .A1(n3441), .B0(n4487), .B1(n3415), .Y(n1460)
         );
  AOI222XLTS U3351 ( .A0(n528), .A1(n3774), .B0(n4129), .B1(n3856), .C0(n6297), 
        .C1(n3844), .Y(n1461) );
  AOI22X1TS U3352 ( .A0(n4382), .A1(n3441), .B0(n4478), .B1(n3415), .Y(n1454)
         );
  AOI222XLTS U3353 ( .A0(n532), .A1(n3775), .B0(n4120), .B1(n3857), .C0(n6298), 
        .C1(n3849), .Y(n1455) );
  AOI22X1TS U3354 ( .A0(n4376), .A1(n3430), .B0(n4470), .B1(n3414), .Y(n1450)
         );
  AOI222XLTS U3355 ( .A0(n536), .A1(n3774), .B0(n4114), .B1(n3858), .C0(n6299), 
        .C1(n734), .Y(n1451) );
  AOI22X1TS U3356 ( .A0(n4352), .A1(n3428), .B0(n4452), .B1(n3412), .Y(n1434)
         );
  AOI222XLTS U3357 ( .A0(n500), .A1(n3776), .B0(n4090), .B1(n3860), .C0(n6300), 
        .C1(n3843), .Y(n1435) );
  AOI22X1TS U3358 ( .A0(n4349), .A1(n3428), .B0(n4447), .B1(n3412), .Y(n1432)
         );
  AOI222XLTS U3359 ( .A0(n502), .A1(n3777), .B0(n4087), .B1(n3860), .C0(n6301), 
        .C1(n3842), .Y(n1433) );
  AOI22X1TS U3360 ( .A0(n4343), .A1(n3428), .B0(n4443), .B1(n3412), .Y(n1428)
         );
  AOI222XLTS U3361 ( .A0(n506), .A1(n3777), .B0(n4081), .B1(n3860), .C0(n6302), 
        .C1(n3842), .Y(n1429) );
  AOI22X1TS U3362 ( .A0(n4358), .A1(n3429), .B0(n4455), .B1(n3413), .Y(n1438)
         );
  AOI222XLTS U3363 ( .A0(n496), .A1(n3776), .B0(n4096), .B1(n3859), .C0(n6312), 
        .C1(n3843), .Y(n1439) );
  AOI22X1TS U3364 ( .A0(n3478), .A1(n42), .B0(n3950), .B1(n3468), .Y(n1904) );
  AOI222XLTS U3365 ( .A0(n2997), .A1(n3894), .B0(n4216), .B1(n3494), .C0(n4054), .C1(n3929), .Y(n1905) );
  AOI22X1TS U3366 ( .A0(n3480), .A1(n33), .B0(n3944), .B1(n3468), .Y(n1900) );
  AOI222XLTS U3367 ( .A0(n3001), .A1(n3903), .B0(n4211), .B1(n3502), .C0(n4048), .C1(n3929), .Y(n1901) );
  AOI22X1TS U3368 ( .A0(n3480), .A1(n27), .B0(n3941), .B1(n3468), .Y(n1898) );
  AOI222XLTS U3369 ( .A0(n3003), .A1(n3903), .B0(n4209), .B1(n3502), .C0(n4045), .C1(n3929), .Y(n1899) );
  AOI22X1TS U3370 ( .A0(n3479), .A1(n23), .B0(n3938), .B1(n3467), .Y(n1896) );
  AOI222XLTS U3371 ( .A0(n3005), .A1(n3903), .B0(n4206), .B1(n3507), .C0(n4042), .C1(n3928), .Y(n1897) );
  AOI22X1TS U3372 ( .A0(n3480), .A1(n18), .B0(n3935), .B1(n3467), .Y(n1894) );
  AOI222XLTS U3373 ( .A0(n3007), .A1(n3904), .B0(n4202), .B1(n3507), .C0(n4039), .C1(n3928), .Y(n1895) );
  AOI22X1TS U3374 ( .A0(n508), .A1(n3481), .B0(n4429), .B1(n3467), .Y(n1548)
         );
  AOI222XLTS U3375 ( .A0(n2935), .A1(n3902), .B0(n4519), .B1(n3504), .C0(n4165), .C1(n3928), .Y(n1549) );
  AOI22X1TS U3376 ( .A0(n478), .A1(n3481), .B0(n4421), .B1(n3470), .Y(n1544)
         );
  AOI222XLTS U3377 ( .A0(n2939), .A1(n3902), .B0(n4515), .B1(n3501), .C0(n4159), .C1(n3927), .Y(n1545) );
  AOI22X1TS U3378 ( .A0(n480), .A1(n3482), .B0(n4418), .B1(n3477), .Y(n1542)
         );
  AOI222XLTS U3379 ( .A0(n2941), .A1(n3901), .B0(n4511), .B1(n3501), .C0(n4156), .C1(n3927), .Y(n1543) );
  AOI22X1TS U3380 ( .A0(n516), .A1(n3485), .B0(n4415), .B1(n1156), .Y(n1540)
         );
  AOI222XLTS U3381 ( .A0(n2943), .A1(n3901), .B0(n4510), .B1(n3501), .C0(n4153), .C1(n3927), .Y(n1541) );
  AOI22X1TS U3382 ( .A0(n518), .A1(n3481), .B0(n4412), .B1(n3473), .Y(n1538)
         );
  AOI222XLTS U3383 ( .A0(n2945), .A1(n3901), .B0(n4506), .B1(n3500), .C0(n4150), .C1(n3930), .Y(n1539) );
  AOI22X1TS U3384 ( .A0(n520), .A1(n3482), .B0(n4409), .B1(n3475), .Y(n1536)
         );
  AOI222XLTS U3385 ( .A0(n2947), .A1(n3901), .B0(n4503), .B1(n3500), .C0(n4147), .C1(n3930), .Y(n1537) );
  AOI22X1TS U3386 ( .A0(n482), .A1(n3482), .B0(n4406), .B1(n3472), .Y(n1534)
         );
  AOI222XLTS U3387 ( .A0(n2949), .A1(n3900), .B0(n4501), .B1(n3500), .C0(n4144), .C1(n3931), .Y(n1535) );
  AOI22X1TS U3388 ( .A0(n528), .A1(n3487), .B0(n4391), .B1(n3466), .Y(n1524)
         );
  AOI222XLTS U3389 ( .A0(n2959), .A1(n3904), .B0(n4485), .B1(n3498), .C0(n4129), .C1(n3926), .Y(n1525) );
  AOI22X1TS U3390 ( .A0(n536), .A1(n3486), .B0(n4376), .B1(n3465), .Y(n1514)
         );
  AOI222XLTS U3391 ( .A0(n2969), .A1(n3899), .B0(n4471), .B1(n3497), .C0(n4114), .C1(n3925), .Y(n1515) );
  AOI22X1TS U3392 ( .A0(n492), .A1(n3483), .B0(n4364), .B1(n3474), .Y(n1506)
         );
  AOI222XLTS U3393 ( .A0(n2977), .A1(n3898), .B0(n4462), .B1(n3496), .C0(n4102), .C1(n3924), .Y(n1507) );
  AOI22X1TS U3394 ( .A0(n496), .A1(n3483), .B0(n4358), .B1(n3464), .Y(n1502)
         );
  AOI222XLTS U3395 ( .A0(n2981), .A1(n3897), .B0(n4456), .B1(n3496), .C0(n4096), .C1(n3924), .Y(n1503) );
  AOI22X1TS U3396 ( .A0(n500), .A1(n3483), .B0(n4352), .B1(n3463), .Y(n1498)
         );
  AOI222XLTS U3397 ( .A0(n2985), .A1(n3897), .B0(n4451), .B1(n3495), .C0(n4090), .C1(n3933), .Y(n1499) );
  AOI22X1TS U3398 ( .A0(n502), .A1(n3484), .B0(n4349), .B1(n3463), .Y(n1496)
         );
  AOI222XLTS U3399 ( .A0(n2987), .A1(n3896), .B0(n4449), .B1(n3495), .C0(n4087), .C1(n722), .Y(n1497) );
  AOI22X1TS U3400 ( .A0(n506), .A1(n3484), .B0(n4343), .B1(n3463), .Y(n1492)
         );
  AOI222XLTS U3401 ( .A0(n2991), .A1(n3896), .B0(n4442), .B1(n3495), .C0(n4081), .C1(n3934), .Y(n1493) );
  AOI22X1TS U3402 ( .A0(n512), .A1(n3489), .B0(n4433), .B1(n3467), .Y(n1550)
         );
  AOI222XLTS U3403 ( .A0(n2933), .A1(n3902), .B0(n4521), .B1(n3510), .C0(n4168), .C1(n3928), .Y(n1551) );
  AOI22X1TS U3404 ( .A0(n514), .A1(n3481), .B0(n4426), .B1(n1156), .Y(n1546)
         );
  AOI222XLTS U3405 ( .A0(n2937), .A1(n3902), .B0(n4516), .B1(n3501), .C0(n4162), .C1(n3927), .Y(n1547) );
  AOI22X1TS U3406 ( .A0(n522), .A1(n3482), .B0(n4403), .B1(n3472), .Y(n1532)
         );
  AOI222XLTS U3407 ( .A0(n2951), .A1(n3900), .B0(n4497), .B1(n3500), .C0(n4141), .C1(n3932), .Y(n1533) );
  AOI22X1TS U3408 ( .A0(n524), .A1(n3486), .B0(n4400), .B1(n3473), .Y(n1530)
         );
  AOI222XLTS U3409 ( .A0(n2953), .A1(n3900), .B0(n4494), .B1(n3499), .C0(n4138), .C1(n3926), .Y(n1531) );
  AOI22X1TS U3410 ( .A0(n484), .A1(n3486), .B0(n4397), .B1(n3475), .Y(n1528)
         );
  AOI222XLTS U3411 ( .A0(n2955), .A1(n3900), .B0(n4493), .B1(n3499), .C0(n4135), .C1(n3926), .Y(n1529) );
  AOI22X1TS U3412 ( .A0(n526), .A1(n3486), .B0(n4394), .B1(n3474), .Y(n1526)
         );
  AOI222XLTS U3413 ( .A0(n2957), .A1(n3908), .B0(n4488), .B1(n3499), .C0(n4132), .C1(n3926), .Y(n1527) );
  AOI22X1TS U3414 ( .A0(n510), .A1(n3488), .B0(n4385), .B1(n3466), .Y(n1520)
         );
  AOI222XLTS U3415 ( .A0(n2963), .A1(n3907), .B0(n4482), .B1(n3498), .C0(n4123), .C1(n3933), .Y(n1521) );
  AOI22X1TS U3416 ( .A0(n486), .A1(n3485), .B0(n4373), .B1(n3465), .Y(n1512)
         );
  AOI222XLTS U3417 ( .A0(n2971), .A1(n3898), .B0(n4467), .B1(n3497), .C0(n4111), .C1(n3925), .Y(n1513) );
  AOI22X1TS U3418 ( .A0(n488), .A1(n3485), .B0(n4370), .B1(n3465), .Y(n1510)
         );
  AOI222XLTS U3419 ( .A0(n2973), .A1(n3898), .B0(n4465), .B1(n3497), .C0(n4108), .C1(n3925), .Y(n1511) );
  AOI22X1TS U3420 ( .A0(n490), .A1(n3484), .B0(n4367), .B1(n3464), .Y(n1508)
         );
  AOI222XLTS U3421 ( .A0(n2975), .A1(n3898), .B0(n4464), .B1(n3496), .C0(n4105), .C1(n3925), .Y(n1509) );
  AOI22X1TS U3422 ( .A0(n494), .A1(n3483), .B0(n4361), .B1(n3464), .Y(n1504)
         );
  AOI222XLTS U3423 ( .A0(n2979), .A1(n3897), .B0(n4457), .B1(n3496), .C0(n4099), .C1(n3924), .Y(n1505) );
  AOI22X1TS U3424 ( .A0(n498), .A1(n3484), .B0(n4355), .B1(n3464), .Y(n1500)
         );
  AOI222XLTS U3425 ( .A0(n2983), .A1(n3897), .B0(n4453), .B1(n3499), .C0(n4093), .C1(n3924), .Y(n1501) );
  AOI22X1TS U3426 ( .A0(n538), .A1(n3491), .B0(n4340), .B1(n3462), .Y(n1490)
         );
  AOI222XLTS U3427 ( .A0(n2993), .A1(n3896), .B0(n4439), .B1(n3494), .C0(n4078), .C1(n3923), .Y(n1491) );
  AOI22X1TS U3428 ( .A0(n540), .A1(n3489), .B0(n4337), .B1(n3462), .Y(n1488)
         );
  AOI222XLTS U3429 ( .A0(n2995), .A1(n3895), .B0(n4438), .B1(n3494), .C0(n4075), .C1(n3923), .Y(n1489) );
  AOI22X1TS U3430 ( .A0(n530), .A1(n3489), .B0(n4388), .B1(n3466), .Y(n1522)
         );
  AOI222XLTS U3431 ( .A0(n2961), .A1(n3907), .B0(n4483), .B1(n3498), .C0(n4126), .C1(n3932), .Y(n1523) );
  AOI22X1TS U3432 ( .A0(n532), .A1(n3490), .B0(n4382), .B1(n3466), .Y(n1518)
         );
  AOI222XLTS U3433 ( .A0(n2965), .A1(n3899), .B0(n4476), .B1(n3498), .C0(n4120), .C1(n722), .Y(n1519) );
  AOI22X1TS U3434 ( .A0(n534), .A1(n3487), .B0(n4379), .B1(n3465), .Y(n1516)
         );
  AOI222XLTS U3435 ( .A0(n2967), .A1(n3899), .B0(n4475), .B1(n3497), .C0(n4117), .C1(n3931), .Y(n1517) );
  AOI22X1TS U3436 ( .A0(n504), .A1(n3488), .B0(n4346), .B1(n3463), .Y(n1494)
         );
  AOI222XLTS U3437 ( .A0(n2989), .A1(n3896), .B0(n4445), .B1(n3495), .C0(n4084), .C1(n3934), .Y(n1495) );
  AOI22X1TS U3438 ( .A0(n3480), .A1(n37), .B0(n3947), .B1(n3468), .Y(n1902) );
  AOI222XLTS U3439 ( .A0(n2999), .A1(n3905), .B0(n4212), .B1(n3502), .C0(n4051), .C1(n3929), .Y(n1903) );
  OAI211X1TS U3440 ( .A0(n3606), .A1(n774), .B0(n1880), .C0(n1881), .Y(n2530)
         );
  AOI22X1TS U3441 ( .A0(n3989), .A1(n3542), .B0(n4050), .B1(n3916), .Y(n1880)
         );
  AOI222XLTS U3442 ( .A0(n4213), .A1(n3584), .B0(n3570), .B1(n39), .C0(n3948), 
        .C1(n3561), .Y(n1881) );
  AOI22X1TS U3443 ( .A0(n4440), .A1(n3642), .B0(n4077), .B1(n3800), .Y(n1619)
         );
  AOI222XLTS U3444 ( .A0(n4340), .A1(n3786), .B0(n537), .B1(n3633), .C0(n4245), 
        .C1(n3616), .Y(n1620) );
  AOI22X1TS U3445 ( .A0(n4436), .A1(n3642), .B0(n4074), .B1(n3807), .Y(n1617)
         );
  AOI222XLTS U3446 ( .A0(n4337), .A1(n3786), .B0(n539), .B1(n3634), .C0(n4242), 
        .C1(n3617), .Y(n1618) );
  AOI22X1TS U3447 ( .A0(n3947), .A1(n3269), .B0(n4050), .B1(n1759), .Y(n1972)
         );
  AOI22X1TS U3448 ( .A0(n3363), .A1(n28), .B0(n3983), .B1(n3357), .Y(n1945) );
  AOI222XLTS U3449 ( .A0(n65), .A1(n3819), .B0(destinationAddressIn_SOUTH[2]), 
        .B1(n3383), .C0(n4045), .C1(n3834), .Y(n1946) );
  AOI22X1TS U3450 ( .A0(n507), .A1(n3364), .B0(n4331), .B1(n3353), .Y(n1420)
         );
  AOI222XLTS U3451 ( .A0(n66), .A1(n3818), .B0(dataIn_SOUTH[30]), .B1(n3382), 
        .C0(n4165), .C1(n3834), .Y(n1421) );
  AOI22X1TS U3452 ( .A0(n513), .A1(n3364), .B0(n4328), .B1(n3352), .Y(n1418)
         );
  AOI222XLTS U3453 ( .A0(n67), .A1(n3818), .B0(dataIn_SOUTH[29]), .B1(n3381), 
        .C0(n4162), .C1(n3840), .Y(n1419) );
  AOI22X1TS U3454 ( .A0(n477), .A1(n3364), .B0(n4325), .B1(n3352), .Y(n1416)
         );
  AOI222XLTS U3455 ( .A0(n68), .A1(n3818), .B0(dataIn_SOUTH[28]), .B1(n3381), 
        .C0(n4159), .C1(n3836), .Y(n1417) );
  AOI22X1TS U3456 ( .A0(n515), .A1(n3367), .B0(n4319), .B1(n3352), .Y(n1412)
         );
  AOI222XLTS U3457 ( .A0(n69), .A1(n3817), .B0(dataIn_SOUTH[26]), .B1(n3381), 
        .C0(n4153), .C1(n736), .Y(n1413) );
  AOI22X1TS U3458 ( .A0(n517), .A1(n3364), .B0(n4316), .B1(n3351), .Y(n1410)
         );
  AOI222XLTS U3459 ( .A0(n70), .A1(n3817), .B0(dataIn_SOUTH[25]), .B1(n3380), 
        .C0(n4150), .C1(n3837), .Y(n1411) );
  AOI22X1TS U3460 ( .A0(n481), .A1(n3365), .B0(n4310), .B1(n3351), .Y(n1406)
         );
  AOI222XLTS U3461 ( .A0(n71), .A1(n3816), .B0(dataIn_SOUTH[23]), .B1(n3380), 
        .C0(n4144), .C1(n3838), .Y(n1407) );
  AOI22X1TS U3462 ( .A0(n523), .A1(n3366), .B0(n4304), .B1(n3350), .Y(n1402)
         );
  AOI222XLTS U3463 ( .A0(n72), .A1(n3816), .B0(dataIn_SOUTH[21]), .B1(n3379), 
        .C0(n4138), .C1(n3833), .Y(n1403) );
  AOI22X1TS U3464 ( .A0(n483), .A1(n3366), .B0(n4301), .B1(n3350), .Y(n1400)
         );
  AOI222XLTS U3465 ( .A0(n73), .A1(n3816), .B0(dataIn_SOUTH[20]), .B1(n3379), 
        .C0(n4135), .C1(n3833), .Y(n1401) );
  AOI22X1TS U3466 ( .A0(n525), .A1(n3366), .B0(n4298), .B1(n3350), .Y(n1398)
         );
  AOI222XLTS U3467 ( .A0(n74), .A1(n3815), .B0(dataIn_SOUTH[19]), .B1(n3379), 
        .C0(n4132), .C1(n3833), .Y(n1399) );
  AOI22X1TS U3468 ( .A0(n527), .A1(n3370), .B0(n4295), .B1(n3349), .Y(n1396)
         );
  AOI222XLTS U3469 ( .A0(n75), .A1(n3815), .B0(dataIn_SOUTH[18]), .B1(n3378), 
        .C0(n4129), .C1(n3833), .Y(n1397) );
  AOI22X1TS U3470 ( .A0(n529), .A1(n3366), .B0(n4292), .B1(n3349), .Y(n1394)
         );
  AOI222XLTS U3471 ( .A0(n76), .A1(n3815), .B0(dataIn_SOUTH[17]), .B1(n3378), 
        .C0(n4126), .C1(n3832), .Y(n1395) );
  AOI22X1TS U3472 ( .A0(n531), .A1(n3367), .B0(n4286), .B1(n3349), .Y(n1390)
         );
  AOI222XLTS U3473 ( .A0(n77), .A1(n3814), .B0(dataIn_SOUTH[15]), .B1(n3378), 
        .C0(n4120), .C1(n3832), .Y(n1391) );
  AOI22X1TS U3474 ( .A0(n533), .A1(n3372), .B0(n4283), .B1(n3348), .Y(n1388)
         );
  AOI222XLTS U3475 ( .A0(n78), .A1(n3814), .B0(dataIn_SOUTH[14]), .B1(n3377), 
        .C0(n4117), .C1(n3832), .Y(n1389) );
  AOI22X1TS U3476 ( .A0(n535), .A1(n3372), .B0(n4280), .B1(n3348), .Y(n1386)
         );
  AOI222XLTS U3477 ( .A0(n79), .A1(n3814), .B0(dataIn_SOUTH[13]), .B1(n3377), 
        .C0(n4114), .C1(n3831), .Y(n1387) );
  AOI22X1TS U3478 ( .A0(n485), .A1(n3367), .B0(n4277), .B1(n3348), .Y(n1384)
         );
  AOI222XLTS U3479 ( .A0(n80), .A1(n3813), .B0(dataIn_SOUTH[12]), .B1(n3377), 
        .C0(n4111), .C1(n3831), .Y(n1385) );
  AOI22X1TS U3480 ( .A0(n487), .A1(n3367), .B0(n4274), .B1(n3348), .Y(n1382)
         );
  AOI222XLTS U3481 ( .A0(n81), .A1(n3813), .B0(dataIn_SOUTH[11]), .B1(n3377), 
        .C0(n4108), .C1(n3831), .Y(n1383) );
  AOI22X1TS U3482 ( .A0(n491), .A1(n3368), .B0(n4268), .B1(n3350), .Y(n1378)
         );
  AOI222XLTS U3483 ( .A0(n82), .A1(n3813), .B0(dataIn_SOUTH[9]), .B1(n3376), 
        .C0(n4102), .C1(n3830), .Y(n1379) );
  AOI22X1TS U3484 ( .A0(n493), .A1(n3368), .B0(n4265), .B1(n3347), .Y(n1376)
         );
  AOI222XLTS U3485 ( .A0(n83), .A1(n3825), .B0(dataIn_SOUTH[8]), .B1(n3376), 
        .C0(n4099), .C1(n3830), .Y(n1377) );
  AOI22X1TS U3486 ( .A0(n495), .A1(n3368), .B0(n4262), .B1(n3347), .Y(n1374)
         );
  AOI222XLTS U3487 ( .A0(n84), .A1(n3825), .B0(dataIn_SOUTH[7]), .B1(n3376), 
        .C0(n4096), .C1(n3830), .Y(n1375) );
  AOI22X1TS U3488 ( .A0(n499), .A1(n3368), .B0(n4256), .B1(n3346), .Y(n1370)
         );
  AOI222XLTS U3489 ( .A0(n85), .A1(n3824), .B0(dataIn_SOUTH[5]), .B1(n3384), 
        .C0(n4090), .C1(n3829), .Y(n1371) );
  AOI22X1TS U3490 ( .A0(n501), .A1(n3371), .B0(n4253), .B1(n3346), .Y(n1368)
         );
  AOI222XLTS U3491 ( .A0(n86), .A1(n3825), .B0(dataIn_SOUTH[4]), .B1(n3388), 
        .C0(n4087), .C1(n3829), .Y(n1369) );
  AOI22X1TS U3492 ( .A0(n503), .A1(n3370), .B0(n4250), .B1(n3346), .Y(n1366)
         );
  AOI222XLTS U3493 ( .A0(n87), .A1(n3822), .B0(dataIn_SOUTH[3]), .B1(n3390), 
        .C0(n4084), .C1(n3829), .Y(n1367) );
  AOI22X1TS U3494 ( .A0(n3361), .A1(n41), .B0(n3992), .B1(n3356), .Y(n1951) );
  AOI222XLTS U3495 ( .A0(n88), .A1(n3812), .B0(destinationAddressIn_SOUTH[5]), 
        .B1(n3375), .C0(n4054), .C1(n3835), .Y(n1952) );
  AOI22X1TS U3496 ( .A0(n3363), .A1(n38), .B0(n3989), .B1(n3357), .Y(n1949) );
  AOI222XLTS U3497 ( .A0(n89), .A1(n3820), .B0(destinationAddressIn_SOUTH[4]), 
        .B1(n3383), .C0(n4051), .C1(n3836), .Y(n1950) );
  AOI22X1TS U3498 ( .A0(n3363), .A1(n34), .B0(n3986), .B1(n3356), .Y(n1947) );
  AOI222XLTS U3499 ( .A0(n90), .A1(n3819), .B0(destinationAddressIn_SOUTH[3]), 
        .B1(n3383), .C0(n4048), .C1(n3837), .Y(n1948) );
  AOI22X1TS U3500 ( .A0(n3362), .A1(n24), .B0(n3980), .B1(n3353), .Y(n1943) );
  AOI222XLTS U3501 ( .A0(n91), .A1(n3819), .B0(destinationAddressIn_SOUTH[1]), 
        .B1(n3382), .C0(n4042), .C1(n3834), .Y(n1944) );
  AOI22X1TS U3502 ( .A0(n3363), .A1(n19), .B0(n3977), .B1(n3353), .Y(n1941) );
  AOI222XLTS U3503 ( .A0(n92), .A1(n3819), .B0(destinationAddressIn_SOUTH[0]), 
        .B1(n3382), .C0(n4039), .C1(n3835), .Y(n1942) );
  AOI22X1TS U3504 ( .A0(n479), .A1(n3365), .B0(n4322), .B1(n3352), .Y(n1414)
         );
  AOI222XLTS U3505 ( .A0(n93), .A1(n3817), .B0(dataIn_SOUTH[27]), .B1(n3381), 
        .C0(n4156), .C1(n3840), .Y(n1415) );
  AOI22X1TS U3506 ( .A0(n489), .A1(n3369), .B0(n4271), .B1(n3347), .Y(n1380)
         );
  AOI222XLTS U3507 ( .A0(n94), .A1(n3813), .B0(dataIn_SOUTH[10]), .B1(n3376), 
        .C0(n4105), .C1(n3831), .Y(n1381) );
  AOI22X1TS U3508 ( .A0(n537), .A1(n3371), .B0(n4244), .B1(n3345), .Y(n1362)
         );
  AOI222XLTS U3509 ( .A0(n95), .A1(n3821), .B0(dataIn_SOUTH[1]), .B1(n3375), 
        .C0(n4078), .C1(n3828), .Y(n1363) );
  AOI22X1TS U3510 ( .A0(n511), .A1(n3370), .B0(n4334), .B1(n3353), .Y(n1422)
         );
  AOI222XLTS U3511 ( .A0(n96), .A1(n3818), .B0(dataIn_SOUTH[31]), .B1(n3382), 
        .C0(n4168), .C1(n3834), .Y(n1423) );
  AOI22X1TS U3512 ( .A0(n519), .A1(n3365), .B0(n4313), .B1(n3351), .Y(n1408)
         );
  AOI222XLTS U3513 ( .A0(n97), .A1(n3817), .B0(dataIn_SOUTH[24]), .B1(n3380), 
        .C0(n4147), .C1(n3839), .Y(n1409) );
  AOI22X1TS U3514 ( .A0(n521), .A1(n3365), .B0(n4307), .B1(n3351), .Y(n1404)
         );
  AOI222XLTS U3515 ( .A0(n98), .A1(n3816), .B0(dataIn_SOUTH[22]), .B1(n3380), 
        .C0(n4141), .C1(n736), .Y(n1405) );
  AOI22X1TS U3516 ( .A0(n509), .A1(n3374), .B0(n4289), .B1(n3349), .Y(n1392)
         );
  AOI222XLTS U3517 ( .A0(n99), .A1(n3815), .B0(dataIn_SOUTH[16]), .B1(n3378), 
        .C0(n4123), .C1(n3832), .Y(n1393) );
  AOI22X1TS U3518 ( .A0(n497), .A1(n3373), .B0(n4259), .B1(n3347), .Y(n1372)
         );
  AOI222XLTS U3519 ( .A0(n3820), .A1(n666), .B0(dataIn_SOUTH[6]), .B1(n3379), 
        .C0(n4093), .C1(n3830), .Y(n1373) );
  AOI22X1TS U3520 ( .A0(n505), .A1(n3373), .B0(n4247), .B1(n3346), .Y(n1364)
         );
  AOI222XLTS U3521 ( .A0(n3826), .A1(n665), .B0(dataIn_SOUTH[2]), .B1(n3391), 
        .C0(n4081), .C1(n3829), .Y(n1365) );
  AOI22X1TS U3522 ( .A0(n539), .A1(n3369), .B0(n4241), .B1(n3345), .Y(n1360)
         );
  AOI222XLTS U3523 ( .A0(n3820), .A1(n664), .B0(dataIn_SOUTH[0]), .B1(n3375), 
        .C0(n4075), .C1(n3828), .Y(n1361) );
  AOI32XLTS U3524 ( .A0(n444), .A1(n1784), .A2(n1785), .B0(n3906), .B1(n710), 
        .Y(n2567) );
  OAI221XLTS U3525 ( .A0(n467), .A1(n132), .B0(n159), .B1(n577), .C0(n1913), 
        .Y(n2507) );
  AOI222XLTS U3526 ( .A0(n4239), .A1(n3492), .B0(n3975), .B1(n3476), .C0(n4016), .C1(n3522), .Y(n1913) );
  NAND2X1TS U3527 ( .A(readIn_SOUTH), .B(n1806), .Y(n1800) );
  AOI21X1TS U3528 ( .A0(n4190), .A1(n754), .B0(n1802), .Y(n1801) );
  NAND2X1TS U3529 ( .A(n4189), .B(n752), .Y(n1814) );
  OAI33XLTS U3530 ( .A0(n4197), .A1(n752), .A2(n443), .B0(n972), .B1(n927), 
        .B2(n1818), .Y(n1817) );
  OAI22X1TS U3531 ( .A0(n1086), .A1(n1087), .B0(n925), .B1(n1088), .Y(n2888)
         );
  OAI22X1TS U3532 ( .A0(n1087), .A1(n1089), .B0(n926), .B1(n1088), .Y(n2887)
         );
  AOI221X1TS U3533 ( .A0(n1078), .A1(n4430), .B0(n2921), .B1(n4163), .C0(n2375), .Y(n2371) );
  OAI22X1TS U3534 ( .A0(n4432), .A1(n3091), .B0(n881), .B1(n3758), .Y(n2375)
         );
  AOI221X1TS U3535 ( .A0(n1078), .A1(n4427), .B0(n2923), .B1(n4160), .C0(n2369), .Y(n2365) );
  OAI22X1TS U3536 ( .A0(n4441), .A1(n3091), .B0(n880), .B1(n3758), .Y(n2369)
         );
  AOI221X1TS U3537 ( .A0(n1078), .A1(n4422), .B0(n2923), .B1(n4157), .C0(n2363), .Y(n2359) );
  OAI22X1TS U3538 ( .A0(n4450), .A1(n3091), .B0(n879), .B1(n3758), .Y(n2363)
         );
  AOI221X1TS U3539 ( .A0(n1079), .A1(n4419), .B0(n2922), .B1(n4154), .C0(n2357), .Y(n2353) );
  OAI22X1TS U3540 ( .A0(n4459), .A1(n3091), .B0(n878), .B1(n3759), .Y(n2357)
         );
  AOI221X1TS U3541 ( .A0(n1079), .A1(n4416), .B0(n2921), .B1(n4151), .C0(n2351), .Y(n2347) );
  OAI22X1TS U3542 ( .A0(n4468), .A1(n3090), .B0(n877), .B1(n3759), .Y(n2351)
         );
  AOI221X1TS U3543 ( .A0(n1079), .A1(n4413), .B0(n2922), .B1(n4148), .C0(n2345), .Y(n2341) );
  OAI22X1TS U3544 ( .A0(n4477), .A1(n3090), .B0(n859), .B1(n3759), .Y(n2345)
         );
  AOI221X1TS U3545 ( .A0(n1079), .A1(n4410), .B0(n2925), .B1(n4145), .C0(n2339), .Y(n2335) );
  OAI22X1TS U3546 ( .A0(n4486), .A1(n3090), .B0(n876), .B1(n3759), .Y(n2339)
         );
  AOI221X1TS U3547 ( .A0(n1080), .A1(n4407), .B0(n2919), .B1(n4142), .C0(n2333), .Y(n2329) );
  OAI22X1TS U3548 ( .A0(n4495), .A1(n3090), .B0(n858), .B1(n3770), .Y(n2333)
         );
  AOI221X1TS U3549 ( .A0(n1080), .A1(n4404), .B0(n2919), .B1(n4139), .C0(n2327), .Y(n2323) );
  OAI22X1TS U3550 ( .A0(n4504), .A1(n3089), .B0(n875), .B1(n3770), .Y(n2327)
         );
  AOI221X1TS U3551 ( .A0(n1080), .A1(n4401), .B0(n2919), .B1(n4136), .C0(n2321), .Y(n2317) );
  OAI22X1TS U3552 ( .A0(n4513), .A1(n3089), .B0(n874), .B1(n3767), .Y(n2321)
         );
  AOI221X1TS U3553 ( .A0(n1080), .A1(n4398), .B0(n2919), .B1(n4133), .C0(n2315), .Y(n2311) );
  OAI22X1TS U3554 ( .A0(n4522), .A1(n3089), .B0(n857), .B1(n3767), .Y(n2315)
         );
  AOI221X1TS U3555 ( .A0(n1081), .A1(n4395), .B0(n2918), .B1(n4130), .C0(n2309), .Y(n2305) );
  OAI22X1TS U3556 ( .A0(n4531), .A1(n3089), .B0(n873), .B1(n3770), .Y(n2309)
         );
  AOI221X1TS U3557 ( .A0(n1081), .A1(n4392), .B0(n2918), .B1(n4127), .C0(n2303), .Y(n2299) );
  OAI22X1TS U3558 ( .A0(n4540), .A1(n3088), .B0(n856), .B1(n3770), .Y(n2303)
         );
  AOI221X1TS U3559 ( .A0(n1081), .A1(n4389), .B0(n2918), .B1(n4124), .C0(n2297), .Y(n2293) );
  OAI22X1TS U3560 ( .A0(n4549), .A1(n3088), .B0(n872), .B1(n3768), .Y(n2297)
         );
  AOI221X1TS U3561 ( .A0(n1081), .A1(n4386), .B0(n2918), .B1(n4121), .C0(n2291), .Y(n2287) );
  OAI22X1TS U3562 ( .A0(n4558), .A1(n3088), .B0(n871), .B1(n3771), .Y(n2291)
         );
  AOI221X1TS U3563 ( .A0(n1082), .A1(n4383), .B0(n2917), .B1(n4118), .C0(n2285), .Y(n2281) );
  OAI22X1TS U3564 ( .A0(n4567), .A1(n3088), .B0(n855), .B1(n3760), .Y(n2285)
         );
  AOI221X1TS U3565 ( .A0(n1082), .A1(n4380), .B0(n2917), .B1(n4115), .C0(n2279), .Y(n2275) );
  OAI22X1TS U3566 ( .A0(n4576), .A1(n3087), .B0(n870), .B1(n3760), .Y(n2279)
         );
  AOI221X1TS U3567 ( .A0(n1082), .A1(n4377), .B0(n2917), .B1(n4112), .C0(n2273), .Y(n2269) );
  OAI22X1TS U3568 ( .A0(n4585), .A1(n3087), .B0(n854), .B1(n3760), .Y(n2273)
         );
  AOI221X1TS U3569 ( .A0(n1082), .A1(n4374), .B0(n2917), .B1(n4109), .C0(n2267), .Y(n2263) );
  OAI22X1TS U3570 ( .A0(n4594), .A1(n3087), .B0(n869), .B1(n3760), .Y(n2267)
         );
  AOI221X1TS U3571 ( .A0(n1084), .A1(n4371), .B0(n2916), .B1(n4106), .C0(n2261), .Y(n2257) );
  OAI22X1TS U3572 ( .A0(n4603), .A1(n3087), .B0(n868), .B1(n3761), .Y(n2261)
         );
  AOI221X1TS U3573 ( .A0(n1084), .A1(n4368), .B0(n2916), .B1(n4103), .C0(n2255), .Y(n2251) );
  OAI22X1TS U3574 ( .A0(n4612), .A1(n3086), .B0(n867), .B1(n3761), .Y(n2255)
         );
  AOI221X1TS U3575 ( .A0(n1084), .A1(n4365), .B0(n2916), .B1(n4100), .C0(n2249), .Y(n2245) );
  OAI22X1TS U3576 ( .A0(n4621), .A1(n3086), .B0(n866), .B1(n3761), .Y(n2249)
         );
  AOI221X1TS U3577 ( .A0(n1084), .A1(n4362), .B0(n2916), .B1(n4097), .C0(n2243), .Y(n2239) );
  OAI22X1TS U3578 ( .A0(n4630), .A1(n3086), .B0(n865), .B1(n3761), .Y(n2243)
         );
  AOI221X1TS U3579 ( .A0(n1085), .A1(n4359), .B0(n2922), .B1(n4094), .C0(n2237), .Y(n2233) );
  OAI22X1TS U3580 ( .A0(n4639), .A1(n3085), .B0(n850), .B1(n3762), .Y(n2237)
         );
  AOI221X1TS U3581 ( .A0(n1085), .A1(n4356), .B0(n2925), .B1(n4091), .C0(n2231), .Y(n2227) );
  OAI22X1TS U3582 ( .A0(n4648), .A1(n3085), .B0(n864), .B1(n3762), .Y(n2231)
         );
  AOI221X1TS U3583 ( .A0(n1085), .A1(n4353), .B0(n2924), .B1(n4088), .C0(n2225), .Y(n2221) );
  OAI22X1TS U3584 ( .A0(n4657), .A1(n3085), .B0(n853), .B1(n3762), .Y(n2225)
         );
  AOI221X1TS U3585 ( .A0(n1085), .A1(n4350), .B0(n2925), .B1(n4085), .C0(n2219), .Y(n2215) );
  OAI22X1TS U3586 ( .A0(n4666), .A1(n3085), .B0(n852), .B1(n3762), .Y(n2219)
         );
  AOI221X1TS U3587 ( .A0(n1091), .A1(n4347), .B0(n2922), .B1(n4082), .C0(n2213), .Y(n2209) );
  OAI22X1TS U3588 ( .A0(n4675), .A1(n3084), .B0(n863), .B1(n3763), .Y(n2213)
         );
  AOI221X1TS U3589 ( .A0(n1091), .A1(n4344), .B0(n2920), .B1(n4079), .C0(n2207), .Y(n2203) );
  OAI22X1TS U3590 ( .A0(n4684), .A1(n3084), .B0(n851), .B1(n3763), .Y(n2207)
         );
  AOI221X1TS U3591 ( .A0(n1091), .A1(n4341), .B0(n2924), .B1(n4076), .C0(n2201), .Y(n2197) );
  OAI22X1TS U3592 ( .A0(n4693), .A1(n3084), .B0(n862), .B1(n3763), .Y(n2201)
         );
  AOI221X1TS U3593 ( .A0(n1091), .A1(n4338), .B0(n2054), .B1(n4073), .C0(n2195), .Y(n2191) );
  OAI22X1TS U3594 ( .A0(n4702), .A1(n3084), .B0(n861), .B1(n3763), .Y(n2195)
         );
  AOI221X1TS U3595 ( .A0(n1134), .A1(n3951), .B0(n2906), .B1(n4052), .C0(n2153), .Y(n2149) );
  OAI22X1TS U3596 ( .A0(n4715), .A1(n3083), .B0(n887), .B1(n3765), .Y(n2153)
         );
  AOI221X1TS U3597 ( .A0(n1134), .A1(n3948), .B0(n2906), .B1(n4049), .C0(n2147), .Y(n2143) );
  OAI22X1TS U3598 ( .A0(n4724), .A1(n3083), .B0(n886), .B1(n3765), .Y(n2147)
         );
  AOI221X1TS U3599 ( .A0(n1151), .A1(n3945), .B0(n2905), .B1(n4046), .C0(n2141), .Y(n2137) );
  OAI22X1TS U3600 ( .A0(n4733), .A1(n3086), .B0(n885), .B1(n3766), .Y(n2141)
         );
  AOI221X1TS U3601 ( .A0(n1151), .A1(n3942), .B0(n2905), .B1(n4043), .C0(n2135), .Y(n2131) );
  OAI22X1TS U3602 ( .A0(n4742), .A1(n3083), .B0(n860), .B1(n3766), .Y(n2135)
         );
  AOI221X1TS U3603 ( .A0(n1151), .A1(n3936), .B0(n2905), .B1(n4037), .C0(n2122), .Y(n2111) );
  OAI22X1TS U3604 ( .A0(n4760), .A1(n3083), .B0(n883), .B1(n3766), .Y(n2122)
         );
  INVX2TS U3605 ( .A(n2051), .Y(n922) );
  OAI221XLTS U3606 ( .A0(n4194), .A1(n2025), .B0(n148), .B1(n2023), .C0(n6253), 
        .Y(n2051) );
  AOI221X1TS U3607 ( .A0(n1078), .A1(n4434), .B0(n2920), .B1(n4166), .C0(n2381), .Y(n2377) );
  OAI22X1TS U3608 ( .A0(n4423), .A1(n3082), .B0(n882), .B1(n3758), .Y(n2381)
         );
  AOI221X1TS U3609 ( .A0(n1107), .A1(n4185), .B0(n2915), .B1(n4070), .C0(n2189), .Y(n2185) );
  OAI22X1TS U3610 ( .A0(n3082), .A1(n4711), .B0(n892), .B1(n3764), .Y(n2189)
         );
  AOI221X1TS U3611 ( .A0(n1107), .A1(n4182), .B0(n2915), .B1(n4067), .C0(n2183), .Y(n2179) );
  OAI22X1TS U3612 ( .A0(n3082), .A1(n4712), .B0(n893), .B1(n3764), .Y(n2183)
         );
  AOI221X1TS U3613 ( .A0(n1107), .A1(n4176), .B0(n2915), .B1(n4061), .C0(n2171), .Y(n2167) );
  OAI22X1TS U3614 ( .A0(n3081), .A1(n4713), .B0(n890), .B1(n3764), .Y(n2171)
         );
  AOI221X1TS U3615 ( .A0(n1134), .A1(n4173), .B0(n2906), .B1(n4058), .C0(n2165), .Y(n2161) );
  OAI22X1TS U3616 ( .A0(n3081), .A1(n4714), .B0(n889), .B1(n3765), .Y(n2165)
         );
  AOI221X1TS U3617 ( .A0(n1151), .A1(n3939), .B0(n2905), .B1(n4040), .C0(n2129), .Y(n2125) );
  OAI22X1TS U3618 ( .A0(n4751), .A1(n3082), .B0(n884), .B1(n3766), .Y(n2129)
         );
  AOI221X1TS U3619 ( .A0(n1107), .A1(n4179), .B0(n2915), .B1(n4064), .C0(n2177), .Y(n2173) );
  OAI22X1TS U3620 ( .A0(n3081), .A1(n4838), .B0(n891), .B1(n3764), .Y(n2177)
         );
  AOI221X1TS U3621 ( .A0(n1134), .A1(n4170), .B0(n2906), .B1(n4055), .C0(n2159), .Y(n2155) );
  OAI22X1TS U3622 ( .A0(n3081), .A1(n4837), .B0(n888), .B1(n3765), .Y(n2159)
         );
  NAND4X1TS U3623 ( .A(n2376), .B(n2377), .C(n2378), .D(n2379), .Y(n2397) );
  AOI222XLTS U3624 ( .A0(n1007), .A1(n700), .B0(n993), .B1(n2934), .C0(n991), 
        .C1(n2933), .Y(n2378) );
  AOI221X1TS U3625 ( .A0(n1064), .A1(n3012), .B0(n1050), .B1(n96), .C0(n2380), 
        .Y(n2379) );
  AOI222XLTS U3626 ( .A0(n3058), .A1(dataIn_SOUTH[31]), .B0(n3066), .B1(n4335), 
        .C0(n2123), .C1(cacheDataOut[31]), .Y(n2376) );
  NAND4X1TS U3627 ( .A(n2370), .B(n2371), .C(n2372), .D(n2373), .Y(n2398) );
  AOI222XLTS U3628 ( .A0(n1007), .A1(n699), .B0(n993), .B1(n2936), .C0(n991), 
        .C1(n2935), .Y(n2372) );
  AOI221X1TS U3629 ( .A0(n1064), .A1(n3013), .B0(n1050), .B1(n66), .C0(n2374), 
        .Y(n2373) );
  AOI222XLTS U3630 ( .A0(n3061), .A1(n4519), .B0(n3073), .B1(n4332), .C0(n2123), .C1(cacheDataOut[30]), .Y(n2370) );
  NAND4X1TS U3631 ( .A(n2364), .B(n2365), .C(n2366), .D(n2367), .Y(n2399) );
  AOI222XLTS U3632 ( .A0(n1007), .A1(n698), .B0(n993), .B1(n2938), .C0(n991), 
        .C1(n2937), .Y(n2366) );
  AOI221X1TS U3633 ( .A0(n1064), .A1(n3014), .B0(n1050), .B1(n67), .C0(n2368), 
        .Y(n2367) );
  AOI222XLTS U3634 ( .A0(n3060), .A1(dataIn_SOUTH[29]), .B0(n3073), .B1(n4329), 
        .C0(n977), .C1(cacheDataOut[29]), .Y(n2364) );
  NAND4X1TS U3635 ( .A(n2358), .B(n2359), .C(n2360), .D(n2361), .Y(n2400) );
  AOI222XLTS U3636 ( .A0(n1007), .A1(n56), .B0(n993), .B1(n2940), .C0(n990), 
        .C1(n2939), .Y(n2360) );
  AOI221X1TS U3637 ( .A0(n1064), .A1(n3015), .B0(n1050), .B1(n68), .C0(n2362), 
        .Y(n2361) );
  AOI222XLTS U3638 ( .A0(n3059), .A1(n4515), .B0(n3073), .B1(n4326), .C0(n976), 
        .C1(cacheDataOut[28]), .Y(n2358) );
  NAND4X1TS U3639 ( .A(n2352), .B(n2353), .C(n2354), .D(n2355), .Y(n2401) );
  AOI222XLTS U3640 ( .A0(n1017), .A1(n57), .B0(n1004), .B1(n2942), .C0(n979), 
        .C1(n2941), .Y(n2354) );
  AOI221X1TS U3641 ( .A0(n1076), .A1(n3016), .B0(n1060), .B1(n93), .C0(n2356), 
        .Y(n2355) );
  AOI222XLTS U3642 ( .A0(n3058), .A1(dataIn_SOUTH[27]), .B0(n3073), .B1(n4323), 
        .C0(n928), .C1(cacheDataOut[27]), .Y(n2352) );
  NAND4X1TS U3643 ( .A(n2346), .B(n2347), .C(n2348), .D(n2349), .Y(n2402) );
  AOI222XLTS U3644 ( .A0(n1017), .A1(n697), .B0(n1005), .B1(n2944), .C0(n979), 
        .C1(n2943), .Y(n2348) );
  AOI221X1TS U3645 ( .A0(n1074), .A1(n3017), .B0(n1060), .B1(n69), .C0(n2350), 
        .Y(n2349) );
  AOI222XLTS U3646 ( .A0(n3057), .A1(n4510), .B0(n3072), .B1(n4320), .C0(n928), 
        .C1(cacheDataOut[26]), .Y(n2346) );
  NAND4X1TS U3647 ( .A(n2340), .B(n2341), .C(n2342), .D(n2343), .Y(n2403) );
  AOI222XLTS U3648 ( .A0(n1016), .A1(n696), .B0(n1006), .B1(n2946), .C0(n979), 
        .C1(n2945), .Y(n2342) );
  AOI221X1TS U3649 ( .A0(n1077), .A1(n3018), .B0(n1061), .B1(n70), .C0(n2344), 
        .Y(n2343) );
  AOI222XLTS U3650 ( .A0(n2040), .A1(dataIn_SOUTH[25]), .B0(n3072), .B1(n4317), 
        .C0(n928), .C1(cacheDataOut[25]), .Y(n2340) );
  NAND4X1TS U3651 ( .A(n2334), .B(n2335), .C(n2336), .D(n2337), .Y(n2404) );
  AOI222XLTS U3652 ( .A0(n1015), .A1(n695), .B0(n1004), .B1(n2948), .C0(n979), 
        .C1(n2947), .Y(n2336) );
  AOI221X1TS U3653 ( .A0(n1075), .A1(n3019), .B0(n1059), .B1(n97), .C0(n2338), 
        .Y(n2337) );
  AOI222XLTS U3654 ( .A0(n3057), .A1(n4503), .B0(n3072), .B1(n4314), .C0(n928), 
        .C1(cacheDataOut[24]), .Y(n2334) );
  NAND4X1TS U3655 ( .A(n2328), .B(n2329), .C(n2330), .D(n2331), .Y(n2405) );
  AOI222XLTS U3656 ( .A0(n1016), .A1(n58), .B0(n2120), .B1(n2950), .C0(n980), 
        .C1(n2949), .Y(n2330) );
  AOI221X1TS U3657 ( .A0(n1073), .A1(n3020), .B0(n1059), .B1(n71), .C0(n2332), 
        .Y(n2331) );
  AOI222XLTS U3658 ( .A0(n3063), .A1(n4501), .B0(n3072), .B1(n4311), .C0(n932), 
        .C1(cacheDataOut[23]), .Y(n2328) );
  NAND4X1TS U3659 ( .A(n2322), .B(n2323), .C(n2324), .D(n2325), .Y(n2406) );
  AOI222XLTS U3660 ( .A0(n1015), .A1(n694), .B0(n1005), .B1(n2952), .C0(n980), 
        .C1(n2951), .Y(n2324) );
  AOI221X1TS U3661 ( .A0(n1076), .A1(n3021), .B0(n1058), .B1(n98), .C0(n2326), 
        .Y(n2325) );
  AOI222XLTS U3662 ( .A0(n3063), .A1(dataIn_SOUTH[22]), .B0(n3071), .B1(n4308), 
        .C0(n932), .C1(cacheDataOut[22]), .Y(n2322) );
  NAND4X1TS U3663 ( .A(n2316), .B(n2317), .C(n2318), .D(n2319), .Y(n2407) );
  AOI222XLTS U3664 ( .A0(n1020), .A1(n693), .B0(n1003), .B1(n2954), .C0(n980), 
        .C1(n2953), .Y(n2318) );
  AOI221X1TS U3665 ( .A0(n2114), .A1(n3022), .B0(n1057), .B1(n72), .C0(n2320), 
        .Y(n2319) );
  AOI222XLTS U3666 ( .A0(n3061), .A1(dataIn_SOUTH[21]), .B0(n3071), .B1(n4305), 
        .C0(n932), .C1(cacheDataOut[21]), .Y(n2316) );
  NAND4X1TS U3667 ( .A(n2310), .B(n2311), .C(n2312), .D(n2313), .Y(n2408) );
  AOI222XLTS U3668 ( .A0(n1019), .A1(n59), .B0(n1005), .B1(n2956), .C0(n980), 
        .C1(n2955), .Y(n2312) );
  AOI221X1TS U3669 ( .A0(n1077), .A1(n3023), .B0(n1060), .B1(n73), .C0(n2314), 
        .Y(n2313) );
  AOI222XLTS U3670 ( .A0(n3062), .A1(n4493), .B0(n3071), .B1(n4302), .C0(n932), 
        .C1(cacheDataOut[20]), .Y(n2310) );
  NAND4X1TS U3671 ( .A(n2304), .B(n2305), .C(n2306), .D(n2307), .Y(n2409) );
  AOI222XLTS U3672 ( .A0(n1019), .A1(n692), .B0(n994), .B1(n2958), .C0(n981), 
        .C1(n2957), .Y(n2306) );
  AOI221X1TS U3673 ( .A0(n1065), .A1(n3024), .B0(n1061), .B1(n74), .C0(n2308), 
        .Y(n2307) );
  AOI222XLTS U3674 ( .A0(n3009), .A1(dataIn_SOUTH[19]), .B0(n3071), .B1(n4299), 
        .C0(n933), .C1(cacheDataOut[19]), .Y(n2304) );
  NAND4X1TS U3675 ( .A(n2298), .B(n2299), .C(n2300), .D(n2301), .Y(n2410) );
  AOI222XLTS U3676 ( .A0(n1018), .A1(n691), .B0(n994), .B1(n2960), .C0(n981), 
        .C1(n2959), .Y(n2300) );
  AOI221X1TS U3677 ( .A0(n1065), .A1(n3025), .B0(n1062), .B1(n75), .C0(n2302), 
        .Y(n2301) );
  AOI222XLTS U3678 ( .A0(n3009), .A1(dataIn_SOUTH[18]), .B0(n3075), .B1(n4296), 
        .C0(n933), .C1(cacheDataOut[18]), .Y(n2298) );
  NAND4X1TS U3679 ( .A(n2292), .B(n2293), .C(n2294), .D(n2295), .Y(n2411) );
  AOI222XLTS U3680 ( .A0(n1019), .A1(n690), .B0(n994), .B1(n2962), .C0(n981), 
        .C1(n2961), .Y(n2294) );
  AOI221X1TS U3681 ( .A0(n1065), .A1(n3026), .B0(n1058), .B1(n76), .C0(n2296), 
        .Y(n2295) );
  AOI222XLTS U3682 ( .A0(n3009), .A1(dataIn_SOUTH[17]), .B0(n3076), .B1(n4293), 
        .C0(n933), .C1(cacheDataOut[17]), .Y(n2292) );
  NAND4X1TS U3683 ( .A(n2286), .B(n2287), .C(n2288), .D(n2289), .Y(n2412) );
  AOI222XLTS U3684 ( .A0(n1018), .A1(n689), .B0(n994), .B1(n2964), .C0(n981), 
        .C1(n2963), .Y(n2288) );
  AOI221X1TS U3685 ( .A0(n1065), .A1(n3027), .B0(n1060), .B1(n99), .C0(n2290), 
        .Y(n2289) );
  AOI222XLTS U3686 ( .A0(n3009), .A1(n4482), .B0(n3077), .B1(n4290), .C0(n933), 
        .C1(cacheDataOut[16]), .Y(n2286) );
  NAND4X1TS U3687 ( .A(n2280), .B(n2281), .C(n2282), .D(n2283), .Y(n2413) );
  AOI222XLTS U3688 ( .A0(n1008), .A1(n688), .B0(n995), .B1(n2966), .C0(n982), 
        .C1(n2965), .Y(n2282) );
  AOI221X1TS U3689 ( .A0(n1066), .A1(n3028), .B0(n1057), .B1(n77), .C0(n2284), 
        .Y(n2283) );
  AOI222XLTS U3690 ( .A0(n3010), .A1(dataIn_SOUTH[15]), .B0(n3074), .B1(n4287), 
        .C0(n976), .C1(cacheDataOut[15]), .Y(n2280) );
  NAND4X1TS U3691 ( .A(n2274), .B(n2275), .C(n2276), .D(n2277), .Y(n2414) );
  AOI222XLTS U3692 ( .A0(n1008), .A1(n687), .B0(n995), .B1(n2968), .C0(n982), 
        .C1(n2967), .Y(n2276) );
  AOI221X1TS U3693 ( .A0(n1066), .A1(n3029), .B0(n1061), .B1(n78), .C0(n2278), 
        .Y(n2277) );
  AOI222XLTS U3694 ( .A0(n3010), .A1(n4475), .B0(n3075), .B1(n4284), .C0(n975), 
        .C1(cacheDataOut[14]), .Y(n2274) );
  NAND4X1TS U3695 ( .A(n2268), .B(n2269), .C(n2270), .D(n2271), .Y(n2415) );
  AOI222XLTS U3696 ( .A0(n1008), .A1(n686), .B0(n995), .B1(n2970), .C0(n982), 
        .C1(n2969), .Y(n2270) );
  AOI221X1TS U3697 ( .A0(n1066), .A1(n3030), .B0(n1062), .B1(n79), .C0(n2272), 
        .Y(n2271) );
  AOI222XLTS U3698 ( .A0(n3010), .A1(n4471), .B0(n3075), .B1(n4281), .C0(n974), 
        .C1(cacheDataOut[13]), .Y(n2268) );
  NAND4X1TS U3699 ( .A(n2262), .B(n2263), .C(n2264), .D(n2265), .Y(n2416) );
  AOI222XLTS U3700 ( .A0(n1008), .A1(n46), .B0(n995), .B1(n2972), .C0(n982), 
        .C1(n2971), .Y(n2264) );
  AOI221X1TS U3701 ( .A0(n1066), .A1(n3031), .B0(n1063), .B1(n80), .C0(n2266), 
        .Y(n2265) );
  AOI222XLTS U3702 ( .A0(n3010), .A1(dataIn_SOUTH[12]), .B0(n3074), .B1(n4278), 
        .C0(n975), .C1(cacheDataOut[12]), .Y(n2262) );
  NAND4X1TS U3703 ( .A(n2256), .B(n2257), .C(n2258), .D(n2259), .Y(n2417) );
  AOI222XLTS U3704 ( .A0(n1009), .A1(n47), .B0(n996), .B1(n2974), .C0(n2121), 
        .C1(n2973), .Y(n2258) );
  AOI221X1TS U3705 ( .A0(n1067), .A1(n3032), .B0(n1051), .B1(n81), .C0(n2260), 
        .Y(n2259) );
  AOI222XLTS U3706 ( .A0(n3011), .A1(dataIn_SOUTH[11]), .B0(n3075), .B1(n4275), 
        .C0(n956), .C1(cacheDataOut[11]), .Y(n2256) );
  NAND4X1TS U3707 ( .A(n2250), .B(n2251), .C(n2252), .D(n2253), .Y(n2418) );
  AOI222XLTS U3708 ( .A0(n1009), .A1(n48), .B0(n996), .B1(n2976), .C0(n990), 
        .C1(n2975), .Y(n2252) );
  AOI221X1TS U3709 ( .A0(n1067), .A1(n3033), .B0(n1051), .B1(n94), .C0(n2254), 
        .Y(n2253) );
  AOI222XLTS U3710 ( .A0(n3011), .A1(n4464), .B0(n3078), .B1(n4272), .C0(n956), 
        .C1(cacheDataOut[10]), .Y(n2250) );
  NAND4X1TS U3711 ( .A(n2244), .B(n2245), .C(n2246), .D(n2247), .Y(n2419) );
  AOI222XLTS U3712 ( .A0(n1009), .A1(n60), .B0(n996), .B1(n2978), .C0(n989), 
        .C1(n2977), .Y(n2246) );
  AOI221X1TS U3713 ( .A0(n1067), .A1(n3034), .B0(n1051), .B1(n82), .C0(n2248), 
        .Y(n2247) );
  AOI222XLTS U3714 ( .A0(n3011), .A1(n4462), .B0(n3078), .B1(n4269), .C0(n956), 
        .C1(cacheDataOut[9]), .Y(n2244) );
  NAND4X1TS U3715 ( .A(n2238), .B(n2239), .C(n2240), .D(n2241), .Y(n2420) );
  AOI222XLTS U3716 ( .A0(n1009), .A1(n49), .B0(n996), .B1(n2980), .C0(n988), 
        .C1(n2979), .Y(n2240) );
  AOI221X1TS U3717 ( .A0(n1067), .A1(n3035), .B0(n1051), .B1(n83), .C0(n2242), 
        .Y(n2241) );
  AOI222XLTS U3718 ( .A0(n3011), .A1(dataIn_SOUTH[8]), .B0(n3076), .B1(n4266), 
        .C0(n956), .C1(cacheDataOut[8]), .Y(n2238) );
  NAND4X1TS U3719 ( .A(n2232), .B(n2233), .C(n2234), .D(n2235), .Y(n2421) );
  AOI222XLTS U3720 ( .A0(n1010), .A1(n50), .B0(n997), .B1(n2982), .C0(n983), 
        .C1(n2981), .Y(n2234) );
  AOI221X1TS U3721 ( .A0(n1068), .A1(n3036), .B0(n1052), .B1(n84), .C0(n2236), 
        .Y(n2235) );
  AOI222XLTS U3722 ( .A0(n3050), .A1(n4456), .B0(n3077), .B1(n4263), .C0(n961), 
        .C1(cacheDataOut[7]), .Y(n2232) );
  NAND4X1TS U3723 ( .A(n2226), .B(n2227), .C(n2228), .D(n2229), .Y(n2422) );
  AOI222XLTS U3724 ( .A0(n1010), .A1(n51), .B0(n997), .B1(n2984), .C0(n983), 
        .C1(n2983), .Y(n2228) );
  AOI221X1TS U3725 ( .A0(n1068), .A1(n3037), .B0(n1052), .B1(n666), .C0(n2230), 
        .Y(n2229) );
  AOI222XLTS U3726 ( .A0(n3050), .A1(dataIn_SOUTH[6]), .B0(n3070), .B1(n4260), 
        .C0(n961), .C1(cacheDataOut[6]), .Y(n2226) );
  NAND4X1TS U3727 ( .A(n2220), .B(n2221), .C(n2222), .D(n2223), .Y(n2423) );
  AOI222XLTS U3728 ( .A0(n1010), .A1(n61), .B0(n997), .B1(n2986), .C0(n983), 
        .C1(n2985), .Y(n2222) );
  AOI221X1TS U3729 ( .A0(n1068), .A1(n3038), .B0(n1052), .B1(n85), .C0(n2224), 
        .Y(n2223) );
  AOI222XLTS U3730 ( .A0(n3050), .A1(dataIn_SOUTH[5]), .B0(n3070), .B1(n4257), 
        .C0(n961), .C1(cacheDataOut[5]), .Y(n2220) );
  NAND4X1TS U3731 ( .A(n2214), .B(n2215), .C(n2216), .D(n2217), .Y(n2424) );
  AOI222XLTS U3732 ( .A0(n1010), .A1(n52), .B0(n997), .B1(n2988), .C0(n983), 
        .C1(n2987), .Y(n2216) );
  AOI221X1TS U3733 ( .A0(n1068), .A1(n3039), .B0(n1052), .B1(n86), .C0(n2218), 
        .Y(n2217) );
  AOI222XLTS U3734 ( .A0(n3050), .A1(n4449), .B0(n3070), .B1(n4254), .C0(n961), 
        .C1(cacheDataOut[4]), .Y(n2214) );
  NAND4X1TS U3735 ( .A(n2208), .B(n2209), .C(n2210), .D(n2211), .Y(n2425) );
  AOI222XLTS U3736 ( .A0(n1011), .A1(n53), .B0(n998), .B1(n2990), .C0(n984), 
        .C1(n2989), .Y(n2210) );
  AOI221X1TS U3737 ( .A0(n1069), .A1(n3040), .B0(n1053), .B1(n87), .C0(n2212), 
        .Y(n2211) );
  AOI222XLTS U3738 ( .A0(n3051), .A1(n4445), .B0(n3069), .B1(n4251), .C0(n962), 
        .C1(cacheDataOut[3]), .Y(n2208) );
  NAND4X1TS U3739 ( .A(n2202), .B(n2203), .C(n2204), .D(n2205), .Y(n2426) );
  AOI222XLTS U3740 ( .A0(n1011), .A1(n62), .B0(n998), .B1(n2992), .C0(n984), 
        .C1(n2991), .Y(n2204) );
  AOI221X1TS U3741 ( .A0(n1069), .A1(n3041), .B0(n1053), .B1(n665), .C0(n2206), 
        .Y(n2205) );
  AOI222XLTS U3742 ( .A0(n3051), .A1(dataIn_SOUTH[2]), .B0(n3069), .B1(n4248), 
        .C0(n962), .C1(cacheDataOut[2]), .Y(n2202) );
  NAND4X1TS U3743 ( .A(n2196), .B(n2197), .C(n2198), .D(n2199), .Y(n2427) );
  AOI222XLTS U3744 ( .A0(n1011), .A1(n63), .B0(n998), .B1(n2994), .C0(n984), 
        .C1(n2993), .Y(n2198) );
  AOI221X1TS U3745 ( .A0(n1069), .A1(n3042), .B0(n1053), .B1(n95), .C0(n2200), 
        .Y(n2199) );
  AOI222XLTS U3746 ( .A0(n3051), .A1(dataIn_SOUTH[1]), .B0(n3069), .B1(n4245), 
        .C0(n962), .C1(cacheDataOut[1]), .Y(n2196) );
  NAND4X1TS U3747 ( .A(n2190), .B(n2191), .C(n2192), .D(n2193), .Y(n2428) );
  AOI222XLTS U3748 ( .A0(n1011), .A1(n64), .B0(n998), .B1(n2996), .C0(n984), 
        .C1(n2995), .Y(n2192) );
  AOI221X1TS U3749 ( .A0(n1069), .A1(n3043), .B0(n1053), .B1(n664), .C0(n2194), 
        .Y(n2193) );
  AOI222XLTS U3750 ( .A0(n3051), .A1(n4438), .B0(n3069), .B1(n4242), .C0(n962), 
        .C1(cacheDataOut[0]), .Y(n2190) );
  NAND4X1TS U3751 ( .A(n2184), .B(n2185), .C(n2186), .D(n2187), .Y(n2429) );
  AOI222XLTS U3752 ( .A0(n1012), .A1(\requesterAddressbuffer[0][5] ), .B0(n999), .B1(\requesterAddressbuffer[6][5] ), .C0(n985), .C1(n2927), .Y(n2186) );
  AOI221X1TS U3753 ( .A0(n1070), .A1(n2909), .B0(n1054), .B1(
        \requesterAddressbuffer[2][5] ), .C0(n2188), .Y(n2187) );
  AOI222XLTS U3754 ( .A0(n3052), .A1(n4538), .B0(n3068), .B1(n4035), .C0(n963), 
        .C1(n41), .Y(n2184) );
  NAND4X1TS U3755 ( .A(n2178), .B(n2179), .C(n2180), .D(n2181), .Y(n2430) );
  AOI222XLTS U3756 ( .A0(n1012), .A1(\requesterAddressbuffer[0][4] ), .B0(n999), .B1(\requesterAddressbuffer[6][4] ), .C0(n985), .C1(n2928), .Y(n2180) );
  AOI221X1TS U3757 ( .A0(n1070), .A1(n2910), .B0(n1054), .B1(
        \requesterAddressbuffer[2][4] ), .C0(n2182), .Y(n2181) );
  AOI222XLTS U3758 ( .A0(n3052), .A1(n4536), .B0(n3068), .B1(n4032), .C0(n963), 
        .C1(readRequesterAddress[4]), .Y(n2178) );
  NAND4X1TS U3759 ( .A(n2166), .B(n2167), .C(n2168), .D(n2169), .Y(n2432) );
  AOI222XLTS U3760 ( .A0(n1012), .A1(\requesterAddressbuffer[0][2] ), .B0(n999), .B1(\requesterAddressbuffer[6][2] ), .C0(n985), .C1(n2929), .Y(n2168) );
  AOI221X1TS U3761 ( .A0(n1070), .A1(n2911), .B0(n1054), .B1(
        \requesterAddressbuffer[2][2] ), .C0(n2170), .Y(n2169) );
  AOI222XLTS U3762 ( .A0(n3052), .A1(requesterAddressIn_SOUTH[2]), .B0(n3068), 
        .B1(n4026), .C0(n963), .C1(readRequesterAddress[2]), .Y(n2166) );
  NAND4X1TS U3763 ( .A(n2160), .B(n2161), .C(n2162), .D(n2163), .Y(n2433) );
  AOI222XLTS U3764 ( .A0(n1013), .A1(\requesterAddressbuffer[0][1] ), .B0(
        n1000), .B1(\requesterAddressbuffer[6][1] ), .C0(n986), .C1(n2930), 
        .Y(n2162) );
  AOI221X1TS U3765 ( .A0(n1071), .A1(n2912), .B0(n1055), .B1(
        \requesterAddressbuffer[2][1] ), .C0(n2164), .Y(n2163) );
  AOI222XLTS U3766 ( .A0(n3053), .A1(n4528), .B0(n3067), .B1(n4023), .C0(n964), 
        .C1(readRequesterAddress[1]), .Y(n2160) );
  NAND4X1TS U3767 ( .A(n2148), .B(n2149), .C(n2150), .D(n2151), .Y(n2435) );
  AOI222XLTS U3768 ( .A0(n1013), .A1(n704), .B0(n1000), .B1(n2998), .C0(n986), 
        .C1(n2997), .Y(n2150) );
  AOI221X1TS U3769 ( .A0(n1071), .A1(n3044), .B0(n1055), .B1(n88), .C0(n2152), 
        .Y(n2151) );
  AOI222XLTS U3770 ( .A0(n3053), .A1(n4216), .B0(n3067), .B1(n3993), .C0(n964), 
        .C1(n14), .Y(n2148) );
  NAND4X1TS U3771 ( .A(n2142), .B(n2143), .C(n2144), .D(n2145), .Y(n2436) );
  AOI222XLTS U3772 ( .A0(n1013), .A1(n54), .B0(n1000), .B1(n3000), .C0(n986), 
        .C1(n2999), .Y(n2144) );
  AOI221X1TS U3773 ( .A0(n1071), .A1(n3045), .B0(n1055), .B1(n89), .C0(n2146), 
        .Y(n2145) );
  AOI222XLTS U3774 ( .A0(n3053), .A1(destinationAddressIn_SOUTH[4]), .B0(n3067), .B1(n3990), .C0(n964), .C1(readRequesterAddress[4]), .Y(n2142) );
  NAND4X1TS U3775 ( .A(n2136), .B(n2137), .C(n2138), .D(n2139), .Y(n2437) );
  AOI222XLTS U3776 ( .A0(n1014), .A1(n703), .B0(n1001), .B1(n3002), .C0(n987), 
        .C1(n3001), .Y(n2138) );
  AOI221X1TS U3777 ( .A0(n1072), .A1(n3046), .B0(n1056), .B1(n90), .C0(n2140), 
        .Y(n2139) );
  AOI222XLTS U3778 ( .A0(n3054), .A1(n4211), .B0(n3070), .B1(n3987), .C0(n965), 
        .C1(readRequesterAddress[3]), .Y(n2136) );
  NAND4X1TS U3779 ( .A(n2130), .B(n2131), .C(n2132), .D(n2133), .Y(n2438) );
  AOI222XLTS U3780 ( .A0(n1014), .A1(n702), .B0(n1001), .B1(n3004), .C0(n987), 
        .C1(n3003), .Y(n2132) );
  AOI221X1TS U3781 ( .A0(n1072), .A1(n3047), .B0(n1056), .B1(n65), .C0(n2134), 
        .Y(n2133) );
  AOI222XLTS U3782 ( .A0(n3054), .A1(n4209), .B0(n3066), .B1(n3984), .C0(n965), 
        .C1(readRequesterAddress[2]), .Y(n2130) );
  NAND4X1TS U3783 ( .A(n2124), .B(n2125), .C(n2126), .D(n2127), .Y(n2439) );
  AOI222XLTS U3784 ( .A0(n1014), .A1(n701), .B0(n1001), .B1(n3006), .C0(n987), 
        .C1(n3005), .Y(n2126) );
  AOI221X1TS U3785 ( .A0(n1072), .A1(n3048), .B0(n1056), .B1(n91), .C0(n2128), 
        .Y(n2127) );
  AOI222XLTS U3786 ( .A0(n3054), .A1(n4206), .B0(n3066), .B1(n3981), .C0(n965), 
        .C1(readRequesterAddress[1]), .Y(n2124) );
  NAND4X1TS U3787 ( .A(n2110), .B(n2111), .C(n2112), .D(n2113), .Y(n2440) );
  AOI222XLTS U3788 ( .A0(n1014), .A1(n55), .B0(n1001), .B1(n3008), .C0(n987), 
        .C1(n3007), .Y(n2112) );
  AOI221X1TS U3789 ( .A0(n1072), .A1(n3049), .B0(n1056), .B1(n92), .C0(n2116), 
        .Y(n2113) );
  AOI222XLTS U3790 ( .A0(n3054), .A1(destinationAddressIn_SOUTH[0]), .B0(n3066), .B1(n3978), .C0(n965), .C1(readRequesterAddress[0]), .Y(n2110) );
  NAND4X1TS U3791 ( .A(n2172), .B(n2173), .C(n2174), .D(n2175), .Y(n2431) );
  AOI222XLTS U3792 ( .A0(n1012), .A1(\requesterAddressbuffer[0][3] ), .B0(n999), .B1(\requesterAddressbuffer[6][3] ), .C0(n985), .C1(n2931), .Y(n2174) );
  AOI221X1TS U3793 ( .A0(n1070), .A1(n2913), .B0(n1054), .B1(
        \requesterAddressbuffer[2][3] ), .C0(n2176), .Y(n2175) );
  AOI222XLTS U3794 ( .A0(n3052), .A1(n4533), .B0(n3068), .B1(n4029), .C0(n963), 
        .C1(readRequesterAddress[3]), .Y(n2172) );
  NAND4X1TS U3795 ( .A(n2154), .B(n2155), .C(n2156), .D(n2157), .Y(n2434) );
  AOI222XLTS U3796 ( .A0(n1013), .A1(\requesterAddressbuffer[0][0] ), .B0(
        n1000), .B1(\requesterAddressbuffer[6][0] ), .C0(n986), .C1(n2932), 
        .Y(n2156) );
  AOI221X1TS U3797 ( .A0(n1071), .A1(n2914), .B0(n1055), .B1(
        \requesterAddressbuffer[2][0] ), .C0(n2158), .Y(n2157) );
  AOI222XLTS U3798 ( .A0(n3053), .A1(n4525), .B0(n3067), .B1(n4020), .C0(n964), 
        .C1(readRequesterAddress[0]), .Y(n2154) );
  OAI21X1TS U3799 ( .A0(n152), .A1(n922), .B0(n652), .Y(n2041) );
  INVX2TS U3800 ( .A(n2042), .Y(n652) );
  OAI33XLTS U3801 ( .A0(n4833), .A1(n960), .A2(n2018), .B0(n2043), .B1(n4539), 
        .B2(n922), .Y(n2042) );
  NOR4XLTS U3802 ( .A(n2044), .B(n2045), .C(n2046), .D(n2047), .Y(n2043) );
  INVX2TS U3803 ( .A(writeIn_NORTH), .Y(n970) );
  OAI32X1TS U3804 ( .A0(n4835), .A1(n960), .A2(n2018), .B0(n2019), .B1(n2020), 
        .Y(n2450) );
  NOR4BX1TS U3805 ( .AN(n2028), .B(n2029), .C(n2030), .D(n2031), .Y(n2019) );
  OAI31X1TS U3806 ( .A0(n2021), .A1(n469), .A2(n2022), .B0(n4542), .Y(n2020)
         );
  OAI22X1TS U3807 ( .A0(n2035), .A1(n710), .B0(n2036), .B1(n650), .Y(n2029) );
  OAI211X1TS U3808 ( .A0(n3976), .A1(n1167), .B0(n2102), .C0(n2103), .Y(n2441)
         );
  AOI22X1TS U3809 ( .A0(n550), .A1(n2104), .B0(n3093), .B1(
        destinationAddressOut[13]), .Y(n2102) );
  AOI222XLTS U3810 ( .A0(n3055), .A1(n4240), .B0(n2109), .B1(
        destinationAddressIn_NORTH[13]), .C0(n3065), .C1(n4017), .Y(n2103) );
  NAND4X1TS U3811 ( .A(n2105), .B(n2106), .C(n2107), .D(n2108), .Y(n2104) );
  OAI211X1TS U3812 ( .A0(n3973), .A1(n1167), .B0(n2095), .C0(n2096), .Y(n2442)
         );
  AOI22X1TS U3813 ( .A0(n551), .A1(n2097), .B0(n3093), .B1(
        destinationAddressOut[12]), .Y(n2095) );
  AOI222XLTS U3814 ( .A0(n3055), .A1(n4237), .B0(n2109), .B1(
        destinationAddressIn_NORTH[12]), .C0(n3065), .C1(n4014), .Y(n2096) );
  NAND4X1TS U3815 ( .A(n2098), .B(n2099), .C(n2100), .D(n2101), .Y(n2097) );
  OAI211X1TS U3816 ( .A0(n3970), .A1(n1167), .B0(n2088), .C0(n2089), .Y(n2443)
         );
  AOI22X1TS U3817 ( .A0(n552), .A1(n2090), .B0(n3093), .B1(
        destinationAddressOut[11]), .Y(n2088) );
  AOI222XLTS U3818 ( .A0(n3055), .A1(n4234), .B0(n2109), .B1(
        destinationAddressIn_NORTH[11]), .C0(n3065), .C1(n4011), .Y(n2089) );
  NAND4X1TS U3819 ( .A(n2091), .B(n2092), .C(n2093), .D(n2094), .Y(n2090) );
  OAI211X1TS U3820 ( .A0(n3967), .A1(n1198), .B0(n2081), .C0(n2082), .Y(n2444)
         );
  AOI22X1TS U3821 ( .A0(n551), .A1(n2083), .B0(n3093), .B1(
        destinationAddressOut[10]), .Y(n2081) );
  AOI222XLTS U3822 ( .A0(n3055), .A1(n4231), .B0(n2109), .B1(
        destinationAddressIn_NORTH[10]), .C0(n3064), .C1(n4008), .Y(n2082) );
  NAND4X1TS U3823 ( .A(n2084), .B(n2085), .C(n2086), .D(n2087), .Y(n2083) );
  OAI211X1TS U3824 ( .A0(n3964), .A1(n1198), .B0(n2074), .C0(n2075), .Y(n2445)
         );
  AOI22X1TS U3825 ( .A0(n552), .A1(n2076), .B0(n3094), .B1(
        destinationAddressOut[9]), .Y(n2074) );
  AOI222XLTS U3826 ( .A0(n3056), .A1(n4228), .B0(n1939), .B1(
        destinationAddressIn_NORTH[9]), .C0(n3065), .C1(n4005), .Y(n2075) );
  NAND4X1TS U3827 ( .A(n2077), .B(n2078), .C(n2079), .D(n2080), .Y(n2076) );
  OAI211X1TS U3828 ( .A0(n3961), .A1(n1198), .B0(n2067), .C0(n2068), .Y(n2446)
         );
  AOI22X1TS U3829 ( .A0(n551), .A1(n2069), .B0(n3094), .B1(
        destinationAddressOut[8]), .Y(n2067) );
  AOI222XLTS U3830 ( .A0(n3056), .A1(n4225), .B0(n1939), .B1(
        destinationAddressIn_NORTH[8]), .C0(n3064), .C1(n4002), .Y(n2068) );
  NAND4X1TS U3831 ( .A(n2070), .B(n2071), .C(n2072), .D(n2073), .Y(n2069) );
  OAI211X1TS U3832 ( .A0(n3958), .A1(n1215), .B0(n2060), .C0(n2061), .Y(n2447)
         );
  AOI22X1TS U3833 ( .A0(n552), .A1(n2062), .B0(n3094), .B1(
        destinationAddressOut[7]), .Y(n2060) );
  AOI222XLTS U3834 ( .A0(n3056), .A1(n4222), .B0(n1939), .B1(
        destinationAddressIn_NORTH[7]), .C0(n3064), .C1(n3999), .Y(n2061) );
  NAND4X1TS U3835 ( .A(n2063), .B(n2064), .C(n2065), .D(n2066), .Y(n2062) );
  OAI211X1TS U3836 ( .A0(n3955), .A1(n1215), .B0(n2052), .C0(n2053), .Y(n2448)
         );
  AOI22X1TS U3837 ( .A0(n551), .A1(n2055), .B0(n3094), .B1(
        destinationAddressOut[6]), .Y(n2052) );
  AOI222XLTS U3838 ( .A0(n3056), .A1(n4219), .B0(n1939), .B1(
        destinationAddressIn_NORTH[6]), .C0(n3064), .C1(n3996), .Y(n2053) );
  NAND4X1TS U3839 ( .A(n2056), .B(n2057), .C(n2058), .D(n2059), .Y(n2055) );
  INVX2TS U3840 ( .A(readIn_SOUTH), .Y(n972) );
  INVX2TS U3841 ( .A(readIn_NORTH), .Y(n969) );
  OAI21X1TS U3842 ( .A0(n114), .A1(n1097), .B0(n3767), .Y(n2884) );
  INVX2TS U3843 ( .A(destinationAddressIn_NORTH[6]), .Y(n968) );
  INVX2TS U3844 ( .A(destinationAddressIn_NORTH[7]), .Y(n967) );
  INVX2TS U3845 ( .A(destinationAddressIn_NORTH[8]), .Y(n966) );
  OAI21X1TS U3846 ( .A0(n6253), .A1(n1095), .B0(n4542), .Y(n1097) );
  NOR2X1TS U3847 ( .A(n1099), .B(n1097), .Y(n2883) );
  AOI21X1TS U3848 ( .A0(n552), .A1(n137), .B0(n100), .Y(n1099) );
  OAI22X1TS U3849 ( .A0(n45), .A1(n153), .B0(n138), .B1(n136), .Y(n2889) );
  CLKBUFX2TS U3850 ( .A(n5323), .Y(n926) );
  XOR2X1TS U3851 ( .A(n5323), .B(n5), .Y(n2908) );
  NAND2X1TS U3852 ( .A(n100), .B(n136), .Y(n1095) );
  NAND2BX1TS U3853 ( .AN(n1095), .B(n913), .Y(n912) );
  INVX2TS U3854 ( .A(n912), .Y(n2037) );
  AOI22X1TS U3855 ( .A0(n457), .A1(n3138), .B0(n473), .B1(n3184), .Y(n2105) );
  AOI22X1TS U3856 ( .A0(n457), .A1(n3139), .B0(n473), .B1(n3183), .Y(n2098) );
  AOI22X1TS U3857 ( .A0(n457), .A1(n3140), .B0(n473), .B1(n3182), .Y(n2091) );
  AOI22X1TS U3858 ( .A0(n457), .A1(n3141), .B0(n473), .B1(n3181), .Y(n2084) );
  AOI22X1TS U3859 ( .A0(n458), .A1(n3142), .B0(n474), .B1(n3180), .Y(n2077) );
  AOI22X1TS U3860 ( .A0(n458), .A1(n3143), .B0(n474), .B1(n3179), .Y(n2070) );
  AOI22X1TS U3861 ( .A0(n458), .A1(n3144), .B0(n474), .B1(n3178), .Y(n2063) );
  AOI22X1TS U3862 ( .A0(n458), .A1(n3145), .B0(n474), .B1(n3177), .Y(n2056) );
  AOI22X1TS U3863 ( .A0(n145), .A1(n3129), .B0(n156), .B1(n3191), .Y(n2108) );
  AOI22X1TS U3864 ( .A0(n146), .A1(n3130), .B0(n711), .B1(n3190), .Y(n2101) );
  AOI22X1TS U3865 ( .A0(n145), .A1(n3131), .B0(n157), .B1(n3189), .Y(n2094) );
  AOI22X1TS U3866 ( .A0(n146), .A1(n3132), .B0(n156), .B1(n3188), .Y(n2087) );
  AOI22X1TS U3867 ( .A0(n145), .A1(n3133), .B0(n711), .B1(n3187), .Y(n2080) );
  AOI22X1TS U3868 ( .A0(n146), .A1(n3134), .B0(n157), .B1(n3186), .Y(n2073) );
  AOI22X1TS U3869 ( .A0(n145), .A1(n3136), .B0(n156), .B1(n3135), .Y(n2066) );
  AOI22X1TS U3870 ( .A0(n146), .A1(n3137), .B0(n711), .B1(n3185), .Y(n2059) );
  AOI22X1TS U3871 ( .A0(n475), .A1(n3162), .B0(n3161), .B1(n2048), .Y(n2106)
         );
  AOI22X1TS U3872 ( .A0(n475), .A1(n3164), .B0(n3163), .B1(n924), .Y(n2099) );
  AOI22X1TS U3873 ( .A0(n475), .A1(n3166), .B0(n3165), .B1(n462), .Y(n2092) );
  AOI22X1TS U3874 ( .A0(n475), .A1(n3168), .B0(n3167), .B1(n462), .Y(n2085) );
  AOI22X1TS U3875 ( .A0(n476), .A1(n3170), .B0(n3169), .B1(n924), .Y(n2078) );
  AOI22X1TS U3876 ( .A0(n476), .A1(n3172), .B0(n3171), .B1(n462), .Y(n2071) );
  AOI22X1TS U3877 ( .A0(n476), .A1(n3174), .B0(n3173), .B1(n2048), .Y(n2064)
         );
  AOI22X1TS U3878 ( .A0(n476), .A1(n3176), .B0(n3175), .B1(n924), .Y(n2057) );
  AOI22X1TS U3879 ( .A0(n168), .A1(n3147), .B0(n142), .B1(n3146), .Y(n2107) );
  AOI22X1TS U3880 ( .A0(n169), .A1(n3149), .B0(n141), .B1(n3148), .Y(n2100) );
  AOI22X1TS U3881 ( .A0(n2037), .A1(n3151), .B0(n142), .B1(n3150), .Y(n2093)
         );
  AOI22X1TS U3882 ( .A0(n168), .A1(n3154), .B0(n141), .B1(n3153), .Y(n2079) );
  AOI22X1TS U3883 ( .A0(n2037), .A1(n3156), .B0(n142), .B1(n3155), .Y(n2072)
         );
  AOI22X1TS U3884 ( .A0(n168), .A1(n3158), .B0(n141), .B1(n3157), .Y(n2065) );
  AOI22X1TS U3885 ( .A0(n169), .A1(n3160), .B0(n142), .B1(n3159), .Y(n2058) );
  OA22X1TS U3886 ( .A0(n2032), .A1(n563), .B0(n167), .B1(n4796), .Y(n2086) );
  AOI221X1TS U3887 ( .A0(n157), .A1(\readOutbuffer[2] ), .B0(n169), .B1(
        readOutbuffer_7), .C0(n6253), .Y(n2028) );
  AOI32XLTS U3888 ( .A0(n453), .A1(n1814), .A2(n1815), .B0(n3259), .B1(n656), 
        .Y(n2563) );
  AOI32XLTS U3889 ( .A0(n104), .A1(n1808), .A2(n1809), .B0(n3340), .B1(n655), 
        .Y(n2564) );
  AOI32XLTS U3890 ( .A0(n447), .A1(n1810), .A2(n4195), .B0(n1811), .B1(n1782), 
        .Y(n1809) );
  AND3X2TS U3891 ( .A(n447), .B(n1810), .C(n1807), .Y(n1204) );
  NOR2XLTS U3892 ( .A(n143), .B(n957), .Y(n2016) );
  NOR2XLTS U3893 ( .A(n1869), .B(n1775), .Y(n1123) );
  OAI33XLTS U3894 ( .A0(n4197), .A1(n452), .A2(n443), .B0(n438), .B1(n927), 
        .B2(n1790), .Y(n1787) );
  NAND3BX1TS U3895 ( .AN(n1803), .B(n103), .C(n1805), .Y(n1182) );
  AOI32XLTS U3896 ( .A0(n103), .A1(n1800), .A2(n1801), .B0(n3820), .B1(n709), 
        .Y(n2565) );
  OAI221XLTS U3897 ( .A0(n164), .A1(n122), .B0(n163), .B1(n763), .C0(n1953), 
        .Y(n2486) );
  OAI221XLTS U3898 ( .A0(n165), .A1(n124), .B0(n162), .B1(n765), .C0(n1954), 
        .Y(n2485) );
  OAI221XLTS U3899 ( .A0(n164), .A1(n131), .B0(n163), .B1(n764), .C0(n1955), 
        .Y(n2484) );
  OAI221XLTS U3900 ( .A0(n165), .A1(n129), .B0(n1757), .B1(n921), .C0(n1956), 
        .Y(n2483) );
  OAI221XLTS U3901 ( .A0(n164), .A1(n134), .B0(n163), .B1(n920), .C0(n1957), 
        .Y(n2482) );
  OAI221XLTS U3902 ( .A0(n165), .A1(n127), .B0(n1757), .B1(n919), .C0(n1958), 
        .Y(n2481) );
  OAI221XLTS U3903 ( .A0(n164), .A1(n125), .B0(n163), .B1(n918), .C0(n1959), 
        .Y(n2480) );
  OAI221XLTS U3904 ( .A0(n165), .A1(n133), .B0(n1757), .B1(n916), .C0(n1960), 
        .Y(n2479) );
  OAI221XLTS U3905 ( .A0(n1756), .A1(n149), .B0(n162), .B1(n910), .C0(n1758), 
        .Y(n2573) );
  NOR2BX1TS U3906 ( .AN(n1799), .B(n1805), .Y(n1187) );
  AOI21XLTS U3907 ( .A0(n4190), .A1(n759), .B0(n440), .Y(n1763) );
  AOI32XLTS U3908 ( .A0(n1765), .A1(n1766), .A2(n1767), .B0(n4196), .B1(n745), 
        .Y(n1764) );
  AOI32XLTS U3909 ( .A0(n439), .A1(n1792), .A2(n1793), .B0(n3849), .B1(n649), 
        .Y(n2566) );
  OAI221XLTS U3910 ( .A0(n451), .A1(n122), .B0(n549), .B1(n570), .C0(n1929), 
        .Y(n2500) );
  OAI221XLTS U3911 ( .A0(n449), .A1(n967), .B0(n548), .B1(n556), .C0(n1930), 
        .Y(n2499) );
  OAI221XLTS U3912 ( .A0(n450), .A1(n131), .B0(n549), .B1(n567), .C0(n1931), 
        .Y(n2498) );
  OAI221XLTS U3913 ( .A0(n451), .A1(n130), .B0(n548), .B1(n568), .C0(n1932), 
        .Y(n2497) );
  OAI221XLTS U3914 ( .A0(n451), .A1(n134), .B0(n549), .B1(n557), .C0(n1933), 
        .Y(n2496) );
  OAI221XLTS U3915 ( .A0(n450), .A1(n128), .B0(n548), .B1(n571), .C0(n1934), 
        .Y(n2495) );
  OAI221XLTS U3916 ( .A0(n450), .A1(n125), .B0(n549), .B1(n569), .C0(n1935), 
        .Y(n2494) );
  OAI221XLTS U3917 ( .A0(n450), .A1(n132), .B0(n548), .B1(n558), .C0(n1936), 
        .Y(n2493) );
  OAI221XLTS U3918 ( .A0(n451), .A1(n149), .B0(n547), .B1(n706), .C0(n1755), 
        .Y(n2574) );
  AOI32XLTS U3919 ( .A0(n1794), .A1(n1795), .A2(n4195), .B0(n1796), .B1(n1797), 
        .Y(n1793) );
  AOI21XLTS U3920 ( .A0(readIn_SOUTH), .A1(n1774), .B0(n1775), .Y(n1770) );
  OAI211XLTS U3921 ( .A0(n721), .A1(n3937), .B0(n1848), .C0(n1849), .Y(n2548)
         );
  OAI211XLTS U3922 ( .A0(n723), .A1(n3940), .B0(n1850), .C0(n1851), .Y(n2547)
         );
  OAI211XLTS U3923 ( .A0(n725), .A1(n3943), .B0(n1852), .C0(n1853), .Y(n2546)
         );
  OAI211XLTS U3924 ( .A0(n721), .A1(n3946), .B0(n1854), .C0(n1855), .Y(n2545)
         );
  OAI211XLTS U3925 ( .A0(n723), .A1(n3949), .B0(n1856), .C0(n1857), .Y(n2544)
         );
  OAI211XLTS U3926 ( .A0(n725), .A1(n3952), .B0(n1858), .C0(n1859), .Y(n2543)
         );
  OAI211XLTS U3927 ( .A0(n4171), .A1(n721), .B0(n1119), .C0(n1120), .Y(n2876)
         );
  OAI211XLTS U3928 ( .A0(n4174), .A1(n721), .B0(n1124), .C0(n1125), .Y(n2875)
         );
  OAI211XLTS U3929 ( .A0(n4177), .A1(n723), .B0(n1126), .C0(n1127), .Y(n2874)
         );
  OAI211XLTS U3930 ( .A0(n4180), .A1(n723), .B0(n1128), .C0(n1129), .Y(n2873)
         );
  OAI211XLTS U3931 ( .A0(n4183), .A1(n725), .B0(n1130), .C0(n1131), .Y(n2872)
         );
  OAI211XLTS U3932 ( .A0(n4186), .A1(n725), .B0(n1132), .C0(n1133), .Y(n2871)
         );
  NOR2BX1TS U3933 ( .AN(n1774), .B(n1775), .Y(n1121) );
  AOI21XLTS U3934 ( .A0(readIn_NORTH), .A1(n1786), .B0(n1787), .Y(n1785) );
  OA22XLTS U3935 ( .A0(n958), .A1(n2901), .B0(n2902), .B1(n2014), .Y(n2449) );
endmodule


module outputPortArbiter_2 ( clk, reset, selectBit_NORTH, 
        destinationAddressIn_NORTH, requesterAddressIn_NORTH, readIn_NORTH, 
        writeIn_NORTH, dataIn_NORTH, selectBit_SOUTH, 
        destinationAddressIn_SOUTH, requesterAddressIn_SOUTH, readIn_SOUTH, 
        writeIn_SOUTH, dataIn_SOUTH, selectBit_EAST, destinationAddressIn_EAST, 
        requesterAddressIn_EAST, readIn_EAST, writeIn_EAST, dataIn_EAST, 
        selectBit_WEST, destinationAddressIn_WEST, requesterAddressIn_WEST, 
        readIn_WEST, writeIn_WEST, dataIn_WEST, readReady, 
        readRequesterAddress, cacheDataOut, destinationAddressOut, 
        requesterAddressOut, readOut, writeOut, dataOut );
  input [13:0] destinationAddressIn_NORTH;
  input [5:0] requesterAddressIn_NORTH;
  input [31:0] dataIn_NORTH;
  input [13:0] destinationAddressIn_SOUTH;
  input [5:0] requesterAddressIn_SOUTH;
  input [31:0] dataIn_SOUTH;
  input [13:0] destinationAddressIn_EAST;
  input [5:0] requesterAddressIn_EAST;
  input [31:0] dataIn_EAST;
  input [13:0] destinationAddressIn_WEST;
  input [5:0] requesterAddressIn_WEST;
  input [31:0] dataIn_WEST;
  input [5:0] readRequesterAddress;
  input [31:0] cacheDataOut;
  output [13:0] destinationAddressOut;
  output [5:0] requesterAddressOut;
  output [31:0] dataOut;
  input clk, reset, selectBit_NORTH, readIn_NORTH, writeIn_NORTH,
         selectBit_SOUTH, readIn_SOUTH, writeIn_SOUTH, selectBit_EAST,
         readIn_EAST, writeIn_EAST, selectBit_WEST, readIn_WEST, writeIn_WEST,
         readReady;
  output readOut, writeOut;
  wire   n2486, n2484, n2482, n2480, n2457, n2455, n2453, n2485, n2483, n2481,
         n2458, n2454, n2451, n2479, n2456, n2452, n2499, n2496, n2493, n2528,
         n2527, n2526, n2525, n2524, n2523, n2522, n2521, n2498, n2497, n2494,
         n2500, n2495, n2511, n2507, n2538, n2536, n2514, n2513, n2512, n2510,
         n2509, n2508, n2703, n2692, n2691, n2689, n2706, n2705, n2700, n2698,
         n2696, n2695, n2694, n2690, n2687, n2686, n2685, n2684, n2677, n2675,
         n2704, n2702, n2701, n2699, n2697, n2693, n2688, n2683, n2682, n2681,
         n2680, n2679, n2678, n2676, n2520, n2519, n2518, n2517, n2515, n2850,
         \requesterAddressbuffer[2][2] , n2849, \requesterAddressbuffer[2][3] ,
         n2847, \requesterAddressbuffer[2][5] , n2840,
         \requesterAddressbuffer[0][0] , n2839, \requesterAddressbuffer[0][1] ,
         n2838, \requesterAddressbuffer[0][2] , n2836,
         \requesterAddressbuffer[0][4] , n2852, \requesterAddressbuffer[2][0] ,
         n2851, \requesterAddressbuffer[2][1] , n2848,
         \requesterAddressbuffer[2][4] , n2837, \requesterAddressbuffer[0][3] ,
         n2835, \requesterAddressbuffer[0][5] , n2566, \readOutbuffer[2] ,
         readOutbuffer_7, n2569, n2568, n2564, n2576, n2573, n2770, n95, n2768,
         n94, n2764, n93, n2754, n92, n2748, n91, n2746, n90, n2739, n89,
         n2834, n57, n2833, n56, n2832, n55, n2829, n54, n2825, n53, n2814,
         n52, n2811, n51, n2807, n50, n2806, n49, n2769, n88, n2760, n87,
         n2743, n86, n2492, n85, n2491, n84, n2489, n83, n2488, n82, n2487,
         n81, n2464, n48, n2460, n4724, n2767, n80, n2766, n79, n2765, n78,
         n2763, n77, n2762, n76, n2761, n75, n2759, n74, n2758, n73, n2757,
         n72, n2756, n71, n2755, n70, n2753, n69, n2752, n68, n2751, n67,
         n2750, n66, n2749, n65, n2747, n64, n2745, n63, n2744, n62, n2742,
         n61, n2741, n60, n2740, n59, n2490, n58, n2831, n4674, n2830, n4663,
         n2828, n4647, n2827, n4638, n2826, n4633, n2824, n4613, n2823, n4600,
         n2822, n4595, n2821, n4588, n2820, n4575, n2819, n4568, n2818, n4557,
         n2817, n4548, n2816, n4539, n2815, n4530, n2813, n4516, n2812, n4501,
         n2810, n4485, n2809, n4476, n2808, n4469, n2805, n4444, n2804, n4433,
         n2803, n4420, n2463, n4748, n2462, n4743, n2461, n4732, n2459, n4712,
         n2571, n2574, n2575, n2570, n2565, n2567, n2889, N4718, n96, n2887,
         n5323, n4829, n2434, n4833, n2431, n4834, n2450, n4831, n2440, n4756,
         n2439, n4747, n2438, n4738, n2437, n4729, n2436, n4720, n2435, n4711,
         n2433, n4710, n2432, n4709, n2430, n4708, n2429, n4707, n2428, n4698,
         n2427, n4689, n2426, n4680, n2425, n4671, n2424, n4662, n2423, n4653,
         n2422, n4644, n2421, n4635, n2420, n4626, n2419, n4617, n2418, n4608,
         n2417, n4599, n2416, n4590, n2415, n4581, n2414, n4572, n2413, n4563,
         n2412, n4554, n2411, n4545, n2410, n4536, n2409, n4527, n2408, n4518,
         n2407, n4509, n2406, n4500, n2405, n4491, n2404, n4482, n2403, n4473,
         n2402, n4464, n2401, n4455, n2400, n4446, n2399, n4437, n2398, n4428,
         n2397, n4419, n2448, n2447, n2446, n2445, n2444, n2443, n2442, n2441,
         n2549, n2472, n2471, n2470, n2469, n2468, n2467, n2466, n2465, n2530,
         n2674, n2672, n2671, n2670, n2669, n2668, n2667, n2666, n2665, n2664,
         n2662, n2661, n2660, n2657, n2656, n2655, n2654, n2653, n2652, n2651,
         n2650, n2649, n2648, n2647, n2646, n2645, n2644, n2534, n2533, n2532,
         n2531, n2529, n2673, n2663, n2659, n2658, n2643, n2558, n2516, n2638,
         n2624, n2802, n2609, n2608, n2607, n2606, n2605, n2604, n2603, n2602,
         n2601, n2600, n2599, n2598, n2594, n2593, n2592, n2591, n2590, n2589,
         n2588, n2587, n2586, n2585, n2584, n2583, n2582, n2581, n2580, n2579,
         n2561, n2560, n2559, n2557, n2642, n2640, n2639, n2637, n2633, n2628,
         n2614, n2612, n2801, n2799, n2798, n2796, n2795, n2793, n2791, n2790,
         n2789, n2788, n2787, n2786, n2785, n2784, n2781, n2779, n2778, n2777,
         n2776, n2774, n2773, n2772, n2771, n2478, n2477, n2476, n2475, n2473,
         n2562, n2641, n2636, n2632, n2548, n2547, n2546, n2545, n2543, n2800,
         n2797, n2794, n2792, n2783, n2782, n2780, n2775, n2544, n2552, n480,
         n2474, n2731, n6313, n2736, n6300, n2734, n6299, n2733, n6298, n2725,
         n6297, n2723, n6296, n2720, n6295, n2718, n6294, n2715, n6293, n2713,
         n6292, n2504, n6291, n2738, n6276, n2737, n6275, n2735, n6274, n2732,
         n6273, n2730, n6272, n2729, n6271, n2728, n6270, n2727, n6269, n2726,
         n6268, n2724, n6267, n2722, n6266, n2721, n6265, n2719, n6264, n2717,
         n6263, n2716, n6262, n2714, n6261, n2712, n6260, n2711, n6259, n2710,
         n6258, n2709, n6257, n2708, n6256, n2707, n6255, n2506, n6254, n2505,
         n6253, n2503, n6252, n2502, n6251, n2501, n6250, n2858,
         \requesterAddressbuffer[3][0] , n2857, \requesterAddressbuffer[3][1] ,
         n2856, \requesterAddressbuffer[3][2] , n2855,
         \requesterAddressbuffer[3][3] , n2853, \requesterAddressbuffer[3][5] ,
         n2854, \requesterAddressbuffer[3][4] , n2875,
         \requesterAddressbuffer[6][1] , n2874, \requesterAddressbuffer[6][2] ,
         n2873, \requesterAddressbuffer[6][3] , n2872,
         \requesterAddressbuffer[6][4] , n2871, \requesterAddressbuffer[6][5] ,
         n2876, \requesterAddressbuffer[6][0] , n2578, n2882, n2881, n2879,
         n2870, n2869, n2868, n2867, n2866, n2865, n2880, n2878, n2877, n2563,
         n2860, n2859, n2864, n2863, n2862, n2861, n2846, n2845, n2844, n2843,
         n2842, n2841, n2541, n2540, n2537, n2535, n2556, n2555, n2554, n2551,
         n2550, n2553, n2542, n2539, n2577, n2572, n2883, n5, n2884, n385,
         n2595, n2596, n2597, n2610, n2611, n2613, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2625, n2626, n2627, n2629, n2630,
         n2631, n2634, n2635, n2885, n6248, n2888, n9, n2886, n6, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n660, n662, n664,
         n665, n667, n668, n669, n670, n671, n675, n678, n679, n681, n682,
         n684, n685, n686, n688, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n939, n942, n943, n944,
         n945, n946, n947, n948, n951, n953, n954, n955, n964, n965, n968,
         n1023, n1078, n1080, n1081, n1082, n1083, n1084, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2449, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
         n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
         n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
         n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
         n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n2999, n3000, n3001, n3002, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n1, n2, n3, n4, n7,
         n8, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n659, n661, n663, n666, n672, n673, n674, n676,
         n677, n680, n683, n687, n689, n701, n913, n914, n938, n940, n941,
         n949, n950, n952, n956, n957, n958, n959, n960, n961, n962, n963,
         n966, n967, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1079, n1085, n1102,
         n1129, n1146, n1162, n1193, n1210, n1611, n1749, n1771, n1807, n1934,
         n1980, n2103, n2377, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n3003, n3004, n3005, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4429, n4430, n4431,
         n4432, n4434, n4435, n4436, n4438, n4439, n4440, n4441, n4442, n4443,
         n4445, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4465, n4466, n4467,
         n4468, n4470, n4471, n4472, n4474, n4475, n4477, n4478, n4479, n4480,
         n4481, n4483, n4484, n4486, n4487, n4488, n4489, n4490, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4510, n4511, n4512, n4513, n4514, n4515, n4517,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4528, n4529,
         n4531, n4532, n4533, n4534, n4535, n4537, n4538, n4540, n4541, n4542,
         n4543, n4544, n4546, n4547, n4549, n4550, n4551, n4552, n4553, n4555,
         n4556, n4558, n4559, n4560, n4561, n4562, n4564, n4565, n4566, n4567,
         n4569, n4570, n4571, n4573, n4574, n4576, n4577, n4578, n4579, n4580,
         n4582, n4583, n4584, n4585, n4586, n4587, n4589, n4591, n4592, n4593,
         n4594, n4596, n4597, n4598, n4601, n4602, n4603, n4604, n4605, n4606;

  DFFNSRX2TS \dataoutbuffer_reg[2][0]  ( .D(n2770), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n95) );
  DFFNSRX2TS \dataoutbuffer_reg[2][2]  ( .D(n2768), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n94) );
  DFFNSRX2TS \dataoutbuffer_reg[2][6]  ( .D(n2764), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n93) );
  DFFNSRX2TS \dataoutbuffer_reg[2][16]  ( .D(n2754), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n92) );
  DFFNSRX2TS \dataoutbuffer_reg[2][1]  ( .D(n2769), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n88) );
  DFFNSRX2TS \dataoutbuffer_reg[2][10]  ( .D(n2760), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n87) );
  DFFNSRX2TS \destinationAddressbuffer_reg[2][3]  ( .D(n2489), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n83) );
  DFFNSRX2TS \destinationAddressbuffer_reg[2][4]  ( .D(n2488), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n82) );
  DFFNSRX2TS \dataoutbuffer_reg[2][3]  ( .D(n2767), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n80) );
  DFFNSRX2TS \dataoutbuffer_reg[2][4]  ( .D(n2766), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n79) );
  DFFNSRX2TS \dataoutbuffer_reg[2][5]  ( .D(n2765), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n78) );
  DFFNSRX2TS \dataoutbuffer_reg[2][7]  ( .D(n2763), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n77) );
  DFFNSRX2TS \dataoutbuffer_reg[2][8]  ( .D(n2762), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n76) );
  DFFNSRX2TS \dataoutbuffer_reg[2][9]  ( .D(n2761), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n75) );
  DFFNSRX2TS \dataoutbuffer_reg[2][11]  ( .D(n2759), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n74) );
  DFFNSRX2TS \dataoutbuffer_reg[2][12]  ( .D(n2758), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n73) );
  DFFNSRX2TS \dataoutbuffer_reg[2][13]  ( .D(n2757), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n72) );
  DFFNSRX2TS \dataoutbuffer_reg[2][14]  ( .D(n2756), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n71) );
  DFFNSRX2TS \dataoutbuffer_reg[2][15]  ( .D(n2755), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n70) );
  DFFNSRX2TS \dataoutbuffer_reg[2][17]  ( .D(n2753), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n69) );
  DFFNSRX2TS \dataoutbuffer_reg[2][18]  ( .D(n2752), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n68) );
  DFFNSRX2TS \dataoutbuffer_reg[2][19]  ( .D(n2751), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n67) );
  DFFNSRX2TS \destinationAddressbuffer_reg[2][2]  ( .D(n2490), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n58) );
  DFFNSRX2TS empty_reg_reg ( .D(n2885), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        n6248), .QN(n486) );
  DFFNSRX2TS \read_reg_reg[1]  ( .D(n2883), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n5), .QN(n475) );
  DFFNSRX2TS \read_reg_reg[2]  ( .D(n2884), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n3), .QN(n385) );
  DFFNSRX2TS \write_reg_reg[1]  ( .D(n2887), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n467), .QN(n5323) );
  DFFNSRX2TS \write_reg_reg[2]  ( .D(n2886), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n6), .QN(n476) );
  DFFNSRX2TS writeOut_reg ( .D(n602), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        writeOut), .QN(n4829) );
  DFFNSRX2TS \requesterAddressOut_reg[0]  ( .D(n2434), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[0]), .QN(n4833) );
  DFFNSRX2TS \requesterAddressOut_reg[3]  ( .D(n2431), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[3]), .QN(n4834) );
  DFFNSRX2TS readOut_reg ( .D(n2450), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        readOut), .QN(n4831) );
  DFFNSRX2TS \destinationAddressOut_reg[0]  ( .D(n2440), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[0]), .QN(n4756) );
  DFFNSRX2TS \destinationAddressOut_reg[1]  ( .D(n2439), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[1]), .QN(n4747) );
  DFFNSRX2TS \destinationAddressOut_reg[2]  ( .D(n2438), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[2]), .QN(n4738) );
  DFFNSRX2TS \destinationAddressOut_reg[3]  ( .D(n2437), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[3]), .QN(n4729) );
  DFFNSRX2TS \destinationAddressOut_reg[4]  ( .D(n2436), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[4]), .QN(n4720) );
  DFFNSRX2TS \destinationAddressOut_reg[5]  ( .D(n2435), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[5]), .QN(n4711) );
  DFFNSRX2TS \requesterAddressOut_reg[1]  ( .D(n2433), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[1]), .QN(n4710) );
  DFFNSRX2TS \requesterAddressOut_reg[2]  ( .D(n2432), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[2]), .QN(n4709) );
  DFFNSRX2TS \requesterAddressOut_reg[4]  ( .D(n2430), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[4]), .QN(n4708) );
  DFFNSRX2TS \requesterAddressOut_reg[5]  ( .D(n2429), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[5]), .QN(n4707) );
  DFFNSRX2TS \dataOut_reg[0]  ( .D(n2428), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[0]), .QN(n4698) );
  DFFNSRX2TS \dataOut_reg[1]  ( .D(n2427), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[1]), .QN(n4689) );
  DFFNSRX2TS \dataOut_reg[2]  ( .D(n2426), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[2]), .QN(n4680) );
  DFFNSRX2TS \dataOut_reg[3]  ( .D(n2425), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[3]), .QN(n4671) );
  DFFNSRX2TS \dataOut_reg[4]  ( .D(n2424), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[4]), .QN(n4662) );
  DFFNSRX2TS \dataOut_reg[5]  ( .D(n2423), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[5]), .QN(n4653) );
  DFFNSRX2TS \dataOut_reg[6]  ( .D(n2422), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[6]), .QN(n4644) );
  DFFNSRX2TS \dataOut_reg[7]  ( .D(n2421), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[7]), .QN(n4635) );
  DFFNSRX2TS \dataOut_reg[8]  ( .D(n2420), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[8]), .QN(n4626) );
  DFFNSRX2TS \dataOut_reg[9]  ( .D(n2419), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[9]), .QN(n4617) );
  DFFNSRX2TS \dataOut_reg[10]  ( .D(n2418), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[10]), .QN(n4608) );
  DFFNSRX2TS \dataOut_reg[11]  ( .D(n2417), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[11]), .QN(n4599) );
  DFFNSRX2TS \dataOut_reg[12]  ( .D(n2416), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[12]), .QN(n4590) );
  DFFNSRX2TS \dataOut_reg[13]  ( .D(n2415), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[13]), .QN(n4581) );
  DFFNSRX2TS \dataOut_reg[14]  ( .D(n2414), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[14]), .QN(n4572) );
  DFFNSRX2TS \dataOut_reg[15]  ( .D(n2413), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[15]), .QN(n4563) );
  DFFNSRX2TS \dataOut_reg[16]  ( .D(n2412), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[16]), .QN(n4554) );
  DFFNSRX2TS \dataOut_reg[17]  ( .D(n2411), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[17]), .QN(n4545) );
  DFFNSRX2TS \dataOut_reg[18]  ( .D(n2410), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[18]), .QN(n4536) );
  DFFNSRX2TS \dataOut_reg[19]  ( .D(n2409), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[19]), .QN(n4527) );
  DFFNSRX2TS \dataOut_reg[20]  ( .D(n2408), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[20]), .QN(n4518) );
  DFFNSRX2TS \dataOut_reg[21]  ( .D(n2407), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[21]), .QN(n4509) );
  DFFNSRX2TS \dataOut_reg[22]  ( .D(n2406), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[22]), .QN(n4500) );
  DFFNSRX2TS \dataOut_reg[23]  ( .D(n2405), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[23]), .QN(n4491) );
  DFFNSRX2TS \dataOut_reg[24]  ( .D(n2404), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[24]), .QN(n4482) );
  DFFNSRX2TS \dataOut_reg[25]  ( .D(n2403), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[25]), .QN(n4473) );
  DFFNSRX2TS \dataOut_reg[26]  ( .D(n2402), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[26]), .QN(n4464) );
  DFFNSRX2TS \dataOut_reg[27]  ( .D(n2401), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[27]), .QN(n4455) );
  DFFNSRX2TS \dataOut_reg[28]  ( .D(n2400), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[28]), .QN(n4446) );
  DFFNSRX2TS \dataOut_reg[29]  ( .D(n2399), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[29]), .QN(n4437) );
  DFFNSRX2TS \dataOut_reg[30]  ( .D(n2398), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[30]), .QN(n4428) );
  DFFNSRX2TS \dataOut_reg[31]  ( .D(n2397), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[31]), .QN(n4419) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][4]  ( .D(n2530), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n711) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][0]  ( .D(n2534), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n739) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][1]  ( .D(n2533), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n740) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][2]  ( .D(n2532), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n741) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][3]  ( .D(n2531), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n742) );
  DFFNSRXLTS \requesterAddressbuffer_reg[5][0]  ( .D(n2870), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n883) );
  DFFNSRXLTS \requesterAddressbuffer_reg[5][1]  ( .D(n2869), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n884) );
  DFFNSRXLTS \requesterAddressbuffer_reg[5][2]  ( .D(n2868), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n885) );
  DFFNSRXLTS \requesterAddressbuffer_reg[5][3]  ( .D(n2867), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n886) );
  DFFNSRXLTS \requesterAddressbuffer_reg[5][4]  ( .D(n2866), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n887) );
  DFFNSRXLTS \requesterAddressbuffer_reg[5][5]  ( .D(n2865), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n888) );
  DFFNSRXLTS \dataoutbuffer_reg[1][0]  ( .D(n2802), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3037), .QN(n752) );
  DFFNSRXLTS \dataoutbuffer_reg[1][1]  ( .D(n2801), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3036), .QN(n793) );
  DFFNSRXLTS \dataoutbuffer_reg[1][3]  ( .D(n2799), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3034), .QN(n794) );
  DFFNSRXLTS \dataoutbuffer_reg[1][4]  ( .D(n2798), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3033), .QN(n795) );
  DFFNSRXLTS \dataoutbuffer_reg[1][6]  ( .D(n2796), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3031), .QN(n796) );
  DFFNSRXLTS \dataoutbuffer_reg[1][7]  ( .D(n2795), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3030), .QN(n797) );
  DFFNSRXLTS \dataoutbuffer_reg[1][9]  ( .D(n2793), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3028), .QN(n798) );
  DFFNSRXLTS \dataoutbuffer_reg[1][11]  ( .D(n2791), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3026), .QN(n799) );
  DFFNSRXLTS \dataoutbuffer_reg[1][12]  ( .D(n2790), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3025), .QN(n800) );
  DFFNSRXLTS \dataoutbuffer_reg[1][13]  ( .D(n2789), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3024), .QN(n801) );
  DFFNSRXLTS \dataoutbuffer_reg[1][14]  ( .D(n2788), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3023), .QN(n802) );
  DFFNSRXLTS \dataoutbuffer_reg[1][15]  ( .D(n2787), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3022), .QN(n803) );
  DFFNSRXLTS \dataoutbuffer_reg[1][16]  ( .D(n2786), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3021), .QN(n804) );
  DFFNSRXLTS \dataoutbuffer_reg[1][17]  ( .D(n2785), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3020), .QN(n805) );
  DFFNSRXLTS \dataoutbuffer_reg[1][18]  ( .D(n2784), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3019), .QN(n806) );
  DFFNSRXLTS \dataoutbuffer_reg[1][21]  ( .D(n2781), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3016), .QN(n807) );
  DFFNSRXLTS \dataoutbuffer_reg[1][23]  ( .D(n2779), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3014), .QN(n808) );
  DFFNSRXLTS \dataoutbuffer_reg[1][24]  ( .D(n2778), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3013), .QN(n809) );
  DFFNSRXLTS \dataoutbuffer_reg[1][25]  ( .D(n2777), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3012), .QN(n810) );
  DFFNSRXLTS \dataoutbuffer_reg[1][26]  ( .D(n2776), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3011), .QN(n811) );
  DFFNSRXLTS \dataoutbuffer_reg[1][28]  ( .D(n2774), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3009), .QN(n812) );
  DFFNSRXLTS \dataoutbuffer_reg[1][29]  ( .D(n2773), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3008), .QN(n813) );
  DFFNSRXLTS \dataoutbuffer_reg[1][30]  ( .D(n2772), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3007), .QN(n814) );
  DFFNSRXLTS \dataoutbuffer_reg[1][31]  ( .D(n2771), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3006), .QN(n815) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][0]  ( .D(n2478), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3043), .QN(n816) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][1]  ( .D(n2477), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3042), .QN(n817) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][2]  ( .D(n2476), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3041), .QN(n818) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][3]  ( .D(n2475), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3040), .QN(n819) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][5]  ( .D(n2473), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3038), .QN(n820) );
  DFFNSRXLTS \dataoutbuffer_reg[1][2]  ( .D(n2800), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3035), .QN(n825) );
  DFFNSRXLTS \dataoutbuffer_reg[1][5]  ( .D(n2797), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3032), .QN(n826) );
  DFFNSRXLTS \dataoutbuffer_reg[1][8]  ( .D(n2794), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3029), .QN(n827) );
  DFFNSRXLTS \dataoutbuffer_reg[1][10]  ( .D(n2792), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3027), .QN(n828) );
  DFFNSRXLTS \dataoutbuffer_reg[1][19]  ( .D(n2783), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3018), .QN(n829) );
  DFFNSRXLTS \dataoutbuffer_reg[1][20]  ( .D(n2782), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3017), .QN(n830) );
  DFFNSRXLTS \dataoutbuffer_reg[1][22]  ( .D(n2780), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3015), .QN(n831) );
  DFFNSRXLTS \dataoutbuffer_reg[1][27]  ( .D(n2775), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3010), .QN(n832) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][0]  ( .D(n2846), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2908), .QN(n893) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][1]  ( .D(n2845), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2906), .QN(n894) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][2]  ( .D(n2844), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2905), .QN(n895) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][3]  ( .D(n2843), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2907), .QN(n896) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][4]  ( .D(n2842), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2904), .QN(n897) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][5]  ( .D(n2841), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2903), .QN(n898) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][4]  ( .D(n2474), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3039), .QN(n834) );
  DFFNSRXLTS \writeOutbuffer_reg[2]  ( .D(n2573), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n604) );
  DFFNSRXLTS \writeOutbuffer_reg[3]  ( .D(n2574), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n644) );
  DFFNSRXLTS \writeOutbuffer_reg[1]  ( .D(n2572), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n912) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][0]  ( .D(n2548), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3002) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][1]  ( .D(n2547), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3000) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][2]  ( .D(n2546), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2998) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][3]  ( .D(n2545), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2996) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][5]  ( .D(n2543), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2992) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][4]  ( .D(n2544), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2994) );
  DFFNSRXLTS \requesterAddressbuffer_reg[6][1]  ( .D(n2875), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][1] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[6][2]  ( .D(n2874), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][2] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[6][3]  ( .D(n2873), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][3] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[6][4]  ( .D(n2872), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][4] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[6][5]  ( .D(n2871), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][5] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[6][0]  ( .D(n2876), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][0] ) );
  DFFNSRXLTS \dataoutbuffer_reg[6][4]  ( .D(n2638), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n2982), .QN(n750) );
  DFFNSRXLTS \dataoutbuffer_reg[6][18]  ( .D(n2624), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2954), .QN(n751) );
  DFFNSRXLTS \dataoutbuffer_reg[6][0]  ( .D(n2642), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n2990), .QN(n785) );
  DFFNSRXLTS \dataoutbuffer_reg[6][2]  ( .D(n2640), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n2986), .QN(n786) );
  DFFNSRXLTS \dataoutbuffer_reg[6][3]  ( .D(n2639), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n2984), .QN(n787) );
  DFFNSRXLTS \dataoutbuffer_reg[6][5]  ( .D(n2637), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n2980), .QN(n788) );
  DFFNSRXLTS \dataoutbuffer_reg[6][9]  ( .D(n2633), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n2972), .QN(n789) );
  DFFNSRXLTS \dataoutbuffer_reg[6][14]  ( .D(n2628), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2962), .QN(n790) );
  DFFNSRXLTS \dataoutbuffer_reg[6][28]  ( .D(n2614), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2934), .QN(n791) );
  DFFNSRXLTS \dataoutbuffer_reg[6][30]  ( .D(n2612), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2930), .QN(n792) );
  DFFNSRXLTS \dataoutbuffer_reg[6][1]  ( .D(n2641), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n2988), .QN(n822) );
  DFFNSRXLTS \dataoutbuffer_reg[6][6]  ( .D(n2636), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n2978), .QN(n823) );
  DFFNSRXLTS \dataoutbuffer_reg[6][10]  ( .D(n2632), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2970), .QN(n824) );
  DFFNSRXLTS \dataoutbuffer_reg[6][31]  ( .D(n2611), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2928), .QN(n919) );
  DFFNSRXLTS \dataoutbuffer_reg[6][29]  ( .D(n2613), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2932), .QN(n920) );
  DFFNSRXLTS \dataoutbuffer_reg[6][27]  ( .D(n2615), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2936), .QN(n921) );
  DFFNSRXLTS \dataoutbuffer_reg[6][26]  ( .D(n2616), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2938), .QN(n922) );
  DFFNSRXLTS \dataoutbuffer_reg[6][25]  ( .D(n2617), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2940), .QN(n923) );
  DFFNSRXLTS \dataoutbuffer_reg[6][24]  ( .D(n2618), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2942), .QN(n924) );
  DFFNSRXLTS \dataoutbuffer_reg[6][23]  ( .D(n2619), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2944), .QN(n925) );
  DFFNSRXLTS \dataoutbuffer_reg[6][22]  ( .D(n2620), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2946), .QN(n926) );
  DFFNSRXLTS \dataoutbuffer_reg[6][21]  ( .D(n2621), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2948), .QN(n927) );
  DFFNSRXLTS \dataoutbuffer_reg[6][20]  ( .D(n2622), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2950), .QN(n928) );
  DFFNSRXLTS \dataoutbuffer_reg[6][19]  ( .D(n2623), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2952), .QN(n929) );
  DFFNSRXLTS \dataoutbuffer_reg[6][17]  ( .D(n2625), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2956), .QN(n930) );
  DFFNSRXLTS \dataoutbuffer_reg[6][16]  ( .D(n2626), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2958), .QN(n931) );
  DFFNSRXLTS \dataoutbuffer_reg[6][15]  ( .D(n2627), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2960), .QN(n932) );
  DFFNSRXLTS \dataoutbuffer_reg[6][13]  ( .D(n2629), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2964), .QN(n933) );
  DFFNSRXLTS \dataoutbuffer_reg[6][12]  ( .D(n2630), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2966), .QN(n934) );
  DFFNSRXLTS \dataoutbuffer_reg[6][11]  ( .D(n2631), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2968), .QN(n935) );
  DFFNSRXLTS \dataoutbuffer_reg[6][8]  ( .D(n2634), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n2974), .QN(n936) );
  DFFNSRXLTS \dataoutbuffer_reg[6][7]  ( .D(n2635), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n2976), .QN(n937) );
  DFFNSRXLTS \requesterAddressbuffer_reg[0][0]  ( .D(n2840), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][0] ), .QN(n592) );
  DFFNSRXLTS \requesterAddressbuffer_reg[0][1]  ( .D(n2839), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][1] ), .QN(n593) );
  DFFNSRXLTS \requesterAddressbuffer_reg[0][2]  ( .D(n2838), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][2] ), .QN(n594) );
  DFFNSRXLTS \requesterAddressbuffer_reg[0][4]  ( .D(n2836), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][4] ), .QN(n595) );
  DFFNSRXLTS \requesterAddressbuffer_reg[0][3]  ( .D(n2837), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][3] ), .QN(n596) );
  DFFNSRXLTS \requesterAddressbuffer_reg[0][5]  ( .D(n2835), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][5] ), .QN(n597) );
  DFFNSRXLTS \dataoutbuffer_reg[0][0]  ( .D(n2834), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n57), .QN(n605) );
  DFFNSRXLTS \dataoutbuffer_reg[0][1]  ( .D(n2833), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n56), .QN(n606) );
  DFFNSRXLTS \dataoutbuffer_reg[0][2]  ( .D(n2832), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n55), .QN(n607) );
  DFFNSRXLTS \dataoutbuffer_reg[0][5]  ( .D(n2829), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n54), .QN(n608) );
  DFFNSRXLTS \dataoutbuffer_reg[0][9]  ( .D(n2825), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n53), .QN(n609) );
  DFFNSRXLTS \dataoutbuffer_reg[0][20]  ( .D(n2814), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n52), .QN(n610) );
  DFFNSRXLTS \dataoutbuffer_reg[0][23]  ( .D(n2811), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n51), .QN(n611) );
  DFFNSRXLTS \dataoutbuffer_reg[0][27]  ( .D(n2807), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n50), .QN(n612) );
  DFFNSRXLTS \dataoutbuffer_reg[0][28]  ( .D(n2806), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n49), .QN(n613) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][0]  ( .D(n2464), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n48), .QN(n614) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][13]  ( .D(n2451), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3177), .QN(n562) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][13]  ( .D(n2479), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3185), .QN(n563) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][13]  ( .D(n2493), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3154), .QN(n568) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][13]  ( .D(n2465), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3123), .QN(n710) );
  DFFNSRXLTS \writeOutbuffer_reg[0]  ( .D(n2571), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n643) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][6]  ( .D(n2486), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3178), .QN(n550) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][8]  ( .D(n2484), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3180), .QN(n551) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][10]  ( .D(n2482), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3182), .QN(n552) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][12]  ( .D(n2480), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3184), .QN(n553) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][7]  ( .D(n2457), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3171), .QN(n554) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][9]  ( .D(n2455), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3173), .QN(n555) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][11]  ( .D(n2453), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3175), .QN(n556) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][7]  ( .D(n2485), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3179), .QN(n557) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][9]  ( .D(n2483), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3181), .QN(n558) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][11]  ( .D(n2481), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3183), .QN(n559) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][6]  ( .D(n2458), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3170), .QN(n560) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][10]  ( .D(n2454), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3174), .QN(n561) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][8]  ( .D(n2456), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3172), .QN(n564) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][12]  ( .D(n2452), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3176), .QN(n565) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][7]  ( .D(n2499), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3166), .QN(n566) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][10]  ( .D(n2496), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3160), .QN(n567) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][8]  ( .D(n2498), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3164), .QN(n577) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][9]  ( .D(n2497), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3162), .QN(n578) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][12]  ( .D(n2494), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3156), .QN(n579) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][6]  ( .D(n2500), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3168), .QN(n580) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][11]  ( .D(n2495), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3158), .QN(n581) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][6]  ( .D(n2472), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3130), .QN(n703) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][7]  ( .D(n2471), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3129), .QN(n704) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][8]  ( .D(n2470), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3128), .QN(n705) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][9]  ( .D(n2469), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3127), .QN(n706) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][10]  ( .D(n2468), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3126), .QN(n707) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][11]  ( .D(n2467), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3125), .QN(n708) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][12]  ( .D(n2466), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3124), .QN(n709) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][5]  ( .D(n2459), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n642), .QN(n4712) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][4]  ( .D(n2460), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n615), .QN(n4724) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][3]  ( .D(n2461), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n641), .QN(n4732) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][2]  ( .D(n2462), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n640), .QN(n4743) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][1]  ( .D(n2463), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n639), .QN(n4748) );
  DFFNSRXLTS \dataoutbuffer_reg[0][31]  ( .D(n2803), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n638), .QN(n4420) );
  DFFNSRXLTS \dataoutbuffer_reg[0][30]  ( .D(n2804), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n637), .QN(n4433) );
  DFFNSRXLTS \dataoutbuffer_reg[0][29]  ( .D(n2805), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n636), .QN(n4444) );
  DFFNSRXLTS \dataoutbuffer_reg[0][26]  ( .D(n2808), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n635), .QN(n4469) );
  DFFNSRXLTS \dataoutbuffer_reg[0][25]  ( .D(n2809), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n634), .QN(n4476) );
  DFFNSRXLTS \dataoutbuffer_reg[0][24]  ( .D(n2810), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n633), .QN(n4485) );
  DFFNSRXLTS \dataoutbuffer_reg[0][22]  ( .D(n2812), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n632), .QN(n4501) );
  DFFNSRXLTS \dataoutbuffer_reg[0][21]  ( .D(n2813), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n631), .QN(n4516) );
  DFFNSRXLTS \dataoutbuffer_reg[0][19]  ( .D(n2815), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n630), .QN(n4530) );
  DFFNSRXLTS \dataoutbuffer_reg[0][18]  ( .D(n2816), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n629), .QN(n4539) );
  DFFNSRXLTS \dataoutbuffer_reg[0][17]  ( .D(n2817), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n628), .QN(n4548) );
  DFFNSRXLTS \dataoutbuffer_reg[0][16]  ( .D(n2818), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n627), .QN(n4557) );
  DFFNSRXLTS \dataoutbuffer_reg[0][15]  ( .D(n2819), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n626), .QN(n4568) );
  DFFNSRXLTS \dataoutbuffer_reg[0][14]  ( .D(n2820), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n625), .QN(n4575) );
  DFFNSRXLTS \dataoutbuffer_reg[0][13]  ( .D(n2821), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n624), .QN(n4588) );
  DFFNSRXLTS \dataoutbuffer_reg[0][12]  ( .D(n2822), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n623), .QN(n4595) );
  DFFNSRXLTS \dataoutbuffer_reg[0][11]  ( .D(n2823), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n622), .QN(n4600) );
  DFFNSRXLTS \dataoutbuffer_reg[0][10]  ( .D(n2824), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n621), .QN(n4613) );
  DFFNSRXLTS \dataoutbuffer_reg[0][8]  ( .D(n2826), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n620), .QN(n4633) );
  DFFNSRXLTS \dataoutbuffer_reg[0][7]  ( .D(n2827), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n619), .QN(n4638) );
  DFFNSRXLTS \dataoutbuffer_reg[0][6]  ( .D(n2828), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n618), .QN(n4647) );
  DFFNSRXLTS \dataoutbuffer_reg[0][4]  ( .D(n2830), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n617), .QN(n4663) );
  DFFNSRXLTS \dataoutbuffer_reg[0][3]  ( .D(n2831), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n616), .QN(n4674) );
  DFFNSRXLTS \read_reg_reg[0]  ( .D(n2889), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n658), .QN(n10) );
  DFFNSRXLTS full_reg_reg ( .D(N4718), .CKN(clk), .SN(1'b1), .RN(1'b1), .QN(
        n96) );
  DFFNSRXLTS \destinationAddressOut_reg[7]  ( .D(n2447), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[7]) );
  DFFNSRXLTS \destinationAddressOut_reg[6]  ( .D(n2448), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[6]) );
  DFFNSRXLTS \destinationAddressOut_reg[9]  ( .D(n2445), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[9]) );
  DFFNSRXLTS \destinationAddressOut_reg[8]  ( .D(n2446), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[8]) );
  DFFNSRXLTS \destinationAddressOut_reg[13]  ( .D(n2441), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[13]) );
  DFFNSRXLTS \destinationAddressOut_reg[12]  ( .D(n2442), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[12]) );
  DFFNSRXLTS \destinationAddressOut_reg[11]  ( .D(n2443), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[11]) );
  DFFNSRXLTS \destinationAddressOut_reg[10]  ( .D(n2444), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[10]) );
  DFFNSRXLTS \write_reg_reg[0]  ( .D(n2888), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n9), .QN(n948) );
  DFFNSRXLTS \readOutbuffer_reg[5]  ( .D(n2568), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n600) );
  DFFNSRXLTS \readOutbuffer_reg[3]  ( .D(n2566), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n598) );
  DFFNSRXLTS \readOutbuffer_reg[6]  ( .D(n2569), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n599) );
  DFFNSRXLTS \readOutbuffer_reg[4]  ( .D(n2567), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n647) );
  DFFNSRXLTS \readOutbuffer_reg[1]  ( .D(n2564), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n601) );
  DFFNSRXLTS \readOutbuffer_reg[7]  ( .D(n2570), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer_7) );
  DFFNSRXLTS \readOutbuffer_reg[0]  ( .D(n2563), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n892) );
  DFFNSRXLTS \readOutbuffer_reg[2]  ( .D(n2565), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\readOutbuffer[2] ), .QN(n646) );
  DFFNSRXLTS \writeOutbuffer_reg[5]  ( .D(n2576), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n603) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][13]  ( .D(n2507), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3131), .QN(n583) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][12]  ( .D(n2508), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3132), .QN(n591) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][11]  ( .D(n2509), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3133), .QN(n590) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][10]  ( .D(n2510), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3134), .QN(n589) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][9]  ( .D(n2511), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3135), .QN(n582) );
  DFFNSRXLTS \writeOutbuffer_reg[4]  ( .D(n2575), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n645) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][8]  ( .D(n2512), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3136), .QN(n588) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][7]  ( .D(n2513), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3137), .QN(n587) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][6]  ( .D(n2514), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3138), .QN(n586) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][5]  ( .D(n2853), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][5] ), .QN(n877) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][4]  ( .D(n2854), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][4] ), .QN(n878) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][3]  ( .D(n2855), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][3] ), .QN(n876) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][2]  ( .D(n2856), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][2] ), .QN(n875) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][1]  ( .D(n2857), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][1] ), .QN(n874) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][0]  ( .D(n2858), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][0] ), .QN(n873) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][5]  ( .D(n2529), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n743) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][13]  ( .D(n2521), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3139), .QN(n576) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][12]  ( .D(n2522), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3141), .QN(n575) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][11]  ( .D(n2523), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3143), .QN(n574) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][10]  ( .D(n2524), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3145), .QN(n573) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][9]  ( .D(n2525), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3146), .QN(n572) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][8]  ( .D(n2526), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3148), .QN(n571) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][7]  ( .D(n2527), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3150), .QN(n570) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][6]  ( .D(n2528), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3152), .QN(n569) );
  DFFNSRXLTS \dataoutbuffer_reg[3][1]  ( .D(n2737), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n6275), .QN(n847) );
  DFFNSRXLTS \dataoutbuffer_reg[3][0]  ( .D(n2738), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n6276), .QN(n846) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][3]  ( .D(n2559), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n783) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][2]  ( .D(n2560), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n782) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][1]  ( .D(n2561), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n781) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][0]  ( .D(n2562), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n821) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][4]  ( .D(n2558), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n749) );
  DFFNSRXLTS \dataoutbuffer_reg[5][31]  ( .D(n2643), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n748) );
  DFFNSRXLTS \dataoutbuffer_reg[5][30]  ( .D(n2644), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n738) );
  DFFNSRXLTS \dataoutbuffer_reg[5][29]  ( .D(n2645), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n737) );
  DFFNSRXLTS \dataoutbuffer_reg[5][28]  ( .D(n2646), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n736) );
  DFFNSRXLTS \dataoutbuffer_reg[5][27]  ( .D(n2647), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n735) );
  DFFNSRXLTS \dataoutbuffer_reg[5][26]  ( .D(n2648), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n734) );
  DFFNSRXLTS \dataoutbuffer_reg[5][25]  ( .D(n2649), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n733) );
  DFFNSRXLTS \dataoutbuffer_reg[5][24]  ( .D(n2650), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n732) );
  DFFNSRXLTS \dataoutbuffer_reg[5][23]  ( .D(n2651), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n731) );
  DFFNSRXLTS \dataoutbuffer_reg[5][22]  ( .D(n2652), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n730) );
  DFFNSRXLTS \dataoutbuffer_reg[5][21]  ( .D(n2653), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n729) );
  DFFNSRXLTS \dataoutbuffer_reg[5][20]  ( .D(n2654), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n728) );
  DFFNSRXLTS \dataoutbuffer_reg[5][19]  ( .D(n2655), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n727) );
  DFFNSRXLTS \dataoutbuffer_reg[5][18]  ( .D(n2656), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n726) );
  DFFNSRXLTS \dataoutbuffer_reg[5][17]  ( .D(n2657), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n725) );
  DFFNSRXLTS \dataoutbuffer_reg[5][16]  ( .D(n2658), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n747) );
  DFFNSRXLTS \dataoutbuffer_reg[5][15]  ( .D(n2659), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n746) );
  DFFNSRXLTS \dataoutbuffer_reg[5][14]  ( .D(n2660), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n724) );
  DFFNSRXLTS \dataoutbuffer_reg[5][13]  ( .D(n2661), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n723) );
  DFFNSRXLTS \dataoutbuffer_reg[5][12]  ( .D(n2662), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n722) );
  DFFNSRXLTS \dataoutbuffer_reg[5][11]  ( .D(n2663), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n745) );
  DFFNSRXLTS \dataoutbuffer_reg[5][10]  ( .D(n2664), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n721) );
  DFFNSRXLTS \dataoutbuffer_reg[5][9]  ( .D(n2665), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n720) );
  DFFNSRXLTS \dataoutbuffer_reg[5][8]  ( .D(n2666), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n719) );
  DFFNSRXLTS \dataoutbuffer_reg[5][7]  ( .D(n2667), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n718) );
  DFFNSRXLTS \dataoutbuffer_reg[5][6]  ( .D(n2668), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n717) );
  DFFNSRXLTS \dataoutbuffer_reg[5][5]  ( .D(n2669), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n716) );
  DFFNSRXLTS \dataoutbuffer_reg[5][4]  ( .D(n2670), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n715) );
  DFFNSRXLTS \dataoutbuffer_reg[5][3]  ( .D(n2671), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n714) );
  DFFNSRXLTS \dataoutbuffer_reg[5][2]  ( .D(n2672), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n713) );
  DFFNSRXLTS \dataoutbuffer_reg[5][1]  ( .D(n2673), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n744) );
  DFFNSRXLTS \dataoutbuffer_reg[5][0]  ( .D(n2674), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n712) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][5]  ( .D(n2501), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n6250), .QN(n872) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][4]  ( .D(n2502), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n6251), .QN(n871) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][3]  ( .D(n2503), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n6252), .QN(n870) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][2]  ( .D(n2504), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n6291), .QN(n845) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][1]  ( .D(n2505), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n6253), .QN(n869) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][0]  ( .D(n2506), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n6254), .QN(n868) );
  DFFNSRXLTS \dataoutbuffer_reg[3][31]  ( .D(n2707), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6255), .QN(n867) );
  DFFNSRXLTS \dataoutbuffer_reg[3][30]  ( .D(n2708), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6256), .QN(n866) );
  DFFNSRXLTS \dataoutbuffer_reg[3][29]  ( .D(n2709), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6257), .QN(n865) );
  DFFNSRXLTS \dataoutbuffer_reg[3][28]  ( .D(n2710), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6258), .QN(n864) );
  DFFNSRXLTS \dataoutbuffer_reg[3][27]  ( .D(n2711), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6259), .QN(n863) );
  DFFNSRXLTS \dataoutbuffer_reg[3][26]  ( .D(n2712), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6260), .QN(n862) );
  DFFNSRXLTS \dataoutbuffer_reg[3][25]  ( .D(n2713), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6292), .QN(n844) );
  DFFNSRXLTS \dataoutbuffer_reg[3][24]  ( .D(n2714), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6261), .QN(n861) );
  DFFNSRXLTS \dataoutbuffer_reg[3][23]  ( .D(n2715), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6293), .QN(n843) );
  DFFNSRXLTS \dataoutbuffer_reg[3][22]  ( .D(n2716), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6262), .QN(n860) );
  DFFNSRXLTS \dataoutbuffer_reg[3][21]  ( .D(n2717), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6263), .QN(n859) );
  DFFNSRXLTS \dataoutbuffer_reg[3][20]  ( .D(n2718), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6294), .QN(n842) );
  DFFNSRXLTS \dataoutbuffer_reg[3][19]  ( .D(n2719), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6264), .QN(n858) );
  DFFNSRXLTS \dataoutbuffer_reg[3][18]  ( .D(n2720), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6295), .QN(n841) );
  DFFNSRXLTS \dataoutbuffer_reg[3][17]  ( .D(n2721), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6265), .QN(n857) );
  DFFNSRXLTS \dataoutbuffer_reg[3][16]  ( .D(n2722), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6266), .QN(n856) );
  DFFNSRXLTS \dataoutbuffer_reg[3][15]  ( .D(n2723), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6296), .QN(n840) );
  DFFNSRXLTS \dataoutbuffer_reg[3][14]  ( .D(n2724), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6267), .QN(n855) );
  DFFNSRXLTS \dataoutbuffer_reg[3][13]  ( .D(n2725), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6297), .QN(n839) );
  DFFNSRXLTS \dataoutbuffer_reg[3][12]  ( .D(n2726), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6268), .QN(n854) );
  DFFNSRXLTS \dataoutbuffer_reg[3][11]  ( .D(n2727), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6269), .QN(n853) );
  DFFNSRXLTS \dataoutbuffer_reg[3][10]  ( .D(n2728), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n6270), .QN(n852) );
  DFFNSRXLTS \dataoutbuffer_reg[3][9]  ( .D(n2729), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n6271), .QN(n851) );
  DFFNSRXLTS \dataoutbuffer_reg[3][8]  ( .D(n2730), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n6272), .QN(n850) );
  DFFNSRXLTS \dataoutbuffer_reg[3][7]  ( .D(n2731), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n6313), .QN(n835) );
  DFFNSRXLTS \dataoutbuffer_reg[3][6]  ( .D(n2732), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n6273), .QN(n849) );
  DFFNSRXLTS \dataoutbuffer_reg[3][5]  ( .D(n2733), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n6298), .QN(n838) );
  DFFNSRXLTS \dataoutbuffer_reg[3][4]  ( .D(n2734), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n6299), .QN(n837) );
  DFFNSRXLTS \dataoutbuffer_reg[3][3]  ( .D(n2735), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n6274), .QN(n848) );
  DFFNSRXLTS \dataoutbuffer_reg[3][2]  ( .D(n2736), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n6300), .QN(n836) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][13]  ( .D(n2549), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3140), .QN(n702) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][12]  ( .D(n2550), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3142), .QN(n907) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][11]  ( .D(n2551), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3144), .QN(n906) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][10]  ( .D(n2552), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n480), .QN(n833) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][9]  ( .D(n2553), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3147), .QN(n908) );
  DFFNSRXLTS \requesterAddressbuffer_reg[7][5]  ( .D(n2877), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n891) );
  DFFNSRXLTS \requesterAddressbuffer_reg[7][4]  ( .D(n2878), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n890) );
  DFFNSRXLTS \requesterAddressbuffer_reg[7][2]  ( .D(n2880), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n889) );
  DFFNSRXLTS \requesterAddressbuffer_reg[7][0]  ( .D(n2882), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n880) );
  DFFNSRXLTS \dataoutbuffer_reg[7][31]  ( .D(n2579), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n780) );
  DFFNSRXLTS \dataoutbuffer_reg[7][30]  ( .D(n2580), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n779) );
  DFFNSRXLTS \dataoutbuffer_reg[7][29]  ( .D(n2581), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n778) );
  DFFNSRXLTS \dataoutbuffer_reg[7][28]  ( .D(n2582), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n777) );
  DFFNSRXLTS \dataoutbuffer_reg[7][27]  ( .D(n2583), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n776) );
  DFFNSRXLTS \dataoutbuffer_reg[7][26]  ( .D(n2584), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n775) );
  DFFNSRXLTS \dataoutbuffer_reg[7][25]  ( .D(n2585), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n774) );
  DFFNSRXLTS \dataoutbuffer_reg[7][24]  ( .D(n2586), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n773) );
  DFFNSRXLTS \dataoutbuffer_reg[7][23]  ( .D(n2587), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n772) );
  DFFNSRXLTS \dataoutbuffer_reg[7][22]  ( .D(n2588), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n771) );
  DFFNSRXLTS \dataoutbuffer_reg[7][21]  ( .D(n2589), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n770) );
  DFFNSRXLTS \dataoutbuffer_reg[7][20]  ( .D(n2590), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n769) );
  DFFNSRXLTS \dataoutbuffer_reg[7][19]  ( .D(n2591), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n768) );
  DFFNSRXLTS \dataoutbuffer_reg[7][18]  ( .D(n2592), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n767) );
  DFFNSRXLTS \dataoutbuffer_reg[7][17]  ( .D(n2593), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n766) );
  DFFNSRXLTS \dataoutbuffer_reg[7][16]  ( .D(n2594), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n765) );
  DFFNSRXLTS \dataoutbuffer_reg[7][15]  ( .D(n2595), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n915) );
  DFFNSRXLTS \dataoutbuffer_reg[7][14]  ( .D(n2596), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n916) );
  DFFNSRXLTS \dataoutbuffer_reg[7][13]  ( .D(n2597), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n917) );
  DFFNSRXLTS \dataoutbuffer_reg[7][12]  ( .D(n2598), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n764) );
  DFFNSRXLTS \dataoutbuffer_reg[7][11]  ( .D(n2599), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n763) );
  DFFNSRXLTS \dataoutbuffer_reg[7][10]  ( .D(n2600), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n762) );
  DFFNSRXLTS \dataoutbuffer_reg[7][9]  ( .D(n2601), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n761) );
  DFFNSRXLTS \dataoutbuffer_reg[7][8]  ( .D(n2602), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n760) );
  DFFNSRXLTS \dataoutbuffer_reg[7][7]  ( .D(n2603), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n759) );
  DFFNSRXLTS \dataoutbuffer_reg[7][6]  ( .D(n2604), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n758) );
  DFFNSRXLTS \dataoutbuffer_reg[7][5]  ( .D(n2605), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n757) );
  DFFNSRXLTS \dataoutbuffer_reg[7][4]  ( .D(n2606), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n756) );
  DFFNSRXLTS \dataoutbuffer_reg[7][3]  ( .D(n2607), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n755) );
  DFFNSRXLTS \dataoutbuffer_reg[7][2]  ( .D(n2608), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n754) );
  DFFNSRXLTS \dataoutbuffer_reg[7][1]  ( .D(n2609), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n753) );
  DFFNSRXLTS \dataoutbuffer_reg[7][0]  ( .D(n2610), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n918) );
  DFFNSRXLTS \requesterAddressbuffer_reg[7][3]  ( .D(n2879), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n882) );
  DFFNSRXLTS \requesterAddressbuffer_reg[7][1]  ( .D(n2881), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n881) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][5]  ( .D(n2557), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n784) );
  DFFNSRXLTS \writeOutbuffer_reg[6]  ( .D(n2577), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n911) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][12]  ( .D(n2536), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3157), .QN(n585) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][11]  ( .D(n2537), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3159), .QN(n901) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][10]  ( .D(n2538), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3161), .QN(n584) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][9]  ( .D(n2539), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3163), .QN(n910) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][8]  ( .D(n2540), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3165), .QN(n900) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][7]  ( .D(n2541), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3167), .QN(n899) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][6]  ( .D(n2542), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3169), .QN(n909) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][13]  ( .D(n2535), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3155), .QN(n902) );
  DFFNSRXLTS \writeOutbuffer_reg[7]  ( .D(n2578), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n879) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][8]  ( .D(n2554), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3149), .QN(n905) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][7]  ( .D(n2555), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3151), .QN(n904) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][6]  ( .D(n2556), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3153), .QN(n903) );
  DFFNSRXLTS \requesterAddressbuffer_reg[4][3]  ( .D(n2861), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2925) );
  DFFNSRXLTS \requesterAddressbuffer_reg[4][2]  ( .D(n2862), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2923) );
  DFFNSRXLTS \requesterAddressbuffer_reg[4][1]  ( .D(n2863), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2924) );
  DFFNSRXLTS \requesterAddressbuffer_reg[4][0]  ( .D(n2864), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2926) );
  DFFNSRXLTS \requesterAddressbuffer_reg[4][5]  ( .D(n2859), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2921) );
  DFFNSRXLTS \requesterAddressbuffer_reg[4][4]  ( .D(n2860), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2922) );
  DFFNSRXLTS \requesterAddressbuffer_reg[2][3]  ( .D(n2849), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][3] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[2][2]  ( .D(n2850), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][2] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[2][1]  ( .D(n2851), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][1] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[2][0]  ( .D(n2852), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][0] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[2][5]  ( .D(n2847), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][5] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[2][4]  ( .D(n2848), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][4] ) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][1]  ( .D(n2519), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2999) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][0]  ( .D(n2520), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3001) );
  DFFNSRXLTS \dataoutbuffer_reg[4][31]  ( .D(n2675), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2927) );
  DFFNSRXLTS \dataoutbuffer_reg[4][30]  ( .D(n2676), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2929) );
  DFFNSRXLTS \dataoutbuffer_reg[4][29]  ( .D(n2677), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2931) );
  DFFNSRXLTS \dataoutbuffer_reg[4][28]  ( .D(n2678), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2933) );
  DFFNSRXLTS \dataoutbuffer_reg[4][27]  ( .D(n2679), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2935) );
  DFFNSRXLTS \dataoutbuffer_reg[4][26]  ( .D(n2680), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2937) );
  DFFNSRXLTS \dataoutbuffer_reg[4][25]  ( .D(n2681), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2939) );
  DFFNSRXLTS \dataoutbuffer_reg[4][24]  ( .D(n2682), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2941) );
  DFFNSRXLTS \dataoutbuffer_reg[4][23]  ( .D(n2683), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2943) );
  DFFNSRXLTS \dataoutbuffer_reg[4][22]  ( .D(n2684), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2945) );
  DFFNSRXLTS \dataoutbuffer_reg[4][21]  ( .D(n2685), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2947) );
  DFFNSRXLTS \dataoutbuffer_reg[4][20]  ( .D(n2686), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2949) );
  DFFNSRXLTS \dataoutbuffer_reg[4][19]  ( .D(n2687), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2951) );
  DFFNSRXLTS \dataoutbuffer_reg[4][18]  ( .D(n2688), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2953) );
  DFFNSRXLTS \dataoutbuffer_reg[4][17]  ( .D(n2689), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2955) );
  DFFNSRXLTS \dataoutbuffer_reg[4][16]  ( .D(n2690), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2957) );
  DFFNSRXLTS \dataoutbuffer_reg[4][15]  ( .D(n2691), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2959) );
  DFFNSRXLTS \dataoutbuffer_reg[4][14]  ( .D(n2692), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2961) );
  DFFNSRXLTS \dataoutbuffer_reg[4][13]  ( .D(n2693), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2963) );
  DFFNSRXLTS \dataoutbuffer_reg[4][12]  ( .D(n2694), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2965) );
  DFFNSRXLTS \dataoutbuffer_reg[4][11]  ( .D(n2695), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2967) );
  DFFNSRXLTS \dataoutbuffer_reg[4][10]  ( .D(n2696), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2969) );
  DFFNSRXLTS \dataoutbuffer_reg[4][9]  ( .D(n2697), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n2971) );
  DFFNSRXLTS \dataoutbuffer_reg[4][8]  ( .D(n2698), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n2973) );
  DFFNSRXLTS \dataoutbuffer_reg[4][7]  ( .D(n2699), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n2975) );
  DFFNSRXLTS \dataoutbuffer_reg[4][6]  ( .D(n2700), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n2977) );
  DFFNSRXLTS \dataoutbuffer_reg[4][5]  ( .D(n2701), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n2979) );
  DFFNSRXLTS \dataoutbuffer_reg[4][4]  ( .D(n2702), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n2981) );
  DFFNSRXLTS \dataoutbuffer_reg[4][3]  ( .D(n2703), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n2983) );
  DFFNSRXLTS \dataoutbuffer_reg[4][2]  ( .D(n2704), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n2985) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][5]  ( .D(n2515), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2991) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][4]  ( .D(n2516), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2993) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][3]  ( .D(n2517), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2995) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][2]  ( .D(n2518), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2997) );
  DFFNSRXLTS \dataoutbuffer_reg[4][1]  ( .D(n2705), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n2987) );
  DFFNSRXLTS \dataoutbuffer_reg[4][0]  ( .D(n2706), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n2989) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][5]  ( .D(n2487), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n81) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][1]  ( .D(n2491), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n84) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][0]  ( .D(n2492), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n85) );
  DFFNSRXLTS \dataoutbuffer_reg[2][31]  ( .D(n2739), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n89) );
  DFFNSRXLTS \dataoutbuffer_reg[2][30]  ( .D(n2740), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n59) );
  DFFNSRXLTS \dataoutbuffer_reg[2][29]  ( .D(n2741), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n60) );
  DFFNSRXLTS \dataoutbuffer_reg[2][28]  ( .D(n2742), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n61) );
  DFFNSRXLTS \dataoutbuffer_reg[2][27]  ( .D(n2743), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n86) );
  DFFNSRXLTS \dataoutbuffer_reg[2][26]  ( .D(n2744), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n62) );
  DFFNSRXLTS \dataoutbuffer_reg[2][25]  ( .D(n2745), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n63) );
  DFFNSRXLTS \dataoutbuffer_reg[2][24]  ( .D(n2746), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n90) );
  DFFNSRXLTS \dataoutbuffer_reg[2][23]  ( .D(n2747), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n64) );
  DFFNSRXLTS \dataoutbuffer_reg[2][22]  ( .D(n2748), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n91) );
  DFFNSRXLTS \dataoutbuffer_reg[2][21]  ( .D(n2749), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n65) );
  DFFNSRXLTS \dataoutbuffer_reg[2][20]  ( .D(n2750), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n66) );
  BUFX3TS U2 ( .A(n1840), .Y(n972) );
  XOR2X2TS U3 ( .A(n2010), .B(n6), .Y(n1840) );
  NAND2X2TS U4 ( .A(n970), .B(n971), .Y(n1957) );
  OAI221XLTS U5 ( .A0(n6), .A1(n688), .B0(n1798), .B1(n1956), .C0(n1800), .Y(
        n1799) );
  INVX2TS U6 ( .A(n3199), .Y(n3122) );
  CLKBUFX2TS U7 ( .A(n3608), .Y(n3606) );
  CLKBUFX2TS U8 ( .A(n3561), .Y(n3559) );
  OAI21X2TS U9 ( .A0(n1827), .A1(n1864), .B0(n3122), .Y(n1770) );
  INVX2TS U10 ( .A(n109), .Y(n110) );
  CLKBUFX2TS U11 ( .A(n3261), .Y(n3258) );
  CLKBUFX2TS U12 ( .A(n3414), .Y(n3402) );
  OAI32X1TS U13 ( .A0(n4214), .A1(n695), .A2(n1798), .B0(n1799), .B1(n964), 
        .Y(n1797) );
  CLKINVX2TS U14 ( .A(selectBit_SOUTH), .Y(n468) );
  CLKINVX2TS U15 ( .A(n914), .Y(n675) );
  INVX2TS U16 ( .A(n941), .Y(n679) );
  CLKINVX2TS U17 ( .A(n1752), .Y(n664) );
  CLKINVX1TS U18 ( .A(n1743), .Y(n940) );
  INVX1TS U19 ( .A(n1840), .Y(n699) );
  AO21X4TS U20 ( .A0(n1839), .A1(n123), .B0(n1782), .Y(n1784) );
  CLKBUFX2TS U21 ( .A(n468), .Y(n1) );
  XOR2X1TS U22 ( .A(n955), .B(selectBit_EAST), .Y(n2902) );
  INVX2TS U23 ( .A(selectBit_NORTH), .Y(n955) );
  OAI21XLTS U24 ( .A0(n960), .A1(n2004), .B0(n110), .Y(n2003) );
  AOI2BB1X4TS U25 ( .A0N(n110), .A1N(n1909), .B0(n1784), .Y(n1780) );
  NAND3X1TS U26 ( .A(n1840), .B(n1866), .C(n1841), .Y(n1863) );
  INVX2TS U27 ( .A(n973), .Y(n974) );
  NOR2X1TS U28 ( .A(selectBit_NORTH), .B(selectBit_SOUTH), .Y(n2379) );
  NOR2X1TS U29 ( .A(n119), .B(n194), .Y(n2008) );
  OAI21X1TS U30 ( .A0(n145), .A1(n1837), .B0(n1838), .Y(n1095) );
  OAI21X1TS U31 ( .A0(n698), .A1(n686), .B0(n678), .Y(n1838) );
  CLKBUFX2TS U32 ( .A(n1095), .Y(n3778) );
  NAND2X1TS U33 ( .A(n967), .B(n2008), .Y(n971) );
  NAND2X1TS U34 ( .A(n2007), .B(n969), .Y(n970) );
  INVX2TS U35 ( .A(n2007), .Y(n967) );
  INVX2TS U36 ( .A(n961), .Y(n670) );
  OA22X1TS U37 ( .A0(n1768), .A1(n180), .B0(n1827), .B1(n1865), .Y(n987) );
  INVX2TS U38 ( .A(n1770), .Y(n671) );
  OR2X2TS U39 ( .A(n978), .B(n468), .Y(n979) );
  NOR2BX1TS U40 ( .AN(n1794), .B(n688), .Y(n1180) );
  CLKBUFX2TS U41 ( .A(n1098), .Y(n3758) );
  CLKBUFX2TS U42 ( .A(n3502), .Y(n3496) );
  AND2X2TS U43 ( .A(n1780), .B(n667), .Y(n1745) );
  OA22X1TS U44 ( .A0(n1780), .A1(n180), .B0(n1865), .B1(n1879), .Y(n1746) );
  NOR2X1TS U45 ( .A(n1023), .B(n1957), .Y(n1841) );
  AND2X2TS U46 ( .A(n1957), .B(selectBit_WEST), .Y(n1888) );
  OA22X1TS U47 ( .A0(n1811), .A1(n178), .B0(n1865), .B1(n128), .Y(n986) );
  NOR3BX1TS U48 ( .AN(n1808), .B(n124), .C(n692), .Y(n1213) );
  NOR2BX1TS U49 ( .AN(n1794), .B(n1800), .Y(n1182) );
  CLKBUFX2TS U50 ( .A(n1213), .Y(n3266) );
  CLKBUFX2TS U51 ( .A(n987), .Y(n3201) );
  OA21XLTS U52 ( .A0(n1933), .A1(n1910), .B0(n1791), .Y(n1932) );
  AOI21X1TS U53 ( .A0(n945), .A1(n700), .B0(n664), .Y(n1794) );
  CLKBUFX2TS U54 ( .A(n3615), .Y(n3608) );
  OA22X1TS U55 ( .A0(n1776), .A1(n179), .B0(n1837), .B1(n130), .Y(n984) );
  CLKBUFX2TS U56 ( .A(n3409), .Y(n3408) );
  CLKBUFX2TS U57 ( .A(n3865), .Y(n3861) );
  CLKBUFX2TS U58 ( .A(n3757), .Y(n3756) );
  CLKBUFX2TS U59 ( .A(n3725), .Y(n3724) );
  CLKBUFX2TS U60 ( .A(n3614), .Y(n3607) );
  CLKBUFX2TS U61 ( .A(n3822), .Y(n3821) );
  CLKBUFX2TS U62 ( .A(n3822), .Y(n3820) );
  CLKBUFX2TS U63 ( .A(n3497), .Y(n3495) );
  CLKBUFX2TS U64 ( .A(n1794), .Y(n102) );
  OAI21X1TS U65 ( .A0(n124), .A1(n1956), .B0(n2002), .Y(n1813) );
  INVX2TS U66 ( .A(n1761), .Y(n698) );
  AOI21X1TS U67 ( .A0(n132), .A1(n684), .B0(n693), .Y(n1806) );
  OAI21X1TS U68 ( .A0(n1864), .A1(n130), .B0(n483), .Y(n1785) );
  NOR2BX1TS U69 ( .AN(n1839), .B(n1798), .Y(n1767) );
  NOR3X1TS U70 ( .A(n1767), .B(n1769), .C(n697), .Y(n1768) );
  AOI21X1TS U71 ( .A0(n1789), .A1(n684), .B0(n696), .Y(n1791) );
  NAND3X1TS U72 ( .A(n1841), .B(n699), .C(n116), .Y(n1790) );
  CLKBUFX2TS U73 ( .A(n3343), .Y(n3341) );
  NAND2X1TS U74 ( .A(n685), .B(n1794), .Y(n1751) );
  CLKBUFX2TS U75 ( .A(n3580), .Y(n3570) );
  CLKBUFX2TS U76 ( .A(n3580), .Y(n3571) );
  AOI222XLTS U77 ( .A0(n4417), .A1(n3859), .B0(n502), .B1(n3652), .C0(n4322), 
        .C1(n3642), .Y(n1653) );
  AOI222XLTS U78 ( .A0(n4422), .A1(n3859), .B0(n524), .B1(n3652), .C0(n4325), 
        .C1(n3642), .Y(n1655) );
  AOI222XLTS U79 ( .A0(n4425), .A1(n3859), .B0(n522), .B1(n3651), .C0(n4328), 
        .C1(n3643), .Y(n1657) );
  AOI222XLTS U80 ( .A0(n4429), .A1(n3859), .B0(n500), .B1(n3651), .C0(n4331), 
        .C1(n3643), .Y(n1659) );
  AOI222XLTS U81 ( .A0(n4432), .A1(n3860), .B0(n520), .B1(n3651), .C0(n4334), 
        .C1(n3643), .Y(n1661) );
  AOI222XLTS U82 ( .A0(n4436), .A1(n3860), .B0(n518), .B1(n3661), .C0(n4337), 
        .C1(n3643), .Y(n1663) );
  AOI222XLTS U83 ( .A0(n4440), .A1(n3860), .B0(n516), .B1(n3654), .C0(n4340), 
        .C1(n3644), .Y(n1665) );
  AOI222XLTS U84 ( .A0(n4443), .A1(n3860), .B0(n498), .B1(n3651), .C0(n4343), 
        .C1(n3644), .Y(n1667) );
  AOI222XLTS U85 ( .A0(n4451), .A1(n3864), .B0(n514), .B1(n3659), .C0(n4349), 
        .C1(n3644), .Y(n1671) );
  AOI222XLTS U86 ( .A0(n4458), .A1(n3864), .B0(n510), .B1(n3657), .C0(n4355), 
        .C1(n3639), .Y(n1675) );
  AOI222XLTS U87 ( .A0(n4454), .A1(n3862), .B0(n512), .B1(n3660), .C0(n4352), 
        .C1(n3649), .Y(n1673) );
  AOI222XLTS U88 ( .A0(n4448), .A1(n3863), .B0(n496), .B1(n3661), .C0(n4346), 
        .C1(n3644), .Y(n1669) );
  AOI222XLTS U89 ( .A0(n4533), .A1(n3336), .B0(n526), .B1(n3324), .C0(n4319), 
        .C1(n3311), .Y(n1330) );
  AOI222XLTS U90 ( .A0(n4499), .A1(n3347), .B0(n544), .B1(n3330), .C0(n4292), 
        .C1(n3309), .Y(n1312) );
  AOI222XLTS U91 ( .A0(n4493), .A1(n3346), .B0(n546), .B1(n3330), .C0(n4286), 
        .C1(n3308), .Y(n1308) );
  AOI222XLTS U92 ( .A0(n4481), .A1(n3347), .B0(n506), .B1(n3326), .C0(n4277), 
        .C1(n3308), .Y(n1302) );
  AOI222XLTS U93 ( .A0(n4470), .A1(n3347), .B0(n508), .B1(n3326), .C0(n4268), 
        .C1(n3307), .Y(n1296) );
  AOI222XLTS U94 ( .A0(n4529), .A1(n3335), .B0(n528), .B1(n3322), .C0(n4316), 
        .C1(n3311), .Y(n1328) );
  AOI222XLTS U95 ( .A0(n4525), .A1(n3335), .B0(n530), .B1(n3324), .C0(n4313), 
        .C1(n3311), .Y(n1326) );
  AOI222XLTS U96 ( .A0(n4522), .A1(n3335), .B0(n532), .B1(n3320), .C0(n4310), 
        .C1(n3311), .Y(n1324) );
  AOI222XLTS U97 ( .A0(n4519), .A1(n3335), .B0(n534), .B1(n3323), .C0(n4307), 
        .C1(n3310), .Y(n1322) );
  AOI222XLTS U98 ( .A0(n4514), .A1(n3346), .B0(n536), .B1(n3322), .C0(n4304), 
        .C1(n3310), .Y(n1320) );
  AOI222XLTS U99 ( .A0(n4511), .A1(n3350), .B0(n538), .B1(n3325), .C0(n4301), 
        .C1(n3310), .Y(n1318) );
  AOI222XLTS U100 ( .A0(n4507), .A1(n1196), .B0(n540), .B1(n3324), .C0(n4298), 
        .C1(n3309), .Y(n1316) );
  AOI222XLTS U101 ( .A0(n4504), .A1(n1196), .B0(n542), .B1(n3331), .C0(n4295), 
        .C1(n3309), .Y(n1314) );
  AOI222XLTS U102 ( .A0(n4496), .A1(n3336), .B0(n504), .B1(n3325), .C0(n4289), 
        .C1(n3309), .Y(n1310) );
  AOI222XLTS U103 ( .A0(n4489), .A1(n3348), .B0(n548), .B1(n3325), .C0(n4283), 
        .C1(n3308), .Y(n1306) );
  AOI222XLTS U104 ( .A0(n4486), .A1(n3348), .B0(n659), .B1(n3325), .C0(n4280), 
        .C1(n3310), .Y(n1304) );
  AOI222XLTS U105 ( .A0(n4478), .A1(n3347), .B0(n663), .B1(n3326), .C0(n4274), 
        .C1(n3308), .Y(n1300) );
  AOI222XLTS U106 ( .A0(n4474), .A1(n3344), .B0(n672), .B1(n3333), .C0(n4271), 
        .C1(n3307), .Y(n1298) );
  AOI222XLTS U107 ( .A0(n4466), .A1(n3334), .B0(n674), .B1(n3326), .C0(n4265), 
        .C1(n3307), .Y(n1294) );
  AOI222XLTS U108 ( .A0(n4462), .A1(n3334), .B0(n677), .B1(n3324), .C0(n4262), 
        .C1(n3307), .Y(n1292) );
  NOR2X1TS U109 ( .A(n1), .B(n2005), .Y(n2001) );
  OAI21X1TS U110 ( .A0(n1932), .A1(n180), .B0(n1923), .Y(n2) );
  AND2X2TS U111 ( .A(n947), .B(n990), .Y(n4) );
  AO21X1TS U112 ( .A0(n943), .A1(n129), .B0(n984), .Y(n7) );
  CLKBUFX2TS U113 ( .A(n670), .Y(n3866) );
  CLKBUFX2TS U114 ( .A(n1166), .Y(n3451) );
  OR2X2TS U115 ( .A(n6248), .B(n4605), .Y(n8) );
  AND2X2TS U116 ( .A(n96), .B(n2045), .Y(n11) );
  INVX1TS U117 ( .A(n1783), .Y(n123) );
  XNOR2X1TS U118 ( .A(n108), .B(n990), .Y(n12) );
  OR2X2TS U119 ( .A(n955), .B(n194), .Y(n13) );
  AND2X2TS U120 ( .A(n6248), .B(n4606), .Y(n14) );
  CLKBUFX2TS U121 ( .A(readIn_NORTH), .Y(n15) );
  INVXLTS U122 ( .A(readRequesterAddress[0]), .Y(n16) );
  INVXLTS U123 ( .A(n16), .Y(n17) );
  INVXLTS U124 ( .A(n16), .Y(n18) );
  INVXLTS U125 ( .A(n16), .Y(n19) );
  INVXLTS U126 ( .A(n16), .Y(n20) );
  INVXLTS U127 ( .A(readRequesterAddress[1]), .Y(n21) );
  INVXLTS U128 ( .A(n21), .Y(n22) );
  INVXLTS U129 ( .A(n21), .Y(n23) );
  INVXLTS U130 ( .A(n21), .Y(n24) );
  INVXLTS U131 ( .A(n21), .Y(n25) );
  INVXLTS U132 ( .A(readRequesterAddress[2]), .Y(n26) );
  INVXLTS U133 ( .A(n26), .Y(n27) );
  INVXLTS U134 ( .A(n26), .Y(n28) );
  INVXLTS U135 ( .A(n26), .Y(n29) );
  INVXLTS U136 ( .A(n26), .Y(n30) );
  INVXLTS U137 ( .A(readRequesterAddress[3]), .Y(n31) );
  INVXLTS U138 ( .A(n31), .Y(n32) );
  INVXLTS U139 ( .A(n31), .Y(n33) );
  INVXLTS U140 ( .A(n31), .Y(n34) );
  INVXLTS U141 ( .A(n31), .Y(n35) );
  INVXLTS U142 ( .A(readRequesterAddress[4]), .Y(n36) );
  INVXLTS U143 ( .A(n36), .Y(n37) );
  INVXLTS U144 ( .A(n36), .Y(n38) );
  INVXLTS U145 ( .A(n36), .Y(n39) );
  INVXLTS U146 ( .A(n36), .Y(n40) );
  INVXLTS U147 ( .A(readRequesterAddress[5]), .Y(n41) );
  INVXLTS U148 ( .A(n41), .Y(n42) );
  INVXLTS U149 ( .A(n41), .Y(n43) );
  INVXLTS U150 ( .A(n41), .Y(n44) );
  INVXLTS U151 ( .A(n41), .Y(n45) );
  INVXLTS U152 ( .A(n121), .Y(n46) );
  INVXLTS U153 ( .A(n5323), .Y(n47) );
  INVXLTS U154 ( .A(n385), .Y(n97) );
  INVXLTS U155 ( .A(n475), .Y(n98) );
  CLKBUFX2TS U156 ( .A(n1782), .Y(n99) );
  NOR3BX1TS U157 ( .AN(n1888), .B(n473), .C(n944), .Y(n1782) );
  CLKBUFX2TS U158 ( .A(n1808), .Y(n100) );
  AND2X2TS U159 ( .A(n1811), .B(n1808), .Y(n1214) );
  CLKBUFX2TS U160 ( .A(n1802), .Y(n101) );
  INVXLTS U161 ( .A(n7), .Y(n103) );
  INVXLTS U162 ( .A(n7), .Y(n104) );
  INVXLTS U163 ( .A(n1081), .Y(n105) );
  INVXLTS U164 ( .A(n105), .Y(n106) );
  CLKINVX2TS U165 ( .A(n13), .Y(n107) );
  INVX1TS U166 ( .A(n13), .Y(n108) );
  INVX1TS U167 ( .A(n1793), .Y(n109) );
  INVXLTS U168 ( .A(n3936), .Y(n111) );
  INVXLTS U169 ( .A(n3936), .Y(n112) );
  INVXLTS U170 ( .A(n182), .Y(n113) );
  INVXLTS U171 ( .A(n113), .Y(n114) );
  INVX2TS U172 ( .A(n944), .Y(n115) );
  INVXLTS U173 ( .A(n115), .Y(n116) );
  INVXLTS U174 ( .A(n2001), .Y(n117) );
  INVX2TS U175 ( .A(n2897), .Y(n118) );
  CLKINVX1TS U176 ( .A(n2897), .Y(n119) );
  INVXLTS U177 ( .A(n2004), .Y(n120) );
  INVXLTS U178 ( .A(n6), .Y(n121) );
  INVXLTS U179 ( .A(n3), .Y(n122) );
  INVXLTS U180 ( .A(n123), .Y(n124) );
  INVXLTS U181 ( .A(n12), .Y(n125) );
  INVXLTS U182 ( .A(n12), .Y(n126) );
  INVXLTS U183 ( .A(n1971), .Y(n127) );
  INVXLTS U184 ( .A(n127), .Y(n128) );
  INVXLTS U185 ( .A(n1879), .Y(n129) );
  INVXLTS U186 ( .A(n129), .Y(n130) );
  INVXLTS U187 ( .A(n1774), .Y(n131) );
  INVXLTS U188 ( .A(n131), .Y(n132) );
  INVXLTS U189 ( .A(n3810), .Y(n133) );
  INVXLTS U190 ( .A(n133), .Y(n134) );
  INVXLTS U191 ( .A(n133), .Y(n135) );
  INVXLTS U192 ( .A(n189), .Y(n136) );
  INVXLTS U193 ( .A(readIn_SOUTH), .Y(n137) );
  INVXLTS U194 ( .A(readIn_SOUTH), .Y(n138) );
  INVXLTS U195 ( .A(n658), .Y(n139) );
  INVXLTS U196 ( .A(n139), .Y(n140) );
  INVXLTS U197 ( .A(n5), .Y(n141) );
  INVXLTS U198 ( .A(n14), .Y(n142) );
  INVXLTS U199 ( .A(n14), .Y(n143) );
  INVXLTS U200 ( .A(n1827), .Y(n144) );
  INVXLTS U201 ( .A(n144), .Y(n145) );
  INVXLTS U202 ( .A(destinationAddressIn_NORTH[7]), .Y(n146) );
  INVXLTS U203 ( .A(destinationAddressIn_NORTH[7]), .Y(n147) );
  INVXLTS U204 ( .A(destinationAddressIn_NORTH[6]), .Y(n148) );
  INVXLTS U205 ( .A(destinationAddressIn_NORTH[6]), .Y(n149) );
  INVXLTS U206 ( .A(destinationAddressIn_NORTH[13]), .Y(n150) );
  INVXLTS U207 ( .A(destinationAddressIn_NORTH[13]), .Y(n151) );
  INVXLTS U208 ( .A(destinationAddressIn_NORTH[11]), .Y(n152) );
  INVXLTS U209 ( .A(destinationAddressIn_NORTH[11]), .Y(n153) );
  INVXLTS U210 ( .A(destinationAddressIn_NORTH[9]), .Y(n154) );
  INVXLTS U211 ( .A(destinationAddressIn_NORTH[9]), .Y(n155) );
  INVXLTS U212 ( .A(destinationAddressIn_NORTH[12]), .Y(n156) );
  INVXLTS U213 ( .A(destinationAddressIn_NORTH[12]), .Y(n157) );
  INVXLTS U214 ( .A(destinationAddressIn_NORTH[10]), .Y(n158) );
  INVXLTS U215 ( .A(destinationAddressIn_NORTH[10]), .Y(n159) );
  INVXLTS U216 ( .A(destinationAddressIn_NORTH[8]), .Y(n160) );
  INVXLTS U217 ( .A(destinationAddressIn_NORTH[8]), .Y(n161) );
  INVXLTS U218 ( .A(n4), .Y(n162) );
  INVXLTS U219 ( .A(n4), .Y(n163) );
  INVXLTS U220 ( .A(n656), .Y(n164) );
  INVXLTS U221 ( .A(n164), .Y(n165) );
  INVXLTS U222 ( .A(n164), .Y(n166) );
  INVXLTS U223 ( .A(n657), .Y(n167) );
  INVXLTS U224 ( .A(n167), .Y(n168) );
  INVXLTS U225 ( .A(n167), .Y(n169) );
  INVXLTS U226 ( .A(n652), .Y(n170) );
  INVXLTS U227 ( .A(n170), .Y(n171) );
  INVXLTS U228 ( .A(n170), .Y(n172) );
  INVXLTS U229 ( .A(n648), .Y(n173) );
  INVXLTS U230 ( .A(n173), .Y(n174) );
  INVXLTS U231 ( .A(n173), .Y(n175) );
  INVX2TS U232 ( .A(n1751), .Y(n662) );
  INVXLTS U233 ( .A(n2043), .Y(n176) );
  INVXLTS U234 ( .A(n2043), .Y(n177) );
  INVXLTS U235 ( .A(n11), .Y(n178) );
  INVXLTS U236 ( .A(n11), .Y(n179) );
  INVXLTS U237 ( .A(n11), .Y(n180) );
  AOI222XLTS U238 ( .A0(n4236), .A1(n3340), .B0(n3327), .B1(n42), .C0(n4009), 
        .C1(n3306), .Y(n1970) );
  INVXLTS U239 ( .A(n8), .Y(n181) );
  INVXLTS U240 ( .A(n8), .Y(n182) );
  INVXLTS U241 ( .A(n8), .Y(n183) );
  INVXLTS U242 ( .A(n8), .Y(n184) );
  INVXLTS U243 ( .A(n3811), .Y(n185) );
  INVXLTS U244 ( .A(n185), .Y(n186) );
  INVXLTS U245 ( .A(n185), .Y(n187) );
  INVXLTS U246 ( .A(n185), .Y(n188) );
  INVXLTS U247 ( .A(n3810), .Y(n189) );
  INVXLTS U248 ( .A(n189), .Y(n190) );
  INVXLTS U249 ( .A(n189), .Y(n191) );
  INVXLTS U250 ( .A(n189), .Y(n192) );
  INVXLTS U251 ( .A(n948), .Y(n193) );
  INVXLTS U252 ( .A(n193), .Y(n194) );
  INVXLTS U253 ( .A(n193), .Y(n195) );
  INVX2TS U523 ( .A(selectBit_EAST), .Y(n968) );
  AOI21X1TS U524 ( .A0(n1839), .A1(n1774), .B0(n694), .Y(n1776) );
  INVX1TS U525 ( .A(n1775), .Y(n694) );
  NAND3X1TS U526 ( .A(n473), .B(n1866), .C(n1888), .Y(n2002) );
  AND3XLTS U527 ( .A(n104), .B(n162), .C(n1776), .Y(n1743) );
  INVX1TS U528 ( .A(n1805), .Y(n693) );
  NAND3X1TS U529 ( .A(n699), .B(n1866), .C(n1841), .Y(n1800) );
  OAI21X1TS U530 ( .A0(n1932), .A1(n179), .B0(n1923), .Y(n466) );
  CLKBUFX2TS U531 ( .A(n136), .Y(n3809) );
  NAND3X1TS U532 ( .A(n947), .B(n47), .C(n691), .Y(n1763) );
  INVX2TS U533 ( .A(n468), .Y(n469) );
  AOI32XLTS U534 ( .A0(n974), .A1(n1), .A2(selectBit_NORTH), .B0(n2902), .B1(
        n469), .Y(n2901) );
  INVX2TS U535 ( .A(n1078), .Y(n470) );
  CLKBUFX2TS U536 ( .A(writeIn_NORTH), .Y(n965) );
  INVX2TS U537 ( .A(n965), .Y(n471) );
  INVX2TS U538 ( .A(n965), .Y(n472) );
  CLKINVX2TS U539 ( .A(n972), .Y(n473) );
  CLKBUFX2TS U540 ( .A(n2378), .Y(n474) );
  NOR2X1TS U541 ( .A(readReady), .B(selectBit_WEST), .Y(n2378) );
  CLKBUFX2TS U542 ( .A(n2030), .Y(n649) );
  INVX2TS U543 ( .A(n649), .Y(n477) );
  INVX2TS U544 ( .A(n649), .Y(n478) );
  CLKAND2X2TS U545 ( .A(n1768), .B(n671), .Y(n1741) );
  CLKINVX2TS U546 ( .A(n1741), .Y(n479) );
  CLKINVX2TS U547 ( .A(n1741), .Y(n481) );
  INVXLTS U548 ( .A(n1741), .Y(n482) );
  INVX2TS U549 ( .A(n1746), .Y(n483) );
  INVXLTS U550 ( .A(n1746), .Y(n484) );
  INVXLTS U551 ( .A(n1746), .Y(n485) );
  CLKBUFX2TS U552 ( .A(n1786), .Y(n487) );
  AND2XLTS U553 ( .A(n696), .B(n1786), .Y(n981) );
  AND3XLTS U554 ( .A(n1791), .B(n110), .C(n1786), .Y(n1166) );
  CLKBUFX2TS U555 ( .A(n1764), .Y(n488) );
  OAI21X1TS U556 ( .A0(n1836), .A1(n145), .B0(n1095), .Y(n1764) );
  INVX2TS U557 ( .A(n953), .Y(n489) );
  NAND2X1TS U558 ( .A(n979), .B(n980), .Y(n2009) );
  OAI2BB1X1TS U559 ( .A0N(n2379), .A1N(selectBit_EAST), .B0(n2901), .Y(n2897)
         );
  INVX2TS U560 ( .A(n1023), .Y(n490) );
  CLKBUFX2TS U561 ( .A(n2031), .Y(n650) );
  INVX2TS U562 ( .A(n650), .Y(n491) );
  INVX2TS U563 ( .A(n650), .Y(n492) );
  CLKBUFX2TS U564 ( .A(n2029), .Y(n651) );
  INVX2TS U565 ( .A(n651), .Y(n493) );
  INVX2TS U566 ( .A(n651), .Y(n494) );
  CLKBUFX2TS U567 ( .A(cacheDataOut[28]), .Y(n495) );
  CLKBUFX2TS U568 ( .A(cacheDataOut[28]), .Y(n496) );
  CLKBUFX2TS U569 ( .A(cacheDataOut[27]), .Y(n497) );
  CLKBUFX2TS U570 ( .A(cacheDataOut[27]), .Y(n498) );
  CLKBUFX2TS U571 ( .A(cacheDataOut[23]), .Y(n499) );
  CLKBUFX2TS U572 ( .A(cacheDataOut[23]), .Y(n500) );
  CLKBUFX2TS U573 ( .A(cacheDataOut[20]), .Y(n501) );
  CLKBUFX2TS U574 ( .A(cacheDataOut[20]), .Y(n502) );
  CLKBUFX2TS U575 ( .A(cacheDataOut[9]), .Y(n503) );
  CLKBUFX2TS U576 ( .A(cacheDataOut[9]), .Y(n504) );
  CLKBUFX2TS U577 ( .A(cacheDataOut[5]), .Y(n505) );
  CLKBUFX2TS U578 ( .A(cacheDataOut[5]), .Y(n506) );
  CLKBUFX2TS U579 ( .A(cacheDataOut[2]), .Y(n507) );
  CLKBUFX2TS U580 ( .A(cacheDataOut[2]), .Y(n508) );
  CLKBUFX2TS U581 ( .A(cacheDataOut[31]), .Y(n509) );
  CLKBUFX2TS U582 ( .A(cacheDataOut[31]), .Y(n510) );
  CLKBUFX2TS U583 ( .A(cacheDataOut[30]), .Y(n511) );
  CLKBUFX2TS U584 ( .A(cacheDataOut[30]), .Y(n512) );
  CLKBUFX2TS U585 ( .A(cacheDataOut[29]), .Y(n513) );
  CLKBUFX2TS U586 ( .A(cacheDataOut[29]), .Y(n514) );
  CLKBUFX2TS U587 ( .A(cacheDataOut[26]), .Y(n515) );
  CLKBUFX2TS U588 ( .A(cacheDataOut[26]), .Y(n516) );
  CLKBUFX2TS U589 ( .A(cacheDataOut[25]), .Y(n517) );
  CLKBUFX2TS U590 ( .A(cacheDataOut[25]), .Y(n518) );
  CLKBUFX2TS U591 ( .A(cacheDataOut[24]), .Y(n519) );
  CLKBUFX2TS U592 ( .A(cacheDataOut[24]), .Y(n520) );
  CLKBUFX2TS U593 ( .A(cacheDataOut[22]), .Y(n521) );
  CLKBUFX2TS U594 ( .A(cacheDataOut[22]), .Y(n522) );
  CLKBUFX2TS U595 ( .A(cacheDataOut[21]), .Y(n523) );
  CLKBUFX2TS U596 ( .A(cacheDataOut[21]), .Y(n524) );
  CLKBUFX2TS U597 ( .A(cacheDataOut[19]), .Y(n525) );
  CLKBUFX2TS U598 ( .A(cacheDataOut[19]), .Y(n526) );
  CLKBUFX2TS U599 ( .A(cacheDataOut[18]), .Y(n527) );
  CLKBUFX2TS U600 ( .A(cacheDataOut[18]), .Y(n528) );
  CLKBUFX2TS U601 ( .A(cacheDataOut[17]), .Y(n529) );
  CLKBUFX2TS U602 ( .A(cacheDataOut[17]), .Y(n530) );
  CLKBUFX2TS U603 ( .A(cacheDataOut[16]), .Y(n531) );
  CLKBUFX2TS U604 ( .A(cacheDataOut[16]), .Y(n532) );
  CLKBUFX2TS U605 ( .A(cacheDataOut[15]), .Y(n533) );
  CLKBUFX2TS U606 ( .A(cacheDataOut[15]), .Y(n534) );
  CLKBUFX2TS U607 ( .A(cacheDataOut[14]), .Y(n535) );
  CLKBUFX2TS U608 ( .A(cacheDataOut[14]), .Y(n536) );
  CLKBUFX2TS U609 ( .A(cacheDataOut[13]), .Y(n537) );
  CLKBUFX2TS U610 ( .A(cacheDataOut[13]), .Y(n538) );
  CLKBUFX2TS U611 ( .A(cacheDataOut[12]), .Y(n539) );
  CLKBUFX2TS U612 ( .A(cacheDataOut[12]), .Y(n540) );
  CLKBUFX2TS U613 ( .A(cacheDataOut[11]), .Y(n541) );
  CLKBUFX2TS U614 ( .A(cacheDataOut[11]), .Y(n542) );
  CLKBUFX2TS U615 ( .A(cacheDataOut[10]), .Y(n543) );
  CLKBUFX2TS U616 ( .A(cacheDataOut[10]), .Y(n544) );
  CLKBUFX2TS U617 ( .A(cacheDataOut[8]), .Y(n545) );
  CLKBUFX2TS U618 ( .A(cacheDataOut[8]), .Y(n546) );
  CLKBUFX2TS U619 ( .A(cacheDataOut[7]), .Y(n547) );
  CLKBUFX2TS U620 ( .A(cacheDataOut[7]), .Y(n548) );
  CLKBUFX2TS U621 ( .A(cacheDataOut[6]), .Y(n549) );
  CLKBUFX2TS U622 ( .A(cacheDataOut[6]), .Y(n659) );
  CLKBUFX2TS U623 ( .A(cacheDataOut[4]), .Y(n661) );
  CLKBUFX2TS U624 ( .A(cacheDataOut[4]), .Y(n663) );
  CLKBUFX2TS U625 ( .A(cacheDataOut[3]), .Y(n666) );
  CLKBUFX2TS U626 ( .A(cacheDataOut[3]), .Y(n672) );
  CLKBUFX2TS U627 ( .A(cacheDataOut[1]), .Y(n673) );
  CLKBUFX2TS U628 ( .A(cacheDataOut[1]), .Y(n674) );
  CLKBUFX2TS U629 ( .A(cacheDataOut[0]), .Y(n676) );
  CLKBUFX2TS U630 ( .A(cacheDataOut[0]), .Y(n677) );
  CLKBUFX2TS U631 ( .A(n976), .Y(n1754) );
  INVX2TS U632 ( .A(n1754), .Y(n680) );
  INVX2TS U633 ( .A(n1754), .Y(n683) );
  INVX2TS U634 ( .A(n1754), .Y(n687) );
  AND3XLTS U635 ( .A(n101), .B(n163), .C(n1806), .Y(n976) );
  AND2X2TS U636 ( .A(n692), .B(n100), .Y(n1756) );
  INVX2TS U637 ( .A(n1756), .Y(n689) );
  INVX2TS U638 ( .A(n1756), .Y(n701) );
  INVX2TS U639 ( .A(n1756), .Y(n913) );
  AOI21X1TS U640 ( .A0(n945), .A1(n127), .B0(n986), .Y(n1808) );
  INVX2TS U641 ( .A(n1743), .Y(n914) );
  INVX2TS U642 ( .A(n1743), .Y(n938) );
  AND2X2TS U643 ( .A(n487), .B(n691), .Y(n1748) );
  INVX2TS U644 ( .A(n1748), .Y(n941) );
  INVX2TS U645 ( .A(n1748), .Y(n949) );
  INVXLTS U646 ( .A(n1748), .Y(n950) );
  AOI21X1TS U647 ( .A0(n943), .A1(n700), .B0(n681), .Y(n1786) );
  INVX2TS U648 ( .A(n1745), .Y(n952) );
  INVX2TS U649 ( .A(n1745), .Y(n956) );
  INVXLTS U650 ( .A(n1745), .Y(n957) );
  INVXLTS U651 ( .A(n3920), .Y(n958) );
  INVXLTS U652 ( .A(n3922), .Y(n959) );
  OAI22X1TS U653 ( .A0(n685), .A1(n179), .B0(n1865), .B1(n1933), .Y(n1752) );
  CLKINVX2TS U654 ( .A(n1799), .Y(n685) );
  CLKBUFX2TS U655 ( .A(n5323), .Y(n960) );
  OAI32X1TS U656 ( .A0(n2011), .A1(n118), .A2(n195), .B0(n989), .B1(n953), .Y(
        n2010) );
  XOR2X1TS U657 ( .A(n2009), .B(n960), .Y(n2007) );
  AND2XLTS U658 ( .A(n1767), .B(n671), .Y(n1113) );
  CLKINVX2TS U659 ( .A(n1113), .Y(n961) );
  INVXLTS U660 ( .A(n1113), .Y(n962) );
  INVXLTS U661 ( .A(n1113), .Y(n963) );
  INVXLTS U662 ( .A(n1113), .Y(n966) );
  INVX2TS U663 ( .A(n2008), .Y(n969) );
  NAND3X1TS U664 ( .A(n944), .B(n972), .C(n1888), .Y(n1775) );
  CLKINVX2TS U665 ( .A(n968), .Y(n973) );
  INVXLTS U666 ( .A(n973), .Y(n975) );
  NAND3XLTS U667 ( .A(n944), .B(n972), .C(n1841), .Y(n1761) );
  CLKBUFX2TS U668 ( .A(n2379), .Y(n977) );
  INVX2TS U669 ( .A(n3548), .Y(n3534) );
  INVX2TS U670 ( .A(n3548), .Y(n3535) );
  INVX2TS U671 ( .A(n3549), .Y(n3536) );
  INVX2TS U672 ( .A(n3549), .Y(n3537) );
  INVX2TS U673 ( .A(n3549), .Y(n3538) );
  INVX2TS U674 ( .A(n3548), .Y(n3540) );
  INVX2TS U675 ( .A(n3548), .Y(n3541) );
  INVX2TS U676 ( .A(n3550), .Y(n3539) );
  INVX1TS U677 ( .A(n1956), .Y(n684) );
  CLKBUFX2TS U678 ( .A(n955), .Y(n978) );
  OR2X1TS U679 ( .A(n2379), .B(n974), .Y(n980) );
  INVX1TS U680 ( .A(n2009), .Y(n953) );
  NAND2XLTS U681 ( .A(n2009), .B(n2900), .Y(n2385) );
  OAI21XLTS U682 ( .A0(n2009), .A1(n2900), .B0(n2385), .Y(n2890) );
  NOR2X1TS U683 ( .A(n489), .B(n467), .Y(n2011) );
  INVX2TS U684 ( .A(n1793), .Y(n691) );
  NAND2XLTS U685 ( .A(n180), .B(n4606), .Y(n1082) );
  NAND2X1TS U686 ( .A(n678), .B(n194), .Y(n1865) );
  NAND3XLTS U687 ( .A(n116), .B(n699), .C(n1888), .Y(n1805) );
  NAND2XLTS U688 ( .A(selectBit_EAST), .B(n1910), .Y(n1956) );
  INVXLTS U689 ( .A(n1923), .Y(n682) );
  AOI21X1TS U690 ( .A0(n943), .A1(n127), .B0(n985), .Y(n1802) );
  NOR3XLTS U691 ( .A(n1783), .B(n1782), .C(n1785), .Y(n1151) );
  NOR2BXLTS U692 ( .AN(n1826), .B(n128), .Y(n1197) );
  NOR2XLTS U693 ( .A(n1863), .B(n1770), .Y(n1118) );
  NOR2BXLTS U694 ( .AN(n1802), .B(n1805), .Y(n1198) );
  NAND2XLTS U695 ( .A(n678), .B(n4606), .Y(n1081) );
  OA22X1TS U696 ( .A0(n1806), .A1(n178), .B0(n1837), .B1(n1971), .Y(n985) );
  NOR2BXLTS U697 ( .AN(n1826), .B(n1827), .Y(n1099) );
  NOR2BXLTS U698 ( .AN(n1826), .B(n130), .Y(n1133) );
  NAND2XLTS U699 ( .A(readReady), .B(n9), .Y(n1836) );
  INVXLTS U700 ( .A(selectBit_WEST), .Y(n1023) );
  XOR2XLTS U701 ( .A(n1078), .B(n490), .Y(n2896) );
  NAND2XLTS U702 ( .A(n470), .B(n195), .Y(n1864) );
  NAND2XLTS U703 ( .A(selectBit_WEST), .B(readReady), .Y(n2898) );
  INVXLTS U704 ( .A(readReady), .Y(n1078) );
  INVXLTS U705 ( .A(n3482), .Y(n3477) );
  INVXLTS U706 ( .A(n3430), .Y(n3425) );
  INVXLTS U707 ( .A(n3481), .Y(n3478) );
  INVXLTS U708 ( .A(n3429), .Y(n3426) );
  INVXLTS U709 ( .A(n3480), .Y(n3479) );
  INVXLTS U710 ( .A(n3428), .Y(n3427) );
  INVXLTS U711 ( .A(n3547), .Y(n3542) );
  INVXLTS U712 ( .A(n3546), .Y(n3543) );
  INVXLTS U713 ( .A(n3545), .Y(n3544) );
  INVX1TS U714 ( .A(n479), .Y(n669) );
  INVXLTS U715 ( .A(n3199), .Y(n3186) );
  INVXLTS U716 ( .A(n3282), .Y(n3279) );
  INVXLTS U717 ( .A(n986), .Y(n3280) );
  CLKBUFX2TS U718 ( .A(n3202), .Y(n3197) );
  CLKBUFX2TS U719 ( .A(n3202), .Y(n3196) );
  CLKBUFX2TS U720 ( .A(n3201), .Y(n3198) );
  CLKBUFX2TS U721 ( .A(n3285), .Y(n3282) );
  CLKBUFX2TS U722 ( .A(n3285), .Y(n3283) );
  AND3XLTS U723 ( .A(n1789), .B(n1790), .C(n1786), .Y(n1165) );
  CLKINVX2TS U724 ( .A(n1801), .Y(n688) );
  INVX1TS U725 ( .A(n1177), .Y(n3434) );
  NAND3BXLTS U726 ( .AN(n1798), .B(n102), .C(n1800), .Y(n1177) );
  CLKBUFX2TS U727 ( .A(n3633), .Y(n3630) );
  CLKBUFX2TS U728 ( .A(n3368), .Y(n3365) );
  CLKBUFX2TS U729 ( .A(n3633), .Y(n3631) );
  CLKBUFX2TS U730 ( .A(n3368), .Y(n3366) );
  INVXLTS U731 ( .A(n1763), .Y(n690) );
  CLKBUFX2TS U732 ( .A(n3120), .Y(n3116) );
  OAI31XLTS U733 ( .A0(n120), .A1(n108), .A2(n943), .B0(n678), .Y(n1837) );
  NAND2XLTS U734 ( .A(n1789), .B(n1839), .Y(n1760) );
  OAI21XLTS U735 ( .A0(n120), .A1(n126), .B0(n162), .Y(n1958) );
  NOR2BXLTS U736 ( .AN(n1802), .B(n162), .Y(n1196) );
  NOR2BXLTS U737 ( .AN(n104), .B(n163), .Y(n1132) );
  NOR2BXLTS U738 ( .AN(n104), .B(n1775), .Y(n1135) );
  NOR2XLTS U739 ( .A(n1763), .B(n1764), .Y(n1098) );
  NOR2XLTS U740 ( .A(n1761), .B(n488), .Y(n1101) );
  NOR3XLTS U741 ( .A(n1784), .B(n946), .C(n1785), .Y(n1149) );
  NOR3BX1TS U742 ( .AN(n1808), .B(n1813), .C(n117), .Y(n1216) );
  OR4XLTS U743 ( .A(n488), .B(n686), .C(n698), .D(n690), .Y(n982) );
  AND3XLTS U744 ( .A(n1774), .B(n1805), .C(n1802), .Y(n1199) );
  CLKINVX2TS U745 ( .A(n2), .Y(n681) );
  AND2XLTS U746 ( .A(n1782), .B(n667), .Y(n983) );
  XNOR2X1TS U747 ( .A(n195), .B(n118), .Y(n1866) );
  NAND3XLTS U748 ( .A(n2378), .B(n974), .C(n2379), .Y(n2045) );
  OAI22XLTS U749 ( .A0(n110), .A1(n964), .B0(n691), .B1(n138), .Y(n1792) );
  NAND2XLTS U750 ( .A(n4206), .B(n696), .Y(n1787) );
  AOI32XLTS U751 ( .A0(n1789), .A1(n1790), .A2(n4212), .B0(n1791), .B1(n1792), 
        .Y(n1788) );
  OAI21XLTS U752 ( .A0(n2378), .A1(n119), .B0(n2898), .Y(n2900) );
  AOI21XLTS U753 ( .A0(n1), .A1(n2005), .B0(n2001), .Y(n1935) );
  AOI32XLTS U754 ( .A0(n101), .A1(n1803), .A2(n1804), .B0(n3367), .B1(n601), 
        .Y(n2564) );
  NAND2XLTS U755 ( .A(n4206), .B(n693), .Y(n1803) );
  AOI32XLTS U756 ( .A0(n132), .A1(n1805), .A2(n4212), .B0(n1806), .B1(n1777), 
        .Y(n1804) );
  AOI32XLTS U757 ( .A0(n104), .A1(n1772), .A2(n1773), .B0(n3630), .B1(n600), 
        .Y(n2568) );
  NAND2XLTS U758 ( .A(n4206), .B(n694), .Y(n1772) );
  AOI32XLTS U759 ( .A0(n1774), .A1(n1775), .A2(n4212), .B0(n1776), .B1(n1777), 
        .Y(n1773) );
  AOI22XLTS U760 ( .A0(n1763), .A1(n964), .B0(n690), .B1(n137), .Y(n1762) );
  NAND2X1TS U761 ( .A(n989), .B(n121), .Y(n1971) );
  NAND2XLTS U762 ( .A(readIn_SOUTH), .B(n1801), .Y(n1795) );
  OAI211XLTS U763 ( .A0(n966), .A1(n3956), .B0(n1844), .C0(n1845), .Y(n2547)
         );
  OAI211XLTS U764 ( .A0(n963), .A1(n3953), .B0(n1842), .C0(n1843), .Y(n2548)
         );
  OAI211XLTS U765 ( .A0(n962), .A1(n3965), .B0(n1850), .C0(n1851), .Y(n2544)
         );
  OAI211XLTS U766 ( .A0(n966), .A1(n3968), .B0(n1852), .C0(n1853), .Y(n2543)
         );
  OAI211XLTS U767 ( .A0(n963), .A1(n3962), .B0(n1848), .C0(n1849), .Y(n2545)
         );
  OAI211XLTS U768 ( .A0(n962), .A1(n3959), .B0(n1846), .C0(n1847), .Y(n2546)
         );
  OAI211XLTS U769 ( .A0(n4199), .A1(n966), .B0(n1125), .C0(n1126), .Y(n2872)
         );
  OAI211XLTS U770 ( .A0(n4196), .A1(n963), .B0(n1123), .C0(n1124), .Y(n2873)
         );
  OAI211XLTS U771 ( .A0(n4193), .A1(n963), .B0(n1121), .C0(n1122), .Y(n2874)
         );
  OAI211XLTS U772 ( .A0(n4190), .A1(n962), .B0(n1119), .C0(n1120), .Y(n2875)
         );
  OAI211XLTS U773 ( .A0(n4187), .A1(n962), .B0(n1114), .C0(n1115), .Y(n2876)
         );
  OAI211XLTS U774 ( .A0(n4202), .A1(n966), .B0(n1127), .C0(n1128), .Y(n2871)
         );
  OAI211XLTS U775 ( .A0(n3618), .A1(n743), .B0(n1877), .C0(n1878), .Y(n2529)
         );
  OAI211XLTS U776 ( .A0(n3187), .A1(n919), .B0(n1674), .C0(n1675), .Y(n2611)
         );
  OAI211XLTS U777 ( .A0(n3187), .A1(n792), .B0(n1672), .C0(n1673), .Y(n2612)
         );
  OAI211XLTS U778 ( .A0(n3353), .A1(n820), .B0(n1969), .C0(n1970), .Y(n2473)
         );
  OAI211XLTS U779 ( .A0(n3353), .A1(n896), .B0(n1204), .C0(n1205), .Y(n2843)
         );
  OAI211XLTS U780 ( .A0(n3353), .A1(n894), .B0(n1200), .C0(n1201), .Y(n2845)
         );
  OAI211XLTS U781 ( .A0(n3270), .A1(n596), .B0(n1221), .C0(n1222), .Y(n2837)
         );
  OAI211XLTS U782 ( .A0(n3270), .A1(n594), .B0(n1219), .C0(n1220), .Y(n2838)
         );
  OAI211XLTS U783 ( .A0(n3270), .A1(n593), .B0(n1217), .C0(n1218), .Y(n2839)
         );
  OAI211XLTS U784 ( .A0(n3618), .A1(n886), .B0(n1140), .C0(n1141), .Y(n2867)
         );
  OAI211XLTS U785 ( .A0(n3618), .A1(n884), .B0(n1136), .C0(n1137), .Y(n2869)
         );
  OAI211XLTS U786 ( .A0(n3543), .A1(n4266), .B0(n1485), .C0(n1486), .Y(n2705)
         );
  OAI211XLTS U787 ( .A0(n3543), .A1(n4263), .B0(n1483), .C0(n1484), .Y(n2706)
         );
  OAI211XLTS U788 ( .A0(n3478), .A1(n4266), .B0(n1421), .C0(n1422), .Y(n2737)
         );
  OAI211XLTS U789 ( .A0(n3478), .A1(n4263), .B0(n1419), .C0(n1420), .Y(n2738)
         );
  OAI211XLTS U790 ( .A0(n3426), .A1(n4362), .B0(n1357), .C0(n1358), .Y(n2769)
         );
  OAI211XLTS U791 ( .A0(n3426), .A1(n4359), .B0(n1355), .C0(n1356), .Y(n2770)
         );
  OAI211XLTS U792 ( .A0(n3274), .A1(n614), .B0(n1981), .C0(n1982), .Y(n2464)
         );
  OAI211XLTS U793 ( .A0(n3534), .A1(n4007), .B0(n1897), .C0(n1898), .Y(n2516)
         );
  OAI211XLTS U794 ( .A0(n3534), .A1(n4010), .B0(n1899), .C0(n1900), .Y(n2515)
         );
  OAI211XLTS U795 ( .A0(n3534), .A1(n4004), .B0(n1895), .C0(n1896), .Y(n2517)
         );
  OAI211XLTS U796 ( .A0(n3534), .A1(n4001), .B0(n1893), .C0(n1894), .Y(n2518)
         );
  OAI211XLTS U797 ( .A0(n3535), .A1(n3998), .B0(n1891), .C0(n1892), .Y(n2519)
         );
  OAI211XLTS U798 ( .A0(n3535), .A1(n3995), .B0(n1889), .C0(n1890), .Y(n2520)
         );
  OAI211XLTS U799 ( .A0(n3535), .A1(n4353), .B0(n1543), .C0(n1544), .Y(n2676)
         );
  OAI211XLTS U800 ( .A0(n3536), .A1(n4347), .B0(n1539), .C0(n1540), .Y(n2678)
         );
  OAI211XLTS U801 ( .A0(n3536), .A1(n4344), .B0(n1537), .C0(n1538), .Y(n2679)
         );
  OAI211XLTS U802 ( .A0(n3536), .A1(n4341), .B0(n1535), .C0(n1536), .Y(n2680)
         );
  OAI211XLTS U803 ( .A0(n3537), .A1(n4338), .B0(n1533), .C0(n1534), .Y(n2681)
         );
  OAI211XLTS U804 ( .A0(n3537), .A1(n4335), .B0(n1531), .C0(n1532), .Y(n2682)
         );
  OAI211XLTS U805 ( .A0(n3537), .A1(n4332), .B0(n1529), .C0(n1530), .Y(n2683)
         );
  OAI211XLTS U806 ( .A0(n3538), .A1(n4317), .B0(n1519), .C0(n1520), .Y(n2688)
         );
  OAI211XLTS U807 ( .A0(n3540), .A1(n4302), .B0(n1509), .C0(n1510), .Y(n2693)
         );
  OAI211XLTS U808 ( .A0(n3541), .A1(n4290), .B0(n1501), .C0(n1502), .Y(n2697)
         );
  OAI211XLTS U809 ( .A0(n3541), .A1(n4284), .B0(n1497), .C0(n1498), .Y(n2699)
         );
  OAI211XLTS U810 ( .A0(n3542), .A1(n4278), .B0(n1493), .C0(n1494), .Y(n2701)
         );
  OAI211XLTS U811 ( .A0(n3542), .A1(n4275), .B0(n1491), .C0(n1492), .Y(n2702)
         );
  OAI211XLTS U812 ( .A0(n3542), .A1(n4269), .B0(n1487), .C0(n1488), .Y(n2704)
         );
  OAI211XLTS U813 ( .A0(n3535), .A1(n4356), .B0(n1545), .C0(n1546), .Y(n2675)
         );
  OAI211XLTS U814 ( .A0(n3536), .A1(n4350), .B0(n1541), .C0(n1542), .Y(n2677)
         );
  OAI211XLTS U815 ( .A0(n3537), .A1(n4329), .B0(n1527), .C0(n1528), .Y(n2684)
         );
  OAI211XLTS U816 ( .A0(n3538), .A1(n4326), .B0(n1525), .C0(n1526), .Y(n2685)
         );
  OAI211XLTS U817 ( .A0(n3538), .A1(n4323), .B0(n1523), .C0(n1524), .Y(n2686)
         );
  OAI211XLTS U818 ( .A0(n3538), .A1(n4320), .B0(n1521), .C0(n1522), .Y(n2687)
         );
  OAI211XLTS U819 ( .A0(n3539), .A1(n4311), .B0(n1515), .C0(n1516), .Y(n2690)
         );
  OAI211XLTS U820 ( .A0(n3540), .A1(n4299), .B0(n1507), .C0(n1508), .Y(n2694)
         );
  OAI211XLTS U821 ( .A0(n3540), .A1(n4296), .B0(n1505), .C0(n1506), .Y(n2695)
         );
  OAI211XLTS U822 ( .A0(n3540), .A1(n4293), .B0(n1503), .C0(n1504), .Y(n2696)
         );
  OAI211XLTS U823 ( .A0(n3541), .A1(n4287), .B0(n1499), .C0(n1500), .Y(n2698)
         );
  OAI211XLTS U824 ( .A0(n3541), .A1(n4281), .B0(n1495), .C0(n1496), .Y(n2700)
         );
  OAI211XLTS U825 ( .A0(n3539), .A1(n4314), .B0(n1517), .C0(n1518), .Y(n2689)
         );
  OAI211XLTS U826 ( .A0(n3539), .A1(n4308), .B0(n1513), .C0(n1514), .Y(n2691)
         );
  OAI211XLTS U827 ( .A0(n3539), .A1(n4305), .B0(n1511), .C0(n1512), .Y(n2692)
         );
  OAI211XLTS U828 ( .A0(n3542), .A1(n4272), .B0(n1489), .C0(n1490), .Y(n2703)
         );
  OAI211XLTS U829 ( .A0(n3470), .A1(n3998), .B0(n1913), .C0(n1914), .Y(n2505)
         );
  OAI211XLTS U830 ( .A0(n3470), .A1(n3995), .B0(n1911), .C0(n1912), .Y(n2506)
         );
  OAI211XLTS U831 ( .A0(n3470), .A1(n4356), .B0(n1481), .C0(n1482), .Y(n2707)
         );
  OAI211XLTS U832 ( .A0(n3470), .A1(n4353), .B0(n1479), .C0(n1480), .Y(n2708)
         );
  OAI211XLTS U833 ( .A0(n3471), .A1(n4350), .B0(n1477), .C0(n1478), .Y(n2709)
         );
  OAI211XLTS U834 ( .A0(n3471), .A1(n4347), .B0(n1475), .C0(n1476), .Y(n2710)
         );
  OAI211XLTS U835 ( .A0(n3471), .A1(n4344), .B0(n1473), .C0(n1474), .Y(n2711)
         );
  OAI211XLTS U836 ( .A0(n3471), .A1(n4341), .B0(n1471), .C0(n1472), .Y(n2712)
         );
  OAI211XLTS U837 ( .A0(n3472), .A1(n4335), .B0(n1467), .C0(n1468), .Y(n2714)
         );
  OAI211XLTS U838 ( .A0(n3472), .A1(n4329), .B0(n1463), .C0(n1464), .Y(n2716)
         );
  OAI211XLTS U839 ( .A0(n3473), .A1(n4326), .B0(n1461), .C0(n1462), .Y(n2717)
         );
  OAI211XLTS U840 ( .A0(n3473), .A1(n4320), .B0(n1457), .C0(n1458), .Y(n2719)
         );
  OAI211XLTS U841 ( .A0(n3474), .A1(n4314), .B0(n1453), .C0(n1454), .Y(n2721)
         );
  OAI211XLTS U842 ( .A0(n3474), .A1(n4311), .B0(n1451), .C0(n1452), .Y(n2722)
         );
  OAI211XLTS U843 ( .A0(n3474), .A1(n4305), .B0(n1447), .C0(n1448), .Y(n2724)
         );
  OAI211XLTS U844 ( .A0(n3475), .A1(n4299), .B0(n1443), .C0(n1444), .Y(n2726)
         );
  OAI211XLTS U845 ( .A0(n3475), .A1(n4296), .B0(n1441), .C0(n1442), .Y(n2727)
         );
  OAI211XLTS U846 ( .A0(n3475), .A1(n4293), .B0(n1439), .C0(n1440), .Y(n2728)
         );
  OAI211XLTS U847 ( .A0(n3476), .A1(n4290), .B0(n1437), .C0(n1438), .Y(n2729)
         );
  OAI211XLTS U848 ( .A0(n3476), .A1(n4287), .B0(n1435), .C0(n1436), .Y(n2730)
         );
  OAI211XLTS U849 ( .A0(n3476), .A1(n4281), .B0(n1431), .C0(n1432), .Y(n2732)
         );
  OAI211XLTS U850 ( .A0(n3477), .A1(n4272), .B0(n1425), .C0(n1426), .Y(n2735)
         );
  OAI211XLTS U851 ( .A0(n3472), .A1(n4338), .B0(n1469), .C0(n1470), .Y(n2713)
         );
  OAI211XLTS U852 ( .A0(n3472), .A1(n4332), .B0(n1465), .C0(n1466), .Y(n2715)
         );
  OAI211XLTS U853 ( .A0(n3473), .A1(n4323), .B0(n1459), .C0(n1460), .Y(n2718)
         );
  OAI211XLTS U854 ( .A0(n3473), .A1(n4317), .B0(n1455), .C0(n1456), .Y(n2720)
         );
  OAI211XLTS U855 ( .A0(n3474), .A1(n4308), .B0(n1449), .C0(n1450), .Y(n2723)
         );
  OAI211XLTS U856 ( .A0(n3475), .A1(n4302), .B0(n1445), .C0(n1446), .Y(n2725)
         );
  OAI211XLTS U857 ( .A0(n3477), .A1(n4278), .B0(n1429), .C0(n1430), .Y(n2733)
         );
  OAI211XLTS U858 ( .A0(n3477), .A1(n4275), .B0(n1427), .C0(n1428), .Y(n2734)
         );
  OAI211XLTS U859 ( .A0(n3477), .A1(n4269), .B0(n1423), .C0(n1424), .Y(n2736)
         );
  OAI211XLTS U860 ( .A0(n3476), .A1(n4284), .B0(n1433), .C0(n1434), .Y(n2731)
         );
  OAI211XLTS U861 ( .A0(n3469), .A1(n4010), .B0(n1921), .C0(n1922), .Y(n2501)
         );
  OAI211XLTS U862 ( .A0(n3469), .A1(n4007), .B0(n1919), .C0(n1920), .Y(n2502)
         );
  OAI211XLTS U863 ( .A0(n3469), .A1(n4004), .B0(n1917), .C0(n1918), .Y(n2503)
         );
  OAI211XLTS U864 ( .A0(n3469), .A1(n4001), .B0(n1915), .C0(n1916), .Y(n2504)
         );
  OAI211XLTS U865 ( .A0(n3417), .A1(n3959), .B0(n1940), .C0(n1941), .Y(n2490)
         );
  OAI211XLTS U866 ( .A0(n3417), .A1(n3965), .B0(n1944), .C0(n1945), .Y(n2488)
         );
  OAI211XLTS U867 ( .A0(n3417), .A1(n3962), .B0(n1942), .C0(n1943), .Y(n2489)
         );
  OAI211XLTS U868 ( .A0(n3417), .A1(n3968), .B0(n1946), .C0(n1947), .Y(n2487)
         );
  OAI211XLTS U869 ( .A0(n3418), .A1(n4457), .B0(n1415), .C0(n1416), .Y(n2740)
         );
  OAI211XLTS U870 ( .A0(n3419), .A1(n4453), .B0(n1413), .C0(n1414), .Y(n2741)
         );
  OAI211XLTS U871 ( .A0(n3419), .A1(n4450), .B0(n1411), .C0(n1412), .Y(n2742)
         );
  OAI211XLTS U872 ( .A0(n3419), .A1(n4442), .B0(n1407), .C0(n1408), .Y(n2744)
         );
  OAI211XLTS U873 ( .A0(n3420), .A1(n4439), .B0(n1405), .C0(n1406), .Y(n2745)
         );
  OAI211XLTS U874 ( .A0(n3420), .A1(n4431), .B0(n1401), .C0(n1402), .Y(n2747)
         );
  OAI211XLTS U875 ( .A0(n3421), .A1(n4424), .B0(n1397), .C0(n1398), .Y(n2749)
         );
  OAI211XLTS U876 ( .A0(n3421), .A1(n4421), .B0(n1395), .C0(n1396), .Y(n2750)
         );
  OAI211XLTS U877 ( .A0(n3421), .A1(n4416), .B0(n1393), .C0(n1394), .Y(n2751)
         );
  OAI211XLTS U878 ( .A0(n3421), .A1(n4413), .B0(n1391), .C0(n1392), .Y(n2752)
         );
  OAI211XLTS U879 ( .A0(n3422), .A1(n4410), .B0(n1389), .C0(n1390), .Y(n2753)
         );
  OAI211XLTS U880 ( .A0(n3422), .A1(n4404), .B0(n1385), .C0(n1386), .Y(n2755)
         );
  OAI211XLTS U881 ( .A0(n3422), .A1(n4401), .B0(n1383), .C0(n1384), .Y(n2756)
         );
  OAI211XLTS U882 ( .A0(n3423), .A1(n4398), .B0(n1381), .C0(n1382), .Y(n2757)
         );
  OAI211XLTS U883 ( .A0(n3423), .A1(n4395), .B0(n1379), .C0(n1380), .Y(n2758)
         );
  OAI211XLTS U884 ( .A0(n3423), .A1(n4392), .B0(n1377), .C0(n1378), .Y(n2759)
         );
  OAI211XLTS U885 ( .A0(n3424), .A1(n4386), .B0(n1373), .C0(n1374), .Y(n2761)
         );
  OAI211XLTS U886 ( .A0(n3424), .A1(n4383), .B0(n1371), .C0(n1372), .Y(n2762)
         );
  OAI211XLTS U887 ( .A0(n3424), .A1(n4380), .B0(n1369), .C0(n1370), .Y(n2763)
         );
  OAI211XLTS U888 ( .A0(n3425), .A1(n4374), .B0(n1365), .C0(n1366), .Y(n2765)
         );
  OAI211XLTS U889 ( .A0(n3425), .A1(n4371), .B0(n1363), .C0(n1364), .Y(n2766)
         );
  OAI211XLTS U890 ( .A0(n3425), .A1(n4368), .B0(n1361), .C0(n1362), .Y(n2767)
         );
  OAI211XLTS U891 ( .A0(n3418), .A1(n3956), .B0(n1938), .C0(n1939), .Y(n2491)
         );
  OAI211XLTS U892 ( .A0(n3418), .A1(n3953), .B0(n1936), .C0(n1937), .Y(n2492)
         );
  OAI211XLTS U893 ( .A0(n3419), .A1(n4447), .B0(n1409), .C0(n1410), .Y(n2743)
         );
  OAI211XLTS U894 ( .A0(n3423), .A1(n4389), .B0(n1375), .C0(n1376), .Y(n2760)
         );
  OAI211XLTS U895 ( .A0(n3418), .A1(n4460), .B0(n1417), .C0(n1418), .Y(n2739)
         );
  OAI211XLTS U896 ( .A0(n3420), .A1(n4435), .B0(n1403), .C0(n1404), .Y(n2746)
         );
  OAI211XLTS U897 ( .A0(n3420), .A1(n4427), .B0(n1399), .C0(n1400), .Y(n2748)
         );
  OAI211XLTS U898 ( .A0(n3422), .A1(n4407), .B0(n1387), .C0(n1388), .Y(n2754)
         );
  OAI211XLTS U899 ( .A0(n3424), .A1(n4377), .B0(n1367), .C0(n1368), .Y(n2764)
         );
  OAI211XLTS U900 ( .A0(n3425), .A1(n4365), .B0(n1359), .C0(n1360), .Y(n2768)
         );
  OAI211XLTS U901 ( .A0(n3624), .A1(n747), .B0(n1579), .C0(n1580), .Y(n2658)
         );
  OAI211XLTS U902 ( .A0(n3623), .A1(n746), .B0(n1577), .C0(n1578), .Y(n2659)
         );
  OAI211XLTS U903 ( .A0(n3622), .A1(n745), .B0(n1569), .C0(n1570), .Y(n2663)
         );
  OAI211XLTS U904 ( .A0(n3620), .A1(n744), .B0(n1549), .C0(n1550), .Y(n2673)
         );
  OAI211XLTS U905 ( .A0(n3626), .A1(n735), .B0(n1601), .C0(n1602), .Y(n2647)
         );
  OAI211XLTS U906 ( .A0(n3626), .A1(n734), .B0(n1599), .C0(n1600), .Y(n2648)
         );
  OAI211XLTS U907 ( .A0(n3626), .A1(n733), .B0(n1597), .C0(n1598), .Y(n2649)
         );
  OAI211XLTS U908 ( .A0(n3626), .A1(n732), .B0(n1595), .C0(n1596), .Y(n2650)
         );
  OAI211XLTS U909 ( .A0(n3625), .A1(n731), .B0(n1593), .C0(n1594), .Y(n2651)
         );
  OAI211XLTS U910 ( .A0(n3625), .A1(n730), .B0(n1591), .C0(n1592), .Y(n2652)
         );
  OAI211XLTS U911 ( .A0(n3625), .A1(n729), .B0(n1589), .C0(n1590), .Y(n2653)
         );
  OAI211XLTS U912 ( .A0(n3625), .A1(n728), .B0(n1587), .C0(n1588), .Y(n2654)
         );
  OAI211XLTS U913 ( .A0(n3624), .A1(n727), .B0(n1585), .C0(n1586), .Y(n2655)
         );
  OAI211XLTS U914 ( .A0(n3624), .A1(n726), .B0(n1583), .C0(n1584), .Y(n2656)
         );
  OAI211XLTS U915 ( .A0(n3624), .A1(n725), .B0(n1581), .C0(n1582), .Y(n2657)
         );
  OAI211XLTS U916 ( .A0(n3623), .A1(n724), .B0(n1575), .C0(n1576), .Y(n2660)
         );
  OAI211XLTS U917 ( .A0(n3623), .A1(n723), .B0(n1573), .C0(n1574), .Y(n2661)
         );
  OAI211XLTS U918 ( .A0(n3622), .A1(n722), .B0(n1571), .C0(n1572), .Y(n2662)
         );
  OAI211XLTS U919 ( .A0(n3622), .A1(n721), .B0(n1567), .C0(n1568), .Y(n2664)
         );
  OAI211XLTS U920 ( .A0(n3622), .A1(n720), .B0(n1565), .C0(n1566), .Y(n2665)
         );
  OAI211XLTS U921 ( .A0(n3621), .A1(n719), .B0(n1563), .C0(n1564), .Y(n2666)
         );
  OAI211XLTS U922 ( .A0(n3621), .A1(n718), .B0(n1561), .C0(n1562), .Y(n2667)
         );
  OAI211XLTS U923 ( .A0(n3621), .A1(n717), .B0(n1559), .C0(n1560), .Y(n2668)
         );
  OAI211XLTS U924 ( .A0(n3621), .A1(n716), .B0(n1557), .C0(n1558), .Y(n2669)
         );
  OAI211XLTS U925 ( .A0(n3620), .A1(n715), .B0(n1555), .C0(n1556), .Y(n2670)
         );
  OAI211XLTS U926 ( .A0(n3620), .A1(n714), .B0(n1553), .C0(n1554), .Y(n2671)
         );
  OAI211XLTS U927 ( .A0(n3620), .A1(n713), .B0(n1551), .C0(n1552), .Y(n2672)
         );
  OAI211XLTS U928 ( .A0(n3619), .A1(n712), .B0(n1547), .C0(n1548), .Y(n2674)
         );
  OAI211XLTS U929 ( .A0(n3193), .A1(n937), .B0(n1626), .C0(n1627), .Y(n2635)
         );
  OAI211XLTS U930 ( .A0(n3193), .A1(n936), .B0(n1628), .C0(n1629), .Y(n2634)
         );
  OAI211XLTS U931 ( .A0(n3192), .A1(n935), .B0(n1634), .C0(n1635), .Y(n2631)
         );
  OAI211XLTS U932 ( .A0(n3192), .A1(n934), .B0(n1636), .C0(n1637), .Y(n2630)
         );
  OAI211XLTS U933 ( .A0(n3192), .A1(n933), .B0(n1638), .C0(n1639), .Y(n2629)
         );
  OAI211XLTS U934 ( .A0(n3191), .A1(n932), .B0(n1642), .C0(n1643), .Y(n2627)
         );
  OAI211XLTS U935 ( .A0(n3191), .A1(n931), .B0(n1644), .C0(n1645), .Y(n2626)
         );
  OAI211XLTS U936 ( .A0(n3191), .A1(n930), .B0(n1646), .C0(n1647), .Y(n2625)
         );
  OAI211XLTS U937 ( .A0(n3190), .A1(n929), .B0(n1650), .C0(n1651), .Y(n2623)
         );
  OAI211XLTS U938 ( .A0(n3190), .A1(n928), .B0(n1652), .C0(n1653), .Y(n2622)
         );
  OAI211XLTS U939 ( .A0(n3190), .A1(n927), .B0(n1654), .C0(n1655), .Y(n2621)
         );
  OAI211XLTS U940 ( .A0(n3189), .A1(n926), .B0(n1656), .C0(n1657), .Y(n2620)
         );
  OAI211XLTS U941 ( .A0(n3189), .A1(n925), .B0(n1658), .C0(n1659), .Y(n2619)
         );
  OAI211XLTS U942 ( .A0(n3189), .A1(n924), .B0(n1660), .C0(n1661), .Y(n2618)
         );
  OAI211XLTS U943 ( .A0(n3189), .A1(n923), .B0(n1662), .C0(n1663), .Y(n2617)
         );
  OAI211XLTS U944 ( .A0(n3188), .A1(n922), .B0(n1664), .C0(n1665), .Y(n2616)
         );
  OAI211XLTS U945 ( .A0(n3188), .A1(n921), .B0(n1666), .C0(n1667), .Y(n2615)
         );
  OAI211XLTS U946 ( .A0(n3188), .A1(n920), .B0(n1670), .C0(n1671), .Y(n2613)
         );
  OAI211XLTS U947 ( .A0(n3192), .A1(n824), .B0(n1632), .C0(n1633), .Y(n2632)
         );
  OAI211XLTS U948 ( .A0(n3193), .A1(n823), .B0(n1624), .C0(n1625), .Y(n2636)
         );
  OAI211XLTS U949 ( .A0(n3188), .A1(n791), .B0(n1668), .C0(n1669), .Y(n2614)
         );
  OAI211XLTS U950 ( .A0(n3191), .A1(n790), .B0(n1640), .C0(n1641), .Y(n2628)
         );
  OAI211XLTS U951 ( .A0(n3193), .A1(n789), .B0(n1630), .C0(n1631), .Y(n2633)
         );
  OAI211XLTS U952 ( .A0(n3194), .A1(n788), .B0(n1622), .C0(n1623), .Y(n2637)
         );
  OAI211XLTS U953 ( .A0(n3190), .A1(n751), .B0(n1648), .C0(n1649), .Y(n2624)
         );
  OAI211XLTS U954 ( .A0(n3194), .A1(n750), .B0(n1620), .C0(n1621), .Y(n2638)
         );
  OAI211XLTS U955 ( .A0(n3194), .A1(n787), .B0(n1618), .C0(n1619), .Y(n2639)
         );
  OAI211XLTS U956 ( .A0(n3194), .A1(n786), .B0(n1616), .C0(n1617), .Y(n2640)
         );
  OAI211XLTS U957 ( .A0(n3361), .A1(n832), .B0(n1345), .C0(n1346), .Y(n2775)
         );
  OAI211XLTS U958 ( .A0(n3360), .A1(n831), .B0(n1335), .C0(n1336), .Y(n2780)
         );
  OAI211XLTS U959 ( .A0(n3360), .A1(n830), .B0(n1331), .C0(n1332), .Y(n2782)
         );
  OAI211XLTS U960 ( .A0(n3359), .A1(n829), .B0(n1329), .C0(n1330), .Y(n2783)
         );
  OAI211XLTS U961 ( .A0(n3357), .A1(n828), .B0(n1311), .C0(n1312), .Y(n2792)
         );
  OAI211XLTS U962 ( .A0(n3356), .A1(n827), .B0(n1307), .C0(n1308), .Y(n2794)
         );
  OAI211XLTS U963 ( .A0(n3356), .A1(n826), .B0(n1301), .C0(n1302), .Y(n2797)
         );
  OAI211XLTS U964 ( .A0(n3355), .A1(n825), .B0(n1295), .C0(n1296), .Y(n2800)
         );
  OAI211XLTS U965 ( .A0(n3362), .A1(n815), .B0(n1353), .C0(n1354), .Y(n2771)
         );
  OAI211XLTS U966 ( .A0(n3362), .A1(n814), .B0(n1351), .C0(n1352), .Y(n2772)
         );
  OAI211XLTS U967 ( .A0(n3362), .A1(n813), .B0(n1349), .C0(n1350), .Y(n2773)
         );
  OAI211XLTS U968 ( .A0(n3362), .A1(n812), .B0(n1347), .C0(n1348), .Y(n2774)
         );
  OAI211XLTS U969 ( .A0(n3361), .A1(n811), .B0(n1343), .C0(n1344), .Y(n2776)
         );
  OAI211XLTS U970 ( .A0(n3361), .A1(n810), .B0(n1341), .C0(n1342), .Y(n2777)
         );
  OAI211XLTS U971 ( .A0(n3361), .A1(n809), .B0(n1339), .C0(n1340), .Y(n2778)
         );
  OAI211XLTS U972 ( .A0(n3360), .A1(n808), .B0(n1337), .C0(n1338), .Y(n2779)
         );
  OAI211XLTS U973 ( .A0(n3360), .A1(n807), .B0(n1333), .C0(n1334), .Y(n2781)
         );
  OAI211XLTS U974 ( .A0(n3359), .A1(n806), .B0(n1327), .C0(n1328), .Y(n2784)
         );
  OAI211XLTS U975 ( .A0(n3359), .A1(n805), .B0(n1325), .C0(n1326), .Y(n2785)
         );
  OAI211XLTS U976 ( .A0(n3359), .A1(n804), .B0(n1323), .C0(n1324), .Y(n2786)
         );
  OAI211XLTS U977 ( .A0(n3358), .A1(n803), .B0(n1321), .C0(n1322), .Y(n2787)
         );
  OAI211XLTS U978 ( .A0(n3358), .A1(n802), .B0(n1319), .C0(n1320), .Y(n2788)
         );
  OAI211XLTS U979 ( .A0(n3358), .A1(n801), .B0(n1317), .C0(n1318), .Y(n2789)
         );
  OAI211XLTS U980 ( .A0(n3357), .A1(n800), .B0(n1315), .C0(n1316), .Y(n2790)
         );
  OAI211XLTS U981 ( .A0(n3357), .A1(n799), .B0(n1313), .C0(n1314), .Y(n2791)
         );
  OAI211XLTS U982 ( .A0(n3357), .A1(n798), .B0(n1309), .C0(n1310), .Y(n2793)
         );
  OAI211XLTS U983 ( .A0(n3356), .A1(n797), .B0(n1305), .C0(n1306), .Y(n2795)
         );
  OAI211XLTS U984 ( .A0(n3356), .A1(n796), .B0(n1303), .C0(n1304), .Y(n2796)
         );
  OAI211XLTS U985 ( .A0(n3355), .A1(n795), .B0(n1299), .C0(n1300), .Y(n2798)
         );
  OAI211XLTS U986 ( .A0(n3355), .A1(n794), .B0(n1297), .C0(n1298), .Y(n2799)
         );
  OAI211XLTS U987 ( .A0(n3355), .A1(n793), .B0(n1293), .C0(n1294), .Y(n2801)
         );
  OAI211XLTS U988 ( .A0(n3354), .A1(n752), .B0(n1291), .C0(n1292), .Y(n2802)
         );
  OAI211XLTS U989 ( .A0(n3354), .A1(n895), .B0(n1202), .C0(n1203), .Y(n2844)
         );
  OAI211XLTS U990 ( .A0(n3354), .A1(n898), .B0(n1208), .C0(n1209), .Y(n2841)
         );
  OAI211XLTS U991 ( .A0(n3354), .A1(n897), .B0(n1206), .C0(n1207), .Y(n2842)
         );
  OAI211XLTS U992 ( .A0(n3358), .A1(n893), .B0(n1194), .C0(n1195), .Y(n2846)
         );
  OAI211XLTS U993 ( .A0(n3272), .A1(n607), .B0(n1231), .C0(n1232), .Y(n2832)
         );
  OAI211XLTS U994 ( .A0(n3271), .A1(n606), .B0(n1229), .C0(n1230), .Y(n2833)
         );
  OAI211XLTS U995 ( .A0(n3273), .A1(n605), .B0(n1227), .C0(n1228), .Y(n2834)
         );
  OAI211XLTS U996 ( .A0(n3273), .A1(n613), .B0(n1283), .C0(n1284), .Y(n2806)
         );
  OAI211XLTS U997 ( .A0(n3273), .A1(n612), .B0(n1281), .C0(n1282), .Y(n2807)
         );
  OAI211XLTS U998 ( .A0(n3273), .A1(n611), .B0(n1273), .C0(n1274), .Y(n2811)
         );
  OAI211XLTS U999 ( .A0(n3272), .A1(n610), .B0(n1267), .C0(n1268), .Y(n2814)
         );
  OAI211XLTS U1000 ( .A0(n3272), .A1(n609), .B0(n1245), .C0(n1246), .Y(n2825)
         );
  OAI211XLTS U1001 ( .A0(n3272), .A1(n608), .B0(n1237), .C0(n1238), .Y(n2829)
         );
  OAI211XLTS U1002 ( .A0(n3271), .A1(n597), .B0(n1225), .C0(n1226), .Y(n2835)
         );
  OAI211XLTS U1003 ( .A0(n3271), .A1(n595), .B0(n1223), .C0(n1224), .Y(n2836)
         );
  OAI211XLTS U1004 ( .A0(n3271), .A1(n592), .B0(n1211), .C0(n1212), .Y(n2840)
         );
  OAI211XLTS U1005 ( .A0(n3619), .A1(n885), .B0(n1138), .C0(n1139), .Y(n2868)
         );
  OAI211XLTS U1006 ( .A0(n3619), .A1(n888), .B0(n1144), .C0(n1145), .Y(n2865)
         );
  OAI211XLTS U1007 ( .A0(n3619), .A1(n887), .B0(n1142), .C0(n1143), .Y(n2866)
         );
  OAI211XLTS U1008 ( .A0(n3623), .A1(n883), .B0(n1130), .C0(n1131), .Y(n2870)
         );
  OAI211XLTS U1009 ( .A0(n3627), .A1(n748), .B0(n1609), .C0(n1610), .Y(n2643)
         );
  OAI211XLTS U1010 ( .A0(n3627), .A1(n738), .B0(n1607), .C0(n1608), .Y(n2644)
         );
  OAI211XLTS U1011 ( .A0(n3627), .A1(n737), .B0(n1605), .C0(n1606), .Y(n2645)
         );
  OAI211XLTS U1012 ( .A0(n3627), .A1(n736), .B0(n1603), .C0(n1604), .Y(n2646)
         );
  OAI211XLTS U1013 ( .A0(n3363), .A1(n819), .B0(n1965), .C0(n1966), .Y(n2475)
         );
  OAI211XLTS U1014 ( .A0(n3363), .A1(n818), .B0(n1963), .C0(n1964), .Y(n2476)
         );
  OAI211XLTS U1015 ( .A0(n3363), .A1(n817), .B0(n1961), .C0(n1962), .Y(n2477)
         );
  OAI211XLTS U1016 ( .A0(n3363), .A1(n816), .B0(n1959), .C0(n1960), .Y(n2478)
         );
  OAI211XLTS U1017 ( .A0(n3628), .A1(n742), .B0(n1873), .C0(n1874), .Y(n2531)
         );
  OAI211XLTS U1018 ( .A0(n3628), .A1(n741), .B0(n1871), .C0(n1872), .Y(n2532)
         );
  OAI211XLTS U1019 ( .A0(n3628), .A1(n740), .B0(n1869), .C0(n1870), .Y(n2533)
         );
  OAI211XLTS U1020 ( .A0(n3628), .A1(n739), .B0(n1867), .C0(n1868), .Y(n2534)
         );
  OAI211XLTS U1021 ( .A0(n3195), .A1(n822), .B0(n1614), .C0(n1615), .Y(n2641)
         );
  OAI211XLTS U1022 ( .A0(n3195), .A1(n785), .B0(n1612), .C0(n1613), .Y(n2642)
         );
  OAI211XLTS U1023 ( .A0(n4052), .A1(n3543), .B0(n1160), .C0(n1161), .Y(n2859)
         );
  OAI211XLTS U1024 ( .A0(n4049), .A1(n3543), .B0(n1158), .C0(n1159), .Y(n2860)
         );
  OAI211XLTS U1025 ( .A0(n4046), .A1(n3544), .B0(n1156), .C0(n1157), .Y(n2861)
         );
  OAI211XLTS U1026 ( .A0(n4043), .A1(n3544), .B0(n1154), .C0(n1155), .Y(n2862)
         );
  OAI211XLTS U1027 ( .A0(n4040), .A1(n3544), .B0(n1152), .C0(n1153), .Y(n2863)
         );
  OAI211XLTS U1028 ( .A0(n4037), .A1(n3544), .B0(n1147), .C0(n1148), .Y(n2864)
         );
  OAI211XLTS U1029 ( .A0(n4046), .A1(n3479), .B0(n1171), .C0(n1172), .Y(n2855)
         );
  OAI211XLTS U1030 ( .A0(n4043), .A1(n3479), .B0(n1169), .C0(n1170), .Y(n2856)
         );
  OAI211XLTS U1031 ( .A0(n4040), .A1(n3479), .B0(n1167), .C0(n1168), .Y(n2857)
         );
  OAI211XLTS U1032 ( .A0(n4037), .A1(n3479), .B0(n1163), .C0(n1164), .Y(n2858)
         );
  OAI211XLTS U1033 ( .A0(n4049), .A1(n3478), .B0(n1173), .C0(n1174), .Y(n2854)
         );
  OAI211XLTS U1034 ( .A0(n4052), .A1(n3478), .B0(n1175), .C0(n1176), .Y(n2853)
         );
  OAI211XLTS U1035 ( .A0(n4202), .A1(n3426), .B0(n1191), .C0(n1192), .Y(n2847)
         );
  OAI211XLTS U1036 ( .A0(n4190), .A1(n3427), .B0(n1183), .C0(n1184), .Y(n2851)
         );
  OAI211XLTS U1037 ( .A0(n4187), .A1(n3427), .B0(n1178), .C0(n1179), .Y(n2852)
         );
  OAI211XLTS U1038 ( .A0(n4196), .A1(n3427), .B0(n1187), .C0(n1188), .Y(n2849)
         );
  OAI211XLTS U1039 ( .A0(n4193), .A1(n3427), .B0(n1185), .C0(n1186), .Y(n2850)
         );
  OAI211XLTS U1040 ( .A0(n4199), .A1(n3426), .B0(n1189), .C0(n1190), .Y(n2848)
         );
  OAI211XLTS U1041 ( .A0(n3364), .A1(n834), .B0(n1967), .C0(n1968), .Y(n2474)
         );
  INVXLTS U1042 ( .A(n3365), .Y(n3364) );
  OAI211XLTS U1043 ( .A0(n3629), .A1(n711), .B0(n1875), .C0(n1876), .Y(n2530)
         );
  INVXLTS U1044 ( .A(n3632), .Y(n3629) );
  OAI211XLTS U1045 ( .A0(n4712), .A1(n3281), .B0(n1991), .C0(n1992), .Y(n2459)
         );
  INVXLTS U1046 ( .A(n986), .Y(n3281) );
  OAI211XLTS U1047 ( .A0(n3773), .A1(n882), .B0(n1107), .C0(n1108), .Y(n2879)
         );
  OAI211XLTS U1048 ( .A0(n3780), .A1(n881), .B0(n1103), .C0(n1104), .Y(n2881)
         );
  OAI211XLTS U1049 ( .A0(n3775), .A1(n784), .B0(n1824), .C0(n1825), .Y(n2557)
         );
  OAI211XLTS U1050 ( .A0(n3772), .A1(n918), .B0(n1676), .C0(n1677), .Y(n2610)
         );
  OAI211XLTS U1051 ( .A0(n3766), .A1(n917), .B0(n1702), .C0(n1703), .Y(n2597)
         );
  OAI211XLTS U1052 ( .A0(n3766), .A1(n916), .B0(n1704), .C0(n1705), .Y(n2596)
         );
  OAI211XLTS U1053 ( .A0(n3767), .A1(n915), .B0(n1706), .C0(n1707), .Y(n2595)
         );
  OAI211XLTS U1054 ( .A0(n3773), .A1(n891), .B0(n1111), .C0(n1112), .Y(n2877)
         );
  OAI211XLTS U1055 ( .A0(n3777), .A1(n890), .B0(n1109), .C0(n1110), .Y(n2878)
         );
  OAI211XLTS U1056 ( .A0(n3774), .A1(n889), .B0(n1105), .C0(n1106), .Y(n2880)
         );
  OAI211XLTS U1057 ( .A0(n3767), .A1(n880), .B0(n1096), .C0(n1097), .Y(n2882)
         );
  OAI211XLTS U1058 ( .A0(n3771), .A1(n780), .B0(n1738), .C0(n1739), .Y(n2579)
         );
  OAI211XLTS U1059 ( .A0(n3771), .A1(n779), .B0(n1736), .C0(n1737), .Y(n2580)
         );
  OAI211XLTS U1060 ( .A0(n3770), .A1(n778), .B0(n1734), .C0(n1735), .Y(n2581)
         );
  OAI211XLTS U1061 ( .A0(n3770), .A1(n777), .B0(n1732), .C0(n1733), .Y(n2582)
         );
  OAI211XLTS U1062 ( .A0(n3770), .A1(n776), .B0(n1730), .C0(n1731), .Y(n2583)
         );
  OAI211XLTS U1063 ( .A0(n3770), .A1(n775), .B0(n1728), .C0(n1729), .Y(n2584)
         );
  OAI211XLTS U1064 ( .A0(n3769), .A1(n774), .B0(n1726), .C0(n1727), .Y(n2585)
         );
  OAI211XLTS U1065 ( .A0(n3769), .A1(n773), .B0(n1724), .C0(n1725), .Y(n2586)
         );
  OAI211XLTS U1066 ( .A0(n3769), .A1(n772), .B0(n1722), .C0(n1723), .Y(n2587)
         );
  OAI211XLTS U1067 ( .A0(n3769), .A1(n771), .B0(n1720), .C0(n1721), .Y(n2588)
         );
  OAI211XLTS U1068 ( .A0(n3768), .A1(n770), .B0(n1718), .C0(n1719), .Y(n2589)
         );
  OAI211XLTS U1069 ( .A0(n3768), .A1(n769), .B0(n1716), .C0(n1717), .Y(n2590)
         );
  OAI211XLTS U1070 ( .A0(n3768), .A1(n768), .B0(n1714), .C0(n1715), .Y(n2591)
         );
  OAI211XLTS U1071 ( .A0(n3768), .A1(n767), .B0(n1712), .C0(n1713), .Y(n2592)
         );
  OAI211XLTS U1072 ( .A0(n3767), .A1(n766), .B0(n1710), .C0(n1711), .Y(n2593)
         );
  OAI211XLTS U1073 ( .A0(n3767), .A1(n765), .B0(n1708), .C0(n1709), .Y(n2594)
         );
  OAI211XLTS U1074 ( .A0(n3766), .A1(n764), .B0(n1700), .C0(n1701), .Y(n2598)
         );
  OAI211XLTS U1075 ( .A0(n3766), .A1(n763), .B0(n1698), .C0(n1699), .Y(n2599)
         );
  OAI211XLTS U1076 ( .A0(n3765), .A1(n762), .B0(n1696), .C0(n1697), .Y(n2600)
         );
  OAI211XLTS U1077 ( .A0(n3765), .A1(n761), .B0(n1694), .C0(n1695), .Y(n2601)
         );
  OAI211XLTS U1078 ( .A0(n3765), .A1(n760), .B0(n1692), .C0(n1693), .Y(n2602)
         );
  OAI211XLTS U1079 ( .A0(n3765), .A1(n759), .B0(n1690), .C0(n1691), .Y(n2603)
         );
  OAI211XLTS U1080 ( .A0(n3779), .A1(n758), .B0(n1688), .C0(n1689), .Y(n2604)
         );
  OAI211XLTS U1081 ( .A0(n3774), .A1(n757), .B0(n1686), .C0(n1687), .Y(n2605)
         );
  OAI211XLTS U1082 ( .A0(n3775), .A1(n756), .B0(n1684), .C0(n1685), .Y(n2606)
         );
  OAI211XLTS U1083 ( .A0(n3776), .A1(n755), .B0(n1682), .C0(n1683), .Y(n2607)
         );
  OAI211XLTS U1084 ( .A0(n3780), .A1(n754), .B0(n1680), .C0(n1681), .Y(n2608)
         );
  OAI211XLTS U1085 ( .A0(n3780), .A1(n753), .B0(n1678), .C0(n1679), .Y(n2609)
         );
  OAI211XLTS U1086 ( .A0(n3771), .A1(n821), .B0(n1814), .C0(n1815), .Y(n2562)
         );
  OAI211XLTS U1087 ( .A0(n3772), .A1(n783), .B0(n1820), .C0(n1821), .Y(n2559)
         );
  OAI211XLTS U1088 ( .A0(n3772), .A1(n782), .B0(n1818), .C0(n1819), .Y(n2560)
         );
  OAI211XLTS U1089 ( .A0(n3771), .A1(n781), .B0(n1816), .C0(n1817), .Y(n2561)
         );
  OAI211XLTS U1090 ( .A0(n3772), .A1(n749), .B0(n1822), .C0(n1823), .Y(n2558)
         );
  OAI211XLTS U1091 ( .A0(n4420), .A1(n3279), .B0(n1289), .C0(n1290), .Y(n2803)
         );
  OAI211XLTS U1092 ( .A0(n4433), .A1(n3279), .B0(n1287), .C0(n1288), .Y(n2804)
         );
  OAI211XLTS U1093 ( .A0(n4444), .A1(n3279), .B0(n1285), .C0(n1286), .Y(n2805)
         );
  OAI211XLTS U1094 ( .A0(n4469), .A1(n3275), .B0(n1279), .C0(n1280), .Y(n2808)
         );
  OAI211XLTS U1095 ( .A0(n4476), .A1(n3274), .B0(n1277), .C0(n1278), .Y(n2809)
         );
  OAI211XLTS U1096 ( .A0(n4485), .A1(n3274), .B0(n1275), .C0(n1276), .Y(n2810)
         );
  OAI211XLTS U1097 ( .A0(n4501), .A1(n3274), .B0(n1271), .C0(n1272), .Y(n2812)
         );
  OAI211XLTS U1098 ( .A0(n4516), .A1(n3275), .B0(n1269), .C0(n1270), .Y(n2813)
         );
  OAI211XLTS U1099 ( .A0(n4530), .A1(n3275), .B0(n1265), .C0(n1266), .Y(n2815)
         );
  OAI211XLTS U1100 ( .A0(n4539), .A1(n3275), .B0(n1263), .C0(n1264), .Y(n2816)
         );
  OAI211XLTS U1101 ( .A0(n4548), .A1(n3276), .B0(n1261), .C0(n1262), .Y(n2817)
         );
  OAI211XLTS U1102 ( .A0(n4557), .A1(n3276), .B0(n1259), .C0(n1260), .Y(n2818)
         );
  OAI211XLTS U1103 ( .A0(n4568), .A1(n3276), .B0(n1257), .C0(n1258), .Y(n2819)
         );
  OAI211XLTS U1104 ( .A0(n4575), .A1(n3276), .B0(n1255), .C0(n1256), .Y(n2820)
         );
  OAI211XLTS U1105 ( .A0(n4588), .A1(n3277), .B0(n1253), .C0(n1254), .Y(n2821)
         );
  OAI211XLTS U1106 ( .A0(n4595), .A1(n3277), .B0(n1251), .C0(n1252), .Y(n2822)
         );
  OAI211XLTS U1107 ( .A0(n4600), .A1(n3277), .B0(n1249), .C0(n1250), .Y(n2823)
         );
  OAI211XLTS U1108 ( .A0(n4613), .A1(n3277), .B0(n1247), .C0(n1248), .Y(n2824)
         );
  OAI211XLTS U1109 ( .A0(n4633), .A1(n3278), .B0(n1243), .C0(n1244), .Y(n2826)
         );
  OAI211XLTS U1110 ( .A0(n4638), .A1(n3278), .B0(n1241), .C0(n1242), .Y(n2827)
         );
  OAI211XLTS U1111 ( .A0(n4647), .A1(n3278), .B0(n1239), .C0(n1240), .Y(n2828)
         );
  OAI211XLTS U1112 ( .A0(n4663), .A1(n3278), .B0(n1235), .C0(n1236), .Y(n2830)
         );
  OAI211XLTS U1113 ( .A0(n4674), .A1(n3279), .B0(n1233), .C0(n1234), .Y(n2831)
         );
  OAI211XLTS U1114 ( .A0(n4732), .A1(n3280), .B0(n1987), .C0(n1988), .Y(n2461)
         );
  OAI211XLTS U1115 ( .A0(n4743), .A1(n3280), .B0(n1985), .C0(n1986), .Y(n2462)
         );
  OAI211XLTS U1116 ( .A0(n4748), .A1(n3280), .B0(n1983), .C0(n1984), .Y(n2463)
         );
  OAI211XLTS U1117 ( .A0(n4724), .A1(n3280), .B0(n1989), .C0(n1990), .Y(n2460)
         );
  NAND2XLTS U1118 ( .A(n2005), .B(n469), .Y(n2004) );
  AOI32XLTS U1119 ( .A0(n100), .A1(n1809), .A2(n1810), .B0(n3284), .B1(n892), 
        .Y(n2563) );
  AOI21XLTS U1120 ( .A0(n15), .A1(n1811), .B0(n1812), .Y(n1810) );
  AOI21XLTS U1121 ( .A0(n15), .A1(n1780), .B0(n1781), .Y(n1779) );
  AOI21XLTS U1122 ( .A0(n4207), .A1(n99), .B0(n1785), .Y(n1778) );
  AOI22XLTS U1123 ( .A0(n1765), .A1(n1766), .B0(n3199), .B1(n599), .Y(n2569)
         );
  AOI21XLTS U1124 ( .A0(readIn_SOUTH), .A1(n1769), .B0(n1770), .Y(n1765) );
  OAI22XLTS U1125 ( .A0(n119), .A1(n2895), .B0(n2896), .B1(n2897), .Y(n2393)
         );
  NAND4XLTS U1126 ( .A(n470), .B(n977), .C(n975), .D(n1023), .Y(n2021) );
  NAND4XLTS U1127 ( .A(n490), .B(n977), .C(n1078), .D(n975), .Y(n2020) );
  NAND4XLTS U1128 ( .A(n469), .B(n474), .C(n975), .D(n978), .Y(n2018) );
  AOI2BB2XLTS U1129 ( .B0(n1758), .B1(n1759), .A0N(n3778), .A1N(
        readOutbuffer_7), .Y(n2570) );
  AOI32XLTS U1130 ( .A0(n1760), .A1(n1761), .A2(n1762), .B0(n4213), .B1(n686), 
        .Y(n1759) );
  AOI21XLTS U1131 ( .A0(n4207), .A1(n698), .B0(n488), .Y(n1758) );
  NAND3XLTS U1132 ( .A(n977), .B(n474), .C(n973), .Y(n2019) );
  NAND2X1TS U1133 ( .A(n46), .B(n47), .Y(n1827) );
  CLKBUFX2TS U1134 ( .A(n5323), .Y(n990) );
  XNOR2X1TS U1135 ( .A(n2892), .B(n2899), .Y(n1089) );
  NAND2X1TS U1136 ( .A(n46), .B(n989), .Y(n1879) );
  NOR2X1TS U1137 ( .A(n141), .B(n10), .Y(n1090) );
  NAND3X1TS U1138 ( .A(n10), .B(n475), .C(n122), .Y(n2029) );
  NAND3X1TS U1139 ( .A(n139), .B(n97), .C(n5), .Y(n2031) );
  NAND3X1TS U1140 ( .A(n141), .B(n658), .C(n385), .Y(n2028) );
  NAND3X1TS U1141 ( .A(n3), .B(n141), .C(n10), .Y(n2030) );
  NAND3X1TS U1142 ( .A(n98), .B(n139), .C(n122), .Y(n2044) );
  NAND2X1TS U1143 ( .A(n1090), .B(n122), .Y(n2026) );
  CLKBUFX2TS U1144 ( .A(n3878), .Y(n3868) );
  CLKBUFX2TS U1145 ( .A(n3877), .Y(n3869) );
  CLKBUFX2TS U1146 ( .A(n3876), .Y(n3871) );
  CLKBUFX2TS U1147 ( .A(n3878), .Y(n3867) );
  CLKBUFX2TS U1148 ( .A(n3877), .Y(n3870) );
  CLKBUFX2TS U1149 ( .A(n3947), .Y(n3940) );
  CLKBUFX2TS U1150 ( .A(n3945), .Y(n3944) );
  CLKBUFX2TS U1151 ( .A(n3946), .Y(n3943) );
  CLKBUFX2TS U1152 ( .A(n3946), .Y(n3942) );
  CLKBUFX2TS U1153 ( .A(n3947), .Y(n3941) );
  CLKBUFX2TS U1154 ( .A(n3948), .Y(n3939) );
  CLKBUFX2TS U1155 ( .A(n3864), .Y(n3859) );
  CLKBUFX2TS U1156 ( .A(n3862), .Y(n3860) );
  CLKBUFX2TS U1157 ( .A(n3862), .Y(n3857) );
  CLKBUFX2TS U1158 ( .A(n3863), .Y(n3856) );
  CLKBUFX2TS U1159 ( .A(n3862), .Y(n3858) );
  CLKBUFX2TS U1160 ( .A(n3863), .Y(n3855) );
  CLKBUFX2TS U1161 ( .A(n3825), .Y(n3812) );
  CLKBUFX2TS U1162 ( .A(n3825), .Y(n3813) );
  CLKBUFX2TS U1163 ( .A(n3824), .Y(n3814) );
  CLKBUFX2TS U1164 ( .A(n3824), .Y(n3815) );
  CLKBUFX2TS U1165 ( .A(n3823), .Y(n3816) );
  CLKBUFX2TS U1166 ( .A(n3823), .Y(n3817) );
  CLKBUFX2TS U1167 ( .A(n3823), .Y(n3819) );
  CLKBUFX2TS U1168 ( .A(n3822), .Y(n3818) );
  CLKBUFX2TS U1169 ( .A(n3876), .Y(n3872) );
  CLKBUFX2TS U1170 ( .A(n3905), .Y(n3895) );
  CLKBUFX2TS U1171 ( .A(n3875), .Y(n3873) );
  CLKBUFX2TS U1172 ( .A(n3908), .Y(n3901) );
  CLKBUFX2TS U1173 ( .A(n3903), .Y(n3900) );
  CLKBUFX2TS U1174 ( .A(n3904), .Y(n3898) );
  CLKBUFX2TS U1175 ( .A(n3904), .Y(n3897) );
  CLKBUFX2TS U1176 ( .A(n3903), .Y(n3899) );
  CLKBUFX2TS U1177 ( .A(n3905), .Y(n3896) );
  CLKBUFX2TS U1178 ( .A(n3875), .Y(n3874) );
  CLKBUFX2TS U1179 ( .A(n3826), .Y(n3825) );
  CLKBUFX2TS U1180 ( .A(n1748), .Y(n3822) );
  CLKBUFX2TS U1181 ( .A(n3826), .Y(n3824) );
  CLKBUFX2TS U1182 ( .A(n679), .Y(n3823) );
  CLKBUFX2TS U1183 ( .A(n3908), .Y(n3902) );
  CLKBUFX2TS U1184 ( .A(n3907), .Y(n3904) );
  CLKBUFX2TS U1185 ( .A(n3908), .Y(n3903) );
  CLKBUFX2TS U1186 ( .A(n3907), .Y(n3905) );
  CLKBUFX2TS U1187 ( .A(n669), .Y(n3875) );
  CLKBUFX2TS U1188 ( .A(n1741), .Y(n3876) );
  CLKBUFX2TS U1189 ( .A(n3879), .Y(n3878) );
  CLKBUFX2TS U1190 ( .A(n3865), .Y(n3862) );
  CLKBUFX2TS U1191 ( .A(n3865), .Y(n3863) );
  CLKBUFX2TS U1192 ( .A(n669), .Y(n3877) );
  CLKBUFX2TS U1193 ( .A(n3950), .Y(n3945) );
  CLKBUFX2TS U1194 ( .A(n3950), .Y(n3946) );
  CLKBUFX2TS U1195 ( .A(n3950), .Y(n3947) );
  CLKBUFX2TS U1196 ( .A(n660), .Y(n3948) );
  CLKBUFX2TS U1197 ( .A(n3466), .Y(n3452) );
  CLKBUFX2TS U1198 ( .A(n3466), .Y(n3453) );
  CLKBUFX2TS U1199 ( .A(n3463), .Y(n3458) );
  CLKBUFX2TS U1200 ( .A(n3463), .Y(n3457) );
  CLKBUFX2TS U1201 ( .A(n3462), .Y(n3459) );
  CLKBUFX2TS U1202 ( .A(n3464), .Y(n3456) );
  CLKBUFX2TS U1203 ( .A(n3464), .Y(n3455) );
  CLKBUFX2TS U1204 ( .A(n3466), .Y(n3454) );
  CLKBUFX2TS U1205 ( .A(n3383), .Y(n3369) );
  CLKBUFX2TS U1206 ( .A(n3949), .Y(n3938) );
  CLKBUFX2TS U1207 ( .A(n1756), .Y(n3949) );
  CLKBUFX2TS U1208 ( .A(n675), .Y(n3828) );
  CLKBUFX2TS U1209 ( .A(n3383), .Y(n3370) );
  CLKBUFX2TS U1210 ( .A(n3848), .Y(n3847) );
  CLKBUFX2TS U1211 ( .A(n3848), .Y(n3846) );
  CLKBUFX2TS U1212 ( .A(n3849), .Y(n3845) );
  CLKBUFX2TS U1213 ( .A(n3849), .Y(n3844) );
  CLKBUFX2TS U1214 ( .A(n3850), .Y(n3843) );
  CLKBUFX2TS U1215 ( .A(n3850), .Y(n3842) );
  CLKBUFX2TS U1216 ( .A(n3852), .Y(n3841) );
  CLKBUFX2TS U1217 ( .A(n3839), .Y(n3835) );
  CLKBUFX2TS U1218 ( .A(n3837), .Y(n3834) );
  CLKBUFX2TS U1219 ( .A(n3837), .Y(n3833) );
  CLKBUFX2TS U1220 ( .A(n3838), .Y(n3832) );
  CLKBUFX2TS U1221 ( .A(n675), .Y(n3831) );
  CLKBUFX2TS U1222 ( .A(n3838), .Y(n3830) );
  CLKBUFX2TS U1223 ( .A(n1743), .Y(n3829) );
  CLKBUFX2TS U1224 ( .A(n3839), .Y(n3836) );
  CLKBUFX2TS U1225 ( .A(n3380), .Y(n3371) );
  CLKBUFX2TS U1226 ( .A(n3378), .Y(n3375) );
  CLKBUFX2TS U1227 ( .A(n3379), .Y(n3373) );
  CLKBUFX2TS U1228 ( .A(n3379), .Y(n3374) );
  CLKBUFX2TS U1229 ( .A(n3380), .Y(n3372) );
  CLKBUFX2TS U1230 ( .A(n3413), .Y(n3400) );
  CLKBUFX2TS U1231 ( .A(n3264), .Y(n3251) );
  CLKBUFX2TS U1232 ( .A(n3264), .Y(n3252) );
  CLKBUFX2TS U1233 ( .A(n3262), .Y(n3256) );
  CLKBUFX2TS U1234 ( .A(n3262), .Y(n3255) );
  CLKBUFX2TS U1235 ( .A(n3263), .Y(n3254) );
  CLKBUFX2TS U1236 ( .A(n3261), .Y(n3257) );
  CLKBUFX2TS U1237 ( .A(n3263), .Y(n3253) );
  CLKBUFX2TS U1238 ( .A(n3413), .Y(n3401) );
  CLKBUFX2TS U1239 ( .A(n3864), .Y(n3854) );
  CLKBUFX2TS U1240 ( .A(n3865), .Y(n3864) );
  CLKBUFX2TS U1241 ( .A(n3412), .Y(n3405) );
  CLKBUFX2TS U1242 ( .A(n3412), .Y(n3404) );
  CLKBUFX2TS U1243 ( .A(n3410), .Y(n3407) );
  CLKBUFX2TS U1244 ( .A(n3415), .Y(n3406) );
  CLKBUFX2TS U1245 ( .A(n3412), .Y(n3403) );
  CLKBUFX2TS U1246 ( .A(n3245), .Y(n3240) );
  CLKBUFX2TS U1247 ( .A(n3247), .Y(n3236) );
  CLKBUFX2TS U1248 ( .A(n3247), .Y(n3237) );
  CLKBUFX2TS U1249 ( .A(n3246), .Y(n3238) );
  CLKBUFX2TS U1250 ( .A(n3246), .Y(n3239) );
  CLKBUFX2TS U1251 ( .A(n3245), .Y(n3241) );
  CLKBUFX2TS U1252 ( .A(n3244), .Y(n3242) );
  CLKBUFX2TS U1253 ( .A(n3462), .Y(n3460) );
  CLKBUFX2TS U1254 ( .A(n3248), .Y(n3234) );
  CLKBUFX2TS U1255 ( .A(n3248), .Y(n3235) );
  CLKBUFX2TS U1256 ( .A(n3378), .Y(n3376) );
  CLKBUFX2TS U1257 ( .A(n3244), .Y(n3243) );
  CLKBUFX2TS U1258 ( .A(n3935), .Y(n3925) );
  CLKBUFX2TS U1259 ( .A(n3933), .Y(n3930) );
  CLKBUFX2TS U1260 ( .A(n3934), .Y(n3928) );
  CLKBUFX2TS U1261 ( .A(n3932), .Y(n3931) );
  CLKBUFX2TS U1262 ( .A(n3933), .Y(n3929) );
  CLKBUFX2TS U1263 ( .A(n3934), .Y(n3927) );
  CLKBUFX2TS U1264 ( .A(n3935), .Y(n3926) );
  CLKBUFX2TS U1265 ( .A(n3906), .Y(n3894) );
  CLKBUFX2TS U1266 ( .A(n3907), .Y(n3906) );
  INVX2TS U1267 ( .A(n4605), .Y(n4606) );
  CLKBUFX2TS U1268 ( .A(n3806), .Y(n3795) );
  CLKBUFX2TS U1269 ( .A(n3806), .Y(n3796) );
  CLKBUFX2TS U1270 ( .A(n3803), .Y(n3802) );
  CLKBUFX2TS U1271 ( .A(n3805), .Y(n3797) );
  CLKBUFX2TS U1272 ( .A(n3804), .Y(n3799) );
  CLKBUFX2TS U1273 ( .A(n3805), .Y(n3798) );
  CLKBUFX2TS U1274 ( .A(n3803), .Y(n3801) );
  CLKBUFX2TS U1275 ( .A(n3804), .Y(n3800) );
  CLKBUFX2TS U1276 ( .A(n3433), .Y(n3428) );
  CLKBUFX2TS U1277 ( .A(n3485), .Y(n3480) );
  CLKBUFX2TS U1278 ( .A(n3485), .Y(n3481) );
  CLKBUFX2TS U1279 ( .A(n3485), .Y(n3482) );
  CLKBUFX2TS U1280 ( .A(n3433), .Y(n3429) );
  CLKBUFX2TS U1281 ( .A(n3433), .Y(n3430) );
  CLKBUFX2TS U1282 ( .A(n3414), .Y(n3412) );
  CLKBUFX2TS U1283 ( .A(n3415), .Y(n3411) );
  CLKBUFX2TS U1284 ( .A(n3415), .Y(n3410) );
  CLKBUFX2TS U1285 ( .A(n3384), .Y(n3381) );
  CLKBUFX2TS U1286 ( .A(n3384), .Y(n3382) );
  CLKBUFX2TS U1287 ( .A(n3384), .Y(n3383) );
  CLKBUFX2TS U1288 ( .A(n3414), .Y(n3413) );
  CLKBUFX2TS U1289 ( .A(n662), .Y(n3932) );
  CLKBUFX2TS U1290 ( .A(n662), .Y(n3933) );
  CLKBUFX2TS U1291 ( .A(n3937), .Y(n3934) );
  CLKBUFX2TS U1292 ( .A(n3937), .Y(n3935) );
  CLKBUFX2TS U1293 ( .A(n3468), .Y(n3463) );
  CLKBUFX2TS U1294 ( .A(n3467), .Y(n3466) );
  CLKBUFX2TS U1295 ( .A(n3468), .Y(n3464) );
  CLKBUFX2TS U1296 ( .A(n3467), .Y(n3465) );
  CLKBUFX2TS U1297 ( .A(n3853), .Y(n3848) );
  CLKBUFX2TS U1298 ( .A(n3853), .Y(n3849) );
  CLKBUFX2TS U1299 ( .A(n3853), .Y(n3850) );
  CLKBUFX2TS U1300 ( .A(n3839), .Y(n3837) );
  CLKBUFX2TS U1301 ( .A(n3265), .Y(n3262) );
  CLKBUFX2TS U1302 ( .A(n3249), .Y(n3247) );
  CLKBUFX2TS U1303 ( .A(n3249), .Y(n3246) );
  CLKBUFX2TS U1304 ( .A(n1214), .Y(n3245) );
  CLKBUFX2TS U1305 ( .A(n3265), .Y(n3263) );
  CLKBUFX2TS U1306 ( .A(n1214), .Y(n3244) );
  CLKBUFX2TS U1307 ( .A(n3265), .Y(n3264) );
  CLKBUFX2TS U1308 ( .A(n3468), .Y(n3462) );
  CLKBUFX2TS U1309 ( .A(n3266), .Y(n3261) );
  CLKBUFX2TS U1310 ( .A(n3249), .Y(n3248) );
  CLKBUFX2TS U1311 ( .A(n3385), .Y(n3379) );
  CLKBUFX2TS U1312 ( .A(n3385), .Y(n3380) );
  CLKBUFX2TS U1313 ( .A(n3385), .Y(n3378) );
  CLKBUFX2TS U1314 ( .A(n679), .Y(n3826) );
  CLKBUFX2TS U1315 ( .A(n665), .Y(n3908) );
  CLKBUFX2TS U1316 ( .A(n665), .Y(n3907) );
  CLKBUFX2TS U1317 ( .A(n669), .Y(n3879) );
  CLKBUFX2TS U1318 ( .A(n660), .Y(n3950) );
  CLKBUFX2TS U1319 ( .A(n670), .Y(n3865) );
  CLKBUFX2TS U1320 ( .A(n3301), .Y(n3286) );
  CLKBUFX2TS U1321 ( .A(n3215), .Y(n3203) );
  CLKBUFX2TS U1322 ( .A(n3301), .Y(n3287) );
  CLKBUFX2TS U1323 ( .A(n3565), .Y(n3551) );
  CLKBUFX2TS U1324 ( .A(n3218), .Y(n3204) );
  CLKBUFX2TS U1325 ( .A(n3679), .Y(n3669) );
  CLKBUFX2TS U1326 ( .A(n3678), .Y(n3670) );
  CLKBUFX2TS U1327 ( .A(n3713), .Y(n3699) );
  CLKBUFX2TS U1328 ( .A(n3298), .Y(n3296) );
  CLKBUFX2TS U1329 ( .A(n3300), .Y(n3295) );
  CLKBUFX2TS U1330 ( .A(n3302), .Y(n3294) );
  CLKBUFX2TS U1331 ( .A(n3299), .Y(n3293) );
  CLKBUFX2TS U1332 ( .A(n1199), .Y(n3291) );
  CLKBUFX2TS U1333 ( .A(n3300), .Y(n3290) );
  CLKBUFX2TS U1334 ( .A(n3299), .Y(n3292) );
  CLKBUFX2TS U1335 ( .A(n3300), .Y(n3289) );
  CLKBUFX2TS U1336 ( .A(n3300), .Y(n3288) );
  CLKBUFX2TS U1337 ( .A(n3678), .Y(n3671) );
  CLKBUFX2TS U1338 ( .A(n3677), .Y(n3667) );
  CLKBUFX2TS U1339 ( .A(n3680), .Y(n3665) );
  CLKBUFX2TS U1340 ( .A(n3709), .Y(n3706) );
  CLKBUFX2TS U1341 ( .A(n3709), .Y(n3705) );
  CLKBUFX2TS U1342 ( .A(n3710), .Y(n3704) );
  CLKBUFX2TS U1343 ( .A(n3710), .Y(n3703) );
  CLKBUFX2TS U1344 ( .A(n3711), .Y(n3702) );
  CLKBUFX2TS U1345 ( .A(n3711), .Y(n3701) );
  CLKBUFX2TS U1346 ( .A(n3713), .Y(n3700) );
  CLKBUFX2TS U1347 ( .A(n3679), .Y(n3668) );
  CLKBUFX2TS U1348 ( .A(n3680), .Y(n3666) );
  CLKBUFX2TS U1349 ( .A(n3562), .Y(n3557) );
  CLKBUFX2TS U1350 ( .A(n3562), .Y(n3556) );
  CLKBUFX2TS U1351 ( .A(n3563), .Y(n3555) );
  CLKBUFX2TS U1352 ( .A(n3564), .Y(n3553) );
  CLKBUFX2TS U1353 ( .A(n3564), .Y(n3552) );
  CLKBUFX2TS U1354 ( .A(n3563), .Y(n3554) );
  CLKBUFX2TS U1355 ( .A(n3561), .Y(n3558) );
  CLKBUFX2TS U1356 ( .A(n3217), .Y(n3205) );
  CLKBUFX2TS U1357 ( .A(n3214), .Y(n3210) );
  CLKBUFX2TS U1358 ( .A(n3215), .Y(n3209) );
  CLKBUFX2TS U1359 ( .A(n3215), .Y(n3208) );
  CLKBUFX2TS U1360 ( .A(n3216), .Y(n3207) );
  CLKBUFX2TS U1361 ( .A(n3216), .Y(n3206) );
  CLKBUFX2TS U1362 ( .A(n3500), .Y(n3486) );
  CLKBUFX2TS U1363 ( .A(n3649), .Y(n3634) );
  CLKBUFX2TS U1364 ( .A(n3449), .Y(n3435) );
  CLKBUFX2TS U1365 ( .A(n3851), .Y(n3840) );
  CLKBUFX2TS U1366 ( .A(n3852), .Y(n3851) );
  CLKBUFX2TS U1367 ( .A(n3838), .Y(n3827) );
  CLKBUFX2TS U1368 ( .A(n675), .Y(n3838) );
  CLKBUFX2TS U1369 ( .A(n3449), .Y(n3436) );
  CLKBUFX2TS U1370 ( .A(n3649), .Y(n3635) );
  CLKBUFX2TS U1371 ( .A(n3500), .Y(n3487) );
  CLKBUFX2TS U1372 ( .A(n3444), .Y(n3441) );
  CLKBUFX2TS U1373 ( .A(n3447), .Y(n3440) );
  CLKBUFX2TS U1374 ( .A(n3447), .Y(n3439) );
  CLKBUFX2TS U1375 ( .A(n3448), .Y(n3437) );
  CLKBUFX2TS U1376 ( .A(n3448), .Y(n3438) );
  CLKBUFX2TS U1377 ( .A(n3648), .Y(n3636) );
  CLKBUFX2TS U1378 ( .A(n3496), .Y(n3493) );
  CLKBUFX2TS U1379 ( .A(n3496), .Y(n3492) );
  CLKBUFX2TS U1380 ( .A(n3499), .Y(n3489) );
  CLKBUFX2TS U1381 ( .A(n3498), .Y(n3491) );
  CLKBUFX2TS U1382 ( .A(n3498), .Y(n3490) );
  CLKBUFX2TS U1383 ( .A(n3499), .Y(n3488) );
  INVX2TS U1384 ( .A(n3693), .Y(n3692) );
  INVX2TS U1385 ( .A(n3695), .Y(n3690) );
  INVX2TS U1386 ( .A(n3694), .Y(n3691) );
  CLKBUFX2TS U1387 ( .A(n3613), .Y(n3599) );
  CLKBUFX2TS U1388 ( .A(n3379), .Y(n3377) );
  CLKBUFX2TS U1389 ( .A(n3348), .Y(n3334) );
  CLKBUFX2TS U1390 ( .A(n3613), .Y(n3600) );
  CLKBUFX2TS U1391 ( .A(n3759), .Y(n3753) );
  CLKBUFX2TS U1392 ( .A(n3715), .Y(n3707) );
  CLKBUFX2TS U1393 ( .A(n3762), .Y(n3747) );
  CLKBUFX2TS U1394 ( .A(n3343), .Y(n3340) );
  CLKBUFX2TS U1395 ( .A(n3344), .Y(n3339) );
  CLKBUFX2TS U1396 ( .A(n3344), .Y(n3338) );
  CLKBUFX2TS U1397 ( .A(n3345), .Y(n3337) );
  CLKBUFX2TS U1398 ( .A(n3346), .Y(n3335) );
  CLKBUFX2TS U1399 ( .A(n3345), .Y(n3336) );
  CLKBUFX2TS U1400 ( .A(n3760), .Y(n3752) );
  CLKBUFX2TS U1401 ( .A(n3760), .Y(n3751) );
  CLKBUFX2TS U1402 ( .A(n3761), .Y(n3750) );
  CLKBUFX2TS U1403 ( .A(n3761), .Y(n3749) );
  CLKBUFX2TS U1404 ( .A(n3762), .Y(n3748) );
  CLKBUFX2TS U1405 ( .A(n3611), .Y(n3604) );
  CLKBUFX2TS U1406 ( .A(n3611), .Y(n3603) );
  CLKBUFX2TS U1407 ( .A(n3610), .Y(n3605) );
  CLKBUFX2TS U1408 ( .A(n3612), .Y(n3602) );
  CLKBUFX2TS U1409 ( .A(n3612), .Y(n3601) );
  CLKBUFX2TS U1410 ( .A(n3298), .Y(n3297) );
  CLKBUFX2TS U1411 ( .A(n3919), .Y(n3917) );
  CLKBUFX2TS U1412 ( .A(n3922), .Y(n3911) );
  CLKBUFX2TS U1413 ( .A(n3920), .Y(n3916) );
  CLKBUFX2TS U1414 ( .A(n3920), .Y(n3915) );
  CLKBUFX2TS U1415 ( .A(n3921), .Y(n3914) );
  CLKBUFX2TS U1416 ( .A(n3921), .Y(n3913) );
  CLKBUFX2TS U1417 ( .A(n3923), .Y(n3910) );
  CLKBUFX2TS U1418 ( .A(n3922), .Y(n3909) );
  CLKBUFX2TS U1419 ( .A(n3922), .Y(n3912) );
  CLKBUFX2TS U1420 ( .A(n3888), .Y(n3886) );
  CLKBUFX2TS U1421 ( .A(n3888), .Y(n3887) );
  CLKBUFX2TS U1422 ( .A(n3889), .Y(n3885) );
  CLKBUFX2TS U1423 ( .A(n3890), .Y(n3882) );
  CLKBUFX2TS U1424 ( .A(n3891), .Y(n3881) );
  CLKBUFX2TS U1425 ( .A(n3889), .Y(n3884) );
  CLKBUFX2TS U1426 ( .A(n3890), .Y(n3883) );
  CLKBUFX2TS U1427 ( .A(n3891), .Y(n3880) );
  CLKBUFX2TS U1428 ( .A(n3677), .Y(n3673) );
  CLKBUFX2TS U1429 ( .A(n3677), .Y(n3672) );
  CLKBUFX2TS U1430 ( .A(n3532), .Y(n3517) );
  CLKBUFX2TS U1431 ( .A(n3532), .Y(n3518) );
  CLKBUFX2TS U1432 ( .A(n3214), .Y(n3211) );
  CLKBUFX2TS U1433 ( .A(n3758), .Y(n3754) );
  CLKBUFX2TS U1434 ( .A(n3676), .Y(n3674) );
  CLKBUFX2TS U1435 ( .A(n3531), .Y(n3519) );
  CLKBUFX2TS U1436 ( .A(n3730), .Y(n3717) );
  CLKBUFX2TS U1437 ( .A(n3728), .Y(n3716) );
  CLKBUFX2TS U1438 ( .A(n3496), .Y(n3494) );
  CLKBUFX2TS U1439 ( .A(n3581), .Y(n3568) );
  CLKBUFX2TS U1440 ( .A(n3581), .Y(n3569) );
  CLKBUFX2TS U1441 ( .A(n3648), .Y(n3637) );
  CLKBUFX2TS U1442 ( .A(n3317), .Y(n3303) );
  CLKBUFX2TS U1443 ( .A(n3317), .Y(n3304) );
  CLKBUFX2TS U1444 ( .A(n3528), .Y(n3526) );
  CLKBUFX2TS U1445 ( .A(n3528), .Y(n3525) );
  CLKBUFX2TS U1446 ( .A(n3530), .Y(n3521) );
  CLKBUFX2TS U1447 ( .A(n3529), .Y(n3524) );
  CLKBUFX2TS U1448 ( .A(n3529), .Y(n3523) );
  CLKBUFX2TS U1449 ( .A(n3530), .Y(n3522) );
  CLKBUFX2TS U1450 ( .A(n3531), .Y(n3520) );
  CLKBUFX2TS U1451 ( .A(n3647), .Y(n3638) );
  CLKBUFX2TS U1452 ( .A(n3463), .Y(n3461) );
  CLKBUFX2TS U1453 ( .A(n3676), .Y(n3675) );
  CLKBUFX2TS U1454 ( .A(n3316), .Y(n3305) );
  CLKBUFX2TS U1455 ( .A(n3316), .Y(n3306) );
  CLKBUFX2TS U1456 ( .A(n3647), .Y(n3639) );
  CLKBUFX2TS U1457 ( .A(n3728), .Y(n3719) );
  CLKBUFX2TS U1458 ( .A(n3726), .Y(n3723) );
  CLKBUFX2TS U1459 ( .A(n3726), .Y(n3722) );
  CLKBUFX2TS U1460 ( .A(n3727), .Y(n3721) );
  CLKBUFX2TS U1461 ( .A(n3727), .Y(n3720) );
  CLKBUFX2TS U1462 ( .A(n3728), .Y(n3718) );
  CLKBUFX2TS U1463 ( .A(n3583), .Y(n3576) );
  CLKBUFX2TS U1464 ( .A(n3578), .Y(n3574) );
  CLKBUFX2TS U1465 ( .A(n3578), .Y(n3575) );
  CLKBUFX2TS U1466 ( .A(n3579), .Y(n3573) );
  CLKBUFX2TS U1467 ( .A(n3579), .Y(n3572) );
  CLKBUFX2TS U1468 ( .A(n3645), .Y(n3643) );
  CLKBUFX2TS U1469 ( .A(n3316), .Y(n3311) );
  CLKBUFX2TS U1470 ( .A(n3314), .Y(n3309) );
  CLKBUFX2TS U1471 ( .A(n3314), .Y(n3310) );
  CLKBUFX2TS U1472 ( .A(n3315), .Y(n3308) );
  CLKBUFX2TS U1473 ( .A(n3646), .Y(n3641) );
  CLKBUFX2TS U1474 ( .A(n3315), .Y(n3307) );
  CLKBUFX2TS U1475 ( .A(n3645), .Y(n3642) );
  CLKBUFX2TS U1476 ( .A(n3646), .Y(n3640) );
  CLKBUFX2TS U1477 ( .A(n3444), .Y(n3442) );
  CLKBUFX2TS U1478 ( .A(n3260), .Y(n3259) );
  CLKBUFX2TS U1479 ( .A(n3936), .Y(n3924) );
  CLKBUFX2TS U1480 ( .A(n3937), .Y(n3936) );
  CLKBUFX2TS U1481 ( .A(n3758), .Y(n3755) );
  CLKBUFX2TS U1482 ( .A(n3919), .Y(n3918) );
  INVX2TS U1483 ( .A(n3483), .Y(n3470) );
  INVX2TS U1484 ( .A(n3483), .Y(n3471) );
  INVX2TS U1485 ( .A(n3483), .Y(n3469) );
  INVX2TS U1486 ( .A(n3484), .Y(n3472) );
  INVX2TS U1487 ( .A(n3484), .Y(n3473) );
  INVX2TS U1488 ( .A(n3483), .Y(n3474) );
  INVX2TS U1489 ( .A(n3484), .Y(n3475) );
  INVX2TS U1490 ( .A(n3484), .Y(n3476) );
  INVX2TS U1491 ( .A(n3431), .Y(n3421) );
  CLKBUFX2TS U1492 ( .A(n3432), .Y(n3431) );
  INVX2TS U1493 ( .A(n3432), .Y(n3417) );
  INVX2TS U1494 ( .A(n3433), .Y(n3419) );
  INVX2TS U1495 ( .A(n3432), .Y(n3423) );
  INVX2TS U1496 ( .A(n3431), .Y(n3418) );
  INVX2TS U1497 ( .A(n3432), .Y(n3420) );
  INVX2TS U1498 ( .A(n3431), .Y(n3422) );
  INVX2TS U1499 ( .A(n3431), .Y(n3424) );
  CLKBUFX2TS U1500 ( .A(n3330), .Y(n3321) );
  CLKBUFX2TS U1501 ( .A(n3331), .Y(n3323) );
  CLKBUFX2TS U1502 ( .A(n3331), .Y(n3322) );
  CLKBUFX2TS U1503 ( .A(n3330), .Y(n3325) );
  CLKBUFX2TS U1504 ( .A(n3329), .Y(n3326) );
  CLKBUFX2TS U1505 ( .A(n3331), .Y(n3324) );
  CLKBUFX2TS U1506 ( .A(n3230), .Y(n3222) );
  CLKBUFX2TS U1507 ( .A(n3230), .Y(n3221) );
  CLKBUFX2TS U1508 ( .A(n3329), .Y(n3327) );
  CLKBUFX2TS U1509 ( .A(n1197), .Y(n3328) );
  CLKBUFX2TS U1510 ( .A(n3229), .Y(n3223) );
  CLKBUFX2TS U1511 ( .A(n3229), .Y(n3224) );
  CLKBUFX2TS U1512 ( .A(n3226), .Y(n3225) );
  CLKBUFX2TS U1513 ( .A(reset), .Y(n4605) );
  CLKBUFX2TS U1514 ( .A(n3807), .Y(n3806) );
  CLKBUFX2TS U1515 ( .A(n3808), .Y(n3805) );
  CLKBUFX2TS U1516 ( .A(n3808), .Y(n3803) );
  CLKBUFX2TS U1517 ( .A(n3808), .Y(n3804) );
  CLKBUFX2TS U1518 ( .A(n3396), .Y(n3388) );
  CLKBUFX2TS U1519 ( .A(n3396), .Y(n3387) );
  CLKBUFX2TS U1520 ( .A(n3395), .Y(n3389) );
  CLKBUFX2TS U1521 ( .A(n3393), .Y(n3391) );
  CLKBUFX2TS U1522 ( .A(n3393), .Y(n3392) );
  CLKBUFX2TS U1523 ( .A(n3395), .Y(n3390) );
  CLKBUFX2TS U1524 ( .A(n1098), .Y(n3759) );
  CLKBUFX2TS U1525 ( .A(n3698), .Y(n3695) );
  CLKBUFX2TS U1526 ( .A(n3698), .Y(n3694) );
  CLKBUFX2TS U1527 ( .A(n3698), .Y(n3693) );
  CLKBUFX2TS U1528 ( .A(n3550), .Y(n3547) );
  CLKBUFX2TS U1529 ( .A(n3550), .Y(n3545) );
  CLKBUFX2TS U1530 ( .A(n3550), .Y(n3546) );
  CLKBUFX2TS U1531 ( .A(n1180), .Y(n3415) );
  CLKBUFX2TS U1532 ( .A(n1180), .Y(n3414) );
  CLKBUFX2TS U1533 ( .A(n1182), .Y(n3384) );
  CLKBUFX2TS U1534 ( .A(n3923), .Y(n3919) );
  CLKBUFX2TS U1535 ( .A(n3923), .Y(n3920) );
  CLKBUFX2TS U1536 ( .A(n3923), .Y(n3921) );
  CLKBUFX2TS U1537 ( .A(n3730), .Y(n3729) );
  CLKBUFX2TS U1538 ( .A(n3731), .Y(n3726) );
  CLKBUFX2TS U1539 ( .A(n3731), .Y(n3727) );
  CLKBUFX2TS U1540 ( .A(n3731), .Y(n3728) );
  CLKBUFX2TS U1541 ( .A(n3583), .Y(n3578) );
  CLKBUFX2TS U1542 ( .A(n3582), .Y(n3579) );
  CLKBUFX2TS U1543 ( .A(n3582), .Y(n3580) );
  CLKBUFX2TS U1544 ( .A(n3582), .Y(n3581) );
  CLKBUFX2TS U1545 ( .A(n3650), .Y(n3649) );
  CLKBUFX2TS U1546 ( .A(n3681), .Y(n3676) );
  CLKBUFX2TS U1547 ( .A(n3650), .Y(n3648) );
  CLKBUFX2TS U1548 ( .A(n3318), .Y(n3316) );
  CLKBUFX2TS U1549 ( .A(n3350), .Y(n3344) );
  CLKBUFX2TS U1550 ( .A(n3319), .Y(n3313) );
  CLKBUFX2TS U1551 ( .A(n3349), .Y(n3346) );
  CLKBUFX2TS U1552 ( .A(n3350), .Y(n3345) );
  CLKBUFX2TS U1553 ( .A(n3302), .Y(n3299) );
  CLKBUFX2TS U1554 ( .A(n3319), .Y(n3314) );
  CLKBUFX2TS U1555 ( .A(n3349), .Y(n3347) );
  CLKBUFX2TS U1556 ( .A(n3302), .Y(n3300) );
  CLKBUFX2TS U1557 ( .A(n3681), .Y(n3678) );
  CLKBUFX2TS U1558 ( .A(n1101), .Y(n3709) );
  CLKBUFX2TS U1559 ( .A(n1101), .Y(n3710) );
  CLKBUFX2TS U1560 ( .A(n3763), .Y(n3760) );
  CLKBUFX2TS U1561 ( .A(n3714), .Y(n3711) );
  CLKBUFX2TS U1562 ( .A(n3763), .Y(n3761) );
  CLKBUFX2TS U1563 ( .A(n3714), .Y(n3712) );
  CLKBUFX2TS U1564 ( .A(n3763), .Y(n3762) );
  CLKBUFX2TS U1565 ( .A(n3714), .Y(n3713) );
  CLKBUFX2TS U1566 ( .A(n3318), .Y(n3315) );
  CLKBUFX2TS U1567 ( .A(n3349), .Y(n3348) );
  CLKBUFX2TS U1568 ( .A(n1199), .Y(n3301) );
  CLKBUFX2TS U1569 ( .A(n3650), .Y(n3645) );
  CLKBUFX2TS U1570 ( .A(n1116), .Y(n3679) );
  CLKBUFX2TS U1571 ( .A(n1118), .Y(n3646) );
  CLKBUFX2TS U1572 ( .A(n1116), .Y(n3680) );
  CLKBUFX2TS U1573 ( .A(n3615), .Y(n3609) );
  CLKBUFX2TS U1574 ( .A(n3567), .Y(n3562) );
  CLKBUFX2TS U1575 ( .A(n3614), .Y(n3611) );
  CLKBUFX2TS U1576 ( .A(n3566), .Y(n3564) );
  CLKBUFX2TS U1577 ( .A(n3615), .Y(n3610) );
  CLKBUFX2TS U1578 ( .A(n3567), .Y(n3563) );
  CLKBUFX2TS U1579 ( .A(n3614), .Y(n3612) );
  CLKBUFX2TS U1580 ( .A(n3566), .Y(n3565) );
  CLKBUFX2TS U1581 ( .A(n3614), .Y(n3613) );
  CLKBUFX2TS U1582 ( .A(n3350), .Y(n3343) );
  CLKBUFX2TS U1583 ( .A(n3318), .Y(n3317) );
  CLKBUFX2TS U1584 ( .A(n3302), .Y(n3298) );
  CLKBUFX2TS U1585 ( .A(n3218), .Y(n3217) );
  CLKBUFX2TS U1586 ( .A(n3219), .Y(n3215) );
  CLKBUFX2TS U1587 ( .A(n3219), .Y(n3216) );
  CLKBUFX2TS U1588 ( .A(n668), .Y(n3888) );
  CLKBUFX2TS U1589 ( .A(n3502), .Y(n3497) );
  CLKBUFX2TS U1590 ( .A(n3533), .Y(n3528) );
  CLKBUFX2TS U1591 ( .A(n3893), .Y(n3892) );
  CLKBUFX2TS U1592 ( .A(n3501), .Y(n3500) );
  CLKBUFX2TS U1593 ( .A(n3893), .Y(n3889) );
  CLKBUFX2TS U1594 ( .A(n1149), .Y(n3529) );
  CLKBUFX2TS U1595 ( .A(n3533), .Y(n3530) );
  CLKBUFX2TS U1596 ( .A(n3893), .Y(n3890) );
  CLKBUFX2TS U1597 ( .A(n3501), .Y(n3498) );
  CLKBUFX2TS U1598 ( .A(n3533), .Y(n3531) );
  CLKBUFX2TS U1599 ( .A(n3893), .Y(n3891) );
  CLKBUFX2TS U1600 ( .A(n3501), .Y(n3499) );
  CLKBUFX2TS U1601 ( .A(n3650), .Y(n3647) );
  CLKBUFX2TS U1602 ( .A(n3681), .Y(n3677) );
  CLKBUFX2TS U1603 ( .A(n3533), .Y(n3532) );
  CLKBUFX2TS U1604 ( .A(n3567), .Y(n3561) );
  CLKBUFX2TS U1605 ( .A(n3219), .Y(n3214) );
  CLKBUFX2TS U1606 ( .A(n3416), .Y(n3409) );
  CLKBUFX2TS U1607 ( .A(n1180), .Y(n3416) );
  CLKBUFX2TS U1608 ( .A(n3451), .Y(n3445) );
  CLKBUFX2TS U1609 ( .A(n3450), .Y(n3449) );
  CLKBUFX2TS U1610 ( .A(n3451), .Y(n3446) );
  CLKBUFX2TS U1611 ( .A(n3450), .Y(n3447) );
  CLKBUFX2TS U1612 ( .A(n3450), .Y(n3448) );
  CLKBUFX2TS U1613 ( .A(n3921), .Y(n3922) );
  CLKBUFX2TS U1614 ( .A(n1214), .Y(n3250) );
  CLKBUFX2TS U1615 ( .A(n3451), .Y(n3444) );
  CLKBUFX2TS U1616 ( .A(n3267), .Y(n3260) );
  CLKBUFX2TS U1617 ( .A(n1213), .Y(n3267) );
  CLKBUFX2TS U1618 ( .A(n1165), .Y(n3467) );
  CLKBUFX2TS U1619 ( .A(n1165), .Y(n3468) );
  CLKBUFX2TS U1620 ( .A(n1213), .Y(n3265) );
  CLKBUFX2TS U1621 ( .A(n1214), .Y(n3249) );
  CLKBUFX2TS U1622 ( .A(n662), .Y(n3937) );
  CLKBUFX2TS U1623 ( .A(n976), .Y(n3853) );
  CLKBUFX2TS U1624 ( .A(n976), .Y(n3852) );
  CLKBUFX2TS U1625 ( .A(n675), .Y(n3839) );
  CLKBUFX2TS U1626 ( .A(n1182), .Y(n3385) );
  INVX2TS U1627 ( .A(n3696), .Y(n3683) );
  CLKBUFX2TS U1628 ( .A(n3697), .Y(n3696) );
  INVX2TS U1629 ( .A(n3696), .Y(n3684) );
  INVX2TS U1630 ( .A(n3698), .Y(n3685) );
  INVX2TS U1631 ( .A(n3697), .Y(n3686) );
  INVX2TS U1632 ( .A(n3696), .Y(n3687) );
  INVX2TS U1633 ( .A(n3697), .Y(n3688) );
  INVX2TS U1634 ( .A(n982), .Y(n3689) );
  INVX2TS U1635 ( .A(n3697), .Y(n3682) );
  INVX2TS U1636 ( .A(n952), .Y(n665) );
  INVX2TS U1637 ( .A(n689), .Y(n660) );
  CLKBUFX2TS U1638 ( .A(n981), .Y(n3483) );
  CLKBUFX2TS U1639 ( .A(n981), .Y(n3484) );
  CLKBUFX2TS U1640 ( .A(n3434), .Y(n3432) );
  CLKBUFX2TS U1641 ( .A(n981), .Y(n3485) );
  CLKBUFX2TS U1642 ( .A(n3434), .Y(n3433) );
  CLKBUFX2TS U1643 ( .A(n3567), .Y(n3560) );
  CLKBUFX2TS U1644 ( .A(n3213), .Y(n3212) );
  CLKBUFX2TS U1645 ( .A(n3532), .Y(n3527) );
  CLKBUFX2TS U1646 ( .A(n3315), .Y(n3312) );
  CLKBUFX2TS U1647 ( .A(n3649), .Y(n3644) );
  CLKBUFX2TS U1648 ( .A(n3584), .Y(n3577) );
  CLKBUFX2TS U1649 ( .A(n3349), .Y(n3342) );
  CLKBUFX2TS U1650 ( .A(n3451), .Y(n3443) );
  CLKBUFX2TS U1651 ( .A(n3549), .Y(n3548) );
  CLKBUFX2TS U1652 ( .A(n3333), .Y(n3330) );
  CLKBUFX2TS U1653 ( .A(n1197), .Y(n3329) );
  CLKBUFX2TS U1654 ( .A(n3333), .Y(n3331) );
  CLKBUFX2TS U1655 ( .A(n3232), .Y(n3229) );
  CLKBUFX2TS U1656 ( .A(n3233), .Y(n3228) );
  CLKBUFX2TS U1657 ( .A(n3233), .Y(n3227) );
  CLKBUFX2TS U1658 ( .A(n3233), .Y(n3226) );
  CLKBUFX2TS U1659 ( .A(n3232), .Y(n3230) );
  INVX2TS U1660 ( .A(n3120), .Y(n3105) );
  INVX2TS U1661 ( .A(n3120), .Y(n3106) );
  INVX2TS U1662 ( .A(n3121), .Y(n3115) );
  INVX2TS U1663 ( .A(n3121), .Y(n3114) );
  INVX2TS U1664 ( .A(n3119), .Y(n3113) );
  INVX2TS U1665 ( .A(n3119), .Y(n3112) );
  INVX2TS U1666 ( .A(n3116), .Y(n3111) );
  INVX2TS U1667 ( .A(n3116), .Y(n3109) );
  INVX2TS U1668 ( .A(n3116), .Y(n3108) );
  INVX2TS U1669 ( .A(n3116), .Y(n3110) );
  INVX2TS U1670 ( .A(n3120), .Y(n3107) );
  CLKBUFX2TS U1671 ( .A(n3332), .Y(n3320) );
  CLKBUFX2TS U1672 ( .A(n3333), .Y(n3332) );
  CLKBUFX2TS U1673 ( .A(n3777), .Y(n3764) );
  CLKBUFX2TS U1674 ( .A(n3660), .Y(n3652) );
  CLKBUFX2TS U1675 ( .A(n3659), .Y(n3654) );
  CLKBUFX2TS U1676 ( .A(n3661), .Y(n3651) );
  CLKBUFX2TS U1677 ( .A(n3659), .Y(n3655) );
  CLKBUFX2TS U1678 ( .A(n3658), .Y(n3657) );
  CLKBUFX2TS U1679 ( .A(n3743), .Y(n3734) );
  CLKBUFX2TS U1680 ( .A(n3743), .Y(n3735) );
  CLKBUFX2TS U1681 ( .A(n3742), .Y(n3736) );
  CLKBUFX2TS U1682 ( .A(n3742), .Y(n3737) );
  CLKBUFX2TS U1683 ( .A(n3739), .Y(n3738) );
  CLKBUFX2TS U1684 ( .A(n3660), .Y(n3653) );
  CLKBUFX2TS U1685 ( .A(n3658), .Y(n3656) );
  CLKBUFX2TS U1686 ( .A(n3597), .Y(n3585) );
  CLKBUFX2TS U1687 ( .A(n3596), .Y(n3587) );
  CLKBUFX2TS U1688 ( .A(n1133), .Y(n3586) );
  CLKBUFX2TS U1689 ( .A(n3595), .Y(n3589) );
  CLKBUFX2TS U1690 ( .A(n3595), .Y(n3590) );
  CLKBUFX2TS U1691 ( .A(n3596), .Y(n3588) );
  CLKBUFX2TS U1692 ( .A(n3595), .Y(n3591) );
  CLKBUFX2TS U1693 ( .A(n3594), .Y(n3592) );
  CLKBUFX2TS U1694 ( .A(n3594), .Y(n3593) );
  CLKBUFX2TS U1695 ( .A(n3231), .Y(n3220) );
  CLKBUFX2TS U1696 ( .A(n3232), .Y(n3231) );
  CLKBUFX2TS U1697 ( .A(n3774), .Y(n3770) );
  CLKBUFX2TS U1698 ( .A(n3774), .Y(n3769) );
  CLKBUFX2TS U1699 ( .A(n3775), .Y(n3768) );
  CLKBUFX2TS U1700 ( .A(n3775), .Y(n3767) );
  CLKBUFX2TS U1701 ( .A(n3776), .Y(n3766) );
  CLKBUFX2TS U1702 ( .A(n3776), .Y(n3765) );
  CLKBUFX2TS U1703 ( .A(n3065), .Y(n3061) );
  CLKBUFX2TS U1704 ( .A(n3065), .Y(n3060) );
  CLKBUFX2TS U1705 ( .A(n3066), .Y(n3059) );
  CLKBUFX2TS U1706 ( .A(n3066), .Y(n3058) );
  CLKBUFX2TS U1707 ( .A(n3067), .Y(n3057) );
  CLKBUFX2TS U1708 ( .A(n3067), .Y(n3056) );
  INVX2TS U1709 ( .A(n3198), .Y(n3187) );
  INVX2TS U1710 ( .A(n3198), .Y(n3189) );
  INVX2TS U1711 ( .A(n3197), .Y(n3192) );
  INVX2TS U1712 ( .A(n3198), .Y(n3188) );
  INVX2TS U1713 ( .A(n3197), .Y(n3191) );
  INVX2TS U1714 ( .A(n3196), .Y(n3193) );
  INVX2TS U1715 ( .A(n3197), .Y(n3190) );
  INVX2TS U1716 ( .A(n3196), .Y(n3194) );
  INVX2TS U1717 ( .A(n3368), .Y(n3361) );
  INVX2TS U1718 ( .A(n3367), .Y(n3360) );
  INVX2TS U1719 ( .A(n3366), .Y(n3359) );
  INVX2TS U1720 ( .A(n3630), .Y(n3626) );
  INVX2TS U1721 ( .A(n3630), .Y(n3625) );
  INVX2TS U1722 ( .A(n3630), .Y(n3624) );
  INVX2TS U1723 ( .A(n3366), .Y(n3353) );
  INVX2TS U1724 ( .A(n3633), .Y(n3618) );
  INVX2TS U1725 ( .A(n3283), .Y(n3270) );
  INVX2TS U1726 ( .A(n3365), .Y(n3358) );
  INVX2TS U1727 ( .A(n3365), .Y(n3357) );
  INVX2TS U1728 ( .A(n3365), .Y(n3356) );
  INVX2TS U1729 ( .A(n3366), .Y(n3355) );
  INVX2TS U1730 ( .A(n3366), .Y(n3354) );
  INVX2TS U1731 ( .A(n3631), .Y(n3623) );
  INVX2TS U1732 ( .A(n3631), .Y(n3622) );
  INVX2TS U1733 ( .A(n3631), .Y(n3621) );
  INVX2TS U1734 ( .A(n984), .Y(n3620) );
  INVX2TS U1735 ( .A(n984), .Y(n3619) );
  INVX2TS U1736 ( .A(n3283), .Y(n3272) );
  INVX2TS U1737 ( .A(n3282), .Y(n3273) );
  INVX2TS U1738 ( .A(n3283), .Y(n3271) );
  INVX2TS U1739 ( .A(n3285), .Y(n3276) );
  INVX2TS U1740 ( .A(n3284), .Y(n3277) );
  INVX2TS U1741 ( .A(n3283), .Y(n3278) );
  INVX2TS U1742 ( .A(n3282), .Y(n3274) );
  INVX2TS U1743 ( .A(n3282), .Y(n3275) );
  INVX2TS U1744 ( .A(n3196), .Y(n3195) );
  INVX2TS U1745 ( .A(n3367), .Y(n3351) );
  INVX2TS U1746 ( .A(n3367), .Y(n3352) );
  INVX2TS U1747 ( .A(n3632), .Y(n3616) );
  INVX2TS U1748 ( .A(n3632), .Y(n3617) );
  INVX2TS U1749 ( .A(n3284), .Y(n3268) );
  INVX2TS U1750 ( .A(n3284), .Y(n3269) );
  CLKBUFX2TS U1751 ( .A(n3399), .Y(n3393) );
  CLKBUFX2TS U1752 ( .A(n3398), .Y(n3395) );
  CLKBUFX2TS U1753 ( .A(n3399), .Y(n3394) );
  CLKBUFX2TS U1754 ( .A(n3398), .Y(n3396) );
  CLKBUFX2TS U1755 ( .A(n682), .Y(n3807) );
  CLKBUFX2TS U1756 ( .A(n682), .Y(n3808) );
  CLKBUFX2TS U1757 ( .A(n3514), .Y(n3503) );
  CLKBUFX2TS U1758 ( .A(n3397), .Y(n3386) );
  CLKBUFX2TS U1759 ( .A(n3398), .Y(n3397) );
  CLKBUFX2TS U1760 ( .A(n3511), .Y(n3507) );
  CLKBUFX2TS U1761 ( .A(n3510), .Y(n3508) );
  CLKBUFX2TS U1762 ( .A(n3512), .Y(n3504) );
  CLKBUFX2TS U1763 ( .A(n3511), .Y(n3506) );
  CLKBUFX2TS U1764 ( .A(n3512), .Y(n3505) );
  CLKBUFX2TS U1765 ( .A(n3510), .Y(n3509) );
  CLKBUFX2TS U1766 ( .A(n3081), .Y(n3080) );
  CLKBUFX2TS U1767 ( .A(n3086), .Y(n3071) );
  CLKBUFX2TS U1768 ( .A(n3086), .Y(n3072) );
  CLKBUFX2TS U1769 ( .A(n3085), .Y(n3073) );
  CLKBUFX2TS U1770 ( .A(n3085), .Y(n3074) );
  CLKBUFX2TS U1771 ( .A(n3083), .Y(n3075) );
  CLKBUFX2TS U1772 ( .A(n3083), .Y(n3076) );
  CLKBUFX2TS U1773 ( .A(n3081), .Y(n3079) );
  CLKBUFX2TS U1774 ( .A(n3082), .Y(n3077) );
  CLKBUFX2TS U1775 ( .A(n3082), .Y(n3078) );
  CLKBUFX2TS U1776 ( .A(n3103), .Y(n3089) );
  CLKBUFX2TS U1777 ( .A(n3103), .Y(n3088) );
  CLKBUFX2TS U1778 ( .A(n3098), .Y(n3097) );
  CLKBUFX2TS U1779 ( .A(n3098), .Y(n3096) );
  CLKBUFX2TS U1780 ( .A(n3099), .Y(n3095) );
  CLKBUFX2TS U1781 ( .A(n3099), .Y(n3094) );
  CLKBUFX2TS U1782 ( .A(n3101), .Y(n3093) );
  CLKBUFX2TS U1783 ( .A(n3102), .Y(n3090) );
  CLKBUFX2TS U1784 ( .A(n3101), .Y(n3092) );
  CLKBUFX2TS U1785 ( .A(n3102), .Y(n3091) );
  INVX2TS U1786 ( .A(n3050), .Y(n3049) );
  INVX2TS U1787 ( .A(n3051), .Y(n3048) );
  INVX2TS U1788 ( .A(n3052), .Y(n3047) );
  CLKBUFX2TS U1789 ( .A(n1074), .Y(n1062) );
  CLKBUFX2TS U1790 ( .A(n1074), .Y(n1063) );
  CLKBUFX2TS U1791 ( .A(n1073), .Y(n1064) );
  CLKBUFX2TS U1792 ( .A(n1075), .Y(n1065) );
  CLKBUFX2TS U1793 ( .A(n1073), .Y(n1066) );
  CLKBUFX2TS U1794 ( .A(n1072), .Y(n1067) );
  CLKBUFX2TS U1795 ( .A(n1071), .Y(n1070) );
  CLKBUFX2TS U1796 ( .A(n1072), .Y(n1068) );
  CLKBUFX2TS U1797 ( .A(n1071), .Y(n1069) );
  CLKBUFX2TS U1798 ( .A(n3793), .Y(n3781) );
  CLKBUFX2TS U1799 ( .A(n3793), .Y(n3782) );
  CLKBUFX2TS U1800 ( .A(n1060), .Y(n1048) );
  CLKBUFX2TS U1801 ( .A(n3792), .Y(n3783) );
  CLKBUFX2TS U1802 ( .A(n1060), .Y(n1049) );
  CLKBUFX2TS U1803 ( .A(n1059), .Y(n1050) );
  CLKBUFX2TS U1804 ( .A(n1061), .Y(n1051) );
  CLKBUFX2TS U1805 ( .A(n3791), .Y(n3784) );
  CLKBUFX2TS U1806 ( .A(n1059), .Y(n1052) );
  CLKBUFX2TS U1807 ( .A(n3791), .Y(n3785) );
  CLKBUFX2TS U1808 ( .A(n1058), .Y(n1053) );
  CLKBUFX2TS U1809 ( .A(n3789), .Y(n3788) );
  CLKBUFX2TS U1810 ( .A(n1057), .Y(n1056) );
  CLKBUFX2TS U1811 ( .A(n3790), .Y(n3786) );
  CLKBUFX2TS U1812 ( .A(n1058), .Y(n1054) );
  CLKBUFX2TS U1813 ( .A(n3790), .Y(n3787) );
  CLKBUFX2TS U1814 ( .A(n1057), .Y(n1055) );
  CLKBUFX2TS U1815 ( .A(n1045), .Y(n1034) );
  CLKBUFX2TS U1816 ( .A(n1043), .Y(n1035) );
  CLKBUFX2TS U1817 ( .A(n1043), .Y(n1036) );
  CLKBUFX2TS U1818 ( .A(n1042), .Y(n1037) );
  CLKBUFX2TS U1819 ( .A(n1041), .Y(n1040) );
  CLKBUFX2TS U1820 ( .A(n1042), .Y(n1038) );
  CLKBUFX2TS U1821 ( .A(n1041), .Y(n1039) );
  CLKBUFX2TS U1822 ( .A(n1002), .Y(n991) );
  CLKBUFX2TS U1823 ( .A(n1017), .Y(n1005) );
  CLKBUFX2TS U1824 ( .A(n2115), .Y(n1006) );
  CLKBUFX2TS U1825 ( .A(n1016), .Y(n1007) );
  CLKBUFX2TS U1826 ( .A(n1016), .Y(n1008) );
  CLKBUFX2TS U1827 ( .A(n1000), .Y(n992) );
  CLKBUFX2TS U1828 ( .A(n1000), .Y(n993) );
  CLKBUFX2TS U1829 ( .A(n1018), .Y(n1009) );
  CLKBUFX2TS U1830 ( .A(n999), .Y(n994) );
  CLKBUFX2TS U1831 ( .A(n1015), .Y(n1010) );
  CLKBUFX2TS U1832 ( .A(n998), .Y(n997) );
  CLKBUFX2TS U1833 ( .A(n1014), .Y(n1013) );
  CLKBUFX2TS U1834 ( .A(n999), .Y(n995) );
  CLKBUFX2TS U1835 ( .A(n1015), .Y(n1011) );
  CLKBUFX2TS U1836 ( .A(n998), .Y(n996) );
  CLKBUFX2TS U1837 ( .A(n1014), .Y(n1012) );
  CLKBUFX2TS U1838 ( .A(n1032), .Y(n1019) );
  CLKBUFX2TS U1839 ( .A(n2917), .Y(n1934) );
  CLKBUFX2TS U1840 ( .A(n2114), .Y(n1020) );
  CLKBUFX2TS U1841 ( .A(n2917), .Y(n1980) );
  CLKBUFX2TS U1842 ( .A(n1031), .Y(n1021) );
  CLKBUFX2TS U1843 ( .A(n2916), .Y(n2103) );
  CLKBUFX2TS U1844 ( .A(n1031), .Y(n1022) );
  CLKBUFX2TS U1845 ( .A(n2918), .Y(n2377) );
  CLKBUFX2TS U1846 ( .A(n1033), .Y(n1024) );
  CLKBUFX2TS U1847 ( .A(n2916), .Y(n2909) );
  CLKBUFX2TS U1848 ( .A(n1030), .Y(n1025) );
  CLKBUFX2TS U1849 ( .A(n2915), .Y(n2910) );
  CLKBUFX2TS U1850 ( .A(n1029), .Y(n1028) );
  CLKBUFX2TS U1851 ( .A(n2914), .Y(n2913) );
  CLKBUFX2TS U1852 ( .A(n1030), .Y(n1026) );
  CLKBUFX2TS U1853 ( .A(n2915), .Y(n2911) );
  CLKBUFX2TS U1854 ( .A(n1029), .Y(n1027) );
  CLKBUFX2TS U1855 ( .A(n2914), .Y(n2912) );
  CLKBUFX2TS U1856 ( .A(n1771), .Y(n1076) );
  CLKBUFX2TS U1857 ( .A(n1771), .Y(n1077) );
  CLKBUFX2TS U1858 ( .A(n1749), .Y(n1079) );
  CLKBUFX2TS U1859 ( .A(n1807), .Y(n1085) );
  CLKBUFX2TS U1860 ( .A(n1749), .Y(n1102) );
  CLKBUFX2TS U1861 ( .A(n1611), .Y(n1129) );
  CLKBUFX2TS U1862 ( .A(n1210), .Y(n1193) );
  CLKBUFX2TS U1863 ( .A(n1611), .Y(n1146) );
  CLKBUFX2TS U1864 ( .A(n1210), .Y(n1162) );
  CLKBUFX2TS U1865 ( .A(n3201), .Y(n3199) );
  CLKBUFX2TS U1866 ( .A(n1100), .Y(n3730) );
  CLKBUFX2TS U1867 ( .A(n664), .Y(n3923) );
  CLKBUFX2TS U1868 ( .A(n1098), .Y(n3757) );
  CLKBUFX2TS U1869 ( .A(n1134), .Y(n3584) );
  CLKBUFX2TS U1870 ( .A(n3219), .Y(n3213) );
  INVX2TS U1871 ( .A(n1760), .Y(n686) );
  CLKBUFX2TS U1872 ( .A(n1151), .Y(n3502) );
  CLKBUFX2TS U1873 ( .A(n1151), .Y(n3501) );
  CLKBUFX2TS U1874 ( .A(n1100), .Y(n3731) );
  CLKBUFX2TS U1875 ( .A(n1101), .Y(n3714) );
  CLKBUFX2TS U1876 ( .A(n1116), .Y(n3681) );
  CLKBUFX2TS U1877 ( .A(n1149), .Y(n3533) );
  CLKBUFX2TS U1878 ( .A(n1098), .Y(n3763) );
  CLKBUFX2TS U1879 ( .A(n1135), .Y(n3566) );
  CLKBUFX2TS U1880 ( .A(n1135), .Y(n3567) );
  CLKBUFX2TS U1881 ( .A(n1216), .Y(n3218) );
  CLKBUFX2TS U1882 ( .A(n1216), .Y(n3219) );
  CLKBUFX2TS U1883 ( .A(n1132), .Y(n3615) );
  CLKBUFX2TS U1884 ( .A(n1198), .Y(n3319) );
  CLKBUFX2TS U1885 ( .A(n1196), .Y(n3349) );
  CLKBUFX2TS U1886 ( .A(n1132), .Y(n3614) );
  CLKBUFX2TS U1887 ( .A(n1196), .Y(n3350) );
  CLKBUFX2TS U1888 ( .A(n1198), .Y(n3318) );
  CLKBUFX2TS U1889 ( .A(n1118), .Y(n3650) );
  CLKBUFX2TS U1890 ( .A(n668), .Y(n3893) );
  CLKBUFX2TS U1891 ( .A(n1134), .Y(n3583) );
  CLKBUFX2TS U1892 ( .A(n1134), .Y(n3582) );
  CLKBUFX2TS U1893 ( .A(n1199), .Y(n3302) );
  INVX2TS U1894 ( .A(n2890), .Y(n951) );
  INVX2TS U1895 ( .A(n1790), .Y(n696) );
  CLKBUFX2TS U1896 ( .A(n1166), .Y(n3450) );
  CLKBUFX2TS U1897 ( .A(n681), .Y(n3810) );
  CLKBUFX2TS U1898 ( .A(n681), .Y(n3811) );
  CLKBUFX2TS U1899 ( .A(n3778), .Y(n3777) );
  CLKBUFX2TS U1900 ( .A(n3732), .Y(n3725) );
  CLKBUFX2TS U1901 ( .A(n1100), .Y(n3732) );
  CLKBUFX2TS U1902 ( .A(n3715), .Y(n3708) );
  CLKBUFX2TS U1903 ( .A(n1101), .Y(n3715) );
  CLKBUFX2TS U1904 ( .A(n982), .Y(n3697) );
  CLKBUFX2TS U1905 ( .A(n983), .Y(n3549) );
  CLKBUFX2TS U1906 ( .A(n982), .Y(n3698) );
  CLKBUFX2TS U1907 ( .A(n983), .Y(n3550) );
  CLKBUFX2TS U1908 ( .A(n3368), .Y(n3367) );
  CLKBUFX2TS U1909 ( .A(n3633), .Y(n3632) );
  CLKBUFX2TS U1910 ( .A(n3285), .Y(n3284) );
  CLKBUFX2TS U1911 ( .A(n3663), .Y(n3661) );
  CLKBUFX2TS U1912 ( .A(n3664), .Y(n3659) );
  CLKBUFX2TS U1913 ( .A(n3745), .Y(n3743) );
  CLKBUFX2TS U1914 ( .A(n3745), .Y(n3742) );
  CLKBUFX2TS U1915 ( .A(n3746), .Y(n3741) );
  CLKBUFX2TS U1916 ( .A(n3746), .Y(n3740) );
  CLKBUFX2TS U1917 ( .A(n3746), .Y(n3739) );
  CLKBUFX2TS U1918 ( .A(n3664), .Y(n3660) );
  CLKBUFX2TS U1919 ( .A(n3664), .Y(n3658) );
  CLKBUFX2TS U1920 ( .A(n3598), .Y(n3595) );
  CLKBUFX2TS U1921 ( .A(n3598), .Y(n3596) );
  CLKBUFX2TS U1922 ( .A(n3598), .Y(n3594) );
  CLKBUFX2TS U1923 ( .A(n3070), .Y(n3065) );
  CLKBUFX2TS U1924 ( .A(n3069), .Y(n3066) );
  CLKBUFX2TS U1925 ( .A(n3069), .Y(n3067) );
  CLKBUFX2TS U1926 ( .A(n3779), .Y(n3774) );
  CLKBUFX2TS U1927 ( .A(n3779), .Y(n3775) );
  CLKBUFX2TS U1928 ( .A(n3779), .Y(n3776) );
  CLKBUFX2TS U1929 ( .A(n1197), .Y(n3333) );
  CLKBUFX2TS U1930 ( .A(n1215), .Y(n3233) );
  CLKBUFX2TS U1931 ( .A(n1215), .Y(n3232) );
  CLKBUFX2TS U1932 ( .A(n3119), .Y(n3117) );
  CLKBUFX2TS U1933 ( .A(n3119), .Y(n3118) );
  CLKBUFX2TS U1934 ( .A(n3744), .Y(n3733) );
  CLKBUFX2TS U1935 ( .A(n3745), .Y(n3744) );
  CLKBUFX2TS U1936 ( .A(n1133), .Y(n3597) );
  CLKBUFX2TS U1937 ( .A(n3202), .Y(n3200) );
  CLKBUFX2TS U1938 ( .A(n3068), .Y(n3055) );
  CLKBUFX2TS U1939 ( .A(n3069), .Y(n3068) );
  CLKBUFX2TS U1940 ( .A(n3773), .Y(n3771) );
  CLKBUFX2TS U1941 ( .A(n3064), .Y(n3063) );
  CLKBUFX2TS U1942 ( .A(n3064), .Y(n3062) );
  CLKBUFX2TS U1943 ( .A(n3773), .Y(n3772) );
  INVX2TS U1944 ( .A(n985), .Y(n3363) );
  INVX2TS U1945 ( .A(n985), .Y(n3362) );
  INVX2TS U1946 ( .A(n3631), .Y(n3628) );
  INVX2TS U1947 ( .A(n3632), .Y(n3627) );
  CLKBUFX2TS U1948 ( .A(n988), .Y(n3050) );
  CLKBUFX2TS U1949 ( .A(n3053), .Y(n3051) );
  CLKBUFX2TS U1950 ( .A(n988), .Y(n3052) );
  CLKBUFX2TS U1951 ( .A(n3663), .Y(n3662) );
  CLKBUFX2TS U1952 ( .A(n3104), .Y(n3103) );
  CLKBUFX2TS U1953 ( .A(n2034), .Y(n3086) );
  CLKBUFX2TS U1954 ( .A(n3104), .Y(n3098) );
  CLKBUFX2TS U1955 ( .A(n2034), .Y(n3085) );
  CLKBUFX2TS U1956 ( .A(n2033), .Y(n3099) );
  CLKBUFX2TS U1957 ( .A(n3081), .Y(n3084) );
  CLKBUFX2TS U1958 ( .A(n3087), .Y(n3083) );
  CLKBUFX2TS U1959 ( .A(n2033), .Y(n3100) );
  CLKBUFX2TS U1960 ( .A(n3087), .Y(n3081) );
  CLKBUFX2TS U1961 ( .A(n3104), .Y(n3101) );
  CLKBUFX2TS U1962 ( .A(n3104), .Y(n3102) );
  CLKBUFX2TS U1963 ( .A(n3087), .Y(n3082) );
  CLKBUFX2TS U1964 ( .A(n3515), .Y(n3514) );
  CLKBUFX2TS U1965 ( .A(n3515), .Y(n3513) );
  CLKBUFX2TS U1966 ( .A(n3516), .Y(n3511) );
  CLKBUFX2TS U1967 ( .A(n3516), .Y(n3512) );
  CLKBUFX2TS U1968 ( .A(n3516), .Y(n3510) );
  CLKBUFX2TS U1969 ( .A(n1181), .Y(n3399) );
  CLKBUFX2TS U1970 ( .A(n1181), .Y(n3398) );
  INVX2TS U1971 ( .A(n1800), .Y(n695) );
  CLKBUFX2TS U1972 ( .A(n4237), .Y(n4239) );
  CLKBUFX2TS U1973 ( .A(n4240), .Y(n4242) );
  INVX2TS U1974 ( .A(n3052), .Y(n2919) );
  INVX2TS U1975 ( .A(n3053), .Y(n2920) );
  CLKBUFX2TS U1976 ( .A(n988), .Y(n3053) );
  INVX2TS U1977 ( .A(n3053), .Y(n3003) );
  INVX2TS U1978 ( .A(n3054), .Y(n3004) );
  INVX2TS U1979 ( .A(n3054), .Y(n3005) );
  INVX2TS U1980 ( .A(n3053), .Y(n3044) );
  INVX2TS U1981 ( .A(n3054), .Y(n3045) );
  INVX2TS U1982 ( .A(n3054), .Y(n3046) );
  CLKBUFX2TS U1983 ( .A(n3794), .Y(n3793) );
  CLKBUFX2TS U1984 ( .A(n1061), .Y(n1060) );
  CLKBUFX2TS U1985 ( .A(n1075), .Y(n1074) );
  CLKBUFX2TS U1986 ( .A(n1093), .Y(n3792) );
  CLKBUFX2TS U1987 ( .A(n2112), .Y(n1059) );
  CLKBUFX2TS U1988 ( .A(n2111), .Y(n1073) );
  CLKBUFX2TS U1989 ( .A(n3794), .Y(n3791) );
  CLKBUFX2TS U1990 ( .A(n3794), .Y(n3789) );
  CLKBUFX2TS U1991 ( .A(n1061), .Y(n1058) );
  CLKBUFX2TS U1992 ( .A(n1075), .Y(n1072) );
  CLKBUFX2TS U1993 ( .A(n3794), .Y(n3790) );
  CLKBUFX2TS U1994 ( .A(n1061), .Y(n1057) );
  CLKBUFX2TS U1995 ( .A(n1075), .Y(n1071) );
  CLKBUFX2TS U1996 ( .A(n1003), .Y(n1002) );
  CLKBUFX2TS U1997 ( .A(n1046), .Y(n1045) );
  CLKBUFX2TS U1998 ( .A(n1807), .Y(n1771) );
  CLKBUFX2TS U1999 ( .A(n2918), .Y(n2917) );
  CLKBUFX2TS U2000 ( .A(n1003), .Y(n1001) );
  CLKBUFX2TS U2001 ( .A(n1018), .Y(n1016) );
  CLKBUFX2TS U2002 ( .A(n1033), .Y(n1031) );
  CLKBUFX2TS U2003 ( .A(n1046), .Y(n1044) );
  CLKBUFX2TS U2004 ( .A(n2109), .Y(n1749) );
  CLKBUFX2TS U2005 ( .A(n2108), .Y(n2916) );
  CLKBUFX2TS U2006 ( .A(n1004), .Y(n1000) );
  CLKBUFX2TS U2007 ( .A(n1047), .Y(n1043) );
  CLKBUFX2TS U2008 ( .A(n1004), .Y(n999) );
  CLKBUFX2TS U2009 ( .A(n1018), .Y(n1015) );
  CLKBUFX2TS U2010 ( .A(n1033), .Y(n1030) );
  CLKBUFX2TS U2011 ( .A(n1047), .Y(n1042) );
  CLKBUFX2TS U2012 ( .A(n1807), .Y(n1611) );
  CLKBUFX2TS U2013 ( .A(n2918), .Y(n2915) );
  CLKBUFX2TS U2014 ( .A(n1004), .Y(n998) );
  CLKBUFX2TS U2015 ( .A(n1018), .Y(n1014) );
  CLKBUFX2TS U2016 ( .A(n1033), .Y(n1029) );
  CLKBUFX2TS U2017 ( .A(n1047), .Y(n1041) );
  CLKBUFX2TS U2018 ( .A(n1807), .Y(n1210) );
  CLKBUFX2TS U2019 ( .A(n2918), .Y(n2914) );
  CLKBUFX2TS U2020 ( .A(n4240), .Y(n4241) );
  CLKBUFX2TS U2021 ( .A(n4237), .Y(n4238) );
  CLKBUFX2TS U2022 ( .A(n2115), .Y(n1017) );
  CLKBUFX2TS U2023 ( .A(n2114), .Y(n1032) );
  INVX2TS U2024 ( .A(n4215), .Y(n4212) );
  NOR2BX1TS U2025 ( .AN(n125), .B(n1935), .Y(n1774) );
  OAI211X1TS U2026 ( .A0(n120), .A1(n125), .B0(n163), .C0(n1935), .Y(n1783) );
  NOR2BX1TS U2027 ( .AN(n1769), .B(n1770), .Y(n1116) );
  AOI2BB1X1TS U2028 ( .A0N(n691), .A1N(n1909), .B0(n1813), .Y(n1811) );
  NOR2X1TS U2029 ( .A(n1760), .B(n1764), .Y(n1100) );
  NOR2X1TS U2030 ( .A(n117), .B(n126), .Y(n1801) );
  NOR2X1TS U2031 ( .A(n125), .B(n1935), .Y(n1789) );
  INVX2TS U2032 ( .A(n1866), .Y(n944) );
  INVX2TS U2033 ( .A(n1785), .Y(n667) );
  NAND2X1TS U2034 ( .A(n951), .B(n2386), .Y(n2388) );
  AND3X2TS U2035 ( .A(n132), .B(n1775), .C(n103), .Y(n1134) );
  NAND2X1TS U2036 ( .A(n700), .B(n1826), .Y(n1923) );
  NAND2X1TS U2037 ( .A(n1935), .B(n1958), .Y(n1798) );
  INVX2TS U2038 ( .A(n2001), .Y(n946) );
  INVX2TS U2039 ( .A(n483), .Y(n668) );
  INVX2TS U2040 ( .A(n1863), .Y(n697) );
  NOR2BX1TS U2041 ( .AN(n1854), .B(n1971), .Y(n1215) );
  NAND2BX1TS U2042 ( .AN(n2385), .B(n2386), .Y(n2384) );
  INVX2TS U2043 ( .A(n2002), .Y(n692) );
  NAND2X1TS U2044 ( .A(n2001), .B(n126), .Y(n1909) );
  CLKBUFX2TS U2045 ( .A(n3121), .Y(n3120) );
  CLKBUFX2TS U2046 ( .A(n3121), .Y(n3119) );
  CLKBUFX2TS U2047 ( .A(n987), .Y(n3202) );
  CLKBUFX2TS U2048 ( .A(n985), .Y(n3368) );
  CLKBUFX2TS U2049 ( .A(n984), .Y(n3633) );
  CLKBUFX2TS U2050 ( .A(n986), .Y(n3285) );
  CLKBUFX2TS U2051 ( .A(n2048), .Y(n3069) );
  CLKBUFX2TS U2052 ( .A(n1095), .Y(n3779) );
  CLKBUFX2TS U2053 ( .A(n1117), .Y(n3663) );
  CLKBUFX2TS U2054 ( .A(n1099), .Y(n3746) );
  CLKBUFX2TS U2055 ( .A(n1117), .Y(n3664) );
  CLKBUFX2TS U2056 ( .A(n1099), .Y(n3745) );
  CLKBUFX2TS U2057 ( .A(n1133), .Y(n3598) );
  CLKBUFX2TS U2058 ( .A(n3070), .Y(n3064) );
  CLKBUFX2TS U2059 ( .A(n2048), .Y(n3070) );
  CLKBUFX2TS U2060 ( .A(n3780), .Y(n3773) );
  CLKBUFX2TS U2061 ( .A(n1095), .Y(n3780) );
  NOR2BX1TS U2062 ( .AN(n1854), .B(n1933), .Y(n1181) );
  INVX2TS U2063 ( .A(n2045), .Y(n954) );
  CLKBUFX2TS U2064 ( .A(destinationAddressIn_SOUTH[7]), .Y(n4240) );
  CLKBUFX2TS U2065 ( .A(destinationAddressIn_SOUTH[6]), .Y(n4237) );
  CLKBUFX2TS U2066 ( .A(n2033), .Y(n3104) );
  CLKBUFX2TS U2067 ( .A(n1150), .Y(n3515) );
  CLKBUFX2TS U2068 ( .A(n1150), .Y(n3516) );
  CLKBUFX2TS U2069 ( .A(n2034), .Y(n3087) );
  CLKBUFX2TS U2070 ( .A(n988), .Y(n3054) );
  INVX2TS U2071 ( .A(n4208), .Y(n4206) );
  CLKBUFX2TS U2072 ( .A(n1093), .Y(n3794) );
  CLKBUFX2TS U2073 ( .A(n2112), .Y(n1061) );
  CLKBUFX2TS U2074 ( .A(n2111), .Y(n1075) );
  CLKBUFX2TS U2075 ( .A(n2117), .Y(n1003) );
  CLKBUFX2TS U2076 ( .A(n2113), .Y(n1046) );
  CLKBUFX2TS U2077 ( .A(n2117), .Y(n1004) );
  CLKBUFX2TS U2078 ( .A(n2115), .Y(n1018) );
  CLKBUFX2TS U2079 ( .A(n2114), .Y(n1033) );
  CLKBUFX2TS U2080 ( .A(n2113), .Y(n1047) );
  CLKBUFX2TS U2081 ( .A(n2109), .Y(n1807) );
  CLKBUFX2TS U2082 ( .A(n2108), .Y(n2918) );
  CLKBUFX2TS U2083 ( .A(n4182), .Y(n4183) );
  CLKBUFX2TS U2084 ( .A(n4137), .Y(n4138) );
  CLKBUFX2TS U2085 ( .A(n4134), .Y(n4135) );
  CLKBUFX2TS U2086 ( .A(n4122), .Y(n4123) );
  CLKBUFX2TS U2087 ( .A(n4092), .Y(n4093) );
  CLKBUFX2TS U2088 ( .A(n4179), .Y(n4180) );
  CLKBUFX2TS U2089 ( .A(n4176), .Y(n4177) );
  CLKBUFX2TS U2090 ( .A(n4173), .Y(n4174) );
  CLKBUFX2TS U2091 ( .A(n4170), .Y(n4171) );
  CLKBUFX2TS U2092 ( .A(n4167), .Y(n4168) );
  CLKBUFX2TS U2093 ( .A(n4164), .Y(n4165) );
  CLKBUFX2TS U2094 ( .A(n4161), .Y(n4162) );
  CLKBUFX2TS U2095 ( .A(n4158), .Y(n4159) );
  CLKBUFX2TS U2096 ( .A(n4155), .Y(n4156) );
  CLKBUFX2TS U2097 ( .A(n4152), .Y(n4153) );
  CLKBUFX2TS U2098 ( .A(n4149), .Y(n4150) );
  CLKBUFX2TS U2099 ( .A(n4146), .Y(n4147) );
  CLKBUFX2TS U2100 ( .A(n4143), .Y(n4144) );
  CLKBUFX2TS U2101 ( .A(n4140), .Y(n4141) );
  CLKBUFX2TS U2102 ( .A(n4131), .Y(n4132) );
  CLKBUFX2TS U2103 ( .A(n4128), .Y(n4129) );
  CLKBUFX2TS U2104 ( .A(n4125), .Y(n4126) );
  CLKBUFX2TS U2105 ( .A(n4119), .Y(n4120) );
  CLKBUFX2TS U2106 ( .A(n4116), .Y(n4117) );
  CLKBUFX2TS U2107 ( .A(n4113), .Y(n4114) );
  CLKBUFX2TS U2108 ( .A(n4110), .Y(n4111) );
  CLKBUFX2TS U2109 ( .A(n4107), .Y(n4108) );
  CLKBUFX2TS U2110 ( .A(n4104), .Y(n4105) );
  CLKBUFX2TS U2111 ( .A(n4101), .Y(n4102) );
  CLKBUFX2TS U2112 ( .A(n4098), .Y(n4099) );
  CLKBUFX2TS U2113 ( .A(n4095), .Y(n4096) );
  CLKBUFX2TS U2114 ( .A(n4089), .Y(n4090) );
  INVX2TS U2115 ( .A(n4001), .Y(n3999) );
  INVX2TS U2116 ( .A(n4353), .Y(n4351) );
  INVX2TS U2117 ( .A(n4350), .Y(n4348) );
  INVX2TS U2118 ( .A(n4341), .Y(n4339) );
  INVX2TS U2119 ( .A(n4338), .Y(n4336) );
  INVX2TS U2120 ( .A(n4326), .Y(n4324) );
  INVX2TS U2121 ( .A(n4320), .Y(n4318) );
  INVX2TS U2122 ( .A(n4317), .Y(n4315) );
  INVX2TS U2123 ( .A(n4314), .Y(n4312) );
  INVX2TS U2124 ( .A(n4308), .Y(n4306) );
  INVX2TS U2125 ( .A(n4305), .Y(n4303) );
  INVX2TS U2126 ( .A(n4302), .Y(n4300) );
  INVX2TS U2127 ( .A(n4299), .Y(n4297) );
  INVX2TS U2128 ( .A(n4296), .Y(n4294) );
  INVX2TS U2129 ( .A(n4287), .Y(n4285) );
  INVX2TS U2130 ( .A(n4284), .Y(n4282) );
  INVX2TS U2131 ( .A(n4275), .Y(n4273) );
  INVX2TS U2132 ( .A(n4272), .Y(n4270) );
  INVX2TS U2133 ( .A(n4010), .Y(n4008) );
  INVX2TS U2134 ( .A(n4007), .Y(n4005) );
  INVX2TS U2135 ( .A(n4004), .Y(n4002) );
  INVX2TS U2136 ( .A(n3998), .Y(n3996) );
  INVX2TS U2137 ( .A(n3995), .Y(n3993) );
  INVX2TS U2138 ( .A(n4293), .Y(n4291) );
  INVX2TS U2139 ( .A(n4347), .Y(n4345) );
  INVX2TS U2140 ( .A(n4344), .Y(n4342) );
  INVX2TS U2141 ( .A(n4332), .Y(n4330) );
  INVX2TS U2142 ( .A(n4323), .Y(n4321) );
  INVX2TS U2143 ( .A(n4290), .Y(n4288) );
  INVX2TS U2144 ( .A(n4278), .Y(n4276) );
  INVX2TS U2145 ( .A(n4266), .Y(n4264) );
  INVX2TS U2146 ( .A(n4356), .Y(n4354) );
  INVX2TS U2147 ( .A(n4335), .Y(n4333) );
  INVX2TS U2148 ( .A(n4329), .Y(n4327) );
  INVX2TS U2149 ( .A(n4311), .Y(n4309) );
  INVX2TS U2150 ( .A(n4281), .Y(n4279) );
  INVX2TS U2151 ( .A(n4269), .Y(n4267) );
  INVX2TS U2152 ( .A(n4263), .Y(n4261) );
  CLKBUFX2TS U2153 ( .A(n4578), .Y(n4579) );
  CLKBUFX2TS U2154 ( .A(n4574), .Y(n4576) );
  CLKBUFX2TS U2155 ( .A(n4570), .Y(n4571) );
  CLKBUFX2TS U2156 ( .A(n4559), .Y(n4560) );
  CLKBUFX2TS U2157 ( .A(n4555), .Y(n4556) );
  CLKBUFX2TS U2158 ( .A(n4551), .Y(n4552) );
  CLKBUFX2TS U2159 ( .A(n4543), .Y(n4544) );
  CLKBUFX2TS U2160 ( .A(n4540), .Y(n4541) );
  CLKBUFX2TS U2161 ( .A(n4532), .Y(n4533) );
  CLKBUFX2TS U2162 ( .A(n4528), .Y(n4529) );
  CLKBUFX2TS U2163 ( .A(n4524), .Y(n4525) );
  CLKBUFX2TS U2164 ( .A(n4521), .Y(n4522) );
  CLKBUFX2TS U2165 ( .A(n4517), .Y(n4519) );
  CLKBUFX2TS U2166 ( .A(n4513), .Y(n4514) );
  CLKBUFX2TS U2167 ( .A(n4510), .Y(n4511) );
  CLKBUFX2TS U2168 ( .A(n4506), .Y(n4507) );
  CLKBUFX2TS U2169 ( .A(n4503), .Y(n4504) );
  CLKBUFX2TS U2170 ( .A(n4498), .Y(n4499) );
  CLKBUFX2TS U2171 ( .A(n4492), .Y(n4493) );
  CLKBUFX2TS U2172 ( .A(n4488), .Y(n4489) );
  CLKBUFX2TS U2173 ( .A(n4484), .Y(n4486) );
  CLKBUFX2TS U2174 ( .A(n4477), .Y(n4478) );
  CLKBUFX2TS U2175 ( .A(n4472), .Y(n4474) );
  CLKBUFX2TS U2176 ( .A(n4566), .Y(n4567) );
  CLKBUFX2TS U2177 ( .A(n4562), .Y(n4564) );
  CLKBUFX2TS U2178 ( .A(n4547), .Y(n4549) );
  CLKBUFX2TS U2179 ( .A(n4535), .Y(n4537) );
  CLKBUFX2TS U2180 ( .A(n4495), .Y(n4496) );
  CLKBUFX2TS U2181 ( .A(n4480), .Y(n4481) );
  CLKBUFX2TS U2182 ( .A(n4468), .Y(n4470) );
  CLKBUFX2TS U2183 ( .A(n4465), .Y(n4466) );
  CLKBUFX2TS U2184 ( .A(n4461), .Y(n4462) );
  INVX2TS U2185 ( .A(n4049), .Y(n4047) );
  INVX2TS U2186 ( .A(n4040), .Y(n4038) );
  INVX2TS U2187 ( .A(n4037), .Y(n4035) );
  INVX2TS U2188 ( .A(n4052), .Y(n4050) );
  INVX2TS U2189 ( .A(n4046), .Y(n4044) );
  INVX2TS U2190 ( .A(n4043), .Y(n4041) );
  CLKBUFX2TS U2191 ( .A(n4068), .Y(n4069) );
  CLKBUFX2TS U2192 ( .A(n4062), .Y(n4063) );
  CLKBUFX2TS U2193 ( .A(n4059), .Y(n4060) );
  CLKBUFX2TS U2194 ( .A(n4056), .Y(n4057) );
  CLKBUFX2TS U2195 ( .A(n4053), .Y(n4054) );
  CLKBUFX2TS U2196 ( .A(n4065), .Y(n4066) );
  CLKBUFX2TS U2197 ( .A(n4083), .Y(n4084) );
  CLKBUFX2TS U2198 ( .A(n4086), .Y(n4087) );
  CLKBUFX2TS U2199 ( .A(n4080), .Y(n4081) );
  CLKBUFX2TS U2200 ( .A(n4077), .Y(n4078) );
  CLKBUFX2TS U2201 ( .A(n4074), .Y(n4075) );
  CLKBUFX2TS U2202 ( .A(n4071), .Y(n4072) );
  INVX2TS U2203 ( .A(n3965), .Y(n3963) );
  INVX2TS U2204 ( .A(n3968), .Y(n3966) );
  INVX2TS U2205 ( .A(n3962), .Y(n3960) );
  INVX2TS U2206 ( .A(n3959), .Y(n3957) );
  INVX2TS U2207 ( .A(n3956), .Y(n3954) );
  INVX2TS U2208 ( .A(n3953), .Y(n3951) );
  INVX2TS U2209 ( .A(n4457), .Y(n4454) );
  INVX2TS U2210 ( .A(n4450), .Y(n4448) );
  INVX2TS U2211 ( .A(n4447), .Y(n4443) );
  INVX2TS U2212 ( .A(n4442), .Y(n4440) );
  INVX2TS U2213 ( .A(n4439), .Y(n4436) );
  INVX2TS U2214 ( .A(n4435), .Y(n4432) );
  INVX2TS U2215 ( .A(n4431), .Y(n4429) );
  INVX2TS U2216 ( .A(n4413), .Y(n4411) );
  INVX2TS U2217 ( .A(n4398), .Y(n4396) );
  INVX2TS U2218 ( .A(n4386), .Y(n4384) );
  INVX2TS U2219 ( .A(n4380), .Y(n4378) );
  INVX2TS U2220 ( .A(n4374), .Y(n4372) );
  INVX2TS U2221 ( .A(n4371), .Y(n4369) );
  INVX2TS U2222 ( .A(n4365), .Y(n4363) );
  INVX2TS U2223 ( .A(n4460), .Y(n4458) );
  INVX2TS U2224 ( .A(n4453), .Y(n4451) );
  INVX2TS U2225 ( .A(n4427), .Y(n4425) );
  INVX2TS U2226 ( .A(n4424), .Y(n4422) );
  INVX2TS U2227 ( .A(n4421), .Y(n4417) );
  INVX2TS U2228 ( .A(n4416), .Y(n4414) );
  INVX2TS U2229 ( .A(n4407), .Y(n4405) );
  INVX2TS U2230 ( .A(n4395), .Y(n4393) );
  INVX2TS U2231 ( .A(n4392), .Y(n4390) );
  INVX2TS U2232 ( .A(n4389), .Y(n4387) );
  INVX2TS U2233 ( .A(n4383), .Y(n4381) );
  INVX2TS U2234 ( .A(n4377), .Y(n4375) );
  INVX2TS U2235 ( .A(n4362), .Y(n4360) );
  INVX2TS U2236 ( .A(n4359), .Y(n4357) );
  INVX2TS U2237 ( .A(n4410), .Y(n4408) );
  INVX2TS U2238 ( .A(n4404), .Y(n4402) );
  INVX2TS U2239 ( .A(n4401), .Y(n4399) );
  INVX2TS U2240 ( .A(n4368), .Y(n4366) );
  CLKBUFX2TS U2241 ( .A(n4234), .Y(n4235) );
  CLKBUFX2TS U2242 ( .A(n4228), .Y(n4229) );
  CLKBUFX2TS U2243 ( .A(n4225), .Y(n4226) );
  CLKBUFX2TS U2244 ( .A(n4222), .Y(n4223) );
  CLKBUFX2TS U2245 ( .A(n4231), .Y(n4232) );
  CLKBUFX2TS U2246 ( .A(n4219), .Y(n4220) );
  CLKBUFX2TS U2247 ( .A(n4602), .Y(n4603) );
  CLKBUFX2TS U2248 ( .A(n4593), .Y(n4594) );
  CLKBUFX2TS U2249 ( .A(n4597), .Y(n4598) );
  CLKBUFX2TS U2250 ( .A(n4589), .Y(n4591) );
  CLKBUFX2TS U2251 ( .A(n4585), .Y(n4586) );
  CLKBUFX2TS U2252 ( .A(n4582), .Y(n4583) );
  INVX2TS U2253 ( .A(n4202), .Y(n4200) );
  INVX2TS U2254 ( .A(n4196), .Y(n4194) );
  INVX2TS U2255 ( .A(n4199), .Y(n4197) );
  INVX2TS U2256 ( .A(n4193), .Y(n4191) );
  INVX2TS U2257 ( .A(n4190), .Y(n4188) );
  INVX2TS U2258 ( .A(n4187), .Y(n4185) );
  INVX2TS U2259 ( .A(n4208), .Y(n4207) );
  CLKBUFX2TS U2260 ( .A(n4252), .Y(n4253) );
  CLKBUFX2TS U2261 ( .A(n4216), .Y(n4217) );
  CLKBUFX2TS U2262 ( .A(n4258), .Y(n4259) );
  CLKBUFX2TS U2263 ( .A(n4246), .Y(n4247) );
  CLKBUFX2TS U2264 ( .A(n4255), .Y(n4256) );
  CLKBUFX2TS U2265 ( .A(n4249), .Y(n4250) );
  CLKBUFX2TS U2266 ( .A(n4243), .Y(n4244) );
  CLKBUFX2TS U2267 ( .A(n4574), .Y(n4577) );
  CLKBUFX2TS U2268 ( .A(n4566), .Y(n4569) );
  CLKBUFX2TS U2269 ( .A(n4562), .Y(n4565) );
  CLKBUFX2TS U2270 ( .A(n4559), .Y(n4561) );
  CLKBUFX2TS U2271 ( .A(n4555), .Y(n4558) );
  CLKBUFX2TS U2272 ( .A(n4551), .Y(n4553) );
  CLKBUFX2TS U2273 ( .A(n4547), .Y(n4550) );
  CLKBUFX2TS U2274 ( .A(n4528), .Y(n4531) );
  CLKBUFX2TS U2275 ( .A(n4510), .Y(n4512) );
  CLKBUFX2TS U2276 ( .A(n4495), .Y(n4497) );
  CLKBUFX2TS U2277 ( .A(n4488), .Y(n4490) );
  CLKBUFX2TS U2278 ( .A(n4480), .Y(n4483) );
  CLKBUFX2TS U2279 ( .A(n4477), .Y(n4479) );
  CLKBUFX2TS U2280 ( .A(n4468), .Y(n4471) );
  CLKBUFX2TS U2281 ( .A(n4578), .Y(n4580) );
  CLKBUFX2TS U2282 ( .A(n4570), .Y(n4573) );
  CLKBUFX2TS U2283 ( .A(n4543), .Y(n4546) );
  CLKBUFX2TS U2284 ( .A(n4540), .Y(n4542) );
  CLKBUFX2TS U2285 ( .A(n4535), .Y(n4538) );
  CLKBUFX2TS U2286 ( .A(n4532), .Y(n4534) );
  CLKBUFX2TS U2287 ( .A(n4521), .Y(n4523) );
  CLKBUFX2TS U2288 ( .A(n4506), .Y(n4508) );
  CLKBUFX2TS U2289 ( .A(n4503), .Y(n4505) );
  CLKBUFX2TS U2290 ( .A(n4498), .Y(n4502) );
  CLKBUFX2TS U2291 ( .A(n4492), .Y(n4494) );
  CLKBUFX2TS U2292 ( .A(n4484), .Y(n4487) );
  CLKBUFX2TS U2293 ( .A(n4465), .Y(n4467) );
  CLKBUFX2TS U2294 ( .A(n4461), .Y(n4463) );
  CLKBUFX2TS U2295 ( .A(n4524), .Y(n4526) );
  CLKBUFX2TS U2296 ( .A(n4517), .Y(n4520) );
  CLKBUFX2TS U2297 ( .A(n4513), .Y(n4515) );
  CLKBUFX2TS U2298 ( .A(n4472), .Y(n4475) );
  CLKBUFX2TS U2299 ( .A(n4231), .Y(n4233) );
  CLKBUFX2TS U2300 ( .A(n4234), .Y(n4236) );
  CLKBUFX2TS U2301 ( .A(n4228), .Y(n4230) );
  CLKBUFX2TS U2302 ( .A(n4225), .Y(n4227) );
  CLKBUFX2TS U2303 ( .A(n4222), .Y(n4224) );
  CLKBUFX2TS U2304 ( .A(n4219), .Y(n4221) );
  CLKBUFX2TS U2305 ( .A(n4597), .Y(n4601) );
  CLKBUFX2TS U2306 ( .A(n4585), .Y(n4587) );
  CLKBUFX2TS U2307 ( .A(n4582), .Y(n4584) );
  CLKBUFX2TS U2308 ( .A(n4602), .Y(n4604) );
  CLKBUFX2TS U2309 ( .A(n4593), .Y(n4596) );
  CLKBUFX2TS U2310 ( .A(n4589), .Y(n4592) );
  CLKBUFX2TS U2311 ( .A(n4255), .Y(n4257) );
  CLKBUFX2TS U2312 ( .A(n4252), .Y(n4254) );
  CLKBUFX2TS U2313 ( .A(n4246), .Y(n4248) );
  CLKBUFX2TS U2314 ( .A(n4243), .Y(n4245) );
  CLKBUFX2TS U2315 ( .A(n4258), .Y(n4260) );
  CLKBUFX2TS U2316 ( .A(n4249), .Y(n4251) );
  CLKBUFX2TS U2317 ( .A(n4216), .Y(n4218) );
  CLKBUFX2TS U2318 ( .A(n4065), .Y(n4067) );
  CLKBUFX2TS U2319 ( .A(n4068), .Y(n4070) );
  CLKBUFX2TS U2320 ( .A(n4062), .Y(n4064) );
  CLKBUFX2TS U2321 ( .A(n4059), .Y(n4061) );
  CLKBUFX2TS U2322 ( .A(n4056), .Y(n4058) );
  CLKBUFX2TS U2323 ( .A(n4053), .Y(n4055) );
  CLKBUFX2TS U2324 ( .A(n4179), .Y(n4181) );
  CLKBUFX2TS U2325 ( .A(n4173), .Y(n4175) );
  CLKBUFX2TS U2326 ( .A(n4170), .Y(n4172) );
  CLKBUFX2TS U2327 ( .A(n4167), .Y(n4169) );
  CLKBUFX2TS U2328 ( .A(n4164), .Y(n4166) );
  CLKBUFX2TS U2329 ( .A(n4161), .Y(n4163) );
  CLKBUFX2TS U2330 ( .A(n4158), .Y(n4160) );
  CLKBUFX2TS U2331 ( .A(n4143), .Y(n4145) );
  CLKBUFX2TS U2332 ( .A(n4128), .Y(n4130) );
  CLKBUFX2TS U2333 ( .A(n4116), .Y(n4118) );
  CLKBUFX2TS U2334 ( .A(n4110), .Y(n4112) );
  CLKBUFX2TS U2335 ( .A(n4104), .Y(n4106) );
  CLKBUFX2TS U2336 ( .A(n4101), .Y(n4103) );
  CLKBUFX2TS U2337 ( .A(n4095), .Y(n4097) );
  CLKBUFX2TS U2338 ( .A(n4182), .Y(n4184) );
  CLKBUFX2TS U2339 ( .A(n4176), .Y(n4178) );
  CLKBUFX2TS U2340 ( .A(n4155), .Y(n4157) );
  CLKBUFX2TS U2341 ( .A(n4152), .Y(n4154) );
  CLKBUFX2TS U2342 ( .A(n4149), .Y(n4151) );
  CLKBUFX2TS U2343 ( .A(n4146), .Y(n4148) );
  CLKBUFX2TS U2344 ( .A(n4137), .Y(n4139) );
  CLKBUFX2TS U2345 ( .A(n4125), .Y(n4127) );
  CLKBUFX2TS U2346 ( .A(n4122), .Y(n4124) );
  CLKBUFX2TS U2347 ( .A(n4119), .Y(n4121) );
  CLKBUFX2TS U2348 ( .A(n4113), .Y(n4115) );
  CLKBUFX2TS U2349 ( .A(n4107), .Y(n4109) );
  CLKBUFX2TS U2350 ( .A(n4092), .Y(n4094) );
  CLKBUFX2TS U2351 ( .A(n4089), .Y(n4091) );
  CLKBUFX2TS U2352 ( .A(n4140), .Y(n4142) );
  CLKBUFX2TS U2353 ( .A(n4134), .Y(n4136) );
  CLKBUFX2TS U2354 ( .A(n4131), .Y(n4133) );
  CLKBUFX2TS U2355 ( .A(n4098), .Y(n4100) );
  CLKBUFX2TS U2356 ( .A(n4083), .Y(n4085) );
  CLKBUFX2TS U2357 ( .A(n4074), .Y(n4076) );
  CLKBUFX2TS U2358 ( .A(n4071), .Y(n4073) );
  CLKBUFX2TS U2359 ( .A(n4086), .Y(n4088) );
  CLKBUFX2TS U2360 ( .A(n4080), .Y(n4082) );
  CLKBUFX2TS U2361 ( .A(n4077), .Y(n4079) );
  CLKBUFX2TS U2362 ( .A(n4215), .Y(n4214) );
  INVX2TS U2363 ( .A(n4010), .Y(n4009) );
  INVX2TS U2364 ( .A(n4004), .Y(n4003) );
  INVX2TS U2365 ( .A(n4001), .Y(n4000) );
  INVX2TS U2366 ( .A(n3998), .Y(n3997) );
  INVX2TS U2367 ( .A(n4007), .Y(n4006) );
  INVX2TS U2368 ( .A(n3995), .Y(n3994) );
  INVX2TS U2369 ( .A(n4052), .Y(n4051) );
  INVX2TS U2370 ( .A(n4046), .Y(n4045) );
  INVX2TS U2371 ( .A(n4049), .Y(n4048) );
  INVX2TS U2372 ( .A(n4043), .Y(n4042) );
  INVX2TS U2373 ( .A(n4040), .Y(n4039) );
  INVX2TS U2374 ( .A(n4037), .Y(n4036) );
  INVX2TS U2375 ( .A(n3986), .Y(n3984) );
  INVX2TS U2376 ( .A(n4205), .Y(n4203) );
  INVX2TS U2377 ( .A(n4013), .Y(n4011) );
  INVX2TS U2378 ( .A(n4016), .Y(n4014) );
  INVX2TS U2379 ( .A(n4211), .Y(n4209) );
  INVX2TS U2380 ( .A(n3992), .Y(n3990) );
  INVX2TS U2381 ( .A(n3980), .Y(n3978) );
  INVX2TS U2382 ( .A(n3974), .Y(n3972) );
  INVX2TS U2383 ( .A(n3989), .Y(n3987) );
  INVX2TS U2384 ( .A(n3983), .Y(n3981) );
  INVX2TS U2385 ( .A(n3977), .Y(n3975) );
  INVX2TS U2386 ( .A(n3971), .Y(n3969) );
  INVX2TS U2387 ( .A(n4460), .Y(n4459) );
  INVX2TS U2388 ( .A(n4457), .Y(n4456) );
  INVX2TS U2389 ( .A(n4453), .Y(n4452) );
  INVX2TS U2390 ( .A(n4442), .Y(n4441) );
  INVX2TS U2391 ( .A(n4439), .Y(n4438) );
  INVX2TS U2392 ( .A(n4435), .Y(n4434) );
  INVX2TS U2393 ( .A(n4427), .Y(n4426) );
  INVX2TS U2394 ( .A(n4424), .Y(n4423) );
  INVX2TS U2395 ( .A(n4416), .Y(n4415) );
  INVX2TS U2396 ( .A(n4413), .Y(n4412) );
  INVX2TS U2397 ( .A(n4410), .Y(n4409) );
  INVX2TS U2398 ( .A(n4407), .Y(n4406) );
  INVX2TS U2399 ( .A(n4404), .Y(n4403) );
  INVX2TS U2400 ( .A(n4401), .Y(n4400) );
  INVX2TS U2401 ( .A(n4398), .Y(n4397) );
  INVX2TS U2402 ( .A(n4395), .Y(n4394) );
  INVX2TS U2403 ( .A(n4392), .Y(n4391) );
  INVX2TS U2404 ( .A(n4389), .Y(n4388) );
  INVX2TS U2405 ( .A(n4383), .Y(n4382) );
  INVX2TS U2406 ( .A(n4380), .Y(n4379) );
  INVX2TS U2407 ( .A(n4377), .Y(n4376) );
  INVX2TS U2408 ( .A(n4371), .Y(n4370) );
  INVX2TS U2409 ( .A(n4368), .Y(n4367) );
  INVX2TS U2410 ( .A(n4450), .Y(n4449) );
  INVX2TS U2411 ( .A(n4447), .Y(n4445) );
  INVX2TS U2412 ( .A(n4431), .Y(n4430) );
  INVX2TS U2413 ( .A(n4421), .Y(n4418) );
  INVX2TS U2414 ( .A(n4386), .Y(n4385) );
  INVX2TS U2415 ( .A(n4374), .Y(n4373) );
  INVX2TS U2416 ( .A(n4365), .Y(n4364) );
  INVX2TS U2417 ( .A(n4362), .Y(n4361) );
  INVX2TS U2418 ( .A(n4359), .Y(n4358) );
  INVX2TS U2419 ( .A(n4211), .Y(n4210) );
  INVX2TS U2420 ( .A(n3989), .Y(n3988) );
  INVX2TS U2421 ( .A(n3986), .Y(n3985) );
  INVX2TS U2422 ( .A(n3980), .Y(n3979) );
  INVX2TS U2423 ( .A(n3977), .Y(n3976) );
  INVX2TS U2424 ( .A(n3971), .Y(n3970) );
  INVX2TS U2425 ( .A(n3992), .Y(n3991) );
  INVX2TS U2426 ( .A(n3983), .Y(n3982) );
  INVX2TS U2427 ( .A(n3974), .Y(n3973) );
  INVX2TS U2428 ( .A(n4205), .Y(n4204) );
  INVX2TS U2429 ( .A(n4016), .Y(n4015) );
  INVX2TS U2430 ( .A(n4013), .Y(n4012) );
  INVX2TS U2431 ( .A(n4356), .Y(n4355) );
  INVX2TS U2432 ( .A(n4353), .Y(n4352) );
  INVX2TS U2433 ( .A(n4350), .Y(n4349) );
  INVX2TS U2434 ( .A(n4347), .Y(n4346) );
  INVX2TS U2435 ( .A(n4344), .Y(n4343) );
  INVX2TS U2436 ( .A(n4341), .Y(n4340) );
  INVX2TS U2437 ( .A(n4338), .Y(n4337) );
  INVX2TS U2438 ( .A(n4335), .Y(n4334) );
  INVX2TS U2439 ( .A(n4332), .Y(n4331) );
  INVX2TS U2440 ( .A(n4329), .Y(n4328) );
  INVX2TS U2441 ( .A(n4326), .Y(n4325) );
  INVX2TS U2442 ( .A(n4323), .Y(n4322) );
  INVX2TS U2443 ( .A(n4320), .Y(n4319) );
  INVX2TS U2444 ( .A(n4317), .Y(n4316) );
  INVX2TS U2445 ( .A(n4314), .Y(n4313) );
  INVX2TS U2446 ( .A(n4311), .Y(n4310) );
  INVX2TS U2447 ( .A(n4308), .Y(n4307) );
  INVX2TS U2448 ( .A(n4305), .Y(n4304) );
  INVX2TS U2449 ( .A(n4302), .Y(n4301) );
  INVX2TS U2450 ( .A(n4299), .Y(n4298) );
  INVX2TS U2451 ( .A(n4296), .Y(n4295) );
  INVX2TS U2452 ( .A(n4293), .Y(n4292) );
  INVX2TS U2453 ( .A(n4290), .Y(n4289) );
  INVX2TS U2454 ( .A(n4287), .Y(n4286) );
  INVX2TS U2455 ( .A(n4284), .Y(n4283) );
  INVX2TS U2456 ( .A(n4281), .Y(n4280) );
  INVX2TS U2457 ( .A(n4278), .Y(n4277) );
  INVX2TS U2458 ( .A(n4275), .Y(n4274) );
  INVX2TS U2459 ( .A(n4272), .Y(n4271) );
  INVX2TS U2460 ( .A(n4269), .Y(n4268) );
  INVX2TS U2461 ( .A(n4266), .Y(n4265) );
  INVX2TS U2462 ( .A(n4263), .Y(n4262) );
  INVX2TS U2463 ( .A(n3968), .Y(n3967) );
  INVX2TS U2464 ( .A(n3965), .Y(n3964) );
  INVX2TS U2465 ( .A(n3962), .Y(n3961) );
  INVX2TS U2466 ( .A(n3959), .Y(n3958) );
  INVX2TS U2467 ( .A(n3956), .Y(n3955) );
  INVX2TS U2468 ( .A(n3953), .Y(n3952) );
  INVX2TS U2469 ( .A(n4202), .Y(n4201) );
  INVX2TS U2470 ( .A(n4199), .Y(n4198) );
  INVX2TS U2471 ( .A(n4193), .Y(n4192) );
  INVX2TS U2472 ( .A(n4190), .Y(n4189) );
  INVX2TS U2473 ( .A(n4196), .Y(n4195) );
  INVX2TS U2474 ( .A(n4187), .Y(n4186) );
  INVX2TS U2475 ( .A(n1933), .Y(n700) );
  INVX2TS U2476 ( .A(n2043), .Y(n653) );
  INVX2TS U2477 ( .A(n2027), .Y(n657) );
  OAI21X1TS U2478 ( .A0(n654), .A1(n2395), .B0(n2396), .Y(n2386) );
  AOI32X1TS U2479 ( .A0(n1091), .A1(n655), .A2(n1087), .B0(n2449), .B1(n2385), 
        .Y(n2396) );
  OAI22X1TS U2480 ( .A0(n1089), .A1(n2890), .B0(n2449), .B1(n2385), .Y(n2395)
         );
  INVX2TS U2481 ( .A(n2894), .Y(n654) );
  INVX2TS U2482 ( .A(n2012), .Y(n3121) );
  NAND4X1TS U2483 ( .A(n2019), .B(n2017), .C(n942), .D(n2376), .Y(n2012) );
  AND3X2TS U2484 ( .A(n2020), .B(n2018), .C(n2021), .Y(n2376) );
  AOI21X1TS U2485 ( .A0(n195), .A1(n978), .B0(n107), .Y(n2005) );
  AOI222XLTS U2486 ( .A0(n4203), .A1(n3482), .B0(n4210), .B1(n3460), .C0(n4218), .C1(n3442), .Y(n1750) );
  AOI222XLTS U2487 ( .A0(n4217), .A1(n3402), .B0(n4204), .B1(n3376), .C0(n4209), .C1(n3430), .Y(n1753) );
  NOR2X1TS U2488 ( .A(n688), .B(n476), .Y(n1769) );
  NOR2X1TS U2489 ( .A(n1910), .B(n974), .Y(n1839) );
  NOR2X1TS U2490 ( .A(n1836), .B(n179), .Y(n1826) );
  NAND2X1TS U2491 ( .A(n2006), .B(n128), .Y(n1793) );
  OAI2BB2XLTS U2492 ( .B0(n108), .B1(n476), .A0N(n145), .A1N(n107), .Y(n2006)
         );
  NAND2X1TS U2493 ( .A(n1763), .B(n2003), .Y(n1910) );
  INVX2TS U2494 ( .A(n2032), .Y(n602) );
  AOI221X1TS U2495 ( .A0(n4204), .A1(n3100), .B0(writeIn_SOUTH), .B1(n3085), 
        .C0(n2035), .Y(n2032) );
  OAI211X1TS U2496 ( .A0(n655), .A1(n951), .B0(n1087), .C0(n2393), .Y(n2894)
         );
  INVX2TS U2497 ( .A(n178), .Y(n678) );
  XOR2X1TS U2498 ( .A(n2394), .B(n2389), .Y(n1083) );
  XOR2X1TS U2499 ( .A(n2388), .B(n989), .Y(n2394) );
  INVX2TS U2500 ( .A(n2004), .Y(n947) );
  OAI221XLTS U2501 ( .A0(n680), .A1(n472), .B0(n3353), .B1(n912), .C0(n1755), 
        .Y(n2572) );
  AOI222XLTS U2502 ( .A0(n4209), .A1(n3297), .B0(n4204), .B1(n3305), .C0(n4218), .C1(n3341), .Y(n1755) );
  OAI221XLTS U2503 ( .A0(n914), .A1(n472), .B0(n3618), .B1(n603), .C0(n1744), 
        .Y(n2576) );
  AOI222XLTS U2504 ( .A0(n4203), .A1(n3559), .B0(n4210), .B1(n3570), .C0(n4218), .C1(n3606), .Y(n1744) );
  OAI221XLTS U2505 ( .A0(n481), .A1(n471), .B0(n3187), .B1(n911), .C0(n1742), 
        .Y(n2577) );
  AOI222XLTS U2506 ( .A0(n4217), .A1(n3672), .B0(n4204), .B1(n3638), .C0(n4209), .C1(n3866), .Y(n1742) );
  OAI221XLTS U2507 ( .A0(n952), .A1(n471), .B0(n483), .B1(n645), .C0(n1747), 
        .Y(n2575) );
  AOI222XLTS U2508 ( .A0(n4217), .A1(n3519), .B0(n4210), .B1(n3494), .C0(n4203), .C1(n3547), .Y(n1747) );
  OAI221XLTS U2509 ( .A0(n3695), .A1(n471), .B0(n3778), .B1(n879), .C0(n1740), 
        .Y(n2578) );
  AOI222XLTS U2510 ( .A0(n4203), .A1(n3707), .B0(n4210), .B1(n3725), .C0(n4218), .C1(n3755), .Y(n1740) );
  NOR2X1TS U2511 ( .A(n2017), .B(n143), .Y(n2048) );
  OAI22XLTS U2512 ( .A0(n964), .A1(n2017), .B0(n138), .B1(n2018), .Y(n2016) );
  NOR2BX1TS U2513 ( .AN(n1854), .B(n145), .Y(n1117) );
  OAI22X1TS U2514 ( .A0(n1084), .A1(n106), .B0(n1082), .B1(n476), .Y(n2886) );
  OAI22X1TS U2515 ( .A0(n1080), .A1(n106), .B0(n1082), .B1(n194), .Y(n2888) );
  XOR2X1TS U2516 ( .A(n2382), .B(n2383), .Y(n1084) );
  OAI2BB2XLTS U2517 ( .B0(n2387), .B1(n47), .A0N(n2388), .A1N(n2389), .Y(n2382) );
  XOR2X1TS U2518 ( .A(n121), .B(n2384), .Y(n2383) );
  NOR2X1TS U2519 ( .A(n2388), .B(n2389), .Y(n2387) );
  NOR2X1TS U2520 ( .A(n1864), .B(n178), .Y(n1854) );
  INVX2TS U2521 ( .A(n1836), .Y(n943) );
  NOR2BX1TS U2522 ( .AN(n1854), .B(n1879), .Y(n1150) );
  NOR2X1TS U2523 ( .A(n2020), .B(n142), .Y(n2033) );
  NOR2X1TS U2524 ( .A(n2018), .B(n142), .Y(n2034) );
  INVX2TS U2525 ( .A(writeIn_EAST), .Y(n4211) );
  INVX2TS U2526 ( .A(n142), .Y(n942) );
  OR2X2TS U2527 ( .A(n2019), .B(n143), .Y(n988) );
  OAI221XLTS U2528 ( .A0(n4214), .A1(n2019), .B0(n4208), .B1(n2020), .C0(n2021), .Y(n2015) );
  INVX2TS U2529 ( .A(n1864), .Y(n945) );
  NOR2BX1TS U2530 ( .AN(n183), .B(n2030), .Y(n2115) );
  NOR2BX1TS U2531 ( .AN(n184), .B(n2031), .Y(n2114) );
  NOR2BX1TS U2532 ( .AN(n114), .B(n2029), .Y(n2113) );
  NOR2BX1TS U2533 ( .AN(n181), .B(n2044), .Y(n2109) );
  NOR2BX1TS U2534 ( .AN(n182), .B(n2028), .Y(n2108) );
  NOR2X1TS U2535 ( .A(n2021), .B(n143), .Y(n2117) );
  OAI22X1TS U2536 ( .A0(n748), .A1(n1072), .B0(n780), .B1(n1058), .Y(n2374) );
  OAI22X1TS U2537 ( .A0(n738), .A1(n1071), .B0(n779), .B1(n1057), .Y(n2368) );
  OAI22X1TS U2538 ( .A0(n737), .A1(n1073), .B0(n778), .B1(n1060), .Y(n2362) );
  OAI22X1TS U2539 ( .A0(n736), .A1(n1074), .B0(n777), .B1(n1059), .Y(n2356) );
  OAI22X1TS U2540 ( .A0(n735), .A1(n1062), .B0(n776), .B1(n1048), .Y(n2350) );
  OAI22X1TS U2541 ( .A0(n734), .A1(n1062), .B0(n775), .B1(n1048), .Y(n2344) );
  OAI22X1TS U2542 ( .A0(n733), .A1(n1062), .B0(n774), .B1(n1048), .Y(n2338) );
  OAI22X1TS U2543 ( .A0(n732), .A1(n1062), .B0(n773), .B1(n1048), .Y(n2332) );
  OAI22X1TS U2544 ( .A0(n731), .A1(n1063), .B0(n772), .B1(n1049), .Y(n2326) );
  OAI22X1TS U2545 ( .A0(n730), .A1(n1063), .B0(n771), .B1(n1049), .Y(n2320) );
  OAI22X1TS U2546 ( .A0(n729), .A1(n1063), .B0(n770), .B1(n1049), .Y(n2314) );
  OAI22X1TS U2547 ( .A0(n728), .A1(n1063), .B0(n769), .B1(n1049), .Y(n2308) );
  OAI22X1TS U2548 ( .A0(n727), .A1(n1064), .B0(n768), .B1(n1050), .Y(n2302) );
  OAI22X1TS U2549 ( .A0(n726), .A1(n1064), .B0(n767), .B1(n1050), .Y(n2296) );
  OAI22X1TS U2550 ( .A0(n725), .A1(n1064), .B0(n766), .B1(n1050), .Y(n2290) );
  OAI22X1TS U2551 ( .A0(n747), .A1(n1064), .B0(n765), .B1(n1050), .Y(n2284) );
  OAI22X1TS U2552 ( .A0(n746), .A1(n1073), .B0(n915), .B1(n1059), .Y(n2278) );
  OAI22X1TS U2553 ( .A0(n724), .A1(n1072), .B0(n916), .B1(n1058), .Y(n2272) );
  OAI22X1TS U2554 ( .A0(n723), .A1(n1071), .B0(n917), .B1(n1057), .Y(n2266) );
  OAI22X1TS U2555 ( .A0(n722), .A1(n1074), .B0(n764), .B1(n1060), .Y(n2260) );
  OAI22X1TS U2556 ( .A0(n745), .A1(n1065), .B0(n763), .B1(n1051), .Y(n2254) );
  OAI22X1TS U2557 ( .A0(n721), .A1(n1065), .B0(n762), .B1(n1051), .Y(n2248) );
  OAI22X1TS U2558 ( .A0(n720), .A1(n1065), .B0(n761), .B1(n1051), .Y(n2242) );
  OAI22X1TS U2559 ( .A0(n719), .A1(n1065), .B0(n760), .B1(n1051), .Y(n2236) );
  OAI22X1TS U2560 ( .A0(n718), .A1(n1066), .B0(n759), .B1(n1052), .Y(n2230) );
  OAI22X1TS U2561 ( .A0(n717), .A1(n1066), .B0(n758), .B1(n1052), .Y(n2224) );
  OAI22X1TS U2562 ( .A0(n716), .A1(n1066), .B0(n757), .B1(n1052), .Y(n2218) );
  OAI22X1TS U2563 ( .A0(n715), .A1(n1066), .B0(n756), .B1(n1052), .Y(n2212) );
  OAI22X1TS U2564 ( .A0(n714), .A1(n1067), .B0(n755), .B1(n1053), .Y(n2206) );
  OAI22X1TS U2565 ( .A0(n713), .A1(n1067), .B0(n754), .B1(n1053), .Y(n2200) );
  OAI22X1TS U2566 ( .A0(n744), .A1(n1067), .B0(n753), .B1(n1053), .Y(n2194) );
  OAI22X1TS U2567 ( .A0(n712), .A1(n1067), .B0(n918), .B1(n1053), .Y(n2188) );
  OAI22X1TS U2568 ( .A0(n888), .A1(n1068), .B0(n891), .B1(n1054), .Y(n2182) );
  OAI22X1TS U2569 ( .A0(n887), .A1(n1068), .B0(n890), .B1(n1054), .Y(n2176) );
  OAI22X1TS U2570 ( .A0(n885), .A1(n1068), .B0(n889), .B1(n1054), .Y(n2164) );
  OAI22X1TS U2571 ( .A0(n884), .A1(n1069), .B0(n881), .B1(n1055), .Y(n2158) );
  OAI22X1TS U2572 ( .A0(n743), .A1(n1069), .B0(n784), .B1(n1055), .Y(n2146) );
  OAI22X1TS U2573 ( .A0(n711), .A1(n1069), .B0(n749), .B1(n1055), .Y(n2140) );
  OAI22X1TS U2574 ( .A0(n742), .A1(n1070), .B0(n783), .B1(n1056), .Y(n2134) );
  OAI22X1TS U2575 ( .A0(n741), .A1(n1070), .B0(n782), .B1(n1056), .Y(n2128) );
  OAI22X1TS U2576 ( .A0(n740), .A1(n1070), .B0(n781), .B1(n1056), .Y(n2122) );
  OAI22X1TS U2577 ( .A0(n739), .A1(n1070), .B0(n821), .B1(n1056), .Y(n2110) );
  OAI22X1TS U2578 ( .A0(n886), .A1(n1068), .B0(n882), .B1(n1054), .Y(n2170) );
  OAI22X1TS U2579 ( .A0(n883), .A1(n1069), .B0(n880), .B1(n1055), .Y(n2152) );
  AOI21X1TS U2580 ( .A0(n184), .A1(n1086), .B0(n105), .Y(n2885) );
  NAND3BX1TS U2581 ( .AN(n1087), .B(n1088), .C(n1089), .Y(n1086) );
  XOR2X1TS U2582 ( .A(n1090), .B(n1091), .Y(n1088) );
  NAND2X1TS U2583 ( .A(n171), .B(n184), .Y(n1093) );
  NAND2X1TS U2584 ( .A(n176), .B(n183), .Y(n2112) );
  NAND2X1TS U2585 ( .A(n168), .B(n181), .Y(n2111) );
  INVX2TS U2586 ( .A(requesterAddressIn_WEST[4]), .Y(n4049) );
  INVX2TS U2587 ( .A(requesterAddressIn_WEST[5]), .Y(n4052) );
  INVX2TS U2588 ( .A(requesterAddressIn_WEST[3]), .Y(n4046) );
  INVX2TS U2589 ( .A(requesterAddressIn_WEST[2]), .Y(n4043) );
  INVX2TS U2590 ( .A(requesterAddressIn_WEST[1]), .Y(n4040) );
  INVX2TS U2591 ( .A(requesterAddressIn_WEST[0]), .Y(n4037) );
  INVX2TS U2592 ( .A(requesterAddressIn_EAST[4]), .Y(n4199) );
  INVX2TS U2593 ( .A(requesterAddressIn_EAST[1]), .Y(n4190) );
  INVX2TS U2594 ( .A(requesterAddressIn_EAST[0]), .Y(n4187) );
  INVX2TS U2595 ( .A(requesterAddressIn_EAST[5]), .Y(n4202) );
  INVX2TS U2596 ( .A(requesterAddressIn_EAST[3]), .Y(n4196) );
  INVX2TS U2597 ( .A(requesterAddressIn_EAST[2]), .Y(n4193) );
  INVX2TS U2598 ( .A(destinationAddressIn_WEST[4]), .Y(n4007) );
  INVX2TS U2599 ( .A(destinationAddressIn_EAST[2]), .Y(n3959) );
  INVX2TS U2600 ( .A(destinationAddressIn_EAST[5]), .Y(n3968) );
  INVX2TS U2601 ( .A(destinationAddressIn_EAST[4]), .Y(n3965) );
  INVX2TS U2602 ( .A(destinationAddressIn_EAST[3]), .Y(n3962) );
  INVX2TS U2603 ( .A(destinationAddressIn_EAST[1]), .Y(n3956) );
  INVX2TS U2604 ( .A(destinationAddressIn_EAST[0]), .Y(n3953) );
  INVX2TS U2605 ( .A(destinationAddressIn_WEST[5]), .Y(n4010) );
  INVX2TS U2606 ( .A(destinationAddressIn_WEST[3]), .Y(n4004) );
  INVX2TS U2607 ( .A(destinationAddressIn_WEST[2]), .Y(n4001) );
  INVX2TS U2608 ( .A(destinationAddressIn_WEST[1]), .Y(n3998) );
  INVX2TS U2609 ( .A(destinationAddressIn_WEST[0]), .Y(n3995) );
  INVX2TS U2610 ( .A(dataIn_WEST[30]), .Y(n4353) );
  INVX2TS U2611 ( .A(dataIn_WEST[28]), .Y(n4347) );
  INVX2TS U2612 ( .A(dataIn_WEST[27]), .Y(n4344) );
  INVX2TS U2613 ( .A(dataIn_WEST[26]), .Y(n4341) );
  INVX2TS U2614 ( .A(dataIn_WEST[25]), .Y(n4338) );
  INVX2TS U2615 ( .A(dataIn_WEST[24]), .Y(n4335) );
  INVX2TS U2616 ( .A(dataIn_WEST[23]), .Y(n4332) );
  INVX2TS U2617 ( .A(dataIn_WEST[18]), .Y(n4317) );
  INVX2TS U2618 ( .A(dataIn_WEST[13]), .Y(n4302) );
  INVX2TS U2619 ( .A(dataIn_WEST[9]), .Y(n4290) );
  INVX2TS U2620 ( .A(dataIn_WEST[7]), .Y(n4284) );
  INVX2TS U2621 ( .A(dataIn_WEST[5]), .Y(n4278) );
  INVX2TS U2622 ( .A(dataIn_WEST[4]), .Y(n4275) );
  INVX2TS U2623 ( .A(dataIn_WEST[2]), .Y(n4269) );
  INVX2TS U2624 ( .A(dataIn_WEST[31]), .Y(n4356) );
  INVX2TS U2625 ( .A(dataIn_WEST[29]), .Y(n4350) );
  INVX2TS U2626 ( .A(dataIn_WEST[22]), .Y(n4329) );
  INVX2TS U2627 ( .A(dataIn_WEST[21]), .Y(n4326) );
  INVX2TS U2628 ( .A(dataIn_WEST[20]), .Y(n4323) );
  INVX2TS U2629 ( .A(dataIn_WEST[19]), .Y(n4320) );
  INVX2TS U2630 ( .A(dataIn_WEST[16]), .Y(n4311) );
  INVX2TS U2631 ( .A(dataIn_WEST[12]), .Y(n4299) );
  INVX2TS U2632 ( .A(dataIn_WEST[11]), .Y(n4296) );
  INVX2TS U2633 ( .A(dataIn_WEST[10]), .Y(n4293) );
  INVX2TS U2634 ( .A(dataIn_WEST[8]), .Y(n4287) );
  INVX2TS U2635 ( .A(dataIn_WEST[6]), .Y(n4281) );
  INVX2TS U2636 ( .A(dataIn_WEST[1]), .Y(n4266) );
  INVX2TS U2637 ( .A(dataIn_WEST[0]), .Y(n4263) );
  INVX2TS U2638 ( .A(dataIn_WEST[17]), .Y(n4314) );
  INVX2TS U2639 ( .A(dataIn_WEST[15]), .Y(n4308) );
  INVX2TS U2640 ( .A(dataIn_WEST[14]), .Y(n4305) );
  INVX2TS U2641 ( .A(dataIn_WEST[3]), .Y(n4272) );
  INVX2TS U2642 ( .A(readIn_WEST), .Y(n4208) );
  INVX2TS U2643 ( .A(destinationAddressIn_EAST[13]), .Y(n3992) );
  INVX2TS U2644 ( .A(destinationAddressIn_EAST[11]), .Y(n3986) );
  INVX2TS U2645 ( .A(destinationAddressIn_EAST[9]), .Y(n3980) );
  INVX2TS U2646 ( .A(destinationAddressIn_EAST[7]), .Y(n3974) );
  INVX2TS U2647 ( .A(destinationAddressIn_EAST[12]), .Y(n3989) );
  INVX2TS U2648 ( .A(destinationAddressIn_EAST[10]), .Y(n3983) );
  INVX2TS U2649 ( .A(destinationAddressIn_EAST[8]), .Y(n3977) );
  INVX2TS U2650 ( .A(destinationAddressIn_EAST[6]), .Y(n3971) );
  INVX2TS U2651 ( .A(dataIn_EAST[30]), .Y(n4457) );
  INVX2TS U2652 ( .A(dataIn_EAST[28]), .Y(n4450) );
  INVX2TS U2653 ( .A(dataIn_EAST[27]), .Y(n4447) );
  INVX2TS U2654 ( .A(dataIn_EAST[26]), .Y(n4442) );
  INVX2TS U2655 ( .A(dataIn_EAST[25]), .Y(n4439) );
  INVX2TS U2656 ( .A(dataIn_EAST[24]), .Y(n4435) );
  INVX2TS U2657 ( .A(dataIn_EAST[23]), .Y(n4431) );
  INVX2TS U2658 ( .A(dataIn_EAST[18]), .Y(n4413) );
  INVX2TS U2659 ( .A(dataIn_EAST[13]), .Y(n4398) );
  INVX2TS U2660 ( .A(dataIn_EAST[9]), .Y(n4386) );
  INVX2TS U2661 ( .A(dataIn_EAST[7]), .Y(n4380) );
  INVX2TS U2662 ( .A(dataIn_EAST[5]), .Y(n4374) );
  INVX2TS U2663 ( .A(dataIn_EAST[4]), .Y(n4371) );
  INVX2TS U2664 ( .A(dataIn_EAST[2]), .Y(n4365) );
  INVX2TS U2665 ( .A(dataIn_EAST[31]), .Y(n4460) );
  INVX2TS U2666 ( .A(dataIn_EAST[29]), .Y(n4453) );
  INVX2TS U2667 ( .A(dataIn_EAST[22]), .Y(n4427) );
  INVX2TS U2668 ( .A(dataIn_EAST[21]), .Y(n4424) );
  INVX2TS U2669 ( .A(dataIn_EAST[20]), .Y(n4421) );
  INVX2TS U2670 ( .A(dataIn_EAST[19]), .Y(n4416) );
  INVX2TS U2671 ( .A(dataIn_EAST[16]), .Y(n4407) );
  INVX2TS U2672 ( .A(dataIn_EAST[12]), .Y(n4395) );
  INVX2TS U2673 ( .A(dataIn_EAST[11]), .Y(n4392) );
  INVX2TS U2674 ( .A(dataIn_EAST[10]), .Y(n4389) );
  INVX2TS U2675 ( .A(dataIn_EAST[8]), .Y(n4383) );
  INVX2TS U2676 ( .A(dataIn_EAST[6]), .Y(n4377) );
  INVX2TS U2677 ( .A(dataIn_EAST[1]), .Y(n4362) );
  INVX2TS U2678 ( .A(dataIn_EAST[0]), .Y(n4359) );
  INVX2TS U2679 ( .A(dataIn_EAST[17]), .Y(n4410) );
  INVX2TS U2680 ( .A(dataIn_EAST[15]), .Y(n4404) );
  INVX2TS U2681 ( .A(dataIn_EAST[14]), .Y(n4401) );
  INVX2TS U2682 ( .A(dataIn_EAST[3]), .Y(n4368) );
  INVX2TS U2683 ( .A(writeIn_WEST), .Y(n4205) );
  INVX2TS U2684 ( .A(destinationAddressIn_WEST[7]), .Y(n4016) );
  INVX2TS U2685 ( .A(destinationAddressIn_WEST[6]), .Y(n4013) );
  CLKBUFX2TS U2686 ( .A(writeIn_SOUTH), .Y(n4216) );
  CLKBUFX2TS U2687 ( .A(destinationAddressIn_SOUTH[13]), .Y(n4258) );
  CLKBUFX2TS U2688 ( .A(destinationAddressIn_SOUTH[11]), .Y(n4252) );
  CLKBUFX2TS U2689 ( .A(destinationAddressIn_SOUTH[9]), .Y(n4246) );
  CLKBUFX2TS U2690 ( .A(destinationAddressIn_SOUTH[12]), .Y(n4255) );
  CLKBUFX2TS U2691 ( .A(destinationAddressIn_SOUTH[10]), .Y(n4249) );
  CLKBUFX2TS U2692 ( .A(destinationAddressIn_SOUTH[8]), .Y(n4243) );
  CLKBUFX2TS U2693 ( .A(destinationAddressIn_SOUTH[4]), .Y(n4231) );
  CLKBUFX2TS U2694 ( .A(destinationAddressIn_NORTH[4]), .Y(n4065) );
  CLKBUFX2TS U2695 ( .A(requesterAddressIn_NORTH[4]), .Y(n4083) );
  CLKBUFX2TS U2696 ( .A(requesterAddressIn_SOUTH[4]), .Y(n4597) );
  CLKBUFX2TS U2697 ( .A(requesterAddressIn_NORTH[1]), .Y(n4074) );
  CLKBUFX2TS U2698 ( .A(requesterAddressIn_SOUTH[1]), .Y(n4585) );
  CLKBUFX2TS U2699 ( .A(requesterAddressIn_NORTH[0]), .Y(n4071) );
  CLKBUFX2TS U2700 ( .A(requesterAddressIn_SOUTH[0]), .Y(n4582) );
  CLKBUFX2TS U2701 ( .A(requesterAddressIn_NORTH[5]), .Y(n4086) );
  CLKBUFX2TS U2702 ( .A(requesterAddressIn_SOUTH[5]), .Y(n4602) );
  CLKBUFX2TS U2703 ( .A(requesterAddressIn_NORTH[3]), .Y(n4080) );
  CLKBUFX2TS U2704 ( .A(requesterAddressIn_SOUTH[3]), .Y(n4593) );
  CLKBUFX2TS U2705 ( .A(requesterAddressIn_NORTH[2]), .Y(n4077) );
  CLKBUFX2TS U2706 ( .A(requesterAddressIn_SOUTH[2]), .Y(n4589) );
  CLKBUFX2TS U2707 ( .A(destinationAddressIn_NORTH[5]), .Y(n4068) );
  CLKBUFX2TS U2708 ( .A(destinationAddressIn_SOUTH[5]), .Y(n4234) );
  CLKBUFX2TS U2709 ( .A(destinationAddressIn_NORTH[3]), .Y(n4062) );
  CLKBUFX2TS U2710 ( .A(destinationAddressIn_SOUTH[3]), .Y(n4228) );
  CLKBUFX2TS U2711 ( .A(destinationAddressIn_NORTH[2]), .Y(n4059) );
  CLKBUFX2TS U2712 ( .A(destinationAddressIn_SOUTH[2]), .Y(n4225) );
  CLKBUFX2TS U2713 ( .A(destinationAddressIn_NORTH[1]), .Y(n4056) );
  CLKBUFX2TS U2714 ( .A(destinationAddressIn_SOUTH[1]), .Y(n4222) );
  CLKBUFX2TS U2715 ( .A(destinationAddressIn_NORTH[0]), .Y(n4053) );
  CLKBUFX2TS U2716 ( .A(destinationAddressIn_SOUTH[0]), .Y(n4219) );
  CLKBUFX2TS U2717 ( .A(dataIn_NORTH[30]), .Y(n4179) );
  CLKBUFX2TS U2718 ( .A(dataIn_SOUTH[30]), .Y(n4574) );
  CLKBUFX2TS U2719 ( .A(dataIn_NORTH[28]), .Y(n4173) );
  CLKBUFX2TS U2720 ( .A(dataIn_SOUTH[28]), .Y(n4566) );
  CLKBUFX2TS U2721 ( .A(dataIn_NORTH[27]), .Y(n4170) );
  CLKBUFX2TS U2722 ( .A(dataIn_SOUTH[27]), .Y(n4562) );
  CLKBUFX2TS U2723 ( .A(dataIn_NORTH[26]), .Y(n4167) );
  CLKBUFX2TS U2724 ( .A(dataIn_SOUTH[26]), .Y(n4559) );
  CLKBUFX2TS U2725 ( .A(dataIn_NORTH[25]), .Y(n4164) );
  CLKBUFX2TS U2726 ( .A(dataIn_SOUTH[25]), .Y(n4555) );
  CLKBUFX2TS U2727 ( .A(dataIn_NORTH[24]), .Y(n4161) );
  CLKBUFX2TS U2728 ( .A(dataIn_SOUTH[24]), .Y(n4551) );
  CLKBUFX2TS U2729 ( .A(dataIn_NORTH[23]), .Y(n4158) );
  CLKBUFX2TS U2730 ( .A(dataIn_SOUTH[23]), .Y(n4547) );
  CLKBUFX2TS U2731 ( .A(dataIn_NORTH[18]), .Y(n4143) );
  CLKBUFX2TS U2732 ( .A(dataIn_SOUTH[18]), .Y(n4528) );
  CLKBUFX2TS U2733 ( .A(dataIn_NORTH[13]), .Y(n4128) );
  CLKBUFX2TS U2734 ( .A(dataIn_SOUTH[13]), .Y(n4510) );
  CLKBUFX2TS U2735 ( .A(dataIn_NORTH[9]), .Y(n4116) );
  CLKBUFX2TS U2736 ( .A(dataIn_SOUTH[9]), .Y(n4495) );
  CLKBUFX2TS U2737 ( .A(dataIn_NORTH[7]), .Y(n4110) );
  CLKBUFX2TS U2738 ( .A(dataIn_SOUTH[7]), .Y(n4488) );
  CLKBUFX2TS U2739 ( .A(dataIn_NORTH[5]), .Y(n4104) );
  CLKBUFX2TS U2740 ( .A(dataIn_SOUTH[5]), .Y(n4480) );
  CLKBUFX2TS U2741 ( .A(dataIn_NORTH[4]), .Y(n4101) );
  CLKBUFX2TS U2742 ( .A(dataIn_SOUTH[4]), .Y(n4477) );
  CLKBUFX2TS U2743 ( .A(dataIn_NORTH[2]), .Y(n4095) );
  CLKBUFX2TS U2744 ( .A(dataIn_SOUTH[2]), .Y(n4468) );
  CLKBUFX2TS U2745 ( .A(dataIn_NORTH[31]), .Y(n4182) );
  CLKBUFX2TS U2746 ( .A(dataIn_SOUTH[31]), .Y(n4578) );
  CLKBUFX2TS U2747 ( .A(dataIn_NORTH[29]), .Y(n4176) );
  CLKBUFX2TS U2748 ( .A(dataIn_SOUTH[29]), .Y(n4570) );
  CLKBUFX2TS U2749 ( .A(dataIn_NORTH[22]), .Y(n4155) );
  CLKBUFX2TS U2750 ( .A(dataIn_SOUTH[22]), .Y(n4543) );
  CLKBUFX2TS U2751 ( .A(dataIn_NORTH[21]), .Y(n4152) );
  CLKBUFX2TS U2752 ( .A(dataIn_SOUTH[21]), .Y(n4540) );
  CLKBUFX2TS U2753 ( .A(dataIn_NORTH[20]), .Y(n4149) );
  CLKBUFX2TS U2754 ( .A(dataIn_SOUTH[20]), .Y(n4535) );
  CLKBUFX2TS U2755 ( .A(dataIn_NORTH[19]), .Y(n4146) );
  CLKBUFX2TS U2756 ( .A(dataIn_SOUTH[19]), .Y(n4532) );
  CLKBUFX2TS U2757 ( .A(dataIn_NORTH[16]), .Y(n4137) );
  CLKBUFX2TS U2758 ( .A(dataIn_SOUTH[16]), .Y(n4521) );
  CLKBUFX2TS U2759 ( .A(dataIn_NORTH[12]), .Y(n4125) );
  CLKBUFX2TS U2760 ( .A(dataIn_SOUTH[12]), .Y(n4506) );
  CLKBUFX2TS U2761 ( .A(dataIn_NORTH[11]), .Y(n4122) );
  CLKBUFX2TS U2762 ( .A(dataIn_SOUTH[11]), .Y(n4503) );
  CLKBUFX2TS U2763 ( .A(dataIn_NORTH[10]), .Y(n4119) );
  CLKBUFX2TS U2764 ( .A(dataIn_SOUTH[10]), .Y(n4498) );
  CLKBUFX2TS U2765 ( .A(dataIn_NORTH[8]), .Y(n4113) );
  CLKBUFX2TS U2766 ( .A(dataIn_SOUTH[8]), .Y(n4492) );
  CLKBUFX2TS U2767 ( .A(dataIn_NORTH[6]), .Y(n4107) );
  CLKBUFX2TS U2768 ( .A(dataIn_SOUTH[6]), .Y(n4484) );
  CLKBUFX2TS U2769 ( .A(dataIn_NORTH[1]), .Y(n4092) );
  CLKBUFX2TS U2770 ( .A(dataIn_SOUTH[1]), .Y(n4465) );
  CLKBUFX2TS U2771 ( .A(dataIn_NORTH[0]), .Y(n4089) );
  CLKBUFX2TS U2772 ( .A(dataIn_SOUTH[0]), .Y(n4461) );
  CLKBUFX2TS U2773 ( .A(dataIn_NORTH[17]), .Y(n4140) );
  CLKBUFX2TS U2774 ( .A(dataIn_SOUTH[17]), .Y(n4524) );
  CLKBUFX2TS U2775 ( .A(dataIn_NORTH[15]), .Y(n4134) );
  CLKBUFX2TS U2776 ( .A(dataIn_SOUTH[15]), .Y(n4517) );
  CLKBUFX2TS U2777 ( .A(dataIn_NORTH[14]), .Y(n4131) );
  CLKBUFX2TS U2778 ( .A(dataIn_SOUTH[14]), .Y(n4513) );
  CLKBUFX2TS U2779 ( .A(dataIn_NORTH[3]), .Y(n4098) );
  CLKBUFX2TS U2780 ( .A(dataIn_SOUTH[3]), .Y(n4472) );
  INVX2TS U2781 ( .A(readIn_EAST), .Y(n4215) );
  INVX2TS U2782 ( .A(n4028), .Y(n4027) );
  INVX2TS U2783 ( .A(n4031), .Y(n4029) );
  INVX2TS U2784 ( .A(n4028), .Y(n4026) );
  INVX2TS U2785 ( .A(n4022), .Y(n4020) );
  INVX2TS U2786 ( .A(n4019), .Y(n4017) );
  INVX2TS U2787 ( .A(n4034), .Y(n4032) );
  INVX2TS U2788 ( .A(n4025), .Y(n4023) );
  INVX2TS U2789 ( .A(n4034), .Y(n4033) );
  INVX2TS U2790 ( .A(n4022), .Y(n4021) );
  INVX2TS U2791 ( .A(n4031), .Y(n4030) );
  INVX2TS U2792 ( .A(n4025), .Y(n4024) );
  INVX2TS U2793 ( .A(n4019), .Y(n4018) );
  AO21X1TS U2794 ( .A0(n486), .A1(n1090), .B0(n4605), .Y(n1092) );
  NOR2X1TS U2795 ( .A(n948), .B(n140), .Y(n2892) );
  XOR2X1TS U2796 ( .A(n1091), .B(n2891), .Y(n2449) );
  AOI21X1TS U2797 ( .A0(n2892), .A1(n475), .B0(n2893), .Y(n2891) );
  AOI2BB1X1TS U2798 ( .A0N(n141), .A1N(n2892), .B0(n990), .Y(n2893) );
  INVX2TS U2799 ( .A(n1089), .Y(n655) );
  NAND2X1TS U2800 ( .A(n467), .B(n121), .Y(n1933) );
  AOI21X1TS U2801 ( .A0(n658), .A1(n948), .B0(n2892), .Y(n1087) );
  OAI22X1TS U2802 ( .A0(n604), .A1(n2044), .B0(n912), .B1(n2028), .Y(n2039) );
  OAI22X1TS U2803 ( .A0(n643), .A1(n2029), .B0(n645), .B1(n2030), .Y(n2042) );
  OAI22X1TS U2804 ( .A0(n2026), .A1(n644), .B0(n911), .B1(n2031), .Y(n2041) );
  OAI22X1TS U2805 ( .A0(n603), .A1(n2027), .B0(n879), .B1(n2043), .Y(n2040) );
  NAND3X1TS U2806 ( .A(n475), .B(n140), .C(n3), .Y(n2027) );
  INVX2TS U2807 ( .A(n2028), .Y(n656) );
  NAND2X1TS U2808 ( .A(n1090), .B(n97), .Y(n2043) );
  INVX2TS U2809 ( .A(n2026), .Y(n652) );
  INVX2TS U2810 ( .A(n2044), .Y(n648) );
  OAI22X1TS U2811 ( .A0(n2026), .A1(n598), .B0(n2027), .B1(n600), .Y(n2025) );
  OAI22X1TS U2812 ( .A0(n2028), .A1(n601), .B0(n2029), .B1(n892), .Y(n2024) );
  AOI222XLTS U2813 ( .A0(n4026), .A1(n3480), .B0(n3985), .B1(n3461), .C0(n4254), .C1(n3443), .Y(n1929) );
  AOI222XLTS U2814 ( .A0(n4011), .A1(n3482), .B0(n3970), .B1(n3460), .C0(n4239), .C1(n3442), .Y(n1924) );
  AOI222XLTS U2815 ( .A0(n4029), .A1(n3480), .B0(n3988), .B1(n3461), .C0(n4257), .C1(n3443), .Y(n1930) );
  AOI222XLTS U2816 ( .A0(n4020), .A1(n3481), .B0(n3979), .B1(n3461), .C0(n4248), .C1(n3443), .Y(n1927) );
  AOI222XLTS U2817 ( .A0(n4017), .A1(n3481), .B0(n3976), .B1(n3460), .C0(n4245), .C1(n3442), .Y(n1926) );
  AOI222XLTS U2818 ( .A0(n4032), .A1(n3480), .B0(n3991), .B1(n3467), .C0(n4260), .C1(n3450), .Y(n1931) );
  AOI222XLTS U2819 ( .A0(n4023), .A1(n3481), .B0(n3982), .B1(n3461), .C0(n4251), .C1(n3443), .Y(n1928) );
  AOI222XLTS U2820 ( .A0(n4014), .A1(n3482), .B0(n3973), .B1(n3460), .C0(n4242), .C1(n3442), .Y(n1925) );
  AOI222XLTS U2821 ( .A0(n4259), .A1(n3400), .B0(n4033), .B1(n3384), .C0(n3990), .C1(n3428), .Y(n1955) );
  AOI222XLTS U2822 ( .A0(n4253), .A1(n3400), .B0(n4027), .B1(n3377), .C0(n3984), .C1(n3428), .Y(n1953) );
  AOI222XLTS U2823 ( .A0(n4247), .A1(n3401), .B0(n4021), .B1(n3377), .C0(n3978), .C1(n3429), .Y(n1951) );
  AOI222XLTS U2824 ( .A0(n4241), .A1(n3401), .B0(n4015), .B1(n3376), .C0(n3972), .C1(n3430), .Y(n1949) );
  AOI222XLTS U2825 ( .A0(n4256), .A1(n3400), .B0(n4030), .B1(n3377), .C0(n3987), .C1(n3428), .Y(n1954) );
  AOI222XLTS U2826 ( .A0(n4250), .A1(n3400), .B0(n4024), .B1(n3377), .C0(n3981), .C1(n3429), .Y(n1952) );
  AOI222XLTS U2827 ( .A0(n4244), .A1(n3401), .B0(n4018), .B1(n3376), .C0(n3975), .C1(n3429), .Y(n1950) );
  AOI222XLTS U2828 ( .A0(n4238), .A1(n3401), .B0(n4012), .B1(n3376), .C0(n3969), .C1(n3430), .Y(n1948) );
  OAI221XLTS U2829 ( .A0(n4211), .A1(n2019), .B0(n471), .B1(n2017), .C0(n6248), 
        .Y(n2036) );
  XOR2X1TS U2830 ( .A(n5), .B(n1083), .Y(n2390) );
  OAI32X1TS U2831 ( .A0(n2380), .A1(n2381), .A2(n1081), .B0(n96), .B1(n142), 
        .Y(N4718) );
  XOR2X1TS U2832 ( .A(n1084), .B(n385), .Y(n2381) );
  NAND2X1TS U2833 ( .A(n2390), .B(n2391), .Y(n2380) );
  XOR2X1TS U2834 ( .A(n140), .B(n1080), .Y(n2391) );
  OAI221XLTS U2835 ( .A0(n680), .A1(n150), .B0(n3351), .B1(n710), .C0(n1979), 
        .Y(n2465) );
  AOI222XLTS U2836 ( .A0(n3990), .A1(n1199), .B0(n4033), .B1(n3303), .C0(n4260), .C1(n3346), .Y(n1979) );
  OAI221XLTS U2837 ( .A0(n680), .A1(n156), .B0(n3351), .B1(n709), .C0(n1978), 
        .Y(n2466) );
  AOI222XLTS U2838 ( .A0(n3987), .A1(n3301), .B0(n4030), .B1(n3303), .C0(n4257), .C1(n3342), .Y(n1978) );
  OAI221XLTS U2839 ( .A0(n687), .A1(n152), .B0(n3351), .B1(n708), .C0(n1977), 
        .Y(n2467) );
  AOI222XLTS U2840 ( .A0(n3984), .A1(n3299), .B0(n4027), .B1(n3303), .C0(n4254), .C1(n3342), .Y(n1977) );
  OAI221XLTS U2841 ( .A0(n683), .A1(n158), .B0(n3351), .B1(n707), .C0(n1976), 
        .Y(n2468) );
  AOI222XLTS U2842 ( .A0(n3981), .A1(n3301), .B0(n4024), .B1(n3303), .C0(n4251), .C1(n3342), .Y(n1976) );
  OAI221XLTS U2843 ( .A0(n687), .A1(n154), .B0(n3352), .B1(n706), .C0(n1975), 
        .Y(n2469) );
  AOI222XLTS U2844 ( .A0(n3978), .A1(n3299), .B0(n4021), .B1(n3304), .C0(n4248), .C1(n3342), .Y(n1975) );
  OAI221XLTS U2845 ( .A0(n683), .A1(n160), .B0(n3352), .B1(n705), .C0(n1974), 
        .Y(n2470) );
  AOI222XLTS U2846 ( .A0(n3975), .A1(n3297), .B0(n4018), .B1(n3304), .C0(n4245), .C1(n3341), .Y(n1974) );
  OAI221XLTS U2847 ( .A0(n687), .A1(n146), .B0(n3352), .B1(n704), .C0(n1973), 
        .Y(n2471) );
  AOI222XLTS U2848 ( .A0(n3972), .A1(n3297), .B0(n4015), .B1(n3304), .C0(n4242), .C1(n3341), .Y(n1973) );
  OAI221XLTS U2849 ( .A0(n683), .A1(n149), .B0(n3352), .B1(n703), .C0(n1972), 
        .Y(n2472) );
  AOI222XLTS U2850 ( .A0(n3969), .A1(n3297), .B0(n4012), .B1(n3304), .C0(n4239), .C1(n3341), .Y(n1972) );
  OAI221XLTS U2851 ( .A0(n479), .A1(n155), .B0(n3186), .B1(n910), .C0(n1858), 
        .Y(n2539) );
  AOI222XLTS U2852 ( .A0(n4247), .A1(n3673), .B0(n4021), .B1(n3637), .C0(n3978), .C1(n3861), .Y(n1858) );
  OAI221XLTS U2853 ( .A0(n481), .A1(n161), .B0(n3186), .B1(n900), .C0(n1857), 
        .Y(n2540) );
  AOI222XLTS U2854 ( .A0(n4244), .A1(n3673), .B0(n4018), .B1(n3638), .C0(n3975), .C1(n3866), .Y(n1857) );
  OAI221XLTS U2855 ( .A0(n482), .A1(n147), .B0(n3186), .B1(n899), .C0(n1856), 
        .Y(n2541) );
  AOI222XLTS U2856 ( .A0(n4241), .A1(n3673), .B0(n4015), .B1(n3637), .C0(n3972), .C1(n3866), .Y(n1856) );
  OAI221XLTS U2857 ( .A0(n481), .A1(n159), .B0(n3186), .B1(n584), .C0(n1859), 
        .Y(n2538) );
  AOI222XLTS U2858 ( .A0(n4250), .A1(n3672), .B0(n4024), .B1(n3638), .C0(n3981), .C1(n3861), .Y(n1859) );
  OAI221XLTS U2859 ( .A0(n940), .A1(n151), .B0(n3616), .B1(n576), .C0(n1887), 
        .Y(n2521) );
  AOI222XLTS U2860 ( .A0(n4032), .A1(n3566), .B0(n3991), .B1(n3568), .C0(n4260), .C1(n3611), .Y(n1887) );
  OAI221XLTS U2861 ( .A0(n938), .A1(n157), .B0(n3616), .B1(n575), .C0(n1886), 
        .Y(n2522) );
  AOI222XLTS U2862 ( .A0(n4029), .A1(n3560), .B0(n3988), .B1(n3568), .C0(n4257), .C1(n3607), .Y(n1886) );
  OAI221XLTS U2863 ( .A0(n940), .A1(n153), .B0(n3616), .B1(n574), .C0(n1885), 
        .Y(n2523) );
  AOI222XLTS U2864 ( .A0(n4026), .A1(n3560), .B0(n3985), .B1(n3568), .C0(n4254), .C1(n3607), .Y(n1885) );
  OAI221XLTS U2865 ( .A0(n938), .A1(n158), .B0(n3616), .B1(n573), .C0(n1884), 
        .Y(n2524) );
  AOI222XLTS U2866 ( .A0(n4023), .A1(n3560), .B0(n3982), .B1(n3568), .C0(n4251), .C1(n3607), .Y(n1884) );
  OAI221XLTS U2867 ( .A0(n940), .A1(n154), .B0(n3617), .B1(n572), .C0(n1883), 
        .Y(n2525) );
  AOI222XLTS U2868 ( .A0(n4020), .A1(n3560), .B0(n3979), .B1(n3569), .C0(n4248), .C1(n3607), .Y(n1883) );
  OAI221XLTS U2869 ( .A0(n938), .A1(n160), .B0(n3617), .B1(n571), .C0(n1882), 
        .Y(n2526) );
  AOI222XLTS U2870 ( .A0(n4017), .A1(n3559), .B0(n3976), .B1(n3569), .C0(n4245), .C1(n3606), .Y(n1882) );
  OAI221XLTS U2871 ( .A0(n940), .A1(n146), .B0(n3617), .B1(n570), .C0(n1881), 
        .Y(n2527) );
  AOI222XLTS U2872 ( .A0(n4014), .A1(n3559), .B0(n3973), .B1(n3569), .C0(n4242), .C1(n3606), .Y(n1881) );
  OAI221XLTS U2873 ( .A0(n938), .A1(n148), .B0(n3617), .B1(n569), .C0(n1880), 
        .Y(n2528) );
  AOI222XLTS U2874 ( .A0(n4011), .A1(n3559), .B0(n3970), .B1(n3569), .C0(n4239), .C1(n3606), .Y(n1880) );
  OAI221XLTS U2875 ( .A0(n689), .A1(n4031), .B0(n3268), .B1(n565), .C0(n1999), 
        .Y(n2452) );
  AOI222XLTS U2876 ( .A0(n4256), .A1(n3212), .B0(
        destinationAddressIn_NORTH[12]), .B1(n3234), .C0(n3987), .C1(n3259), 
        .Y(n1999) );
  OAI221XLTS U2877 ( .A0(n913), .A1(n4019), .B0(n3269), .B1(n564), .C0(n1995), 
        .Y(n2456) );
  AOI222XLTS U2878 ( .A0(n4244), .A1(n3211), .B0(destinationAddressIn_NORTH[8]), .B1(n3235), .C0(n3975), .C1(n3258), .Y(n1995) );
  OAI221XLTS U2879 ( .A0(n701), .A1(n4034), .B0(n3268), .B1(n562), .C0(n2000), 
        .Y(n2451) );
  AOI222XLTS U2880 ( .A0(n4259), .A1(n3218), .B0(
        destinationAddressIn_NORTH[13]), .B1(n3234), .C0(n3990), .C1(n3266), 
        .Y(n2000) );
  OAI221XLTS U2881 ( .A0(n913), .A1(n4025), .B0(n3268), .B1(n561), .C0(n1997), 
        .Y(n2454) );
  AOI222XLTS U2882 ( .A0(n4250), .A1(n3212), .B0(
        destinationAddressIn_NORTH[10]), .B1(n3234), .C0(n3981), .C1(n3259), 
        .Y(n1997) );
  OAI221XLTS U2883 ( .A0(n701), .A1(n4013), .B0(n3269), .B1(n560), .C0(n1993), 
        .Y(n2458) );
  AOI222XLTS U2884 ( .A0(n4238), .A1(n3211), .B0(destinationAddressIn_NORTH[6]), .B1(n3235), .C0(n3969), .C1(n3258), .Y(n1993) );
  OAI221XLTS U2885 ( .A0(n913), .A1(n4028), .B0(n3268), .B1(n556), .C0(n1998), 
        .Y(n2453) );
  AOI222XLTS U2886 ( .A0(n4253), .A1(n3212), .B0(
        destinationAddressIn_NORTH[11]), .B1(n3234), .C0(n3984), .C1(n3259), 
        .Y(n1998) );
  OAI221XLTS U2887 ( .A0(n701), .A1(n4022), .B0(n3269), .B1(n555), .C0(n1996), 
        .Y(n2455) );
  AOI222XLTS U2888 ( .A0(n4247), .A1(n3212), .B0(destinationAddressIn_NORTH[9]), .B1(n3235), .C0(n3978), .C1(n3259), .Y(n1996) );
  OAI221XLTS U2889 ( .A0(n913), .A1(n4016), .B0(n3269), .B1(n554), .C0(n1994), 
        .Y(n2457) );
  AOI222XLTS U2890 ( .A0(n4241), .A1(n3211), .B0(destinationAddressIn_NORTH[7]), .B1(n3235), .C0(n3972), .C1(n3258), .Y(n1994) );
  OAI221XLTS U2891 ( .A0(n482), .A1(n148), .B0(n3187), .B1(n909), .C0(n1855), 
        .Y(n2542) );
  AOI222XLTS U2892 ( .A0(n4238), .A1(n3672), .B0(n4012), .B1(n3639), .C0(n3969), .C1(n3866), .Y(n1855) );
  OAI221XLTS U2893 ( .A0(n701), .A1(n4205), .B0(n3270), .B1(n643), .C0(n1757), 
        .Y(n2571) );
  AOI222XLTS U2894 ( .A0(n4217), .A1(n3211), .B0(writeIn_NORTH), .B1(n3237), 
        .C0(n4209), .C1(n3258), .Y(n1757) );
  OAI221XLTS U2895 ( .A0(n956), .A1(n156), .B0(n485), .B1(n591), .C0(n1907), 
        .Y(n2508) );
  AOI222XLTS U2896 ( .A0(n4256), .A1(n3517), .B0(n3988), .B1(n3495), .C0(n4029), .C1(n3545), .Y(n1907) );
  OAI221XLTS U2897 ( .A0(n957), .A1(n152), .B0(n484), .B1(n590), .C0(n1906), 
        .Y(n2509) );
  AOI222XLTS U2898 ( .A0(n4253), .A1(n3517), .B0(n3985), .B1(n3495), .C0(n4026), .C1(n3545), .Y(n1906) );
  OAI221XLTS U2899 ( .A0(n956), .A1(n158), .B0(n485), .B1(n589), .C0(n1905), 
        .Y(n2510) );
  AOI222XLTS U2900 ( .A0(n4250), .A1(n3517), .B0(n3982), .B1(n3495), .C0(n4023), .C1(n3546), .Y(n1905) );
  OAI221XLTS U2901 ( .A0(n957), .A1(n161), .B0(n484), .B1(n588), .C0(n1903), 
        .Y(n2512) );
  AOI222XLTS U2902 ( .A0(n4244), .A1(n3518), .B0(n3976), .B1(n3494), .C0(n4017), .C1(n3546), .Y(n1903) );
  OAI221XLTS U2903 ( .A0(n956), .A1(n147), .B0(n485), .B1(n587), .C0(n1902), 
        .Y(n2513) );
  AOI222XLTS U2904 ( .A0(n4241), .A1(n3518), .B0(n3973), .B1(n3494), .C0(n4014), .C1(n3547), .Y(n1902) );
  OAI221XLTS U2905 ( .A0(n957), .A1(n149), .B0(n484), .B1(n586), .C0(n1901), 
        .Y(n2514) );
  AOI222XLTS U2906 ( .A0(n4238), .A1(n3518), .B0(n3970), .B1(n3494), .C0(n4011), .C1(n3547), .Y(n1901) );
  OAI221XLTS U2907 ( .A0(n957), .A1(n150), .B0(n484), .B1(n583), .C0(n1908), 
        .Y(n2507) );
  AOI222XLTS U2908 ( .A0(n4259), .A1(n3517), .B0(n3991), .B1(n3501), .C0(n4032), .C1(n3545), .Y(n1908) );
  OAI221XLTS U2909 ( .A0(n956), .A1(n154), .B0(n485), .B1(n582), .C0(n1904), 
        .Y(n2511) );
  AOI222XLTS U2910 ( .A0(n4247), .A1(n3518), .B0(n3979), .B1(n3495), .C0(n4020), .C1(n3546), .Y(n1904) );
  OAI221XLTS U2911 ( .A0(n482), .A1(n150), .B0(n3122), .B1(n902), .C0(n1862), 
        .Y(n2535) );
  AOI222XLTS U2912 ( .A0(n4259), .A1(n3672), .B0(n4033), .B1(n3637), .C0(n3990), .C1(n3863), .Y(n1862) );
  OAI221XLTS U2913 ( .A0(n482), .A1(n152), .B0(n3122), .B1(n901), .C0(n1860), 
        .Y(n2537) );
  AOI222XLTS U2914 ( .A0(n4253), .A1(n3674), .B0(n4027), .B1(n3637), .C0(n3984), .C1(n3861), .Y(n1860) );
  OAI221XLTS U2915 ( .A0(n481), .A1(n156), .B0(n3122), .B1(n585), .C0(n1861), 
        .Y(n2536) );
  AOI222XLTS U2916 ( .A0(n4256), .A1(n3673), .B0(n4030), .B1(n3638), .C0(n3987), .C1(n3861), .Y(n1861) );
  OAI221XLTS U2917 ( .A0(n3694), .A1(n155), .B0(n3764), .B1(n908), .C0(n1831), 
        .Y(n2553) );
  AOI222XLTS U2918 ( .A0(n4020), .A1(n3708), .B0(n3979), .B1(n3717), .C0(
        destinationAddressIn_SOUTH[9]), .C1(n3756), .Y(n1831) );
  OAI221XLTS U2919 ( .A0(n3693), .A1(n153), .B0(n3764), .B1(n906), .C0(n1833), 
        .Y(n2551) );
  AOI222XLTS U2920 ( .A0(n4026), .A1(n3708), .B0(n3985), .B1(n3716), .C0(
        destinationAddressIn_SOUTH[11]), .C1(n3756), .Y(n1833) );
  OAI221XLTS U2921 ( .A0(n3694), .A1(n160), .B0(n3764), .B1(n905), .C0(n1830), 
        .Y(n2554) );
  AOI222XLTS U2922 ( .A0(n4017), .A1(n3707), .B0(n3976), .B1(n3717), .C0(
        destinationAddressIn_SOUTH[8]), .C1(n3755), .Y(n1830) );
  OAI221XLTS U2923 ( .A0(n3695), .A1(n146), .B0(n3777), .B1(n904), .C0(n1829), 
        .Y(n2555) );
  AOI222XLTS U2924 ( .A0(n4014), .A1(n3707), .B0(n3973), .B1(n3717), .C0(n4240), .C1(n3755), .Y(n1829) );
  OAI221XLTS U2925 ( .A0(n3695), .A1(n148), .B0(n3777), .B1(n903), .C0(n1828), 
        .Y(n2556) );
  AOI222XLTS U2926 ( .A0(n4011), .A1(n3707), .B0(n3970), .B1(n3717), .C0(n4237), .C1(n3755), .Y(n1828) );
  OAI221XLTS U2927 ( .A0(n3694), .A1(n159), .B0(n3764), .B1(n833), .C0(n1832), 
        .Y(n2552) );
  AOI222XLTS U2928 ( .A0(n4023), .A1(n3708), .B0(n3982), .B1(n3716), .C0(
        destinationAddressIn_SOUTH[10]), .C1(n3756), .Y(n1832) );
  OAI221XLTS U2929 ( .A0(n3693), .A1(n157), .B0(n3776), .B1(n907), .C0(n1834), 
        .Y(n2550) );
  AOI222XLTS U2930 ( .A0(n4029), .A1(n3708), .B0(n3988), .B1(n3716), .C0(
        destinationAddressIn_SOUTH[12]), .C1(n3756), .Y(n1834) );
  OAI221XLTS U2931 ( .A0(n3693), .A1(n151), .B0(n3778), .B1(n702), .C0(n1835), 
        .Y(n2549) );
  AOI222XLTS U2932 ( .A0(n4032), .A1(n3714), .B0(n3991), .B1(n3716), .C0(
        destinationAddressIn_SOUTH[13]), .C1(n3763), .Y(n1835) );
  AOI22X1TS U2933 ( .A0(n3551), .A1(n4050), .B0(n3828), .B1(n4087), .Y(n1144)
         );
  AOI222XLTS U2934 ( .A0(n3600), .A1(n4604), .B0(n3592), .B1(n43), .C0(n3571), 
        .C1(n4201), .Y(n1145) );
  AOI22X1TS U2935 ( .A0(n3565), .A1(n4047), .B0(n3828), .B1(n4084), .Y(n1142)
         );
  AOI222XLTS U2936 ( .A0(n3599), .A1(n4601), .B0(n3592), .B1(n37), .C0(n3571), 
        .C1(n4198), .Y(n1143) );
  AOI22X1TS U2937 ( .A0(n3562), .A1(n4044), .B0(n3827), .B1(n4081), .Y(n1140)
         );
  AOI222XLTS U2938 ( .A0(n3599), .A1(n4596), .B0(n3591), .B1(n32), .C0(n3570), 
        .C1(n4195), .Y(n1141) );
  AOI22X1TS U2939 ( .A0(n3563), .A1(n4041), .B0(n3827), .B1(n4078), .Y(n1138)
         );
  AOI222XLTS U2940 ( .A0(n3599), .A1(n4592), .B0(n3591), .B1(n27), .C0(n3570), 
        .C1(n4192), .Y(n1139) );
  AOI22X1TS U2941 ( .A0(n3564), .A1(n4038), .B0(n3827), .B1(n4075), .Y(n1136)
         );
  AOI222XLTS U2942 ( .A0(n3599), .A1(n4587), .B0(n3591), .B1(n22), .C0(n3570), 
        .C1(n4189), .Y(n1137) );
  AOI22X1TS U2943 ( .A0(n3551), .A1(n4035), .B0(n3827), .B1(n4072), .Y(n1130)
         );
  AOI222XLTS U2944 ( .A0(n3600), .A1(n4584), .B0(n3592), .B1(n17), .C0(n3571), 
        .C1(n4186), .Y(n1131) );
  AOI222XLTS U2945 ( .A0(n4233), .A1(n3340), .B0(n3328), .B1(n38), .C0(n4006), 
        .C1(n3314), .Y(n1968) );
  AOI22X1TS U2946 ( .A0(n3287), .A1(n4200), .B0(n3850), .B1(n4087), .Y(n1208)
         );
  AOI222XLTS U2947 ( .A0(n3334), .A1(n4604), .B0(n3332), .B1(n44), .C0(n3306), 
        .C1(n4051), .Y(n1209) );
  AOI22X1TS U2948 ( .A0(n3286), .A1(n4197), .B0(n3851), .B1(n4084), .Y(n1206)
         );
  AOI222XLTS U2949 ( .A0(n3345), .A1(n4601), .B0(n3329), .B1(n39), .C0(n3306), 
        .C1(n4048), .Y(n1207) );
  AOI22X1TS U2950 ( .A0(n3286), .A1(n4194), .B0(n3840), .B1(n4081), .Y(n1204)
         );
  AOI222XLTS U2951 ( .A0(n3344), .A1(n4596), .B0(n3327), .B1(n33), .C0(n3305), 
        .C1(n4045), .Y(n1205) );
  AOI22X1TS U2952 ( .A0(n3286), .A1(n4191), .B0(n3840), .B1(n4078), .Y(n1202)
         );
  AOI222XLTS U2953 ( .A0(n3348), .A1(n4592), .B0(n3327), .B1(n28), .C0(n3305), 
        .C1(n4042), .Y(n1203) );
  AOI22X1TS U2954 ( .A0(n3286), .A1(n4188), .B0(n3840), .B1(n4075), .Y(n1200)
         );
  AOI222XLTS U2955 ( .A0(n3345), .A1(n4587), .B0(n3327), .B1(n23), .C0(n3305), 
        .C1(n4039), .Y(n1201) );
  AOI22X1TS U2956 ( .A0(n3287), .A1(n4185), .B0(n3840), .B1(n4072), .Y(n1194)
         );
  AOI222XLTS U2957 ( .A0(n3334), .A1(n4584), .B0(n3329), .B1(n18), .C0(n3306), 
        .C1(n4036), .Y(n1195) );
  AOI22X1TS U2958 ( .A0(n3966), .A1(n3459), .B0(n4235), .B1(n3441), .Y(n1921)
         );
  AOI222XLTS U2959 ( .A0(n3808), .A1(n45), .B0(n4070), .B1(n3822), .C0(n6250), 
        .C1(n186), .Y(n1922) );
  AOI22X1TS U2960 ( .A0(n3963), .A1(n3459), .B0(n4232), .B1(n3441), .Y(n1919)
         );
  AOI222XLTS U2961 ( .A0(n3796), .A1(n40), .B0(n4067), .B1(n3823), .C0(n6251), 
        .C1(n190), .Y(n1920) );
  AOI22X1TS U2962 ( .A0(n3960), .A1(n3459), .B0(n4229), .B1(n3441), .Y(n1917)
         );
  AOI222XLTS U2963 ( .A0(n3796), .A1(n35), .B0(n4064), .B1(n679), .C0(n6252), 
        .C1(n136), .Y(n1918) );
  AOI22X1TS U2964 ( .A0(n3954), .A1(n3458), .B0(n4223), .B1(n3445), .Y(n1913)
         );
  AOI222XLTS U2965 ( .A0(n3795), .A1(n25), .B0(n4058), .B1(n3812), .C0(n6253), 
        .C1(n187), .Y(n1914) );
  AOI22X1TS U2966 ( .A0(n3951), .A1(n3458), .B0(n4220), .B1(n3449), .Y(n1911)
         );
  AOI222XLTS U2967 ( .A0(n3796), .A1(n20), .B0(n4055), .B1(n3812), .C0(n6254), 
        .C1(n3810), .Y(n1912) );
  AOI22X1TS U2968 ( .A0(n3957), .A1(n3459), .B0(n4226), .B1(n3441), .Y(n1915)
         );
  AOI222XLTS U2969 ( .A0(n3796), .A1(n30), .B0(n4061), .B1(n679), .C0(n6291), 
        .C1(n188), .Y(n1916) );
  AOI22X1TS U2970 ( .A0(n3658), .A1(n38), .B0(n3634), .B1(n4047), .Y(n1125) );
  AOI222XLTS U2971 ( .A0(\requesterAddressbuffer[6][4] ), .A1(n3199), .B0(
        n3678), .B1(n4597), .C0(n3872), .C1(n4085), .Y(n1126) );
  AOI22X1TS U2972 ( .A0(n3663), .A1(n28), .B0(n3634), .B1(n4041), .Y(n1121) );
  AOI222XLTS U2973 ( .A0(\requesterAddressbuffer[6][2] ), .A1(n3197), .B0(
        n3681), .B1(n4589), .C0(n3872), .C1(n4079), .Y(n1122) );
  AOI22X1TS U2974 ( .A0(n3664), .A1(n23), .B0(n3635), .B1(n4038), .Y(n1119) );
  AOI222XLTS U2975 ( .A0(\requesterAddressbuffer[6][1] ), .A1(n3196), .B0(
        n3679), .B1(n4585), .C0(n3872), .C1(n4076), .Y(n1120) );
  AOI22X1TS U2976 ( .A0(n3662), .A1(n43), .B0(n4008), .B1(n3635), .Y(n1852) );
  AOI222XLTS U2977 ( .A0(n2992), .A1(n3198), .B0(n4236), .B1(n3674), .C0(n4069), .C1(n3874), .Y(n1853) );
  AOI22X1TS U2978 ( .A0(n4235), .A1(n3210), .B0(n4009), .B1(n3944), .Y(n1991)
         );
  AOI222XLTS U2979 ( .A0(n3966), .A1(n3257), .B0(n4070), .B1(n3236), .C0(n3220), .C1(n44), .Y(n1992) );
  AOI22X1TS U2980 ( .A0(n3662), .A1(n38), .B0(n4005), .B1(n3636), .Y(n1850) );
  AOI222XLTS U2981 ( .A0(n2994), .A1(n3201), .B0(n4233), .B1(n3675), .C0(n4066), .C1(n3874), .Y(n1851) );
  AOI22X1TS U2982 ( .A0(n3663), .A1(n33), .B0(n4002), .B1(n3636), .Y(n1848) );
  AOI222XLTS U2983 ( .A0(n2996), .A1(n3201), .B0(n4230), .B1(n3675), .C0(n4063), .C1(n3874), .Y(n1849) );
  AOI22X1TS U2984 ( .A0(n3660), .A1(n29), .B0(n3999), .B1(n3635), .Y(n1846) );
  AOI222XLTS U2985 ( .A0(n2998), .A1(n987), .B0(n4227), .B1(n3675), .C0(n4060), 
        .C1(n3874), .Y(n1847) );
  AOI22X1TS U2986 ( .A0(n3662), .A1(n22), .B0(n3996), .B1(n3636), .Y(n1844) );
  AOI222XLTS U2987 ( .A0(n3000), .A1(n3202), .B0(n4224), .B1(n3674), .C0(n4057), .C1(n3873), .Y(n1845) );
  AOI22X1TS U2988 ( .A0(n3659), .A1(n17), .B0(n3993), .B1(n3636), .Y(n1842) );
  AOI222XLTS U2989 ( .A0(n3002), .A1(n3200), .B0(n4221), .B1(n3674), .C0(n4054), .C1(n3873), .Y(n1843) );
  AOI22X1TS U2990 ( .A0(n4229), .A1(n3210), .B0(n4003), .B1(n3944), .Y(n1987)
         );
  AOI222XLTS U2991 ( .A0(n3960), .A1(n3257), .B0(n4064), .B1(n3236), .C0(n3222), .C1(n34), .Y(n1988) );
  AOI22X1TS U2992 ( .A0(n4226), .A1(n3210), .B0(n4000), .B1(n3944), .Y(n1985)
         );
  AOI222XLTS U2993 ( .A0(n3957), .A1(n3257), .B0(n4061), .B1(n3236), .C0(n3222), .C1(n29), .Y(n1986) );
  AOI22X1TS U2994 ( .A0(n4223), .A1(n3209), .B0(n3997), .B1(n3945), .Y(n1983)
         );
  AOI222XLTS U2995 ( .A0(n3954), .A1(n3267), .B0(n4058), .B1(n3237), .C0(n3221), .C1(n24), .Y(n1984) );
  AOI22X1TS U2996 ( .A0(n4579), .A1(n3209), .B0(n4354), .B1(n3945), .Y(n1289)
         );
  AOI222XLTS U2997 ( .A0(n4459), .A1(n3264), .B0(n4184), .B1(n3237), .C0(n510), 
        .C1(n3225), .Y(n1290) );
  AOI22X1TS U2998 ( .A0(n4576), .A1(n3209), .B0(n4351), .B1(n3946), .Y(n1287)
         );
  AOI222XLTS U2999 ( .A0(n4456), .A1(n1213), .B0(n4181), .B1(n3238), .C0(n512), 
        .C1(n3223), .Y(n1288) );
  AOI22X1TS U3000 ( .A0(n4571), .A1(n3208), .B0(n4348), .B1(n3943), .Y(n1285)
         );
  AOI222XLTS U3001 ( .A0(n4452), .A1(n3262), .B0(n4178), .B1(n3238), .C0(n514), 
        .C1(n3223), .Y(n1286) );
  AOI22X1TS U3002 ( .A0(n4560), .A1(n3208), .B0(n4339), .B1(n3943), .Y(n1279)
         );
  AOI222XLTS U3003 ( .A0(n4441), .A1(n3263), .B0(n4169), .B1(n3239), .C0(n516), 
        .C1(n3227), .Y(n1280) );
  AOI22X1TS U3004 ( .A0(n4556), .A1(n3207), .B0(n4336), .B1(n3942), .Y(n1277)
         );
  AOI222XLTS U3005 ( .A0(n4438), .A1(n3267), .B0(n4166), .B1(n3239), .C0(n518), 
        .C1(n3223), .Y(n1278) );
  AOI22X1TS U3006 ( .A0(n4552), .A1(n3207), .B0(n4333), .B1(n3942), .Y(n1275)
         );
  AOI222XLTS U3007 ( .A0(n4434), .A1(n3266), .B0(n4163), .B1(n3239), .C0(n520), 
        .C1(n3224), .Y(n1276) );
  AOI22X1TS U3008 ( .A0(n4544), .A1(n3207), .B0(n4327), .B1(n3942), .Y(n1271)
         );
  AOI222XLTS U3009 ( .A0(n4426), .A1(n3264), .B0(n4157), .B1(n3250), .C0(n522), 
        .C1(n3224), .Y(n1272) );
  AOI22X1TS U3010 ( .A0(n4541), .A1(n3206), .B0(n4324), .B1(n3941), .Y(n1269)
         );
  AOI222XLTS U3011 ( .A0(n4423), .A1(n3267), .B0(n4154), .B1(n3250), .C0(n524), 
        .C1(n3228), .Y(n1270) );
  AOI22X1TS U3012 ( .A0(n4533), .A1(n3206), .B0(n4318), .B1(n3941), .Y(n1265)
         );
  AOI222XLTS U3013 ( .A0(n4415), .A1(n3261), .B0(n4148), .B1(n3245), .C0(n526), 
        .C1(n3228), .Y(n1266) );
  AOI22X1TS U3014 ( .A0(n4529), .A1(n3205), .B0(n4315), .B1(n3941), .Y(n1263)
         );
  AOI222XLTS U3015 ( .A0(n4412), .A1(n3256), .B0(n4145), .B1(n3244), .C0(n528), 
        .C1(n3228), .Y(n1264) );
  AOI22X1TS U3016 ( .A0(n4525), .A1(n3205), .B0(n4312), .B1(n3940), .Y(n1261)
         );
  AOI222XLTS U3017 ( .A0(n4409), .A1(n3256), .B0(n4142), .B1(n3244), .C0(n530), 
        .C1(n3232), .Y(n1262) );
  AOI22X1TS U3018 ( .A0(n4522), .A1(n3205), .B0(n4309), .B1(n3940), .Y(n1259)
         );
  AOI222XLTS U3019 ( .A0(n4406), .A1(n3256), .B0(n4139), .B1(n3245), .C0(n532), 
        .C1(n3228), .Y(n1260) );
  AOI22X1TS U3020 ( .A0(n4519), .A1(n3205), .B0(n4306), .B1(n3940), .Y(n1257)
         );
  AOI222XLTS U3021 ( .A0(n4403), .A1(n3256), .B0(n4136), .B1(n3246), .C0(n534), 
        .C1(n3227), .Y(n1258) );
  AOI22X1TS U3022 ( .A0(n4514), .A1(n3217), .B0(n4303), .B1(n3940), .Y(n1255)
         );
  AOI222XLTS U3023 ( .A0(n4400), .A1(n3255), .B0(n4133), .B1(n3240), .C0(n536), 
        .C1(n3229), .Y(n1256) );
  AOI22X1TS U3024 ( .A0(n4511), .A1(n3213), .B0(n4300), .B1(n3949), .Y(n1253)
         );
  AOI222XLTS U3025 ( .A0(n4397), .A1(n3255), .B0(n4130), .B1(n3240), .C0(n538), 
        .C1(n3226), .Y(n1254) );
  AOI22X1TS U3026 ( .A0(n4507), .A1(n3214), .B0(n4297), .B1(n3948), .Y(n1251)
         );
  AOI222XLTS U3027 ( .A0(n4394), .A1(n3255), .B0(n4127), .B1(n3240), .C0(n540), 
        .C1(n3233), .Y(n1252) );
  AOI22X1TS U3028 ( .A0(n4504), .A1(n3213), .B0(n4294), .B1(n3949), .Y(n1249)
         );
  AOI222XLTS U3029 ( .A0(n4391), .A1(n3255), .B0(n4124), .B1(n3240), .C0(n542), 
        .C1(n3229), .Y(n1250) );
  AOI22X1TS U3030 ( .A0(n4499), .A1(n3218), .B0(n4291), .B1(n660), .Y(n1247)
         );
  AOI222XLTS U3031 ( .A0(n4388), .A1(n3254), .B0(n4121), .B1(n3241), .C0(n544), 
        .C1(n3225), .Y(n1248) );
  AOI22X1TS U3032 ( .A0(n4493), .A1(n3217), .B0(n4285), .B1(n3939), .Y(n1243)
         );
  AOI222XLTS U3033 ( .A0(n4382), .A1(n3254), .B0(n4115), .B1(n3241), .C0(n546), 
        .C1(n3227), .Y(n1244) );
  AOI22X1TS U3034 ( .A0(n4489), .A1(n3215), .B0(n4282), .B1(n3939), .Y(n1241)
         );
  AOI222XLTS U3035 ( .A0(n4379), .A1(n3254), .B0(n4112), .B1(n3241), .C0(n548), 
        .C1(n3226), .Y(n1242) );
  AOI22X1TS U3036 ( .A0(n4486), .A1(n3216), .B0(n4279), .B1(n3939), .Y(n1239)
         );
  AOI222XLTS U3037 ( .A0(n4376), .A1(n3254), .B0(n4109), .B1(n3242), .C0(n659), 
        .C1(n3230), .Y(n1240) );
  AOI22X1TS U3038 ( .A0(n4478), .A1(n3213), .B0(n4273), .B1(n3949), .Y(n1235)
         );
  AOI222XLTS U3039 ( .A0(n4370), .A1(n3253), .B0(n4103), .B1(n3242), .C0(n663), 
        .C1(n3231), .Y(n1236) );
  AOI22X1TS U3040 ( .A0(n4474), .A1(n3216), .B0(n4270), .B1(n3948), .Y(n1233)
         );
  AOI222XLTS U3041 ( .A0(n4367), .A1(n3253), .B0(n4100), .B1(n3242), .C0(n672), 
        .C1(n3225), .Y(n1234) );
  AOI22X1TS U3042 ( .A0(n4232), .A1(n3210), .B0(n4006), .B1(n3944), .Y(n1989)
         );
  AOI222XLTS U3043 ( .A0(n3963), .A1(n3257), .B0(n4067), .B1(n3236), .C0(n3222), .C1(n39), .Y(n1990) );
  AOI22X1TS U3044 ( .A0(n3515), .A1(n35), .B0(n3486), .B1(n4194), .Y(n1156) );
  AOI222XLTS U3045 ( .A0(n2925), .A1(n3892), .B0(n3527), .B1(n4596), .C0(n3894), .C1(n4082), .Y(n1157) );
  AOI22X1TS U3046 ( .A0(n3516), .A1(n30), .B0(n3486), .B1(n4191), .Y(n1154) );
  AOI222XLTS U3047 ( .A0(n2923), .A1(n3888), .B0(n3527), .B1(n4592), .C0(n3894), .C1(n4079), .Y(n1155) );
  AOI22X1TS U3048 ( .A0(n3515), .A1(n25), .B0(n3486), .B1(n4188), .Y(n1152) );
  AOI222XLTS U3049 ( .A0(n2924), .A1(n3892), .B0(n3527), .B1(n4587), .C0(n3894), .C1(n4076), .Y(n1153) );
  AOI22X1TS U3050 ( .A0(n3503), .A1(n20), .B0(n3487), .B1(n4185), .Y(n1147) );
  AOI222XLTS U3051 ( .A0(n2926), .A1(n3883), .B0(n3527), .B1(n4584), .C0(n3894), .C1(n4073), .Y(n1148) );
  AOI22X1TS U3052 ( .A0(n3452), .A1(n4194), .B0(n3435), .B1(n4594), .Y(n1171)
         );
  AOI222XLTS U3053 ( .A0(n3806), .A1(n34), .B0(n3821), .B1(n4081), .C0(
        \requesterAddressbuffer[3][3] ), .C1(n135), .Y(n1172) );
  AOI22X1TS U3054 ( .A0(n3452), .A1(n4191), .B0(n3435), .B1(n4591), .Y(n1169)
         );
  AOI222XLTS U3055 ( .A0(n3807), .A1(n29), .B0(n3821), .B1(n4078), .C0(
        \requesterAddressbuffer[3][2] ), .C1(n3810), .Y(n1170) );
  AOI22X1TS U3056 ( .A0(n3452), .A1(n4188), .B0(n3435), .B1(n4586), .Y(n1167)
         );
  AOI222XLTS U3057 ( .A0(n3807), .A1(n24), .B0(n3821), .B1(n4075), .C0(
        \requesterAddressbuffer[3][1] ), .C1(n186), .Y(n1168) );
  AOI22X1TS U3058 ( .A0(n3453), .A1(n4185), .B0(n3436), .B1(n4583), .Y(n1163)
         );
  AOI222XLTS U3059 ( .A0(n3795), .A1(n19), .B0(n3821), .B1(n4072), .C0(
        \requesterAddressbuffer[3][0] ), .C1(n190), .Y(n1164) );
  AOI22X1TS U3060 ( .A0(n3503), .A1(n45), .B0(n3487), .B1(n4200), .Y(n1160) );
  AOI222XLTS U3061 ( .A0(n2921), .A1(n3888), .B0(n3530), .B1(n4604), .C0(n3895), .C1(n4088), .Y(n1161) );
  AOI22X1TS U3062 ( .A0(n3503), .A1(n40), .B0(n3486), .B1(n4197), .Y(n1158) );
  AOI222XLTS U3063 ( .A0(n2922), .A1(n3889), .B0(n3532), .B1(n4601), .C0(n3895), .C1(n4085), .Y(n1159) );
  AOI22X1TS U3064 ( .A0(n3452), .A1(n4197), .B0(n3435), .B1(n4598), .Y(n1173)
         );
  AOI222XLTS U3065 ( .A0(n3795), .A1(n39), .B0(n3820), .B1(n4084), .C0(
        \requesterAddressbuffer[3][4] ), .C1(n134), .Y(n1174) );
  AOI22X1TS U3066 ( .A0(n3453), .A1(n4200), .B0(n3436), .B1(n4603), .Y(n1175)
         );
  AOI222XLTS U3067 ( .A0(n3795), .A1(n44), .B0(n3820), .B1(n4087), .C0(
        \requesterAddressbuffer[3][5] ), .C1(n3811), .Y(n1176) );
  AOI22X1TS U3068 ( .A0(n3387), .A1(n37), .B0(n3369), .B1(n4047), .Y(n1189) );
  AOI222XLTS U3069 ( .A0(\requesterAddressbuffer[2][4] ), .A1(n3918), .B0(
        n3409), .B1(n4601), .C0(n3925), .C1(n4085), .Y(n1190) );
  AOI22X1TS U3070 ( .A0(n3386), .A1(n22), .B0(n3369), .B1(n4038), .Y(n1183) );
  AOI222XLTS U3071 ( .A0(\requesterAddressbuffer[2][1] ), .A1(n3919), .B0(
        n3408), .B1(n4587), .C0(n3924), .C1(n4076), .Y(n1184) );
  AOI22X1TS U3072 ( .A0(n3387), .A1(n17), .B0(n3370), .B1(n4035), .Y(n1178) );
  AOI222XLTS U3073 ( .A0(\requesterAddressbuffer[2][0] ), .A1(n3912), .B0(
        n3408), .B1(n4584), .C0(n3924), .C1(n4073), .Y(n1179) );
  AOI22X1TS U3074 ( .A0(n3387), .A1(n42), .B0(n3370), .B1(n4050), .Y(n1191) );
  AOI222XLTS U3075 ( .A0(\requesterAddressbuffer[2][5] ), .A1(n3918), .B0(
        n3412), .B1(n4604), .C0(n3925), .C1(n4088), .Y(n1192) );
  AOI22X1TS U3076 ( .A0(n3386), .A1(n32), .B0(n3369), .B1(n4044), .Y(n1187) );
  AOI222XLTS U3077 ( .A0(\requesterAddressbuffer[2][3] ), .A1(n3919), .B0(
        n3408), .B1(n4596), .C0(n3924), .C1(n4082), .Y(n1188) );
  AOI22X1TS U3078 ( .A0(n3386), .A1(n27), .B0(n3369), .B1(n4041), .Y(n1185) );
  AOI222XLTS U3079 ( .A0(\requesterAddressbuffer[2][2] ), .A1(n664), .B0(n3408), .B1(n4592), .C0(n3924), .C1(n4079), .Y(n1186) );
  AOI22X1TS U3080 ( .A0(n3661), .A1(n18), .B0(n3634), .B1(n4035), .Y(n1114) );
  AOI222XLTS U3081 ( .A0(\requesterAddressbuffer[6][0] ), .A1(n3200), .B0(
        n1116), .B1(n4582), .C0(n3873), .C1(n4073), .Y(n1115) );
  AOI22X1TS U3082 ( .A0(n3658), .A1(n43), .B0(n3635), .B1(n4050), .Y(n1127) );
  AOI222XLTS U3083 ( .A0(\requesterAddressbuffer[6][5] ), .A1(n3200), .B0(
        n3675), .B1(n4602), .C0(n3873), .C1(n4088), .Y(n1128) );
  AOI22X1TS U3084 ( .A0(n3662), .A1(n33), .B0(n3634), .B1(n4044), .Y(n1123) );
  AOI222XLTS U3085 ( .A0(\requesterAddressbuffer[6][3] ), .A1(n3200), .B0(
        n3678), .B1(n4593), .C0(n3872), .C1(n4082), .Y(n1124) );
  AOI22X1TS U3086 ( .A0(n4261), .A1(n3700), .B0(n4090), .B1(n3691), .Y(n1676)
         );
  AOI222XLTS U3087 ( .A0(n4463), .A1(n3748), .B0(n677), .B1(n3738), .C0(n4358), 
        .C1(n3728), .Y(n1677) );
  AOI22X1TS U3088 ( .A0(n4300), .A1(n3701), .B0(n4129), .B1(n3688), .Y(n1702)
         );
  AOI222XLTS U3089 ( .A0(n4512), .A1(n3751), .B0(n538), .B1(n3741), .C0(n4397), 
        .C1(n3719), .Y(n1703) );
  AOI22X1TS U3090 ( .A0(n4303), .A1(n3701), .B0(n4132), .B1(n3687), .Y(n1704)
         );
  AOI222XLTS U3091 ( .A0(n4515), .A1(n3751), .B0(n536), .B1(n3741), .C0(n4400), 
        .C1(n3719), .Y(n1705) );
  AOI22X1TS U3092 ( .A0(n4306), .A1(n3702), .B0(n4135), .B1(n3687), .Y(n1706)
         );
  AOI222XLTS U3093 ( .A0(n4520), .A1(n3752), .B0(n534), .B1(n3744), .C0(n4403), 
        .C1(n3719), .Y(n1707) );
  AOI22X1TS U3094 ( .A0(n4050), .A1(n3700), .B0(n4087), .B1(n3691), .Y(n1111)
         );
  AOI222XLTS U3095 ( .A0(n4603), .A1(n3748), .B0(n42), .B1(n3738), .C0(n4201), 
        .C1(n3726), .Y(n1112) );
  AOI22X1TS U3096 ( .A0(n4047), .A1(n3699), .B0(n4084), .B1(n3691), .Y(n1109)
         );
  AOI222XLTS U3097 ( .A0(n4598), .A1(n3747), .B0(n37), .B1(n3738), .C0(n4198), 
        .C1(n3729), .Y(n1110) );
  AOI22X1TS U3098 ( .A0(n4041), .A1(n3699), .B0(n4078), .B1(n3692), .Y(n1105)
         );
  AOI222XLTS U3099 ( .A0(n4591), .A1(n3747), .B0(n27), .B1(n3739), .C0(n4192), 
        .C1(n3729), .Y(n1106) );
  AOI22X1TS U3100 ( .A0(n4044), .A1(n3699), .B0(n4081), .B1(n3692), .Y(n1107)
         );
  AOI222XLTS U3101 ( .A0(n4594), .A1(n3747), .B0(n32), .B1(n3744), .C0(n4195), 
        .C1(n3729), .Y(n1108) );
  AOI22X1TS U3102 ( .A0(n4038), .A1(n3699), .B0(n4075), .B1(n3692), .Y(n1103)
         );
  AOI222XLTS U3103 ( .A0(n4586), .A1(n3747), .B0(n22), .B1(n3739), .C0(n4189), 
        .C1(n3729), .Y(n1104) );
  AOI22X1TS U3104 ( .A0(n4035), .A1(n3703), .B0(n4072), .B1(n3692), .Y(n1096)
         );
  AOI222XLTS U3105 ( .A0(n4583), .A1(n3759), .B0(n17), .B1(n3744), .C0(n4186), 
        .C1(n3719), .Y(n1097) );
  AOI22X1TS U3106 ( .A0(n3993), .A1(n3706), .B0(n4054), .B1(n3683), .Y(n1814)
         );
  AOI222XLTS U3107 ( .A0(n4220), .A1(n3753), .B0(n18), .B1(n3734), .C0(n3952), 
        .C1(n3724), .Y(n1815) );
  AOI22X1TS U3108 ( .A0(n4008), .A1(n3709), .B0(n4069), .B1(n3682), .Y(n1824)
         );
  AOI222XLTS U3109 ( .A0(n4235), .A1(n3754), .B0(n43), .B1(n3733), .C0(n3967), 
        .C1(n3727), .Y(n1825) );
  AOI22X1TS U3110 ( .A0(n4002), .A1(n3710), .B0(n4063), .B1(n3682), .Y(n1820)
         );
  AOI222XLTS U3111 ( .A0(n4229), .A1(n3754), .B0(n33), .B1(n3733), .C0(n3961), 
        .C1(n3724), .Y(n1821) );
  AOI22X1TS U3112 ( .A0(n3999), .A1(n3709), .B0(n4060), .B1(n3682), .Y(n1818)
         );
  AOI222XLTS U3113 ( .A0(n4226), .A1(n3754), .B0(n28), .B1(n3733), .C0(n3958), 
        .C1(n3724), .Y(n1819) );
  AOI22X1TS U3114 ( .A0(n3996), .A1(n3706), .B0(n4057), .B1(n3683), .Y(n1816)
         );
  AOI222XLTS U3115 ( .A0(n4223), .A1(n3753), .B0(n23), .B1(n3734), .C0(n3955), 
        .C1(n3724), .Y(n1817) );
  AOI22X1TS U3116 ( .A0(n4354), .A1(n3706), .B0(n4183), .B1(n3683), .Y(n1738)
         );
  AOI222XLTS U3117 ( .A0(n4580), .A1(n3753), .B0(n510), .B1(n3734), .C0(n4459), 
        .C1(n3723), .Y(n1739) );
  AOI22X1TS U3118 ( .A0(n4351), .A1(n3706), .B0(n4180), .B1(n3683), .Y(n1736)
         );
  AOI222XLTS U3119 ( .A0(n4577), .A1(n3753), .B0(n512), .B1(n3734), .C0(n4456), 
        .C1(n3723), .Y(n1737) );
  AOI22X1TS U3120 ( .A0(n4348), .A1(n3705), .B0(n4177), .B1(n3684), .Y(n1734)
         );
  AOI222XLTS U3121 ( .A0(n4573), .A1(n3759), .B0(n514), .B1(n3735), .C0(n4452), 
        .C1(n3723), .Y(n1735) );
  AOI22X1TS U3122 ( .A0(n4345), .A1(n3705), .B0(n4174), .B1(n3684), .Y(n1732)
         );
  AOI222XLTS U3123 ( .A0(n4569), .A1(n3757), .B0(n496), .B1(n3735), .C0(n4449), 
        .C1(n3723), .Y(n1733) );
  AOI22X1TS U3124 ( .A0(n4342), .A1(n3705), .B0(n4171), .B1(n3684), .Y(n1730)
         );
  AOI222XLTS U3125 ( .A0(n4565), .A1(n3757), .B0(n498), .B1(n3735), .C0(n4445), 
        .C1(n3722), .Y(n1731) );
  AOI22X1TS U3126 ( .A0(n4339), .A1(n3705), .B0(n4168), .B1(n3684), .Y(n1728)
         );
  AOI222XLTS U3127 ( .A0(n4561), .A1(n3757), .B0(n516), .B1(n3735), .C0(n4441), 
        .C1(n3722), .Y(n1729) );
  AOI22X1TS U3128 ( .A0(n4336), .A1(n3704), .B0(n4165), .B1(n3685), .Y(n1726)
         );
  AOI222XLTS U3129 ( .A0(n4558), .A1(n3762), .B0(n518), .B1(n3736), .C0(n4438), 
        .C1(n3722), .Y(n1727) );
  AOI22X1TS U3130 ( .A0(n4333), .A1(n3704), .B0(n4162), .B1(n3685), .Y(n1724)
         );
  AOI222XLTS U3131 ( .A0(n4553), .A1(n3760), .B0(n520), .B1(n3736), .C0(n4434), 
        .C1(n3722), .Y(n1725) );
  AOI22X1TS U3132 ( .A0(n4330), .A1(n3704), .B0(n4159), .B1(n3685), .Y(n1722)
         );
  AOI222XLTS U3133 ( .A0(n4550), .A1(n3761), .B0(n500), .B1(n3736), .C0(n4430), 
        .C1(n3721), .Y(n1723) );
  AOI22X1TS U3134 ( .A0(n4327), .A1(n3704), .B0(n4156), .B1(n3685), .Y(n1720)
         );
  AOI222XLTS U3135 ( .A0(n4546), .A1(n3758), .B0(n522), .B1(n3736), .C0(n4426), 
        .C1(n3721), .Y(n1721) );
  AOI22X1TS U3136 ( .A0(n4324), .A1(n3703), .B0(n4153), .B1(n3686), .Y(n1718)
         );
  AOI222XLTS U3137 ( .A0(n4542), .A1(n3759), .B0(n524), .B1(n3737), .C0(n4423), 
        .C1(n3721), .Y(n1719) );
  AOI22X1TS U3138 ( .A0(n4321), .A1(n3703), .B0(n4150), .B1(n3686), .Y(n1716)
         );
  AOI222XLTS U3139 ( .A0(n4538), .A1(n3758), .B0(n502), .B1(n3737), .C0(n4418), 
        .C1(n3721), .Y(n1717) );
  AOI22X1TS U3140 ( .A0(n4318), .A1(n3703), .B0(n4147), .B1(n3686), .Y(n1714)
         );
  AOI222XLTS U3141 ( .A0(n4534), .A1(n3762), .B0(n526), .B1(n3737), .C0(n4415), 
        .C1(n3720), .Y(n1715) );
  AOI22X1TS U3142 ( .A0(n4315), .A1(n3702), .B0(n4144), .B1(n3686), .Y(n1712)
         );
  AOI222XLTS U3143 ( .A0(n4531), .A1(n3752), .B0(n528), .B1(n3737), .C0(n4412), 
        .C1(n3720), .Y(n1713) );
  AOI22X1TS U3144 ( .A0(n4312), .A1(n3702), .B0(n4141), .B1(n3687), .Y(n1710)
         );
  AOI222XLTS U3145 ( .A0(n4526), .A1(n3752), .B0(n530), .B1(n3745), .C0(n4409), 
        .C1(n3720), .Y(n1711) );
  AOI22X1TS U3146 ( .A0(n4309), .A1(n3702), .B0(n4138), .B1(n3687), .Y(n1708)
         );
  AOI222XLTS U3147 ( .A0(n4523), .A1(n3752), .B0(n532), .B1(n3739), .C0(n4406), 
        .C1(n3720), .Y(n1709) );
  AOI22X1TS U3148 ( .A0(n4297), .A1(n3701), .B0(n4126), .B1(n3688), .Y(n1700)
         );
  AOI222XLTS U3149 ( .A0(n4508), .A1(n3751), .B0(n540), .B1(n3741), .C0(n4394), 
        .C1(n3718), .Y(n1701) );
  AOI22X1TS U3150 ( .A0(n4294), .A1(n3701), .B0(n4123), .B1(n3688), .Y(n1698)
         );
  AOI222XLTS U3151 ( .A0(n4505), .A1(n3751), .B0(n542), .B1(n3743), .C0(n4391), 
        .C1(n3718), .Y(n1699) );
  AOI22X1TS U3152 ( .A0(n4291), .A1(n3712), .B0(n4120), .B1(n3688), .Y(n1696)
         );
  AOI222XLTS U3153 ( .A0(n4502), .A1(n3750), .B0(n544), .B1(n3746), .C0(n4388), 
        .C1(n3718), .Y(n1697) );
  AOI22X1TS U3154 ( .A0(n4288), .A1(n3712), .B0(n4117), .B1(n3689), .Y(n1694)
         );
  AOI222XLTS U3155 ( .A0(n4497), .A1(n3750), .B0(n504), .B1(n3740), .C0(n4385), 
        .C1(n3718), .Y(n1695) );
  AOI22X1TS U3156 ( .A0(n4285), .A1(n3711), .B0(n4114), .B1(n3689), .Y(n1692)
         );
  AOI222XLTS U3157 ( .A0(n4494), .A1(n3750), .B0(n546), .B1(n3740), .C0(n4382), 
        .C1(n3726), .Y(n1693) );
  AOI22X1TS U3158 ( .A0(n4282), .A1(n3713), .B0(n4111), .B1(n3689), .Y(n1690)
         );
  AOI222XLTS U3159 ( .A0(n4490), .A1(n3750), .B0(n548), .B1(n3742), .C0(n4379), 
        .C1(n3730), .Y(n1691) );
  AOI22X1TS U3160 ( .A0(n4279), .A1(n3712), .B0(n4108), .B1(n3689), .Y(n1688)
         );
  AOI222XLTS U3161 ( .A0(n4487), .A1(n3749), .B0(n659), .B1(n3742), .C0(n4376), 
        .C1(n3730), .Y(n1689) );
  AOI22X1TS U3162 ( .A0(n4276), .A1(n3711), .B0(n4105), .B1(n3690), .Y(n1686)
         );
  AOI222XLTS U3163 ( .A0(n4483), .A1(n3749), .B0(n506), .B1(n3740), .C0(n4373), 
        .C1(n3731), .Y(n1687) );
  AOI22X1TS U3164 ( .A0(n4273), .A1(n3713), .B0(n4102), .B1(n3690), .Y(n1684)
         );
  AOI222XLTS U3165 ( .A0(n4479), .A1(n3749), .B0(n663), .B1(n3740), .C0(n4370), 
        .C1(n3732), .Y(n1685) );
  AOI22X1TS U3166 ( .A0(n4270), .A1(n3712), .B0(n4099), .B1(n3690), .Y(n1682)
         );
  AOI222XLTS U3167 ( .A0(n4475), .A1(n3749), .B0(n672), .B1(n3743), .C0(n4367), 
        .C1(n3727), .Y(n1683) );
  AOI22X1TS U3168 ( .A0(n4267), .A1(n3700), .B0(n4096), .B1(n3690), .Y(n1680)
         );
  AOI222XLTS U3169 ( .A0(n4471), .A1(n3748), .B0(n508), .B1(n3741), .C0(n4364), 
        .C1(n3725), .Y(n1681) );
  AOI22X1TS U3170 ( .A0(n4264), .A1(n3700), .B0(n4093), .B1(n3691), .Y(n1678)
         );
  AOI222XLTS U3171 ( .A0(n4467), .A1(n3748), .B0(n674), .B1(n3738), .C0(n4361), 
        .C1(n3732), .Y(n1679) );
  AOI22X1TS U3172 ( .A0(n4005), .A1(n3710), .B0(n4066), .B1(n3682), .Y(n1822)
         );
  AOI222XLTS U3173 ( .A0(n4232), .A1(n3754), .B0(n38), .B1(n3733), .C0(n3964), 
        .C1(n3725), .Y(n1823) );
  AOI22X1TS U3174 ( .A0(n4354), .A1(n3557), .B0(n4183), .B1(n3835), .Y(n1609)
         );
  AOI222XLTS U3175 ( .A0(n4580), .A1(n3609), .B0(n509), .B1(n3585), .C0(n4459), 
        .C1(n3578), .Y(n1610) );
  AOI22X1TS U3176 ( .A0(n4309), .A1(n3553), .B0(n4138), .B1(n3831), .Y(n1579)
         );
  AOI222XLTS U3177 ( .A0(n4523), .A1(n3604), .B0(n531), .B1(n3597), .C0(n4406), 
        .C1(n3584), .Y(n1580) );
  AOI22X1TS U3178 ( .A0(n4306), .A1(n3553), .B0(n4135), .B1(n3831), .Y(n1577)
         );
  AOI222XLTS U3179 ( .A0(n4520), .A1(n3604), .B0(n533), .B1(n3587), .C0(n4403), 
        .C1(n3575), .Y(n1578) );
  AOI22X1TS U3180 ( .A0(n4294), .A1(n3552), .B0(n4123), .B1(n3838), .Y(n1569)
         );
  AOI222XLTS U3181 ( .A0(n4505), .A1(n3603), .B0(n541), .B1(n3589), .C0(n4391), 
        .C1(n3574), .Y(n1570) );
  AOI22X1TS U3182 ( .A0(n4264), .A1(n3551), .B0(n4093), .B1(n3828), .Y(n1549)
         );
  AOI222XLTS U3183 ( .A0(n4467), .A1(n3600), .B0(n673), .B1(n3590), .C0(n4361), 
        .C1(n3572), .Y(n1550) );
  AOI22X1TS U3184 ( .A0(n4008), .A1(n3558), .B0(n4069), .B1(n3836), .Y(n1877)
         );
  AOI222XLTS U3185 ( .A0(n4235), .A1(n3608), .B0(n3591), .B1(n45), .C0(n3967), 
        .C1(n3571), .Y(n1878) );
  AOI22X1TS U3186 ( .A0(n4351), .A1(n3557), .B0(n4180), .B1(n3835), .Y(n1607)
         );
  AOI222XLTS U3187 ( .A0(n4577), .A1(n3611), .B0(n511), .B1(n3597), .C0(n4456), 
        .C1(n3580), .Y(n1608) );
  AOI22X1TS U3188 ( .A0(n4348), .A1(n3556), .B0(n4177), .B1(n3834), .Y(n1605)
         );
  AOI222XLTS U3189 ( .A0(n4573), .A1(n3609), .B0(n513), .B1(n3585), .C0(n4452), 
        .C1(n1134), .Y(n1606) );
  AOI22X1TS U3190 ( .A0(n4345), .A1(n3556), .B0(n4174), .B1(n3834), .Y(n1603)
         );
  AOI222XLTS U3191 ( .A0(n4569), .A1(n3609), .B0(n495), .B1(n3597), .C0(n4449), 
        .C1(n3579), .Y(n1604) );
  AOI22X1TS U3192 ( .A0(n4342), .A1(n3556), .B0(n4171), .B1(n3834), .Y(n1601)
         );
  AOI222XLTS U3193 ( .A0(n4565), .A1(n3612), .B0(n497), .B1(n3594), .C0(n4445), 
        .C1(n3576), .Y(n1602) );
  AOI22X1TS U3194 ( .A0(n4339), .A1(n3556), .B0(n4168), .B1(n3834), .Y(n1599)
         );
  AOI222XLTS U3195 ( .A0(n4561), .A1(n3613), .B0(n515), .B1(n3586), .C0(n4441), 
        .C1(n3576), .Y(n1600) );
  AOI22X1TS U3196 ( .A0(n4336), .A1(n3555), .B0(n4165), .B1(n3833), .Y(n1597)
         );
  AOI222XLTS U3197 ( .A0(n4558), .A1(n3610), .B0(n517), .B1(n3586), .C0(n4438), 
        .C1(n3576), .Y(n1598) );
  AOI22X1TS U3198 ( .A0(n4333), .A1(n3555), .B0(n4162), .B1(n3833), .Y(n1595)
         );
  AOI222XLTS U3199 ( .A0(n4553), .A1(n3610), .B0(n519), .B1(n3585), .C0(n4434), 
        .C1(n3576), .Y(n1596) );
  AOI22X1TS U3200 ( .A0(n4330), .A1(n3555), .B0(n4159), .B1(n3833), .Y(n1593)
         );
  AOI222XLTS U3201 ( .A0(n4550), .A1(n3609), .B0(n499), .B1(n3587), .C0(n4430), 
        .C1(n3583), .Y(n1594) );
  AOI22X1TS U3202 ( .A0(n4327), .A1(n3555), .B0(n4156), .B1(n3833), .Y(n1591)
         );
  AOI222XLTS U3203 ( .A0(n4546), .A1(n3610), .B0(n521), .B1(n3587), .C0(n4426), 
        .C1(n3583), .Y(n1592) );
  AOI22X1TS U3204 ( .A0(n4324), .A1(n3554), .B0(n4153), .B1(n3832), .Y(n1589)
         );
  AOI222XLTS U3205 ( .A0(n4542), .A1(n3605), .B0(n523), .B1(n3585), .C0(n4423), 
        .C1(n3579), .Y(n1590) );
  AOI22X1TS U3206 ( .A0(n4321), .A1(n3554), .B0(n4150), .B1(n3832), .Y(n1587)
         );
  AOI222XLTS U3207 ( .A0(n4538), .A1(n3605), .B0(n501), .B1(n3587), .C0(n4418), 
        .C1(n3581), .Y(n1588) );
  AOI22X1TS U3208 ( .A0(n4318), .A1(n3554), .B0(n4147), .B1(n3832), .Y(n1585)
         );
  AOI222XLTS U3209 ( .A0(n4534), .A1(n3605), .B0(n525), .B1(n3588), .C0(n4415), 
        .C1(n3584), .Y(n1586) );
  AOI22X1TS U3210 ( .A0(n4315), .A1(n3553), .B0(n4144), .B1(n3832), .Y(n1583)
         );
  AOI222XLTS U3211 ( .A0(n4531), .A1(n3604), .B0(n527), .B1(n3586), .C0(n4412), 
        .C1(n3581), .Y(n1584) );
  AOI22X1TS U3212 ( .A0(n4312), .A1(n3553), .B0(n4141), .B1(n3831), .Y(n1581)
         );
  AOI222XLTS U3213 ( .A0(n4526), .A1(n3604), .B0(n529), .B1(n3588), .C0(n4409), 
        .C1(n3580), .Y(n1582) );
  AOI22X1TS U3214 ( .A0(n4303), .A1(n3552), .B0(n4132), .B1(n3831), .Y(n1575)
         );
  AOI222XLTS U3215 ( .A0(n4515), .A1(n3603), .B0(n535), .B1(n3586), .C0(n4400), 
        .C1(n3575), .Y(n1576) );
  AOI22X1TS U3216 ( .A0(n4300), .A1(n3552), .B0(n4129), .B1(n3839), .Y(n1573)
         );
  AOI222XLTS U3217 ( .A0(n4512), .A1(n3603), .B0(n537), .B1(n3595), .C0(n4397), 
        .C1(n3575), .Y(n1574) );
  AOI22X1TS U3218 ( .A0(n4297), .A1(n3552), .B0(n4126), .B1(n3837), .Y(n1571)
         );
  AOI222XLTS U3219 ( .A0(n4508), .A1(n3603), .B0(n539), .B1(n3588), .C0(n4394), 
        .C1(n3574), .Y(n1572) );
  AOI22X1TS U3220 ( .A0(n4291), .A1(n3563), .B0(n4120), .B1(n3837), .Y(n1567)
         );
  AOI222XLTS U3221 ( .A0(n4502), .A1(n3602), .B0(n543), .B1(n3589), .C0(n4388), 
        .C1(n3574), .Y(n1568) );
  AOI22X1TS U3222 ( .A0(n4288), .A1(n3554), .B0(n4117), .B1(n3830), .Y(n1565)
         );
  AOI222XLTS U3223 ( .A0(n4497), .A1(n3605), .B0(n503), .B1(n3594), .C0(n4385), 
        .C1(n3574), .Y(n1566) );
  AOI22X1TS U3224 ( .A0(n4285), .A1(n3565), .B0(n4114), .B1(n3830), .Y(n1563)
         );
  AOI222XLTS U3225 ( .A0(n4494), .A1(n3602), .B0(n545), .B1(n3589), .C0(n4382), 
        .C1(n3573), .Y(n1564) );
  AOI22X1TS U3226 ( .A0(n4282), .A1(n3561), .B0(n4111), .B1(n3830), .Y(n1561)
         );
  AOI222XLTS U3227 ( .A0(n4490), .A1(n3602), .B0(n547), .B1(n3598), .C0(n4379), 
        .C1(n3573), .Y(n1562) );
  AOI22X1TS U3228 ( .A0(n4279), .A1(n1135), .B0(n4108), .B1(n3830), .Y(n1559)
         );
  AOI222XLTS U3229 ( .A0(n4487), .A1(n3602), .B0(n549), .B1(n3596), .C0(n4376), 
        .C1(n3575), .Y(n1560) );
  AOI22X1TS U3230 ( .A0(n4276), .A1(n3564), .B0(n4105), .B1(n3829), .Y(n1557)
         );
  AOI222XLTS U3231 ( .A0(n4483), .A1(n3601), .B0(n505), .B1(n3590), .C0(n4373), 
        .C1(n3573), .Y(n1558) );
  AOI22X1TS U3232 ( .A0(n4273), .A1(n3565), .B0(n4102), .B1(n3829), .Y(n1555)
         );
  AOI222XLTS U3233 ( .A0(n4479), .A1(n3601), .B0(n661), .B1(n3590), .C0(n4370), 
        .C1(n3573), .Y(n1556) );
  AOI22X1TS U3234 ( .A0(n4270), .A1(n3566), .B0(n4099), .B1(n3829), .Y(n1553)
         );
  AOI222XLTS U3235 ( .A0(n4475), .A1(n3601), .B0(n666), .B1(n3589), .C0(n4367), 
        .C1(n3572), .Y(n1554) );
  AOI22X1TS U3236 ( .A0(n4267), .A1(n3562), .B0(n4096), .B1(n3829), .Y(n1551)
         );
  AOI222XLTS U3237 ( .A0(n4471), .A1(n3601), .B0(n507), .B1(n3590), .C0(n4364), 
        .C1(n3572), .Y(n1552) );
  AOI22X1TS U3238 ( .A0(n4261), .A1(n3551), .B0(n4090), .B1(n3828), .Y(n1547)
         );
  AOI222XLTS U3239 ( .A0(n4463), .A1(n3600), .B0(n676), .B1(n3588), .C0(n4358), 
        .C1(n3572), .Y(n1548) );
  AOI22X1TS U3240 ( .A0(n4489), .A1(n3666), .B0(n4111), .B1(n3869), .Y(n1626)
         );
  AOI222XLTS U3241 ( .A0(n4378), .A1(n3855), .B0(n547), .B1(n3655), .C0(n4283), 
        .C1(n3641), .Y(n1627) );
  AOI22X1TS U3242 ( .A0(n4493), .A1(n3667), .B0(n4114), .B1(n3869), .Y(n1628)
         );
  AOI222XLTS U3243 ( .A0(n4381), .A1(n3856), .B0(n545), .B1(n3655), .C0(n4286), 
        .C1(n3641), .Y(n1629) );
  AOI22X1TS U3244 ( .A0(n4504), .A1(n3667), .B0(n4123), .B1(n3870), .Y(n1634)
         );
  AOI222XLTS U3245 ( .A0(n4390), .A1(n3856), .B0(n541), .B1(n3654), .C0(n4295), 
        .C1(n1118), .Y(n1635) );
  AOI22X1TS U3246 ( .A0(n4507), .A1(n3680), .B0(n4126), .B1(n3870), .Y(n1636)
         );
  AOI222XLTS U3247 ( .A0(n4393), .A1(n3857), .B0(n539), .B1(n3654), .C0(n4298), 
        .C1(n3647), .Y(n1637) );
  AOI22X1TS U3248 ( .A0(n4511), .A1(n3680), .B0(n4129), .B1(n3877), .Y(n1638)
         );
  AOI222XLTS U3249 ( .A0(n4396), .A1(n3857), .B0(n537), .B1(n3653), .C0(n4301), 
        .C1(n1118), .Y(n1639) );
  AOI22X1TS U3250 ( .A0(n4519), .A1(n3677), .B0(n4135), .B1(n3868), .Y(n1642)
         );
  AOI222XLTS U3251 ( .A0(n4402), .A1(n3857), .B0(n533), .B1(n3654), .C0(n4307), 
        .C1(n3645), .Y(n1643) );
  AOI22X1TS U3252 ( .A0(n4522), .A1(n3668), .B0(n4138), .B1(n3879), .Y(n1644)
         );
  AOI222XLTS U3253 ( .A0(n4405), .A1(n3858), .B0(n531), .B1(n3653), .C0(n4310), 
        .C1(n3648), .Y(n1645) );
  AOI22X1TS U3254 ( .A0(n4525), .A1(n3668), .B0(n4141), .B1(n3878), .Y(n1646)
         );
  AOI222XLTS U3255 ( .A0(n4408), .A1(n3858), .B0(n529), .B1(n3652), .C0(n4313), 
        .C1(n3648), .Y(n1647) );
  AOI22X1TS U3256 ( .A0(n4533), .A1(n3668), .B0(n4147), .B1(n3868), .Y(n1650)
         );
  AOI222XLTS U3257 ( .A0(n4414), .A1(n3858), .B0(n525), .B1(n3652), .C0(n4319), 
        .C1(n3642), .Y(n1651) );
  AOI22X1TS U3258 ( .A0(n4537), .A1(n3669), .B0(n4150), .B1(n3877), .Y(n1652)
         );
  AOI22X1TS U3259 ( .A0(n4541), .A1(n3669), .B0(n4153), .B1(n3878), .Y(n1654)
         );
  AOI22X1TS U3260 ( .A0(n4544), .A1(n3669), .B0(n4156), .B1(n3867), .Y(n1656)
         );
  AOI22X1TS U3261 ( .A0(n4549), .A1(n3669), .B0(n4159), .B1(n3876), .Y(n1658)
         );
  AOI22X1TS U3262 ( .A0(n4552), .A1(n3670), .B0(n4162), .B1(n3876), .Y(n1660)
         );
  AOI22X1TS U3263 ( .A0(n4556), .A1(n3670), .B0(n4165), .B1(n3867), .Y(n1662)
         );
  AOI22X1TS U3264 ( .A0(n4560), .A1(n3670), .B0(n4168), .B1(n3868), .Y(n1664)
         );
  AOI22X1TS U3265 ( .A0(n4564), .A1(n3670), .B0(n4171), .B1(n3868), .Y(n1666)
         );
  AOI22X1TS U3266 ( .A0(n4571), .A1(n3671), .B0(n4177), .B1(n3875), .Y(n1670)
         );
  AOI22X1TS U3267 ( .A0(n4579), .A1(n3671), .B0(n4183), .B1(n3879), .Y(n1674)
         );
  AOI22X1TS U3268 ( .A0(n4443), .A1(n3294), .B0(n4171), .B1(n3845), .Y(n1345)
         );
  AOI222XLTS U3269 ( .A0(n4564), .A1(n3338), .B0(n497), .B1(n3320), .C0(n4343), 
        .C1(n3316), .Y(n1346) );
  AOI22X1TS U3270 ( .A0(n4425), .A1(n3293), .B0(n4156), .B1(n3844), .Y(n1335)
         );
  AOI222XLTS U3271 ( .A0(n4544), .A1(n3337), .B0(n521), .B1(n3323), .C0(n4328), 
        .C1(n3317), .Y(n1336) );
  AOI22X1TS U3272 ( .A0(n4417), .A1(n3292), .B0(n4150), .B1(n3843), .Y(n1331)
         );
  AOI222XLTS U3273 ( .A0(n4537), .A1(n3336), .B0(n501), .B1(n3323), .C0(n4322), 
        .C1(n3318), .Y(n1332) );
  AOI22X1TS U3274 ( .A0(n4414), .A1(n3292), .B0(n4147), .B1(n3843), .Y(n1329)
         );
  AOI22X1TS U3275 ( .A0(n4387), .A1(n3289), .B0(n4120), .B1(n3848), .Y(n1311)
         );
  AOI22X1TS U3276 ( .A0(n4381), .A1(n3289), .B0(n4114), .B1(n3853), .Y(n1307)
         );
  AOI22X1TS U3277 ( .A0(n4372), .A1(n3288), .B0(n4105), .B1(n3841), .Y(n1301)
         );
  AOI22X1TS U3278 ( .A0(n4363), .A1(n3288), .B0(n4096), .B1(n3841), .Y(n1295)
         );
  AOI22X1TS U3279 ( .A0(n4499), .A1(n3667), .B0(n4120), .B1(n3869), .Y(n1632)
         );
  AOI222XLTS U3280 ( .A0(n4387), .A1(n3856), .B0(n543), .B1(n3657), .C0(n4292), 
        .C1(n3641), .Y(n1633) );
  AOI22X1TS U3281 ( .A0(n4486), .A1(n3666), .B0(n4108), .B1(n3871), .Y(n1624)
         );
  AOI222XLTS U3282 ( .A0(n4375), .A1(n3855), .B0(n549), .B1(n3656), .C0(n4280), 
        .C1(n3647), .Y(n1625) );
  AOI22X1TS U3283 ( .A0(n3966), .A1(n3296), .B0(n4069), .B1(n3847), .Y(n1969)
         );
  AOI22X1TS U3284 ( .A0(n3960), .A1(n3296), .B0(n4063), .B1(n3847), .Y(n1965)
         );
  AOI222XLTS U3285 ( .A0(n4230), .A1(n3340), .B0(n3328), .B1(n34), .C0(n4003), 
        .C1(n3312), .Y(n1966) );
  AOI22X1TS U3286 ( .A0(n3957), .A1(n3296), .B0(n4060), .B1(n3847), .Y(n1963)
         );
  AOI222XLTS U3287 ( .A0(n4227), .A1(n3340), .B0(n3328), .B1(n29), .C0(n4000), 
        .C1(n3312), .Y(n1964) );
  AOI22X1TS U3288 ( .A0(n3954), .A1(n3295), .B0(n4057), .B1(n3846), .Y(n1961)
         );
  AOI222XLTS U3289 ( .A0(n4224), .A1(n3339), .B0(n3328), .B1(n24), .C0(n3997), 
        .C1(n3312), .Y(n1962) );
  AOI22X1TS U3290 ( .A0(n3951), .A1(n3295), .B0(n4054), .B1(n3846), .Y(n1959)
         );
  AOI222XLTS U3291 ( .A0(n4221), .A1(n3339), .B0(n3332), .B1(n19), .C0(n3994), 
        .C1(n3312), .Y(n1960) );
  AOI22X1TS U3292 ( .A0(n4458), .A1(n3295), .B0(n4183), .B1(n3846), .Y(n1353)
         );
  AOI222XLTS U3293 ( .A0(n4579), .A1(n3339), .B0(n509), .B1(n3321), .C0(n4355), 
        .C1(n3314), .Y(n1354) );
  AOI22X1TS U3294 ( .A0(n4454), .A1(n3295), .B0(n4180), .B1(n3846), .Y(n1351)
         );
  AOI222XLTS U3295 ( .A0(n4576), .A1(n3339), .B0(n511), .B1(n3320), .C0(n4352), 
        .C1(n3313), .Y(n1352) );
  AOI22X1TS U3296 ( .A0(n4451), .A1(n3294), .B0(n4177), .B1(n3845), .Y(n1349)
         );
  AOI222XLTS U3297 ( .A0(n4571), .A1(n3338), .B0(n513), .B1(n3321), .C0(n4349), 
        .C1(n3319), .Y(n1350) );
  AOI22X1TS U3298 ( .A0(n4448), .A1(n3294), .B0(n4174), .B1(n3845), .Y(n1347)
         );
  AOI222XLTS U3299 ( .A0(n4567), .A1(n3338), .B0(n495), .B1(n3320), .C0(n4346), 
        .C1(n3315), .Y(n1348) );
  AOI22X1TS U3300 ( .A0(n4440), .A1(n3294), .B0(n4168), .B1(n3845), .Y(n1343)
         );
  AOI222XLTS U3301 ( .A0(n4560), .A1(n3338), .B0(n515), .B1(n3322), .C0(n4340), 
        .C1(n3313), .Y(n1344) );
  AOI22X1TS U3302 ( .A0(n4436), .A1(n3293), .B0(n4165), .B1(n3844), .Y(n1341)
         );
  AOI222XLTS U3303 ( .A0(n4556), .A1(n3337), .B0(n517), .B1(n3322), .C0(n4337), 
        .C1(n3313), .Y(n1342) );
  AOI22X1TS U3304 ( .A0(n4432), .A1(n3293), .B0(n4162), .B1(n3844), .Y(n1339)
         );
  AOI222XLTS U3305 ( .A0(n4552), .A1(n3337), .B0(n519), .B1(n3321), .C0(n4334), 
        .C1(n3313), .Y(n1340) );
  AOI22X1TS U3306 ( .A0(n4429), .A1(n3293), .B0(n4159), .B1(n3844), .Y(n1337)
         );
  AOI222XLTS U3307 ( .A0(n4549), .A1(n3337), .B0(n499), .B1(n3323), .C0(n4331), 
        .C1(n3317), .Y(n1338) );
  AOI22X1TS U3308 ( .A0(n4422), .A1(n3292), .B0(n4153), .B1(n3843), .Y(n1333)
         );
  AOI222XLTS U3309 ( .A0(n4541), .A1(n3336), .B0(n523), .B1(n3321), .C0(n4325), 
        .C1(n3319), .Y(n1334) );
  AOI22X1TS U3310 ( .A0(n4411), .A1(n3291), .B0(n4144), .B1(n3843), .Y(n1327)
         );
  AOI22X1TS U3311 ( .A0(n4408), .A1(n3291), .B0(n4141), .B1(n3842), .Y(n1325)
         );
  AOI22X1TS U3312 ( .A0(n4405), .A1(n3291), .B0(n4138), .B1(n3842), .Y(n1323)
         );
  AOI22X1TS U3313 ( .A0(n4402), .A1(n3291), .B0(n4135), .B1(n3842), .Y(n1321)
         );
  AOI22X1TS U3314 ( .A0(n4399), .A1(n3290), .B0(n4132), .B1(n3842), .Y(n1319)
         );
  AOI22X1TS U3315 ( .A0(n4396), .A1(n3290), .B0(n4129), .B1(n3849), .Y(n1317)
         );
  AOI22X1TS U3316 ( .A0(n4393), .A1(n3290), .B0(n4126), .B1(n3850), .Y(n1315)
         );
  AOI22X1TS U3317 ( .A0(n4390), .A1(n3290), .B0(n4123), .B1(n3848), .Y(n1313)
         );
  AOI22X1TS U3318 ( .A0(n4384), .A1(n3292), .B0(n4117), .B1(n3849), .Y(n1309)
         );
  AOI22X1TS U3319 ( .A0(n4378), .A1(n3289), .B0(n4111), .B1(n3851), .Y(n1305)
         );
  AOI22X1TS U3320 ( .A0(n4375), .A1(n3289), .B0(n4108), .B1(n3852), .Y(n1303)
         );
  AOI22X1TS U3321 ( .A0(n4369), .A1(n3288), .B0(n4102), .B1(n3841), .Y(n1299)
         );
  AOI22X1TS U3322 ( .A0(n4366), .A1(n3288), .B0(n4099), .B1(n3841), .Y(n1297)
         );
  AOI22X1TS U3323 ( .A0(n4360), .A1(n3287), .B0(n4093), .B1(n1754), .Y(n1293)
         );
  AOI22X1TS U3324 ( .A0(n4576), .A1(n3671), .B0(n4180), .B1(n3867), .Y(n1672)
         );
  AOI22X1TS U3325 ( .A0(n4567), .A1(n3671), .B0(n4174), .B1(n3879), .Y(n1668)
         );
  AOI22X1TS U3326 ( .A0(n4514), .A1(n3679), .B0(n4132), .B1(n3869), .Y(n1640)
         );
  AOI222XLTS U3327 ( .A0(n4399), .A1(n3857), .B0(n535), .B1(n3653), .C0(n4304), 
        .C1(n3646), .Y(n1641) );
  AOI22X1TS U3328 ( .A0(n4496), .A1(n3667), .B0(n4117), .B1(n3870), .Y(n1630)
         );
  AOI222XLTS U3329 ( .A0(n4384), .A1(n3856), .B0(n503), .B1(n3655), .C0(n4289), 
        .C1(n3641), .Y(n1631) );
  AOI22X1TS U3330 ( .A0(n4481), .A1(n3666), .B0(n4105), .B1(n3871), .Y(n1622)
         );
  AOI222XLTS U3331 ( .A0(n4372), .A1(n3855), .B0(n505), .B1(n3655), .C0(n4277), 
        .C1(n3640), .Y(n1623) );
  AOI22X1TS U3332 ( .A0(n4474), .A1(n3665), .B0(n4099), .B1(n3871), .Y(n1618)
         );
  AOI222XLTS U3333 ( .A0(n4366), .A1(n3854), .B0(n666), .B1(n3657), .C0(n4271), 
        .C1(n3640), .Y(n1619) );
  AOI22X1TS U3334 ( .A0(n4470), .A1(n3665), .B0(n4096), .B1(n3871), .Y(n1616)
         );
  AOI222XLTS U3335 ( .A0(n4363), .A1(n3854), .B0(n507), .B1(n3656), .C0(n4268), 
        .C1(n3639), .Y(n1617) );
  AOI22X1TS U3336 ( .A0(n4357), .A1(n3287), .B0(n4090), .B1(n3851), .Y(n1291)
         );
  AOI22X1TS U3337 ( .A0(n4529), .A1(n3668), .B0(n4144), .B1(n669), .Y(n1648)
         );
  AOI222XLTS U3338 ( .A0(n4411), .A1(n3858), .B0(n527), .B1(n3653), .C0(n4316), 
        .C1(n3642), .Y(n1649) );
  AOI22X1TS U3339 ( .A0(n4478), .A1(n3666), .B0(n4102), .B1(n3870), .Y(n1620)
         );
  AOI222XLTS U3340 ( .A0(n4369), .A1(n3855), .B0(n661), .B1(n3656), .C0(n4274), 
        .C1(n3640), .Y(n1621) );
  AOI22X1TS U3341 ( .A0(n4002), .A1(n3558), .B0(n4063), .B1(n3836), .Y(n1873)
         );
  AOI222XLTS U3342 ( .A0(n4229), .A1(n3615), .B0(n3593), .B1(n35), .C0(n3961), 
        .C1(n3577), .Y(n1874) );
  AOI22X1TS U3343 ( .A0(n3999), .A1(n3558), .B0(n4060), .B1(n3836), .Y(n1871)
         );
  AOI222XLTS U3344 ( .A0(n4226), .A1(n1132), .B0(n3593), .B1(n30), .C0(n3958), 
        .C1(n3577), .Y(n1872) );
  AOI22X1TS U3345 ( .A0(n3996), .A1(n3557), .B0(n4057), .B1(n3835), .Y(n1869)
         );
  AOI222XLTS U3346 ( .A0(n4223), .A1(n3612), .B0(n3593), .B1(n25), .C0(n3955), 
        .C1(n3577), .Y(n1870) );
  AOI22X1TS U3347 ( .A0(n3993), .A1(n3557), .B0(n4054), .B1(n3835), .Y(n1867)
         );
  AOI222XLTS U3348 ( .A0(n4220), .A1(n3613), .B0(n3592), .B1(n20), .C0(n3952), 
        .C1(n3577), .Y(n1868) );
  AOI22X1TS U3349 ( .A0(n4220), .A1(n3209), .B0(n3994), .B1(n3947), .Y(n1981)
         );
  AOI222XLTS U3350 ( .A0(n3951), .A1(n3266), .B0(n4055), .B1(n3237), .C0(n3222), .C1(n19), .Y(n1982) );
  AOI22X1TS U3351 ( .A0(n4567), .A1(n3208), .B0(n4345), .B1(n3943), .Y(n1283)
         );
  AOI222XLTS U3352 ( .A0(n4449), .A1(n3261), .B0(n4175), .B1(n3238), .C0(n496), 
        .C1(n3223), .Y(n1284) );
  AOI22X1TS U3353 ( .A0(n4564), .A1(n3208), .B0(n4342), .B1(n3943), .Y(n1281)
         );
  AOI222XLTS U3354 ( .A0(n4445), .A1(n3265), .B0(n4172), .B1(n3238), .C0(n498), 
        .C1(n3224), .Y(n1282) );
  AOI22X1TS U3355 ( .A0(n4549), .A1(n3207), .B0(n4330), .B1(n3942), .Y(n1273)
         );
  AOI222XLTS U3356 ( .A0(n4430), .A1(n3260), .B0(n4160), .B1(n3239), .C0(n500), 
        .C1(n3224), .Y(n1274) );
  AOI22X1TS U3357 ( .A0(n4537), .A1(n3206), .B0(n4321), .B1(n3941), .Y(n1267)
         );
  AOI222XLTS U3358 ( .A0(n4418), .A1(n3262), .B0(n4151), .B1(n3247), .C0(n502), 
        .C1(n3226), .Y(n1268) );
  AOI22X1TS U3359 ( .A0(n4496), .A1(n3206), .B0(n4288), .B1(n3939), .Y(n1245)
         );
  AOI222XLTS U3360 ( .A0(n4385), .A1(n3263), .B0(n4118), .B1(n3241), .C0(n504), 
        .C1(n3230), .Y(n1246) );
  AOI22X1TS U3361 ( .A0(n4481), .A1(n3217), .B0(n4276), .B1(n660), .Y(n1237)
         );
  AOI222XLTS U3362 ( .A0(n4373), .A1(n3253), .B0(n4106), .B1(n3242), .C0(n506), 
        .C1(n3227), .Y(n1238) );
  AOI22X1TS U3363 ( .A0(n4470), .A1(n3214), .B0(n4267), .B1(n3950), .Y(n1231)
         );
  AOI222XLTS U3364 ( .A0(n4364), .A1(n3253), .B0(n4097), .B1(n3243), .C0(n508), 
        .C1(n3231), .Y(n1232) );
  AOI22X1TS U3365 ( .A0(n4466), .A1(n3204), .B0(n4264), .B1(n3948), .Y(n1229)
         );
  AOI222XLTS U3366 ( .A0(n4361), .A1(n3252), .B0(n4094), .B1(n3243), .C0(n674), 
        .C1(n3231), .Y(n1230) );
  AOI22X1TS U3367 ( .A0(n4462), .A1(n3204), .B0(n4261), .B1(n3945), .Y(n1227)
         );
  AOI222XLTS U3368 ( .A0(n4358), .A1(n3252), .B0(n4091), .B1(n3243), .C0(n677), 
        .C1(n3225), .Y(n1228) );
  AOI22X1TS U3369 ( .A0(n3204), .A1(n4603), .B0(n3946), .B1(n4051), .Y(n1225)
         );
  AOI222XLTS U3370 ( .A0(n3252), .A1(n4200), .B0(n3243), .B1(n4088), .C0(n3221), .C1(n45), .Y(n1226) );
  AOI22X1TS U3371 ( .A0(n3203), .A1(n4594), .B0(n3938), .B1(n4045), .Y(n1221)
         );
  AOI222XLTS U3372 ( .A0(n3251), .A1(n4194), .B0(n3250), .B1(n4082), .C0(n3220), .C1(n35), .Y(n1222) );
  AOI22X1TS U3373 ( .A0(n3203), .A1(n4598), .B0(n3947), .B1(n4048), .Y(n1223)
         );
  AOI222XLTS U3374 ( .A0(n3251), .A1(n4197), .B0(n3248), .B1(n4085), .C0(n3221), .C1(n40), .Y(n1224) );
  AOI22X1TS U3375 ( .A0(n3203), .A1(n4591), .B0(n3938), .B1(n4042), .Y(n1219)
         );
  AOI222XLTS U3376 ( .A0(n3251), .A1(n4191), .B0(n3246), .B1(n4079), .C0(n3220), .C1(n30), .Y(n1220) );
  AOI22X1TS U3377 ( .A0(n3203), .A1(n4586), .B0(n3938), .B1(n4039), .Y(n1217)
         );
  AOI222XLTS U3378 ( .A0(n3251), .A1(n4188), .B0(n3248), .B1(n4076), .C0(n3220), .C1(n25), .Y(n1218) );
  AOI22X1TS U3379 ( .A0(n3204), .A1(n4583), .B0(n3938), .B1(n4036), .Y(n1211)
         );
  AOI222XLTS U3380 ( .A0(n3252), .A1(n4185), .B0(n3250), .B1(n4073), .C0(n3221), .C1(n20), .Y(n1212) );
  AOI22X1TS U3381 ( .A0(n4458), .A1(n3458), .B0(n4579), .B1(n3444), .Y(n1481)
         );
  AOI222XLTS U3382 ( .A0(n509), .A1(n3802), .B0(n4184), .B1(n3812), .C0(n6255), 
        .C1(n192), .Y(n1482) );
  AOI22X1TS U3383 ( .A0(n4454), .A1(n3458), .B0(n4576), .B1(n1166), .Y(n1479)
         );
  AOI222XLTS U3384 ( .A0(n511), .A1(n3806), .B0(n4181), .B1(n3812), .C0(n6256), 
        .C1(n135), .Y(n1480) );
  AOI22X1TS U3385 ( .A0(n4451), .A1(n3457), .B0(n4571), .B1(n3445), .Y(n1477)
         );
  AOI222XLTS U3386 ( .A0(n513), .A1(n3807), .B0(n4178), .B1(n3813), .C0(n6257), 
        .C1(n190), .Y(n1478) );
  AOI22X1TS U3387 ( .A0(n4448), .A1(n3457), .B0(n4567), .B1(n3445), .Y(n1475)
         );
  AOI222XLTS U3388 ( .A0(n495), .A1(n3803), .B0(n4175), .B1(n3813), .C0(n6258), 
        .C1(n3809), .Y(n1476) );
  AOI22X1TS U3389 ( .A0(n4443), .A1(n3457), .B0(n4564), .B1(n3448), .Y(n1473)
         );
  AOI222XLTS U3390 ( .A0(n497), .A1(n3805), .B0(n4172), .B1(n3813), .C0(n6259), 
        .C1(n192), .Y(n1474) );
  AOI22X1TS U3391 ( .A0(n4440), .A1(n3457), .B0(n4560), .B1(n3447), .Y(n1471)
         );
  AOI222XLTS U3392 ( .A0(n515), .A1(n3799), .B0(n4169), .B1(n3813), .C0(n6260), 
        .C1(n134), .Y(n1472) );
  AOI22X1TS U3393 ( .A0(n4432), .A1(n3456), .B0(n4552), .B1(n3446), .Y(n1467)
         );
  AOI222XLTS U3394 ( .A0(n519), .A1(n3804), .B0(n4163), .B1(n3814), .C0(n6261), 
        .C1(n191), .Y(n1468) );
  AOI22X1TS U3395 ( .A0(n4425), .A1(n3456), .B0(n4544), .B1(n3446), .Y(n1463)
         );
  AOI222XLTS U3396 ( .A0(n521), .A1(n3803), .B0(n4157), .B1(n3814), .C0(n6262), 
        .C1(n192), .Y(n1464) );
  AOI22X1TS U3397 ( .A0(n4422), .A1(n3455), .B0(n4541), .B1(n3446), .Y(n1461)
         );
  AOI222XLTS U3398 ( .A0(n523), .A1(n3797), .B0(n4154), .B1(n3815), .C0(n6263), 
        .C1(n135), .Y(n1462) );
  AOI22X1TS U3399 ( .A0(n4414), .A1(n3455), .B0(n4533), .B1(n3446), .Y(n1457)
         );
  AOI222XLTS U3400 ( .A0(n525), .A1(n3797), .B0(n4148), .B1(n3815), .C0(n6264), 
        .C1(n191), .Y(n1458) );
  AOI22X1TS U3401 ( .A0(n4408), .A1(n3465), .B0(n4525), .B1(n3440), .Y(n1453)
         );
  AOI222XLTS U3402 ( .A0(n529), .A1(n3797), .B0(n4142), .B1(n3816), .C0(n6265), 
        .C1(n681), .Y(n1454) );
  AOI22X1TS U3403 ( .A0(n4405), .A1(n3463), .B0(n4522), .B1(n3440), .Y(n1451)
         );
  AOI222XLTS U3404 ( .A0(n531), .A1(n3798), .B0(n4139), .B1(n3816), .C0(n6266), 
        .C1(n3811), .Y(n1452) );
  AOI22X1TS U3405 ( .A0(n4399), .A1(n3465), .B0(n4514), .B1(n3439), .Y(n1447)
         );
  AOI222XLTS U3406 ( .A0(n535), .A1(n3798), .B0(n4133), .B1(n3816), .C0(n6267), 
        .C1(n188), .Y(n1448) );
  AOI22X1TS U3407 ( .A0(n4393), .A1(n3465), .B0(n4507), .B1(n3439), .Y(n1443)
         );
  AOI222XLTS U3408 ( .A0(n539), .A1(n3799), .B0(n4127), .B1(n3817), .C0(n6268), 
        .C1(n136), .Y(n1444) );
  AOI22X1TS U3409 ( .A0(n4390), .A1(n3467), .B0(n4504), .B1(n3439), .Y(n1441)
         );
  AOI222XLTS U3410 ( .A0(n541), .A1(n3799), .B0(n4124), .B1(n3817), .C0(n6269), 
        .C1(n186), .Y(n1442) );
  AOI22X1TS U3411 ( .A0(n4387), .A1(n3454), .B0(n4499), .B1(n3438), .Y(n1439)
         );
  AOI222XLTS U3412 ( .A0(n543), .A1(n3802), .B0(n4121), .B1(n3817), .C0(n6270), 
        .C1(n191), .Y(n1440) );
  AOI22X1TS U3413 ( .A0(n4384), .A1(n3455), .B0(n4496), .B1(n3445), .Y(n1437)
         );
  AOI222XLTS U3414 ( .A0(n503), .A1(n3800), .B0(n4118), .B1(n3818), .C0(n6271), 
        .C1(n136), .Y(n1438) );
  AOI22X1TS U3415 ( .A0(n4381), .A1(n3454), .B0(n4493), .B1(n3438), .Y(n1435)
         );
  AOI222XLTS U3416 ( .A0(n545), .A1(n3800), .B0(n4115), .B1(n3818), .C0(n6272), 
        .C1(n192), .Y(n1436) );
  AOI22X1TS U3417 ( .A0(n4375), .A1(n3454), .B0(n4486), .B1(n3438), .Y(n1431)
         );
  AOI222XLTS U3418 ( .A0(n549), .A1(n3801), .B0(n4109), .B1(n3818), .C0(n6273), 
        .C1(n187), .Y(n1432) );
  AOI22X1TS U3419 ( .A0(n4366), .A1(n3464), .B0(n4474), .B1(n3437), .Y(n1425)
         );
  AOI222XLTS U3420 ( .A0(n666), .A1(n3802), .B0(n4100), .B1(n3819), .C0(n6274), 
        .C1(n3809), .Y(n1426) );
  AOI22X1TS U3421 ( .A0(n4360), .A1(n3453), .B0(n4466), .B1(n3436), .Y(n1421)
         );
  AOI222XLTS U3422 ( .A0(n673), .A1(n3801), .B0(n4094), .B1(n3820), .C0(n6275), 
        .C1(n187), .Y(n1422) );
  AOI22X1TS U3423 ( .A0(n4357), .A1(n3453), .B0(n4462), .B1(n3436), .Y(n1419)
         );
  AOI222XLTS U3424 ( .A0(n676), .A1(n3802), .B0(n4091), .B1(n3820), .C0(n6276), 
        .C1(n135), .Y(n1420) );
  AOI22X1TS U3425 ( .A0(n4436), .A1(n3456), .B0(n4556), .B1(n3447), .Y(n1469)
         );
  AOI222XLTS U3426 ( .A0(n517), .A1(n3804), .B0(n4166), .B1(n3814), .C0(n6292), 
        .C1(n186), .Y(n1470) );
  AOI22X1TS U3427 ( .A0(n4429), .A1(n3456), .B0(n4549), .B1(n3449), .Y(n1465)
         );
  AOI222XLTS U3428 ( .A0(n499), .A1(n3805), .B0(n4160), .B1(n3814), .C0(n6293), 
        .C1(n190), .Y(n1466) );
  AOI22X1TS U3429 ( .A0(n4417), .A1(n3455), .B0(n4537), .B1(n3448), .Y(n1459)
         );
  AOI222XLTS U3430 ( .A0(n501), .A1(n3797), .B0(n4151), .B1(n3815), .C0(n6294), 
        .C1(n188), .Y(n1460) );
  AOI22X1TS U3431 ( .A0(n4411), .A1(n3468), .B0(n4529), .B1(n3440), .Y(n1455)
         );
  AOI222XLTS U3432 ( .A0(n527), .A1(n3798), .B0(n4145), .B1(n3815), .C0(n6295), 
        .C1(n134), .Y(n1456) );
  AOI22X1TS U3433 ( .A0(n4402), .A1(n1165), .B0(n4519), .B1(n3440), .Y(n1449)
         );
  AOI222XLTS U3434 ( .A0(n533), .A1(n3799), .B0(n4136), .B1(n3816), .C0(n6296), 
        .C1(n191), .Y(n1450) );
  AOI22X1TS U3435 ( .A0(n4396), .A1(n3462), .B0(n4511), .B1(n3439), .Y(n1445)
         );
  AOI222XLTS U3436 ( .A0(n537), .A1(n3798), .B0(n4130), .B1(n3817), .C0(n6297), 
        .C1(n187), .Y(n1446) );
  AOI22X1TS U3437 ( .A0(n4372), .A1(n3466), .B0(n4481), .B1(n3437), .Y(n1429)
         );
  AOI222XLTS U3438 ( .A0(n505), .A1(n3800), .B0(n4106), .B1(n3819), .C0(n6298), 
        .C1(n3811), .Y(n1430) );
  AOI22X1TS U3439 ( .A0(n4369), .A1(n3464), .B0(n4478), .B1(n3437), .Y(n1427)
         );
  AOI222XLTS U3440 ( .A0(n661), .A1(n3801), .B0(n4103), .B1(n3819), .C0(n6299), 
        .C1(n3809), .Y(n1428) );
  AOI22X1TS U3441 ( .A0(n4363), .A1(n3465), .B0(n4470), .B1(n3437), .Y(n1423)
         );
  AOI222XLTS U3442 ( .A0(n507), .A1(n3801), .B0(n4097), .B1(n3819), .C0(n6300), 
        .C1(n188), .Y(n1424) );
  AOI22X1TS U3443 ( .A0(n4378), .A1(n3454), .B0(n4489), .B1(n3438), .Y(n1433)
         );
  AOI222XLTS U3444 ( .A0(n547), .A1(n3800), .B0(n4112), .B1(n3818), .C0(n6313), 
        .C1(n134), .Y(n1434) );
  AOI22X1TS U3445 ( .A0(n3510), .A1(n39), .B0(n3963), .B1(n3493), .Y(n1897) );
  AOI222XLTS U3446 ( .A0(n2993), .A1(n3890), .B0(n4233), .B1(n1149), .C0(n4067), .C1(n3902), .Y(n1898) );
  AOI22X1TS U3447 ( .A0(n3388), .A1(n27), .B0(n3999), .B1(n3375), .Y(n1940) );
  AOI222XLTS U3448 ( .A0(n58), .A1(n3917), .B0(n4225), .B1(n3410), .C0(n4061), 
        .C1(n3933), .Y(n1941) );
  AOI22X1TS U3449 ( .A0(n512), .A1(n3389), .B0(n4351), .B1(n3374), .Y(n1415)
         );
  AOI222XLTS U3450 ( .A0(n59), .A1(n3916), .B0(n4574), .B1(n3407), .C0(n4181), 
        .C1(n3931), .Y(n1416) );
  AOI22X1TS U3451 ( .A0(n514), .A1(n3389), .B0(n4348), .B1(n3373), .Y(n1413)
         );
  AOI222XLTS U3452 ( .A0(n60), .A1(n3916), .B0(n4570), .B1(n3411), .C0(n4178), 
        .C1(n3932), .Y(n1414) );
  AOI22X1TS U3453 ( .A0(n496), .A1(n3389), .B0(n4345), .B1(n3373), .Y(n1411)
         );
  AOI222XLTS U3454 ( .A0(n61), .A1(n3916), .B0(n4566), .B1(n3411), .C0(n4175), 
        .C1(n3935), .Y(n1412) );
  AOI22X1TS U3455 ( .A0(n516), .A1(n3391), .B0(n4339), .B1(n3373), .Y(n1407)
         );
  AOI222XLTS U3456 ( .A0(n62), .A1(n3915), .B0(n4559), .B1(n3411), .C0(n4169), 
        .C1(n3935), .Y(n1408) );
  AOI22X1TS U3457 ( .A0(n518), .A1(n3389), .B0(n4336), .B1(n3372), .Y(n1405)
         );
  AOI222XLTS U3458 ( .A0(n63), .A1(n3915), .B0(n4555), .B1(n3409), .C0(n4166), 
        .C1(n3932), .Y(n1406) );
  AOI22X1TS U3459 ( .A0(n500), .A1(n3390), .B0(n4330), .B1(n3372), .Y(n1401)
         );
  AOI222XLTS U3460 ( .A0(n64), .A1(n3914), .B0(n4547), .B1(n3416), .C0(n4160), 
        .C1(n3933), .Y(n1402) );
  AOI22X1TS U3461 ( .A0(n524), .A1(n3396), .B0(n4324), .B1(n3371), .Y(n1397)
         );
  AOI222XLTS U3462 ( .A0(n65), .A1(n3914), .B0(n4540), .B1(n3406), .C0(n4154), 
        .C1(n3930), .Y(n1398) );
  AOI22X1TS U3463 ( .A0(n502), .A1(n3393), .B0(n4321), .B1(n3371), .Y(n1395)
         );
  AOI222XLTS U3464 ( .A0(n66), .A1(n3914), .B0(n4535), .B1(n3406), .C0(n4151), 
        .C1(n3930), .Y(n1396) );
  AOI22X1TS U3465 ( .A0(n526), .A1(n3394), .B0(n4318), .B1(n3371), .Y(n1393)
         );
  AOI222XLTS U3466 ( .A0(n67), .A1(n3913), .B0(n4532), .B1(n3406), .C0(n4148), 
        .C1(n3930), .Y(n1394) );
  AOI22X1TS U3467 ( .A0(n528), .A1(n3394), .B0(n4315), .B1(n3381), .Y(n1391)
         );
  AOI222XLTS U3468 ( .A0(n68), .A1(n3913), .B0(n4528), .B1(n3413), .C0(n4145), 
        .C1(n3930), .Y(n1392) );
  AOI22X1TS U3469 ( .A0(n530), .A1(n3394), .B0(n4312), .B1(n3381), .Y(n1389)
         );
  AOI222XLTS U3470 ( .A0(n69), .A1(n3913), .B0(n4524), .B1(n3413), .C0(n4142), 
        .C1(n3929), .Y(n1390) );
  AOI22X1TS U3471 ( .A0(n534), .A1(n3391), .B0(n4306), .B1(n3383), .Y(n1385)
         );
  AOI222XLTS U3472 ( .A0(n70), .A1(n3912), .B0(n4517), .B1(n3409), .C0(n4136), 
        .C1(n3929), .Y(n1386) );
  AOI22X1TS U3473 ( .A0(n536), .A1(n3399), .B0(n4303), .B1(n3381), .Y(n1383)
         );
  AOI222XLTS U3474 ( .A0(n71), .A1(n3912), .B0(n4513), .B1(n3405), .C0(n4133), 
        .C1(n3929), .Y(n1384) );
  AOI22X1TS U3475 ( .A0(n538), .A1(n3393), .B0(n4300), .B1(n3379), .Y(n1381)
         );
  AOI222XLTS U3476 ( .A0(n72), .A1(n3912), .B0(n4510), .B1(n3405), .C0(n4130), 
        .C1(n3928), .Y(n1382) );
  AOI22X1TS U3477 ( .A0(n540), .A1(n3391), .B0(n4297), .B1(n3385), .Y(n1379)
         );
  AOI222XLTS U3478 ( .A0(n73), .A1(n3911), .B0(n4506), .B1(n3405), .C0(n4127), 
        .C1(n3928), .Y(n1380) );
  AOI22X1TS U3479 ( .A0(n542), .A1(n3391), .B0(n4294), .B1(n1182), .Y(n1377)
         );
  AOI222XLTS U3480 ( .A0(n74), .A1(n3911), .B0(n4503), .B1(n3405), .C0(n4124), 
        .C1(n3928), .Y(n1378) );
  AOI22X1TS U3481 ( .A0(n504), .A1(n3392), .B0(n4288), .B1(n3371), .Y(n1373)
         );
  AOI222XLTS U3482 ( .A0(n75), .A1(n3911), .B0(n4495), .B1(n3404), .C0(n4118), 
        .C1(n3927), .Y(n1374) );
  AOI22X1TS U3483 ( .A0(n546), .A1(n3392), .B0(n4285), .B1(n3382), .Y(n1371)
         );
  AOI222XLTS U3484 ( .A0(n76), .A1(n3910), .B0(n4492), .B1(n3404), .C0(n4115), 
        .C1(n3927), .Y(n1372) );
  AOI22X1TS U3485 ( .A0(n548), .A1(n3392), .B0(n4282), .B1(n3382), .Y(n1369)
         );
  AOI222XLTS U3486 ( .A0(n77), .A1(n3910), .B0(n4488), .B1(n3404), .C0(n4112), 
        .C1(n3927), .Y(n1370) );
  AOI22X1TS U3487 ( .A0(n506), .A1(n3392), .B0(n4276), .B1(n3380), .Y(n1365)
         );
  AOI222XLTS U3488 ( .A0(n78), .A1(n3910), .B0(n4480), .B1(n3403), .C0(n4106), 
        .C1(n3926), .Y(n1366) );
  AOI22X1TS U3489 ( .A0(n663), .A1(n3395), .B0(n4273), .B1(n3382), .Y(n1363)
         );
  AOI222XLTS U3490 ( .A0(n79), .A1(n3909), .B0(n4477), .B1(n3403), .C0(n4103), 
        .C1(n3926), .Y(n1364) );
  AOI22X1TS U3491 ( .A0(n672), .A1(n3397), .B0(n4270), .B1(n3380), .Y(n1361)
         );
  AOI222XLTS U3492 ( .A0(n80), .A1(n3909), .B0(n4472), .B1(n3403), .C0(n4100), 
        .C1(n3926), .Y(n1362) );
  AOI22X1TS U3493 ( .A0(n3386), .A1(n44), .B0(n4008), .B1(n3375), .Y(n1946) );
  AOI222XLTS U3494 ( .A0(n81), .A1(n3921), .B0(n4234), .B1(n3402), .C0(n4070), 
        .C1(n3932), .Y(n1947) );
  AOI22X1TS U3495 ( .A0(n3388), .A1(n37), .B0(n4005), .B1(n3375), .Y(n1944) );
  AOI222XLTS U3496 ( .A0(n82), .A1(n3918), .B0(n4231), .B1(n3410), .C0(n4067), 
        .C1(n3936), .Y(n1945) );
  AOI22X1TS U3497 ( .A0(n3388), .A1(n32), .B0(n4002), .B1(n3375), .Y(n1942) );
  AOI222XLTS U3498 ( .A0(n83), .A1(n3917), .B0(n4228), .B1(n3410), .C0(n4064), 
        .C1(n662), .Y(n1943) );
  AOI22X1TS U3499 ( .A0(n3387), .A1(n23), .B0(n3996), .B1(n3374), .Y(n1938) );
  AOI222XLTS U3500 ( .A0(n84), .A1(n3917), .B0(n4222), .B1(n3407), .C0(n4058), 
        .C1(n3931), .Y(n1939) );
  AOI22X1TS U3501 ( .A0(n3388), .A1(n18), .B0(n3993), .B1(n3374), .Y(n1936) );
  AOI222XLTS U3502 ( .A0(n85), .A1(n3917), .B0(n4219), .B1(n3407), .C0(n4055), 
        .C1(n3931), .Y(n1937) );
  AOI22X1TS U3503 ( .A0(n498), .A1(n3390), .B0(n4342), .B1(n3373), .Y(n1409)
         );
  AOI222XLTS U3504 ( .A0(n86), .A1(n3915), .B0(n4562), .B1(n3415), .C0(n4172), 
        .C1(n3934), .Y(n1410) );
  AOI22X1TS U3505 ( .A0(n544), .A1(n3397), .B0(n4291), .B1(n3381), .Y(n1375)
         );
  AOI222XLTS U3506 ( .A0(n87), .A1(n3911), .B0(n4498), .B1(n3404), .C0(n4121), 
        .C1(n3928), .Y(n1376) );
  AOI22X1TS U3507 ( .A0(n674), .A1(n3398), .B0(n4264), .B1(n3370), .Y(n1357)
         );
  AOI222XLTS U3508 ( .A0(n88), .A1(n3909), .B0(n4465), .B1(n3402), .C0(n4094), 
        .C1(n3925), .Y(n1358) );
  AOI22X1TS U3509 ( .A0(n510), .A1(n3397), .B0(n4354), .B1(n3374), .Y(n1417)
         );
  AOI222XLTS U3510 ( .A0(n89), .A1(n3916), .B0(n4578), .B1(n3407), .C0(n4184), 
        .C1(n3931), .Y(n1418) );
  AOI22X1TS U3511 ( .A0(n520), .A1(n3390), .B0(n4333), .B1(n3372), .Y(n1403)
         );
  AOI222XLTS U3512 ( .A0(n90), .A1(n3915), .B0(n4551), .B1(n3416), .C0(n4163), 
        .C1(n3937), .Y(n1404) );
  AOI22X1TS U3513 ( .A0(n522), .A1(n3390), .B0(n4327), .B1(n3372), .Y(n1399)
         );
  AOI222XLTS U3514 ( .A0(n91), .A1(n3914), .B0(n4543), .B1(n3411), .C0(n4157), 
        .C1(n3934), .Y(n1400) );
  AOI22X1TS U3515 ( .A0(n532), .A1(n3394), .B0(n4309), .B1(n3378), .Y(n1387)
         );
  AOI222XLTS U3516 ( .A0(n92), .A1(n3913), .B0(n4521), .B1(n3416), .C0(n4139), 
        .C1(n3929), .Y(n1388) );
  AOI22X1TS U3517 ( .A0(n659), .A1(n3399), .B0(n4279), .B1(n3383), .Y(n1367)
         );
  AOI222XLTS U3518 ( .A0(n93), .A1(n3910), .B0(n4484), .B1(n3406), .C0(n4109), 
        .C1(n3927), .Y(n1368) );
  AOI22X1TS U3519 ( .A0(n508), .A1(n3396), .B0(n4267), .B1(n3382), .Y(n1359)
         );
  AOI222XLTS U3520 ( .A0(n94), .A1(n3909), .B0(n4468), .B1(n3403), .C0(n4097), 
        .C1(n3926), .Y(n1360) );
  AOI22X1TS U3521 ( .A0(n677), .A1(n3395), .B0(n4261), .B1(n3370), .Y(n1355)
         );
  AOI222XLTS U3522 ( .A0(n95), .A1(n3920), .B0(n4461), .B1(n3402), .C0(n4091), 
        .C1(n3925), .Y(n1356) );
  AOI22X1TS U3523 ( .A0(n3514), .A1(n42), .B0(n3966), .B1(n3493), .Y(n1899) );
  AOI222XLTS U3524 ( .A0(n2991), .A1(n3890), .B0(n4236), .B1(n3519), .C0(n4070), .C1(n3903), .Y(n1900) );
  AOI22X1TS U3525 ( .A0(n3511), .A1(n34), .B0(n3960), .B1(n3493), .Y(n1895) );
  AOI222XLTS U3526 ( .A0(n2995), .A1(n3891), .B0(n4230), .B1(n3528), .C0(n4064), .C1(n3902), .Y(n1896) );
  AOI22X1TS U3527 ( .A0(n3512), .A1(n28), .B0(n3957), .B1(n3493), .Y(n1893) );
  AOI222XLTS U3528 ( .A0(n2997), .A1(n668), .B0(n4227), .B1(n1149), .C0(n4061), 
        .C1(n3902), .Y(n1894) );
  AOI22X1TS U3529 ( .A0(n3503), .A1(n24), .B0(n3954), .B1(n3500), .Y(n1891) );
  AOI222XLTS U3530 ( .A0(n2999), .A1(n668), .B0(n4224), .B1(n3529), .C0(n4058), 
        .C1(n3904), .Y(n1892) );
  AOI22X1TS U3531 ( .A0(n3514), .A1(n19), .B0(n3951), .B1(n3500), .Y(n1889) );
  AOI222XLTS U3532 ( .A0(n3001), .A1(n3892), .B0(n4221), .B1(n3530), .C0(n4055), .C1(n3902), .Y(n1890) );
  AOI22X1TS U3533 ( .A0(n511), .A1(n3513), .B0(n4454), .B1(n3498), .Y(n1543)
         );
  AOI222XLTS U3534 ( .A0(n2929), .A1(n3887), .B0(n4577), .B1(n3531), .C0(n4181), .C1(n3905), .Y(n1544) );
  AOI22X1TS U3535 ( .A0(n495), .A1(n3513), .B0(n4448), .B1(n3496), .Y(n1539)
         );
  AOI222XLTS U3536 ( .A0(n2933), .A1(n3887), .B0(n4569), .B1(n3526), .C0(n4175), .C1(n3906), .Y(n1540) );
  AOI22X1TS U3537 ( .A0(n497), .A1(n3513), .B0(n4443), .B1(n3502), .Y(n1537)
         );
  AOI222XLTS U3538 ( .A0(n2935), .A1(n3886), .B0(n4565), .B1(n3526), .C0(n4172), .C1(n3906), .Y(n1538) );
  AOI22X1TS U3539 ( .A0(n515), .A1(n3506), .B0(n4440), .B1(n3498), .Y(n1535)
         );
  AOI222XLTS U3540 ( .A0(n2937), .A1(n3886), .B0(n4561), .B1(n3526), .C0(n4169), .C1(n3906), .Y(n1536) );
  AOI22X1TS U3541 ( .A0(n517), .A1(n3514), .B0(n4436), .B1(n1151), .Y(n1533)
         );
  AOI222XLTS U3542 ( .A0(n2939), .A1(n3886), .B0(n4558), .B1(n3525), .C0(n4166), .C1(n3901), .Y(n1534) );
  AOI22X1TS U3543 ( .A0(n519), .A1(n3510), .B0(n4432), .B1(n3497), .Y(n1531)
         );
  AOI222XLTS U3544 ( .A0(n2941), .A1(n3886), .B0(n4553), .B1(n3525), .C0(n4163), .C1(n3901), .Y(n1532) );
  AOI22X1TS U3545 ( .A0(n499), .A1(n3511), .B0(n4429), .B1(n3497), .Y(n1529)
         );
  AOI222XLTS U3546 ( .A0(n2943), .A1(n3885), .B0(n4550), .B1(n3525), .C0(n4160), .C1(n3901), .Y(n1530) );
  AOI22X1TS U3547 ( .A0(n527), .A1(n3505), .B0(n4411), .B1(n3491), .Y(n1519)
         );
  AOI222XLTS U3548 ( .A0(n2953), .A1(n3884), .B0(n4531), .B1(n3523), .C0(n4145), .C1(n3900), .Y(n1520) );
  AOI22X1TS U3549 ( .A0(n537), .A1(n3505), .B0(n4396), .B1(n3490), .Y(n1509)
         );
  AOI222XLTS U3550 ( .A0(n2963), .A1(n3883), .B0(n4512), .B1(n3522), .C0(n4130), .C1(n3898), .Y(n1510) );
  AOI22X1TS U3551 ( .A0(n503), .A1(n3507), .B0(n4384), .B1(n3492), .Y(n1501)
         );
  AOI222XLTS U3552 ( .A0(n2971), .A1(n3882), .B0(n4497), .B1(n3521), .C0(n4118), .C1(n3897), .Y(n1502) );
  AOI22X1TS U3553 ( .A0(n547), .A1(n3507), .B0(n4378), .B1(n3489), .Y(n1497)
         );
  AOI222XLTS U3554 ( .A0(n2975), .A1(n3881), .B0(n4490), .B1(n3521), .C0(n4112), .C1(n3897), .Y(n1498) );
  AOI22X1TS U3555 ( .A0(n505), .A1(n3507), .B0(n4372), .B1(n3488), .Y(n1493)
         );
  AOI222XLTS U3556 ( .A0(n2979), .A1(n3881), .B0(n4483), .B1(n3520), .C0(n4106), .C1(n3896), .Y(n1494) );
  AOI22X1TS U3557 ( .A0(n661), .A1(n3508), .B0(n4369), .B1(n3488), .Y(n1491)
         );
  AOI222XLTS U3558 ( .A0(n2981), .A1(n3880), .B0(n4479), .B1(n3520), .C0(n4103), .C1(n3896), .Y(n1492) );
  AOI22X1TS U3559 ( .A0(n507), .A1(n3508), .B0(n4363), .B1(n3488), .Y(n1487)
         );
  AOI222XLTS U3560 ( .A0(n2985), .A1(n3880), .B0(n4471), .B1(n3520), .C0(n4097), .C1(n3896), .Y(n1488) );
  AOI22X1TS U3561 ( .A0(n509), .A1(n3509), .B0(n4458), .B1(n3499), .Y(n1545)
         );
  AOI222XLTS U3562 ( .A0(n2927), .A1(n3887), .B0(n4580), .B1(n3531), .C0(n4184), .C1(n3907), .Y(n1546) );
  AOI22X1TS U3563 ( .A0(n513), .A1(n3513), .B0(n4451), .B1(n3499), .Y(n1541)
         );
  AOI222XLTS U3564 ( .A0(n2931), .A1(n3887), .B0(n4573), .B1(n3526), .C0(n4178), .C1(n3908), .Y(n1542) );
  AOI22X1TS U3565 ( .A0(n521), .A1(n3512), .B0(n4425), .B1(n3502), .Y(n1527)
         );
  AOI222XLTS U3566 ( .A0(n2945), .A1(n3885), .B0(n4546), .B1(n3525), .C0(n4157), .C1(n3901), .Y(n1528) );
  AOI22X1TS U3567 ( .A0(n523), .A1(n3504), .B0(n4422), .B1(n3492), .Y(n1525)
         );
  AOI222XLTS U3568 ( .A0(n2947), .A1(n3885), .B0(n4542), .B1(n3524), .C0(n4154), .C1(n3900), .Y(n1526) );
  AOI22X1TS U3569 ( .A0(n501), .A1(n3504), .B0(n4417), .B1(n3492), .Y(n1523)
         );
  AOI222XLTS U3570 ( .A0(n2949), .A1(n3885), .B0(n4538), .B1(n3524), .C0(n4151), .C1(n3900), .Y(n1524) );
  AOI22X1TS U3571 ( .A0(n525), .A1(n3504), .B0(n4414), .B1(n3492), .Y(n1521)
         );
  AOI222XLTS U3572 ( .A0(n2951), .A1(n3884), .B0(n4534), .B1(n3524), .C0(n4148), .C1(n3900), .Y(n1522) );
  AOI22X1TS U3573 ( .A0(n531), .A1(n3505), .B0(n4405), .B1(n3491), .Y(n1515)
         );
  AOI222XLTS U3574 ( .A0(n2957), .A1(n3884), .B0(n4523), .B1(n3523), .C0(n4139), .C1(n3899), .Y(n1516) );
  AOI22X1TS U3575 ( .A0(n539), .A1(n3506), .B0(n4393), .B1(n3490), .Y(n1507)
         );
  AOI222XLTS U3576 ( .A0(n2965), .A1(n3882), .B0(n4508), .B1(n3522), .C0(n4127), .C1(n3898), .Y(n1508) );
  AOI22X1TS U3577 ( .A0(n541), .A1(n3506), .B0(n4390), .B1(n3490), .Y(n1505)
         );
  AOI222XLTS U3578 ( .A0(n2967), .A1(n3882), .B0(n4505), .B1(n3522), .C0(n4124), .C1(n3898), .Y(n1506) );
  AOI22X1TS U3579 ( .A0(n543), .A1(n3509), .B0(n4387), .B1(n3489), .Y(n1503)
         );
  AOI222XLTS U3580 ( .A0(n2969), .A1(n3882), .B0(n4502), .B1(n3521), .C0(n4121), .C1(n3898), .Y(n1504) );
  AOI22X1TS U3581 ( .A0(n545), .A1(n3507), .B0(n4381), .B1(n3489), .Y(n1499)
         );
  AOI222XLTS U3582 ( .A0(n2973), .A1(n3881), .B0(n4494), .B1(n3521), .C0(n4115), .C1(n3897), .Y(n1500) );
  AOI22X1TS U3583 ( .A0(n549), .A1(n3508), .B0(n4375), .B1(n3489), .Y(n1495)
         );
  AOI222XLTS U3584 ( .A0(n2977), .A1(n3881), .B0(n4487), .B1(n3524), .C0(n4109), .C1(n3897), .Y(n1496) );
  AOI22X1TS U3585 ( .A0(n673), .A1(n3508), .B0(n4360), .B1(n3487), .Y(n1485)
         );
  AOI222XLTS U3586 ( .A0(n2987), .A1(n3880), .B0(n4467), .B1(n3519), .C0(n4094), .C1(n3895), .Y(n1486) );
  AOI22X1TS U3587 ( .A0(n676), .A1(n3509), .B0(n4357), .B1(n3487), .Y(n1483)
         );
  AOI222XLTS U3588 ( .A0(n2989), .A1(n3892), .B0(n4463), .B1(n3519), .C0(n4091), .C1(n3895), .Y(n1484) );
  AOI22X1TS U3589 ( .A0(n529), .A1(n3504), .B0(n4408), .B1(n3491), .Y(n1517)
         );
  AOI222XLTS U3590 ( .A0(n2955), .A1(n3884), .B0(n4526), .B1(n3523), .C0(n4142), .C1(n3899), .Y(n1518) );
  AOI22X1TS U3591 ( .A0(n533), .A1(n3506), .B0(n4402), .B1(n3491), .Y(n1513)
         );
  AOI222XLTS U3592 ( .A0(n2959), .A1(n3883), .B0(n4520), .B1(n3523), .C0(n4136), .C1(n3899), .Y(n1514) );
  AOI22X1TS U3593 ( .A0(n535), .A1(n3505), .B0(n4399), .B1(n3490), .Y(n1511)
         );
  AOI222XLTS U3594 ( .A0(n2961), .A1(n3883), .B0(n4515), .B1(n3522), .C0(n4133), .C1(n3899), .Y(n1512) );
  AOI22X1TS U3595 ( .A0(n666), .A1(n3509), .B0(n4366), .B1(n3488), .Y(n1489)
         );
  AOI222XLTS U3596 ( .A0(n2983), .A1(n3880), .B0(n4475), .B1(n3520), .C0(n4100), .C1(n3896), .Y(n1490) );
  AOI22X1TS U3597 ( .A0(n3963), .A1(n3296), .B0(n4066), .B1(n3847), .Y(n1967)
         );
  AOI22X1TS U3598 ( .A0(n4466), .A1(n3665), .B0(n4093), .B1(n3875), .Y(n1614)
         );
  AOI222XLTS U3599 ( .A0(n4360), .A1(n3854), .B0(n673), .B1(n3656), .C0(n4265), 
        .C1(n3639), .Y(n1615) );
  AOI22X1TS U3600 ( .A0(n4462), .A1(n3665), .B0(n4090), .B1(n3867), .Y(n1612)
         );
  AOI222XLTS U3601 ( .A0(n4357), .A1(n3854), .B0(n676), .B1(n3657), .C0(n4262), 
        .C1(n3640), .Y(n1613) );
  AOI22X1TS U3602 ( .A0(n4005), .A1(n3558), .B0(n4066), .B1(n3836), .Y(n1875)
         );
  AOI222XLTS U3603 ( .A0(n4232), .A1(n1132), .B0(n3593), .B1(n40), .C0(n3964), 
        .C1(n3584), .Y(n1876) );
  AO21X1TS U3604 ( .A0(n942), .A1(n2036), .B0(n2037), .Y(n2035) );
  OAI33XLTS U3605 ( .A0(n4829), .A1(n954), .A2(n2012), .B0(n2038), .B1(n4605), 
        .B2(n939), .Y(n2037) );
  NOR4XLTS U3606 ( .A(n2039), .B(n2040), .C(n2041), .D(n2042), .Y(n2038) );
  INVX2TS U3607 ( .A(n2036), .Y(n939) );
  NOR2BX1TS U3608 ( .AN(n2898), .B(n2378), .Y(n2895) );
  AOI21X1TS U3609 ( .A0(n4207), .A1(n695), .B0(n1797), .Y(n1796) );
  NAND3X1TS U3610 ( .A(n2386), .B(n2393), .C(n9), .Y(n2389) );
  AOI221X1TS U3611 ( .A0(n2919), .A1(n4456), .B0(n3063), .B1(n4179), .C0(n2369), .Y(n2365) );
  OAI22X1TS U3612 ( .A0(n4428), .A1(n3115), .B0(n866), .B1(n3781), .Y(n2369)
         );
  AOI221X1TS U3613 ( .A0(n2919), .A1(n4452), .B0(n3063), .B1(n4176), .C0(n2363), .Y(n2359) );
  OAI22X1TS U3614 ( .A0(n4437), .A1(n3115), .B0(n865), .B1(n3781), .Y(n2363)
         );
  AOI221X1TS U3615 ( .A0(n2919), .A1(n4449), .B0(n3063), .B1(n4173), .C0(n2357), .Y(n2353) );
  OAI22X1TS U3616 ( .A0(n4446), .A1(n3115), .B0(n864), .B1(n3781), .Y(n2357)
         );
  AOI221X1TS U3617 ( .A0(n2920), .A1(n4445), .B0(n3062), .B1(n4170), .C0(n2351), .Y(n2347) );
  OAI22X1TS U3618 ( .A0(n4455), .A1(n3115), .B0(n863), .B1(n3782), .Y(n2351)
         );
  AOI221X1TS U3619 ( .A0(n2920), .A1(n4441), .B0(n3062), .B1(n4167), .C0(n2345), .Y(n2341) );
  OAI22X1TS U3620 ( .A0(n4464), .A1(n3114), .B0(n862), .B1(n3782), .Y(n2345)
         );
  AOI221X1TS U3621 ( .A0(n2920), .A1(n4438), .B0(n3062), .B1(n4164), .C0(n2339), .Y(n2335) );
  OAI22X1TS U3622 ( .A0(n4473), .A1(n3114), .B0(n844), .B1(n3782), .Y(n2339)
         );
  AOI221X1TS U3623 ( .A0(n2920), .A1(n4434), .B0(n3062), .B1(n4161), .C0(n2333), .Y(n2329) );
  OAI22X1TS U3624 ( .A0(n4482), .A1(n3114), .B0(n861), .B1(n3782), .Y(n2333)
         );
  AOI221X1TS U3625 ( .A0(n3003), .A1(n4430), .B0(n3067), .B1(n4158), .C0(n2327), .Y(n2323) );
  OAI22X1TS U3626 ( .A0(n4491), .A1(n3114), .B0(n843), .B1(n3783), .Y(n2327)
         );
  AOI221X1TS U3627 ( .A0(n3003), .A1(n4426), .B0(n3064), .B1(n4155), .C0(n2321), .Y(n2317) );
  OAI22X1TS U3628 ( .A0(n4500), .A1(n3113), .B0(n860), .B1(n3783), .Y(n2321)
         );
  AOI221X1TS U3629 ( .A0(n3003), .A1(n4423), .B0(n3067), .B1(n4152), .C0(n2315), .Y(n2311) );
  OAI22X1TS U3630 ( .A0(n4509), .A1(n3113), .B0(n859), .B1(n3783), .Y(n2315)
         );
  AOI221X1TS U3631 ( .A0(n3003), .A1(n4418), .B0(n3068), .B1(n4149), .C0(n2309), .Y(n2305) );
  OAI22X1TS U3632 ( .A0(n4518), .A1(n3113), .B0(n842), .B1(n3783), .Y(n2309)
         );
  AOI221X1TS U3633 ( .A0(n3004), .A1(n4415), .B0(n3064), .B1(n4146), .C0(n2303), .Y(n2299) );
  OAI22X1TS U3634 ( .A0(n4527), .A1(n3113), .B0(n858), .B1(n3792), .Y(n2303)
         );
  AOI221X1TS U3635 ( .A0(n3004), .A1(n4412), .B0(n3070), .B1(n4143), .C0(n2297), .Y(n2293) );
  OAI22X1TS U3636 ( .A0(n4536), .A1(n3112), .B0(n841), .B1(n3793), .Y(n2297)
         );
  AOI221X1TS U3637 ( .A0(n3004), .A1(n4409), .B0(n3065), .B1(n4140), .C0(n2291), .Y(n2287) );
  OAI22X1TS U3638 ( .A0(n4545), .A1(n3112), .B0(n857), .B1(n3791), .Y(n2291)
         );
  AOI221X1TS U3639 ( .A0(n3004), .A1(n4406), .B0(n3070), .B1(n4137), .C0(n2285), .Y(n2281) );
  OAI22X1TS U3640 ( .A0(n4554), .A1(n3112), .B0(n856), .B1(n1093), .Y(n2285)
         );
  AOI221X1TS U3641 ( .A0(n3005), .A1(n4403), .B0(n3061), .B1(n4134), .C0(n2279), .Y(n2275) );
  OAI22X1TS U3642 ( .A0(n4563), .A1(n3112), .B0(n840), .B1(n3790), .Y(n2279)
         );
  AOI221X1TS U3643 ( .A0(n3005), .A1(n4400), .B0(n3061), .B1(n4131), .C0(n2273), .Y(n2269) );
  OAI22X1TS U3644 ( .A0(n4572), .A1(n3111), .B0(n855), .B1(n3792), .Y(n2273)
         );
  AOI221X1TS U3645 ( .A0(n3005), .A1(n4397), .B0(n3061), .B1(n4128), .C0(n2267), .Y(n2263) );
  OAI22X1TS U3646 ( .A0(n4581), .A1(n3111), .B0(n839), .B1(n3793), .Y(n2267)
         );
  AOI221X1TS U3647 ( .A0(n3005), .A1(n4394), .B0(n3061), .B1(n4125), .C0(n2261), .Y(n2257) );
  OAI22X1TS U3648 ( .A0(n4590), .A1(n3111), .B0(n854), .B1(n3791), .Y(n2261)
         );
  AOI221X1TS U3649 ( .A0(n3044), .A1(n4391), .B0(n3060), .B1(n4122), .C0(n2255), .Y(n2251) );
  OAI22X1TS U3650 ( .A0(n4599), .A1(n3111), .B0(n853), .B1(n3789), .Y(n2255)
         );
  AOI221X1TS U3651 ( .A0(n3044), .A1(n4388), .B0(n3060), .B1(n4119), .C0(n2249), .Y(n2245) );
  OAI22X1TS U3652 ( .A0(n4608), .A1(n3110), .B0(n852), .B1(n3790), .Y(n2249)
         );
  AOI221X1TS U3653 ( .A0(n3044), .A1(n4385), .B0(n3060), .B1(n4116), .C0(n2243), .Y(n2239) );
  OAI22X1TS U3654 ( .A0(n4617), .A1(n3110), .B0(n851), .B1(n3792), .Y(n2243)
         );
  AOI221X1TS U3655 ( .A0(n3044), .A1(n4382), .B0(n3060), .B1(n4113), .C0(n2237), .Y(n2233) );
  OAI22X1TS U3656 ( .A0(n4626), .A1(n3110), .B0(n850), .B1(n3789), .Y(n2237)
         );
  AOI221X1TS U3657 ( .A0(n3045), .A1(n4379), .B0(n3059), .B1(n4110), .C0(n2231), .Y(n2227) );
  OAI22X1TS U3658 ( .A0(n4635), .A1(n3109), .B0(n835), .B1(n3784), .Y(n2231)
         );
  AOI221X1TS U3659 ( .A0(n3045), .A1(n4376), .B0(n3059), .B1(n4107), .C0(n2225), .Y(n2221) );
  OAI22X1TS U3660 ( .A0(n4644), .A1(n3109), .B0(n849), .B1(n3784), .Y(n2225)
         );
  AOI221X1TS U3661 ( .A0(n3045), .A1(n4373), .B0(n3059), .B1(n4104), .C0(n2219), .Y(n2215) );
  OAI22X1TS U3662 ( .A0(n4653), .A1(n3109), .B0(n838), .B1(n3784), .Y(n2219)
         );
  AOI221X1TS U3663 ( .A0(n3045), .A1(n4370), .B0(n3059), .B1(n4101), .C0(n2213), .Y(n2209) );
  OAI22X1TS U3664 ( .A0(n4662), .A1(n3109), .B0(n837), .B1(n3784), .Y(n2213)
         );
  AOI221X1TS U3665 ( .A0(n3046), .A1(n4367), .B0(n3058), .B1(n4098), .C0(n2207), .Y(n2203) );
  OAI22X1TS U3666 ( .A0(n4671), .A1(n3108), .B0(n848), .B1(n3785), .Y(n2207)
         );
  AOI221X1TS U3667 ( .A0(n3046), .A1(n4364), .B0(n3058), .B1(n4095), .C0(n2201), .Y(n2197) );
  OAI22X1TS U3668 ( .A0(n4680), .A1(n3108), .B0(n836), .B1(n3785), .Y(n2201)
         );
  AOI221X1TS U3669 ( .A0(n3046), .A1(n4361), .B0(n3058), .B1(n4092), .C0(n2195), .Y(n2191) );
  OAI22X1TS U3670 ( .A0(n4689), .A1(n3108), .B0(n847), .B1(n3785), .Y(n2195)
         );
  AOI221X1TS U3671 ( .A0(n3046), .A1(n4358), .B0(n3058), .B1(n4089), .C0(n2189), .Y(n2185) );
  OAI22X1TS U3672 ( .A0(n4698), .A1(n3108), .B0(n846), .B1(n3785), .Y(n2189)
         );
  AOI221X1TS U3673 ( .A0(n3048), .A1(n3967), .B0(n3056), .B1(n4068), .C0(n2147), .Y(n2143) );
  OAI22X1TS U3674 ( .A0(n4711), .A1(n3107), .B0(n872), .B1(n3787), .Y(n2147)
         );
  AOI221X1TS U3675 ( .A0(n3048), .A1(n3964), .B0(n3056), .B1(n4065), .C0(n2141), .Y(n2137) );
  OAI22X1TS U3676 ( .A0(n4720), .A1(n3107), .B0(n871), .B1(n3787), .Y(n2141)
         );
  AOI221X1TS U3677 ( .A0(n3049), .A1(n3961), .B0(n3066), .B1(n4062), .C0(n2135), .Y(n2131) );
  OAI22X1TS U3678 ( .A0(n4729), .A1(n3110), .B0(n870), .B1(n3788), .Y(n2135)
         );
  AOI221X1TS U3679 ( .A0(n3049), .A1(n3958), .B0(n3066), .B1(n4059), .C0(n2129), .Y(n2125) );
  OAI22X1TS U3680 ( .A0(n4738), .A1(n3107), .B0(n845), .B1(n3788), .Y(n2129)
         );
  AOI221X1TS U3681 ( .A0(n3049), .A1(n3952), .B0(n3065), .B1(n4053), .C0(n2116), .Y(n2105) );
  OAI22X1TS U3682 ( .A0(n4756), .A1(n3107), .B0(n868), .B1(n3788), .Y(n2116)
         );
  OAI22X1TS U3683 ( .A0(n1081), .A1(n1083), .B0(n960), .B1(n1082), .Y(n2887)
         );
  CLKBUFX2TS U3684 ( .A(n5323), .Y(n989) );
  AOI22X1TS U3685 ( .A0(n1778), .A1(n1779), .B0(n3891), .B1(n647), .Y(n2567)
         );
  OAI33XLTS U3686 ( .A0(n4215), .A1(n99), .A2(n124), .B0(n138), .B1(n117), 
        .B2(n1784), .Y(n1781) );
  AOI222XLTS U3687 ( .A0(n4212), .A1(n1767), .B0(readIn_NORTH), .B1(n1768), 
        .C0(n4207), .C1(n697), .Y(n1766) );
  AOI221X1TS U3688 ( .A0(n2919), .A1(n4459), .B0(n3063), .B1(n4182), .C0(n2375), .Y(n2371) );
  OAI22X1TS U3689 ( .A0(n4419), .A1(n3106), .B0(n867), .B1(n3781), .Y(n2375)
         );
  AOI221X1TS U3690 ( .A0(n3047), .A1(n4201), .B0(n3057), .B1(n4086), .C0(n2183), .Y(n2179) );
  OAI22X1TS U3691 ( .A0(n3106), .A1(n4707), .B0(n877), .B1(n3786), .Y(n2183)
         );
  AOI221X1TS U3692 ( .A0(n3047), .A1(n4198), .B0(n3057), .B1(n4083), .C0(n2177), .Y(n2173) );
  OAI22X1TS U3693 ( .A0(n3106), .A1(n4708), .B0(n878), .B1(n3786), .Y(n2177)
         );
  AOI221X1TS U3694 ( .A0(n3047), .A1(n4192), .B0(n3057), .B1(n4077), .C0(n2165), .Y(n2161) );
  OAI22X1TS U3695 ( .A0(n3105), .A1(n4709), .B0(n875), .B1(n3786), .Y(n2165)
         );
  AOI221X1TS U3696 ( .A0(n3048), .A1(n4189), .B0(n3056), .B1(n4074), .C0(n2159), .Y(n2155) );
  OAI22X1TS U3697 ( .A0(n3105), .A1(n4710), .B0(n874), .B1(n3787), .Y(n2159)
         );
  AOI221X1TS U3698 ( .A0(n3049), .A1(n3955), .B0(n3068), .B1(n4056), .C0(n2123), .Y(n2119) );
  OAI22X1TS U3699 ( .A0(n4747), .A1(n3106), .B0(n869), .B1(n3788), .Y(n2123)
         );
  AOI221X1TS U3700 ( .A0(n3047), .A1(n4195), .B0(n3057), .B1(n4080), .C0(n2171), .Y(n2167) );
  OAI22X1TS U3701 ( .A0(n3105), .A1(n4834), .B0(n876), .B1(n3786), .Y(n2171)
         );
  AOI221X1TS U3702 ( .A0(n3048), .A1(n4186), .B0(n3056), .B1(n4071), .C0(n2153), .Y(n2149) );
  OAI22X1TS U3703 ( .A0(n3105), .A1(n4833), .B0(n873), .B1(n3787), .Y(n2153)
         );
  XOR2X1TS U3704 ( .A(n2392), .B(n9), .Y(n1080) );
  NAND2X1TS U3705 ( .A(n2393), .B(n2386), .Y(n2392) );
  NAND4X1TS U3706 ( .A(n2370), .B(n2371), .C(n2372), .D(n2373), .Y(n2397) );
  AOI221X1TS U3707 ( .A0(n2108), .A1(n3006), .B0(n2109), .B1(n89), .C0(n2374), 
        .Y(n2373) );
  AOI222XLTS U3708 ( .A0(n1046), .A1(n638), .B0(n1032), .B1(n2928), .C0(n1017), 
        .C1(n2927), .Y(n2372) );
  AOI222XLTS U3709 ( .A0(n3071), .A1(n4580), .B0(n3090), .B1(n4355), .C0(n1003), .C1(cacheDataOut[31]), .Y(n2370) );
  NAND4X1TS U3710 ( .A(n2364), .B(n2365), .C(n2366), .D(n2367), .Y(n2398) );
  AOI221X1TS U3711 ( .A0(n2108), .A1(n3007), .B0(n2109), .B1(n59), .C0(n2368), 
        .Y(n2367) );
  AOI222XLTS U3712 ( .A0(n1046), .A1(n637), .B0(n1032), .B1(n2930), .C0(n1017), 
        .C1(n2929), .Y(n2366) );
  AOI222XLTS U3713 ( .A0(n3071), .A1(n4577), .B0(n3099), .B1(n4352), .C0(n1003), .C1(cacheDataOut[30]), .Y(n2364) );
  NAND4X1TS U3714 ( .A(n2358), .B(n2359), .C(n2360), .D(n2361), .Y(n2399) );
  AOI221X1TS U3715 ( .A0(n2916), .A1(n3008), .B0(n1749), .B1(n60), .C0(n2362), 
        .Y(n2361) );
  AOI222XLTS U3716 ( .A0(n1047), .A1(n636), .B0(n1032), .B1(n2932), .C0(n1017), 
        .C1(n2931), .Y(n2360) );
  AOI222XLTS U3717 ( .A0(n3071), .A1(n4573), .B0(n3100), .B1(n4349), .C0(n1004), .C1(cacheDataOut[29]), .Y(n2358) );
  NAND4X1TS U3718 ( .A(n2352), .B(n2353), .C(n2354), .D(n2355), .Y(n2400) );
  AOI221X1TS U3719 ( .A0(n2915), .A1(n3009), .B0(n1611), .B1(n61), .C0(n2356), 
        .Y(n2355) );
  AOI222XLTS U3720 ( .A0(n2113), .A1(n49), .B0(n2114), .B1(n2934), .C0(n1016), 
        .C1(n2933), .Y(n2354) );
  AOI222XLTS U3721 ( .A0(n3071), .A1(n4569), .B0(n3099), .B1(n4346), .C0(n2117), .C1(cacheDataOut[28]), .Y(n2352) );
  NAND4X1TS U3722 ( .A(n2346), .B(n2347), .C(n2348), .D(n2349), .Y(n2401) );
  AOI221X1TS U3723 ( .A0(n1934), .A1(n3010), .B0(n1076), .B1(n86), .C0(n2350), 
        .Y(n2349) );
  AOI222XLTS U3724 ( .A0(n1034), .A1(n50), .B0(n1019), .B1(n2936), .C0(n1005), 
        .C1(n2935), .Y(n2348) );
  AOI222XLTS U3725 ( .A0(n3072), .A1(n4565), .B0(n3103), .B1(n4343), .C0(n991), 
        .C1(cacheDataOut[27]), .Y(n2346) );
  NAND4X1TS U3726 ( .A(n2340), .B(n2341), .C(n2342), .D(n2343), .Y(n2402) );
  AOI221X1TS U3727 ( .A0(n1934), .A1(n3011), .B0(n1076), .B1(n62), .C0(n2344), 
        .Y(n2343) );
  AOI222XLTS U3728 ( .A0(n1034), .A1(n635), .B0(n1019), .B1(n2938), .C0(n1005), 
        .C1(n2937), .Y(n2342) );
  AOI222XLTS U3729 ( .A0(n3072), .A1(n4561), .B0(n3097), .B1(n4340), .C0(n991), 
        .C1(cacheDataOut[26]), .Y(n2340) );
  NAND4X1TS U3730 ( .A(n2334), .B(n2335), .C(n2336), .D(n2337), .Y(n2403) );
  AOI221X1TS U3731 ( .A0(n1934), .A1(n3012), .B0(n1076), .B1(n63), .C0(n2338), 
        .Y(n2337) );
  AOI222XLTS U3732 ( .A0(n1034), .A1(n634), .B0(n1019), .B1(n2940), .C0(n1005), 
        .C1(n2939), .Y(n2336) );
  AOI222XLTS U3733 ( .A0(n3072), .A1(n4558), .B0(n3097), .B1(n4337), .C0(n991), 
        .C1(cacheDataOut[25]), .Y(n2334) );
  NAND4X1TS U3734 ( .A(n2328), .B(n2329), .C(n2330), .D(n2331), .Y(n2404) );
  AOI221X1TS U3735 ( .A0(n1934), .A1(n3013), .B0(n1076), .B1(n90), .C0(n2332), 
        .Y(n2331) );
  AOI222XLTS U3736 ( .A0(n1034), .A1(n633), .B0(n1019), .B1(n2942), .C0(n1005), 
        .C1(n2941), .Y(n2330) );
  AOI222XLTS U3737 ( .A0(n3072), .A1(n4553), .B0(n3097), .B1(n4334), .C0(n991), 
        .C1(cacheDataOut[24]), .Y(n2328) );
  NAND4X1TS U3738 ( .A(n2322), .B(n2323), .C(n2324), .D(n2325), .Y(n2405) );
  AOI221X1TS U3739 ( .A0(n1980), .A1(n3014), .B0(n1077), .B1(n64), .C0(n2326), 
        .Y(n2325) );
  AOI222XLTS U3740 ( .A0(n1045), .A1(n51), .B0(n1020), .B1(n2944), .C0(n1006), 
        .C1(n2943), .Y(n2324) );
  AOI222XLTS U3741 ( .A0(n3073), .A1(n4550), .B0(n3097), .B1(n4331), .C0(n1002), .C1(cacheDataOut[23]), .Y(n2322) );
  NAND4X1TS U3742 ( .A(n2316), .B(n2317), .C(n2318), .D(n2319), .Y(n2406) );
  AOI221X1TS U3743 ( .A0(n1980), .A1(n3015), .B0(n1077), .B1(n91), .C0(n2320), 
        .Y(n2319) );
  AOI222XLTS U3744 ( .A0(n1043), .A1(n632), .B0(n1020), .B1(n2946), .C0(n1006), 
        .C1(n2945), .Y(n2318) );
  AOI222XLTS U3745 ( .A0(n3073), .A1(n4546), .B0(n3096), .B1(n4328), .C0(n1002), .C1(cacheDataOut[22]), .Y(n2316) );
  NAND4X1TS U3746 ( .A(n2310), .B(n2311), .C(n2312), .D(n2313), .Y(n2407) );
  AOI221X1TS U3747 ( .A0(n1980), .A1(n3016), .B0(n1077), .B1(n65), .C0(n2314), 
        .Y(n2313) );
  AOI222XLTS U3748 ( .A0(n1042), .A1(n631), .B0(n1020), .B1(n2948), .C0(n1006), 
        .C1(n2947), .Y(n2312) );
  AOI222XLTS U3749 ( .A0(n3073), .A1(n4542), .B0(n3096), .B1(n4325), .C0(n2117), .C1(cacheDataOut[21]), .Y(n2310) );
  NAND4X1TS U3750 ( .A(n2304), .B(n2305), .C(n2306), .D(n2307), .Y(n2408) );
  AOI221X1TS U3751 ( .A0(n1980), .A1(n3017), .B0(n1077), .B1(n66), .C0(n2308), 
        .Y(n2307) );
  AOI222XLTS U3752 ( .A0(n1041), .A1(n52), .B0(n1020), .B1(n2950), .C0(n1006), 
        .C1(n2949), .Y(n2306) );
  AOI222XLTS U3753 ( .A0(n3073), .A1(n4538), .B0(n3096), .B1(n4322), .C0(n1000), .C1(cacheDataOut[20]), .Y(n2304) );
  NAND4X1TS U3754 ( .A(n2298), .B(n2299), .C(n2300), .D(n2301), .Y(n2409) );
  AOI221X1TS U3755 ( .A0(n2103), .A1(n3018), .B0(n1079), .B1(n67), .C0(n2302), 
        .Y(n2301) );
  AOI222XLTS U3756 ( .A0(n1044), .A1(n630), .B0(n1021), .B1(n2952), .C0(n1007), 
        .C1(n2951), .Y(n2300) );
  AOI222XLTS U3757 ( .A0(n3074), .A1(n4534), .B0(n3096), .B1(n4319), .C0(n1001), .C1(cacheDataOut[19]), .Y(n2298) );
  NAND4X1TS U3758 ( .A(n2292), .B(n2293), .C(n2294), .D(n2295), .Y(n2410) );
  AOI221X1TS U3759 ( .A0(n2103), .A1(n3019), .B0(n1079), .B1(n68), .C0(n2296), 
        .Y(n2295) );
  AOI222XLTS U3760 ( .A0(n1044), .A1(n629), .B0(n1021), .B1(n2954), .C0(n1007), 
        .C1(n2953), .Y(n2294) );
  AOI222XLTS U3761 ( .A0(n3074), .A1(n4531), .B0(n3095), .B1(n4316), .C0(n1001), .C1(cacheDataOut[18]), .Y(n2292) );
  NAND4X1TS U3762 ( .A(n2286), .B(n2287), .C(n2288), .D(n2289), .Y(n2411) );
  AOI221X1TS U3763 ( .A0(n2103), .A1(n3020), .B0(n1079), .B1(n69), .C0(n2290), 
        .Y(n2289) );
  AOI222XLTS U3764 ( .A0(n1044), .A1(n628), .B0(n1021), .B1(n2956), .C0(n1007), 
        .C1(n2955), .Y(n2288) );
  AOI222XLTS U3765 ( .A0(n3074), .A1(n4526), .B0(n3095), .B1(n4313), .C0(n998), 
        .C1(cacheDataOut[17]), .Y(n2286) );
  NAND4X1TS U3766 ( .A(n2280), .B(n2281), .C(n2282), .D(n2283), .Y(n2412) );
  AOI221X1TS U3767 ( .A0(n2103), .A1(n3021), .B0(n1079), .B1(n92), .C0(n2284), 
        .Y(n2283) );
  AOI222XLTS U3768 ( .A0(n1045), .A1(n627), .B0(n1021), .B1(n2958), .C0(n1007), 
        .C1(n2957), .Y(n2282) );
  AOI222XLTS U3769 ( .A0(n3074), .A1(n4523), .B0(n3095), .B1(n4310), .C0(n1002), .C1(cacheDataOut[16]), .Y(n2280) );
  NAND4X1TS U3770 ( .A(n2274), .B(n2275), .C(n2276), .D(n2277), .Y(n2413) );
  AOI221X1TS U3771 ( .A0(n2916), .A1(n3022), .B0(n1749), .B1(n70), .C0(n2278), 
        .Y(n2277) );
  AOI222XLTS U3772 ( .A0(n1044), .A1(n626), .B0(n1022), .B1(n2960), .C0(n1008), 
        .C1(n2959), .Y(n2276) );
  AOI222XLTS U3773 ( .A0(n3084), .A1(n4520), .B0(n3095), .B1(n4307), .C0(n1001), .C1(cacheDataOut[15]), .Y(n2274) );
  NAND4X1TS U3774 ( .A(n2268), .B(n2269), .C(n2270), .D(n2271), .Y(n2414) );
  AOI221X1TS U3775 ( .A0(n2914), .A1(n3023), .B0(n1210), .B1(n71), .C0(n2272), 
        .Y(n2271) );
  AOI222XLTS U3776 ( .A0(n1043), .A1(n625), .B0(n1022), .B1(n2962), .C0(n1008), 
        .C1(n2961), .Y(n2270) );
  AOI222XLTS U3777 ( .A0(n3084), .A1(n4515), .B0(n3094), .B1(n4304), .C0(n1001), .C1(cacheDataOut[14]), .Y(n2268) );
  NAND4X1TS U3778 ( .A(n2262), .B(n2263), .C(n2264), .D(n2265), .Y(n2415) );
  AOI221X1TS U3779 ( .A0(n2917), .A1(n3024), .B0(n1771), .B1(n72), .C0(n2266), 
        .Y(n2265) );
  AOI222XLTS U3780 ( .A0(n1042), .A1(n624), .B0(n1022), .B1(n2964), .C0(n1008), 
        .C1(n2963), .Y(n2264) );
  AOI222XLTS U3781 ( .A0(n3084), .A1(n4512), .B0(n3094), .B1(n4301), .C0(n1000), .C1(cacheDataOut[13]), .Y(n2262) );
  NAND4X1TS U3782 ( .A(n2256), .B(n2257), .C(n2258), .D(n2259), .Y(n2416) );
  AOI221X1TS U3783 ( .A0(n2914), .A1(n3025), .B0(n1210), .B1(n73), .C0(n2260), 
        .Y(n2259) );
  AOI222XLTS U3784 ( .A0(n1041), .A1(n623), .B0(n1022), .B1(n2966), .C0(n1008), 
        .C1(n2965), .Y(n2258) );
  AOI222XLTS U3785 ( .A0(n3084), .A1(n4508), .B0(n3094), .B1(n4298), .C0(n999), 
        .C1(cacheDataOut[12]), .Y(n2256) );
  NAND4X1TS U3786 ( .A(n2250), .B(n2251), .C(n2252), .D(n2253), .Y(n2417) );
  AOI221X1TS U3787 ( .A0(n2377), .A1(n3026), .B0(n1085), .B1(n74), .C0(n2254), 
        .Y(n2253) );
  AOI222XLTS U3788 ( .A0(n1035), .A1(n622), .B0(n1031), .B1(n2968), .C0(n2115), 
        .C1(n2967), .Y(n2252) );
  AOI222XLTS U3789 ( .A0(n3083), .A1(n4505), .B0(n3094), .B1(n4295), .C0(n992), 
        .C1(cacheDataOut[11]), .Y(n2250) );
  NAND4X1TS U3790 ( .A(n2244), .B(n2245), .C(n2246), .D(n2247), .Y(n2418) );
  AOI221X1TS U3791 ( .A0(n2377), .A1(n3027), .B0(n1085), .B1(n87), .C0(n2248), 
        .Y(n2247) );
  AOI222XLTS U3792 ( .A0(n1035), .A1(n621), .B0(n1031), .B1(n2970), .C0(n1016), 
        .C1(n2969), .Y(n2246) );
  AOI222XLTS U3793 ( .A0(n3082), .A1(n4502), .B0(n3100), .B1(n4292), .C0(n992), 
        .C1(cacheDataOut[10]), .Y(n2244) );
  NAND4X1TS U3794 ( .A(n2238), .B(n2239), .C(n2240), .D(n2241), .Y(n2419) );
  AOI221X1TS U3795 ( .A0(n2377), .A1(n3028), .B0(n1085), .B1(n75), .C0(n2242), 
        .Y(n2241) );
  AOI222XLTS U3796 ( .A0(n1035), .A1(n53), .B0(n1030), .B1(n2972), .C0(n1015), 
        .C1(n2971), .Y(n2240) );
  AOI222XLTS U3797 ( .A0(n3083), .A1(n4497), .B0(n3103), .B1(n4289), .C0(n992), 
        .C1(cacheDataOut[9]), .Y(n2238) );
  NAND4X1TS U3798 ( .A(n2232), .B(n2233), .C(n2234), .D(n2235), .Y(n2420) );
  AOI221X1TS U3799 ( .A0(n2377), .A1(n3029), .B0(n1085), .B1(n76), .C0(n2236), 
        .Y(n2235) );
  AOI222XLTS U3800 ( .A0(n1035), .A1(n620), .B0(n1029), .B1(n2974), .C0(n1014), 
        .C1(n2973), .Y(n2234) );
  AOI222XLTS U3801 ( .A0(n3082), .A1(n4494), .B0(n3098), .B1(n4286), .C0(n992), 
        .C1(cacheDataOut[8]), .Y(n2232) );
  NAND4X1TS U3802 ( .A(n2226), .B(n2227), .C(n2228), .D(n2229), .Y(n2421) );
  AOI221X1TS U3803 ( .A0(n2909), .A1(n3030), .B0(n1102), .B1(n77), .C0(n2230), 
        .Y(n2229) );
  AOI222XLTS U3804 ( .A0(n1036), .A1(n619), .B0(n1024), .B1(n2976), .C0(n1009), 
        .C1(n2975), .Y(n2228) );
  AOI222XLTS U3805 ( .A0(n3075), .A1(n4490), .B0(n3101), .B1(n4283), .C0(n993), 
        .C1(cacheDataOut[7]), .Y(n2226) );
  NAND4X1TS U3806 ( .A(n2220), .B(n2221), .C(n2222), .D(n2223), .Y(n2422) );
  AOI221X1TS U3807 ( .A0(n2909), .A1(n3031), .B0(n1102), .B1(n93), .C0(n2224), 
        .Y(n2223) );
  AOI222XLTS U3808 ( .A0(n1036), .A1(n618), .B0(n1024), .B1(n2978), .C0(n1009), 
        .C1(n2977), .Y(n2222) );
  AOI222XLTS U3809 ( .A0(n3075), .A1(n4487), .B0(n3100), .B1(n4280), .C0(n993), 
        .C1(cacheDataOut[6]), .Y(n2220) );
  NAND4X1TS U3810 ( .A(n2214), .B(n2215), .C(n2216), .D(n2217), .Y(n2423) );
  AOI221X1TS U3811 ( .A0(n2909), .A1(n3032), .B0(n1102), .B1(n78), .C0(n2218), 
        .Y(n2217) );
  AOI222XLTS U3812 ( .A0(n1036), .A1(n54), .B0(n1024), .B1(n2980), .C0(n1009), 
        .C1(n2979), .Y(n2216) );
  AOI222XLTS U3813 ( .A0(n3075), .A1(n4483), .B0(n3098), .B1(n4277), .C0(n993), 
        .C1(cacheDataOut[5]), .Y(n2214) );
  NAND4X1TS U3814 ( .A(n2208), .B(n2209), .C(n2210), .D(n2211), .Y(n2424) );
  AOI221X1TS U3815 ( .A0(n2909), .A1(n3033), .B0(n1102), .B1(n79), .C0(n2212), 
        .Y(n2211) );
  AOI222XLTS U3816 ( .A0(n1036), .A1(n617), .B0(n1024), .B1(n2982), .C0(n1009), 
        .C1(n2981), .Y(n2210) );
  AOI222XLTS U3817 ( .A0(n3075), .A1(n4479), .B0(n3101), .B1(n4274), .C0(n993), 
        .C1(cacheDataOut[4]), .Y(n2208) );
  NAND4X1TS U3818 ( .A(n2202), .B(n2203), .C(n2204), .D(n2205), .Y(n2425) );
  AOI221X1TS U3819 ( .A0(n2910), .A1(n3034), .B0(n1129), .B1(n80), .C0(n2206), 
        .Y(n2205) );
  AOI222XLTS U3820 ( .A0(n1037), .A1(n616), .B0(n1025), .B1(n2984), .C0(n1010), 
        .C1(n2983), .Y(n2204) );
  AOI222XLTS U3821 ( .A0(n3076), .A1(n4475), .B0(n3093), .B1(n4271), .C0(n994), 
        .C1(cacheDataOut[3]), .Y(n2202) );
  NAND4X1TS U3822 ( .A(n2196), .B(n2197), .C(n2198), .D(n2199), .Y(n2426) );
  AOI221X1TS U3823 ( .A0(n2910), .A1(n3035), .B0(n1129), .B1(n94), .C0(n2200), 
        .Y(n2199) );
  AOI222XLTS U3824 ( .A0(n1037), .A1(n55), .B0(n1025), .B1(n2986), .C0(n1010), 
        .C1(n2985), .Y(n2198) );
  AOI222XLTS U3825 ( .A0(n3076), .A1(n4471), .B0(n3093), .B1(n4268), .C0(n994), 
        .C1(cacheDataOut[2]), .Y(n2196) );
  NAND4X1TS U3826 ( .A(n2190), .B(n2191), .C(n2192), .D(n2193), .Y(n2427) );
  AOI221X1TS U3827 ( .A0(n2910), .A1(n3036), .B0(n1129), .B1(n88), .C0(n2194), 
        .Y(n2193) );
  AOI222XLTS U3828 ( .A0(n1037), .A1(n56), .B0(n1025), .B1(n2988), .C0(n1010), 
        .C1(n2987), .Y(n2192) );
  AOI222XLTS U3829 ( .A0(n3076), .A1(n4467), .B0(n3093), .B1(n4265), .C0(n994), 
        .C1(cacheDataOut[1]), .Y(n2190) );
  NAND4X1TS U3830 ( .A(n2184), .B(n2185), .C(n2186), .D(n2187), .Y(n2428) );
  AOI221X1TS U3831 ( .A0(n2910), .A1(n3037), .B0(n1129), .B1(n95), .C0(n2188), 
        .Y(n2187) );
  AOI222XLTS U3832 ( .A0(n1037), .A1(n57), .B0(n1025), .B1(n2990), .C0(n1010), 
        .C1(n2989), .Y(n2186) );
  AOI222XLTS U3833 ( .A0(n3076), .A1(n4463), .B0(n3093), .B1(n4262), .C0(n994), 
        .C1(cacheDataOut[0]), .Y(n2184) );
  NAND4X1TS U3834 ( .A(n2178), .B(n2179), .C(n2180), .D(n2181), .Y(n2429) );
  AOI221X1TS U3835 ( .A0(n2911), .A1(n2903), .B0(n1146), .B1(
        \requesterAddressbuffer[2][5] ), .C0(n2182), .Y(n2181) );
  AOI222XLTS U3836 ( .A0(n1038), .A1(\requesterAddressbuffer[0][5] ), .B0(
        n1026), .B1(\requesterAddressbuffer[6][5] ), .C0(n1011), .C1(n2921), 
        .Y(n2180) );
  AOI222XLTS U3837 ( .A0(n3077), .A1(n4603), .B0(n3092), .B1(n4051), .C0(n995), 
        .C1(readRequesterAddress[5]), .Y(n2178) );
  NAND4X1TS U3838 ( .A(n2172), .B(n2173), .C(n2174), .D(n2175), .Y(n2430) );
  AOI221X1TS U3839 ( .A0(n2911), .A1(n2904), .B0(n1146), .B1(
        \requesterAddressbuffer[2][4] ), .C0(n2176), .Y(n2175) );
  AOI222XLTS U3840 ( .A0(n1038), .A1(\requesterAddressbuffer[0][4] ), .B0(
        n1026), .B1(\requesterAddressbuffer[6][4] ), .C0(n1011), .C1(n2922), 
        .Y(n2174) );
  AOI222XLTS U3841 ( .A0(n3077), .A1(n4598), .B0(n3092), .B1(n4048), .C0(n995), 
        .C1(readRequesterAddress[4]), .Y(n2172) );
  NAND4X1TS U3842 ( .A(n2160), .B(n2161), .C(n2162), .D(n2163), .Y(n2432) );
  AOI221X1TS U3843 ( .A0(n2911), .A1(n2905), .B0(n1146), .B1(
        \requesterAddressbuffer[2][2] ), .C0(n2164), .Y(n2163) );
  AOI222XLTS U3844 ( .A0(n1038), .A1(\requesterAddressbuffer[0][2] ), .B0(
        n1026), .B1(\requesterAddressbuffer[6][2] ), .C0(n1011), .C1(n2923), 
        .Y(n2162) );
  AOI222XLTS U3845 ( .A0(n3077), .A1(n4591), .B0(n3092), .B1(n4042), .C0(n995), 
        .C1(readRequesterAddress[2]), .Y(n2160) );
  NAND4X1TS U3846 ( .A(n2154), .B(n2155), .C(n2156), .D(n2157), .Y(n2433) );
  AOI221X1TS U3847 ( .A0(n2912), .A1(n2906), .B0(n1162), .B1(
        \requesterAddressbuffer[2][1] ), .C0(n2158), .Y(n2157) );
  AOI222XLTS U3848 ( .A0(n1039), .A1(\requesterAddressbuffer[0][1] ), .B0(
        n1027), .B1(\requesterAddressbuffer[6][1] ), .C0(n1012), .C1(n2924), 
        .Y(n2156) );
  AOI222XLTS U3849 ( .A0(n3078), .A1(n4586), .B0(n3091), .B1(n4039), .C0(n996), 
        .C1(readRequesterAddress[1]), .Y(n2154) );
  NAND4X1TS U3850 ( .A(n2142), .B(n2143), .C(n2144), .D(n2145), .Y(n2435) );
  AOI221X1TS U3851 ( .A0(n2912), .A1(n3038), .B0(n1162), .B1(n81), .C0(n2146), 
        .Y(n2145) );
  AOI222XLTS U3852 ( .A0(n1039), .A1(n642), .B0(n1027), .B1(n2992), .C0(n1012), 
        .C1(n2991), .Y(n2144) );
  AOI222XLTS U3853 ( .A0(n3078), .A1(n4236), .B0(n3091), .B1(n4009), .C0(n996), 
        .C1(readRequesterAddress[5]), .Y(n2142) );
  NAND4X1TS U3854 ( .A(n2136), .B(n2137), .C(n2138), .D(n2139), .Y(n2436) );
  AOI221X1TS U3855 ( .A0(n2912), .A1(n3039), .B0(n1162), .B1(n82), .C0(n2140), 
        .Y(n2139) );
  AOI222XLTS U3856 ( .A0(n1039), .A1(n615), .B0(n1027), .B1(n2994), .C0(n1012), 
        .C1(n2993), .Y(n2138) );
  AOI222XLTS U3857 ( .A0(n3078), .A1(n4233), .B0(n3091), .B1(n4006), .C0(n996), 
        .C1(readRequesterAddress[4]), .Y(n2136) );
  NAND4X1TS U3858 ( .A(n2130), .B(n2131), .C(n2132), .D(n2133), .Y(n2437) );
  AOI221X1TS U3859 ( .A0(n2913), .A1(n3040), .B0(n1193), .B1(n83), .C0(n2134), 
        .Y(n2133) );
  AOI222XLTS U3860 ( .A0(n1040), .A1(n641), .B0(n1028), .B1(n2996), .C0(n1013), 
        .C1(n2995), .Y(n2132) );
  AOI222XLTS U3861 ( .A0(n3079), .A1(n4230), .B0(n3102), .B1(n4003), .C0(n997), 
        .C1(readRequesterAddress[3]), .Y(n2130) );
  NAND4X1TS U3862 ( .A(n2124), .B(n2125), .C(n2126), .D(n2127), .Y(n2438) );
  AOI221X1TS U3863 ( .A0(n2913), .A1(n3041), .B0(n1193), .B1(n58), .C0(n2128), 
        .Y(n2127) );
  AOI222XLTS U3864 ( .A0(n1040), .A1(n640), .B0(n1028), .B1(n2998), .C0(n1013), 
        .C1(n2997), .Y(n2126) );
  AOI222XLTS U3865 ( .A0(n3079), .A1(n4227), .B0(n3090), .B1(n4000), .C0(n997), 
        .C1(readRequesterAddress[2]), .Y(n2124) );
  NAND4X1TS U3866 ( .A(n2118), .B(n2119), .C(n2120), .D(n2121), .Y(n2439) );
  AOI221X1TS U3867 ( .A0(n2913), .A1(n3042), .B0(n1193), .B1(n84), .C0(n2122), 
        .Y(n2121) );
  AOI222XLTS U3868 ( .A0(n1040), .A1(n639), .B0(n1028), .B1(n3000), .C0(n1013), 
        .C1(n2999), .Y(n2120) );
  AOI222XLTS U3869 ( .A0(n3079), .A1(n4224), .B0(n3090), .B1(n3997), .C0(n997), 
        .C1(readRequesterAddress[1]), .Y(n2118) );
  NAND4X1TS U3870 ( .A(n2104), .B(n2105), .C(n2106), .D(n2107), .Y(n2440) );
  AOI221X1TS U3871 ( .A0(n2913), .A1(n3043), .B0(n1193), .B1(n85), .C0(n2110), 
        .Y(n2107) );
  AOI222XLTS U3872 ( .A0(n1040), .A1(n48), .B0(n1028), .B1(n3002), .C0(n1013), 
        .C1(n3001), .Y(n2106) );
  AOI222XLTS U3873 ( .A0(n3079), .A1(n4221), .B0(n3090), .B1(n3994), .C0(n997), 
        .C1(readRequesterAddress[0]), .Y(n2104) );
  NAND4X1TS U3874 ( .A(n2166), .B(n2167), .C(n2168), .D(n2169), .Y(n2431) );
  AOI221X1TS U3875 ( .A0(n2911), .A1(n2907), .B0(n1146), .B1(
        \requesterAddressbuffer[2][3] ), .C0(n2170), .Y(n2169) );
  AOI222XLTS U3876 ( .A0(n1038), .A1(\requesterAddressbuffer[0][3] ), .B0(
        n1026), .B1(\requesterAddressbuffer[6][3] ), .C0(n1011), .C1(n2925), 
        .Y(n2168) );
  AOI222XLTS U3877 ( .A0(n3077), .A1(n4594), .B0(n3092), .B1(n4045), .C0(n995), 
        .C1(readRequesterAddress[3]), .Y(n2166) );
  NAND4X1TS U3878 ( .A(n2148), .B(n2149), .C(n2150), .D(n2151), .Y(n2434) );
  AOI221X1TS U3879 ( .A0(n2912), .A1(n2908), .B0(n1162), .B1(
        \requesterAddressbuffer[2][0] ), .C0(n2152), .Y(n2151) );
  AOI222XLTS U3880 ( .A0(n1039), .A1(\requesterAddressbuffer[0][0] ), .B0(
        n1027), .B1(\requesterAddressbuffer[6][0] ), .C0(n1012), .C1(n2926), 
        .Y(n2150) );
  AOI222XLTS U3881 ( .A0(n3078), .A1(n4583), .B0(n3091), .B1(n4036), .C0(n996), 
        .C1(readRequesterAddress[0]), .Y(n2148) );
  INVX2TS U3882 ( .A(n4214), .Y(n4213) );
  OAI32X1TS U3883 ( .A0(n4831), .A1(n954), .A2(n2012), .B0(n2013), .B1(n2014), 
        .Y(n2450) );
  NOR4BX1TS U3884 ( .AN(n2022), .B(n2023), .C(n2024), .D(n2025), .Y(n2013) );
  OAI31X1TS U3885 ( .A0(n2015), .A1(n486), .A2(n2016), .B0(n4606), .Y(n2014)
         );
  OAI22X1TS U3886 ( .A0(n2030), .A1(n647), .B0(n2031), .B1(n599), .Y(n2023) );
  OAI211X1TS U3887 ( .A0(n3992), .A1(n3050), .B0(n2096), .C0(n2097), .Y(n2441)
         );
  AOI22X1TS U3888 ( .A0(n114), .A1(n2098), .B0(n3117), .B1(
        destinationAddressOut[13]), .Y(n2096) );
  AOI222XLTS U3889 ( .A0(n3080), .A1(n4260), .B0(n3069), .B1(
        destinationAddressIn_NORTH[13]), .C0(n3089), .C1(n4033), .Y(n2097) );
  NAND4X1TS U3890 ( .A(n2099), .B(n2100), .C(n2101), .D(n2102), .Y(n2098) );
  OAI211X1TS U3891 ( .A0(n3989), .A1(n3050), .B0(n2089), .C0(n2090), .Y(n2442)
         );
  AOI22X1TS U3892 ( .A0(n182), .A1(n2091), .B0(n3117), .B1(
        destinationAddressOut[12]), .Y(n2089) );
  AOI222XLTS U3893 ( .A0(n3080), .A1(n4257), .B0(n2048), .B1(
        destinationAddressIn_NORTH[12]), .C0(n3089), .C1(n4030), .Y(n2090) );
  NAND4X1TS U3894 ( .A(n2092), .B(n2093), .C(n2094), .D(n2095), .Y(n2091) );
  OAI211X1TS U3895 ( .A0(n3986), .A1(n3050), .B0(n2082), .C0(n2083), .Y(n2443)
         );
  AOI22X1TS U3896 ( .A0(n184), .A1(n2084), .B0(n3117), .B1(
        destinationAddressOut[11]), .Y(n2082) );
  AOI222XLTS U3897 ( .A0(n3080), .A1(n4254), .B0(n2048), .B1(
        destinationAddressIn_NORTH[11]), .C0(n3089), .C1(n4027), .Y(n2083) );
  NAND4X1TS U3898 ( .A(n2085), .B(n2086), .C(n2087), .D(n2088), .Y(n2084) );
  OAI211X1TS U3899 ( .A0(n3983), .A1(n3051), .B0(n2075), .C0(n2076), .Y(n2444)
         );
  AOI22X1TS U3900 ( .A0(n182), .A1(n2077), .B0(n3117), .B1(
        destinationAddressOut[10]), .Y(n2075) );
  AOI222XLTS U3901 ( .A0(n3080), .A1(n4251), .B0(n3068), .B1(
        destinationAddressIn_NORTH[10]), .C0(n3088), .C1(n4024), .Y(n2076) );
  NAND4X1TS U3902 ( .A(n2078), .B(n2079), .C(n2080), .D(n2081), .Y(n2077) );
  OAI211X1TS U3903 ( .A0(n3980), .A1(n3051), .B0(n2068), .C0(n2069), .Y(n2445)
         );
  AOI22X1TS U3904 ( .A0(n114), .A1(n2070), .B0(n3118), .B1(
        destinationAddressOut[9]), .Y(n2068) );
  AOI222XLTS U3905 ( .A0(n3086), .A1(n4248), .B0(n3055), .B1(
        destinationAddressIn_NORTH[9]), .C0(n3089), .C1(n4021), .Y(n2069) );
  NAND4X1TS U3906 ( .A(n2071), .B(n2072), .C(n2073), .D(n2074), .Y(n2070) );
  OAI211X1TS U3907 ( .A0(n3977), .A1(n3051), .B0(n2061), .C0(n2062), .Y(n2446)
         );
  AOI22X1TS U3908 ( .A0(n183), .A1(n2063), .B0(n3118), .B1(
        destinationAddressOut[8]), .Y(n2061) );
  AOI222XLTS U3909 ( .A0(n3085), .A1(n4245), .B0(n3055), .B1(
        destinationAddressIn_NORTH[8]), .C0(n3088), .C1(n4018), .Y(n2062) );
  NAND4X1TS U3910 ( .A(n2064), .B(n2065), .C(n2066), .D(n2067), .Y(n2063) );
  OAI211X1TS U3911 ( .A0(n3974), .A1(n3052), .B0(n2054), .C0(n2055), .Y(n2447)
         );
  AOI22X1TS U3912 ( .A0(n181), .A1(n2056), .B0(n3118), .B1(
        destinationAddressOut[7]), .Y(n2054) );
  AOI222XLTS U3913 ( .A0(n3086), .A1(n4242), .B0(n3055), .B1(
        destinationAddressIn_NORTH[7]), .C0(n3088), .C1(n4015), .Y(n2055) );
  NAND4X1TS U3914 ( .A(n2057), .B(n2058), .C(n2059), .D(n2060), .Y(n2056) );
  OAI211X1TS U3915 ( .A0(n3971), .A1(n3052), .B0(n2046), .C0(n2047), .Y(n2448)
         );
  AOI22X1TS U3916 ( .A0(n183), .A1(n2049), .B0(n3118), .B1(
        destinationAddressOut[6]), .Y(n2046) );
  AOI222XLTS U3917 ( .A0(n3087), .A1(n4239), .B0(n3055), .B1(
        destinationAddressIn_NORTH[6]), .C0(n3088), .C1(n4012), .Y(n2047) );
  NAND4X1TS U3918 ( .A(n2050), .B(n2051), .C(n2052), .D(n2053), .Y(n2049) );
  NAND2X1TS U3919 ( .A(n4206), .B(n692), .Y(n1809) );
  OAI33XLTS U3920 ( .A0(n4215), .A1(n692), .A2(n1783), .B0(n137), .B1(n946), 
        .B2(n1813), .Y(n1812) );
  OAI2BB2XLTS U3921 ( .B0(n163), .B1(n137), .A0N(n162), .A1N(readIn_NORTH), 
        .Y(n1777) );
  INVX2TS U3922 ( .A(readIn_NORTH), .Y(n964) );
  INVX2TS U3923 ( .A(destinationAddressIn_WEST[13]), .Y(n4034) );
  INVX2TS U3924 ( .A(destinationAddressIn_WEST[11]), .Y(n4028) );
  INVX2TS U3925 ( .A(destinationAddressIn_WEST[9]), .Y(n4022) );
  INVX2TS U3926 ( .A(destinationAddressIn_WEST[12]), .Y(n4031) );
  INVX2TS U3927 ( .A(destinationAddressIn_WEST[10]), .Y(n4025) );
  INVX2TS U3928 ( .A(destinationAddressIn_WEST[8]), .Y(n4019) );
  OAI21X1TS U3929 ( .A0(n122), .A1(n1092), .B0(n3789), .Y(n2884) );
  NOR2X1TS U3930 ( .A(n1094), .B(n1092), .Y(n2883) );
  AOI21X1TS U3931 ( .A0(n114), .A1(n140), .B0(n98), .Y(n1094) );
  AO22X1TS U3932 ( .A0(n658), .A1(n942), .B0(n181), .B1(n10), .Y(n2889) );
  XOR2X1TS U3933 ( .A(n960), .B(n98), .Y(n2899) );
  XNOR2X1TS U3934 ( .A(n97), .B(n46), .Y(n1091) );
  AOI22X1TS U3935 ( .A0(n477), .A1(n3131), .B0(n493), .B1(n3177), .Y(n2099) );
  AOI22X1TS U3936 ( .A0(n477), .A1(n3132), .B0(n493), .B1(n3176), .Y(n2092) );
  AOI22X1TS U3937 ( .A0(n477), .A1(n3133), .B0(n493), .B1(n3175), .Y(n2085) );
  AOI22X1TS U3938 ( .A0(n477), .A1(n3134), .B0(n493), .B1(n3174), .Y(n2078) );
  AOI22X1TS U3939 ( .A0(n478), .A1(n3135), .B0(n494), .B1(n3173), .Y(n2071) );
  AOI22X1TS U3940 ( .A0(n478), .A1(n3136), .B0(n494), .B1(n3172), .Y(n2064) );
  AOI22X1TS U3941 ( .A0(n478), .A1(n3137), .B0(n494), .B1(n3171), .Y(n2057) );
  AOI22X1TS U3942 ( .A0(n478), .A1(n3138), .B0(n494), .B1(n3170), .Y(n2050) );
  AOI22X1TS U3943 ( .A0(n165), .A1(n3123), .B0(n174), .B1(n3185), .Y(n2102) );
  AOI22X1TS U3944 ( .A0(n166), .A1(n3124), .B0(n648), .B1(n3184), .Y(n2095) );
  AOI22X1TS U3945 ( .A0(n165), .A1(n3125), .B0(n175), .B1(n3183), .Y(n2088) );
  AOI22X1TS U3946 ( .A0(n166), .A1(n3126), .B0(n174), .B1(n3182), .Y(n2081) );
  AOI22X1TS U3947 ( .A0(n165), .A1(n3127), .B0(n648), .B1(n3181), .Y(n2074) );
  AOI22X1TS U3948 ( .A0(n166), .A1(n3128), .B0(n175), .B1(n3180), .Y(n2067) );
  AOI22X1TS U3949 ( .A0(n165), .A1(n3129), .B0(n174), .B1(n3179), .Y(n2060) );
  AOI22X1TS U3950 ( .A0(n166), .A1(n3130), .B0(n648), .B1(n3178), .Y(n2053) );
  AOI22X1TS U3951 ( .A0(n491), .A1(n3155), .B0(n3154), .B1(n172), .Y(n2100) );
  AOI22X1TS U3952 ( .A0(n491), .A1(n3157), .B0(n3156), .B1(n172), .Y(n2093) );
  AOI22X1TS U3953 ( .A0(n491), .A1(n3159), .B0(n3158), .B1(n171), .Y(n2086) );
  AOI22X1TS U3954 ( .A0(n491), .A1(n3161), .B0(n3160), .B1(n172), .Y(n2079) );
  AOI22X1TS U3955 ( .A0(n492), .A1(n3163), .B0(n3162), .B1(n652), .Y(n2072) );
  AOI22X1TS U3956 ( .A0(n492), .A1(n3165), .B0(n3164), .B1(n171), .Y(n2065) );
  AOI22X1TS U3957 ( .A0(n492), .A1(n3167), .B0(n3166), .B1(n172), .Y(n2058) );
  AOI22X1TS U3958 ( .A0(n492), .A1(n3169), .B0(n3168), .B1(n652), .Y(n2051) );
  AOI22X1TS U3959 ( .A0(n653), .A1(n3140), .B0(n169), .B1(n3139), .Y(n2101) );
  AOI22X1TS U3960 ( .A0(n176), .A1(n3142), .B0(n169), .B1(n3141), .Y(n2094) );
  AOI22X1TS U3961 ( .A0(n177), .A1(n3144), .B0(n168), .B1(n3143), .Y(n2087) );
  AOI22X1TS U3962 ( .A0(n177), .A1(n480), .B0(n169), .B1(n3145), .Y(n2080) );
  AOI22X1TS U3963 ( .A0(n176), .A1(n3147), .B0(n657), .B1(n3146), .Y(n2073) );
  AOI22X1TS U3964 ( .A0(n177), .A1(n3149), .B0(n168), .B1(n3148), .Y(n2066) );
  AOI22X1TS U3965 ( .A0(n653), .A1(n3151), .B0(n169), .B1(n3150), .Y(n2059) );
  AOI22X1TS U3966 ( .A0(n176), .A1(n3153), .B0(n657), .B1(n3152), .Y(n2052) );
  AOI221X1TS U3967 ( .A0(n175), .A1(\readOutbuffer[2] ), .B0(n177), .B1(
        readOutbuffer_7), .C0(n6248), .Y(n2022) );
  AOI32XLTS U3968 ( .A0(n487), .A1(n1787), .A2(n1788), .B0(n3809), .B1(n598), 
        .Y(n2566) );
  OAI221XLTS U3969 ( .A0(n950), .A1(n149), .B0(n2), .B1(n580), .C0(n1924), .Y(
        n2500) );
  OAI221XLTS U3970 ( .A0(n949), .A1(n147), .B0(n466), .B1(n566), .C0(n1925), 
        .Y(n2499) );
  OAI221XLTS U3971 ( .A0(n950), .A1(n161), .B0(n2), .B1(n577), .C0(n1926), .Y(
        n2498) );
  OAI221XLTS U3972 ( .A0(n949), .A1(n154), .B0(n466), .B1(n578), .C0(n1927), 
        .Y(n2497) );
  OAI221XLTS U3973 ( .A0(n950), .A1(n158), .B0(n185), .B1(n567), .C0(n1928), 
        .Y(n2496) );
  OAI221XLTS U3974 ( .A0(n949), .A1(n152), .B0(n466), .B1(n581), .C0(n1929), 
        .Y(n2495) );
  OAI221XLTS U3975 ( .A0(n950), .A1(n156), .B0(n133), .B1(n579), .C0(n1930), 
        .Y(n2494) );
  OAI221XLTS U3976 ( .A0(n949), .A1(n151), .B0(n133), .B1(n568), .C0(n1931), 
        .Y(n2493) );
  OAI221XLTS U3977 ( .A0(n941), .A1(n472), .B0(n466), .B1(n644), .C0(n1750), 
        .Y(n2574) );
  NAND4XLTS U3978 ( .A(selectBit_NORTH), .B(n474), .C(n975), .D(n1), .Y(n2017)
         );
  AOI32XLTS U3979 ( .A0(n102), .A1(n1795), .A2(n1796), .B0(n3918), .B1(n646), 
        .Y(n2565) );
  OAI221XLTS U3980 ( .A0(n112), .A1(n148), .B0(n959), .B1(n550), .C0(n1948), 
        .Y(n2486) );
  OAI221XLTS U3981 ( .A0(n111), .A1(n146), .B0(n958), .B1(n557), .C0(n1949), 
        .Y(n2485) );
  OAI221XLTS U3982 ( .A0(n112), .A1(n160), .B0(n959), .B1(n551), .C0(n1950), 
        .Y(n2484) );
  OAI221XLTS U3983 ( .A0(n111), .A1(n155), .B0(n958), .B1(n558), .C0(n1951), 
        .Y(n2483) );
  OAI221XLTS U3984 ( .A0(n112), .A1(n159), .B0(n959), .B1(n552), .C0(n1952), 
        .Y(n2482) );
  OAI221XLTS U3985 ( .A0(n1751), .A1(n153), .B0(n958), .B1(n559), .C0(n1953), 
        .Y(n2481) );
  OAI221XLTS U3986 ( .A0(n1751), .A1(n157), .B0(n959), .B1(n553), .C0(n1954), 
        .Y(n2480) );
  OAI221XLTS U3987 ( .A0(n111), .A1(n150), .B0(n958), .B1(n563), .C0(n1955), 
        .Y(n2479) );
  OAI221XLTS U3988 ( .A0(n1751), .A1(n472), .B0(n1752), .B1(n604), .C0(n1753), 
        .Y(n2573) );
endmodule


module outputPortArbiter_1 ( clk, reset, selectBit_NORTH, 
        destinationAddressIn_NORTH, requesterAddressIn_NORTH, readIn_NORTH, 
        writeIn_NORTH, dataIn_NORTH, selectBit_SOUTH, 
        destinationAddressIn_SOUTH, requesterAddressIn_SOUTH, readIn_SOUTH, 
        writeIn_SOUTH, dataIn_SOUTH, selectBit_EAST, destinationAddressIn_EAST, 
        requesterAddressIn_EAST, readIn_EAST, writeIn_EAST, dataIn_EAST, 
        selectBit_WEST, destinationAddressIn_WEST, requesterAddressIn_WEST, 
        readIn_WEST, writeIn_WEST, dataIn_WEST, readReady, 
        readRequesterAddress, cacheDataOut, destinationAddressOut, 
        requesterAddressOut, readOut, writeOut, dataOut );
  input [13:0] destinationAddressIn_NORTH;
  input [5:0] requesterAddressIn_NORTH;
  input [31:0] dataIn_NORTH;
  input [13:0] destinationAddressIn_SOUTH;
  input [5:0] requesterAddressIn_SOUTH;
  input [31:0] dataIn_SOUTH;
  input [13:0] destinationAddressIn_EAST;
  input [5:0] requesterAddressIn_EAST;
  input [31:0] dataIn_EAST;
  input [13:0] destinationAddressIn_WEST;
  input [5:0] requesterAddressIn_WEST;
  input [31:0] dataIn_WEST;
  input [5:0] readRequesterAddress;
  input [31:0] cacheDataOut;
  output [13:0] destinationAddressOut;
  output [5:0] requesterAddressOut;
  output [31:0] dataOut;
  input clk, reset, selectBit_NORTH, readIn_NORTH, writeIn_NORTH,
         selectBit_SOUTH, readIn_SOUTH, writeIn_SOUTH, selectBit_EAST,
         readIn_EAST, writeIn_EAST, selectBit_WEST, readIn_WEST, writeIn_WEST,
         readReady;
  output readOut, writeOut;
  wire   n2486, n2484, n2482, n2480, n2457, n2455, n2453, n2485, n2483, n2481,
         n2458, n2454, n2451, n2479, n2456, n2452, n2499, n2496, n2493, n2498,
         n2497, n2494, n2500, n2495, n2541, n2540, n2537, n2535, n2511, n2507,
         n2556, n2555, n2554, n2552, n567, n2551, n2550, n2549, n2472, n2471,
         n2470, n2469, n2468, n2467, n2466, n2465, n2553, n2542, n2539, n2538,
         n2536, n2510, n2509, n2508, n2638, n2624, n2617, n2610, n2609, n2608,
         n2607, n2606, n2605, n2604, n2603, n2602, n2601, n2600, n2599, n2598,
         n2597, n2596, n2595, n2594, n2593, n2592, n2591, n2590, n2589, n2588,
         n2587, n2586, n2585, n2584, n2583, n2582, n2581, n2580, n2579, n2561,
         n2560, n2559, n2557, n2642, n2640, n2639, n2637, n2635, n2634, n2633,
         n2631, n2628, n2627, n2626, n2625, n2623, n2620, n2618, n2616, n2615,
         n2614, n2612, n2611, n2562, n2558, n2641, n2636, n2632, n2630, n2629,
         n2622, n2621, n2619, n2613, n2543, n2850,
         \requesterAddressbuffer[2][2] , n2849, \requesterAddressbuffer[2][3] ,
         n2847, \requesterAddressbuffer[2][5] , n2840,
         \requesterAddressbuffer[0][0] , n2839, \requesterAddressbuffer[0][1] ,
         n2838, \requesterAddressbuffer[0][2] , n2836,
         \requesterAddressbuffer[0][4] , n2852, \requesterAddressbuffer[2][0] ,
         n2851, \requesterAddressbuffer[2][1] , n2848,
         \requesterAddressbuffer[2][4] , n2837, \requesterAddressbuffer[0][3] ,
         n2835, \requesterAddressbuffer[0][5] , n2566, \readOutbuffer[2] ,
         readOutbuffer_7, n2569, n2578, n2568, n2564, n2563, n2882, n2881,
         n2879, n2880, n2878, n2877, n2572, n2573, n2731, n4654, n2768, n2754,
         n2748, n2746, n2739, n2834, n2833, n2832, n2829, n2825, n2814, n2811,
         n2807, n2806, n2736, n99, n2734, n98, n2733, n97, n2725, n96, n2723,
         n95, n2720, n94, n2718, n93, n2715, n92, n2713, n91, n2504, n90,
         n2492, n2491, n2464, n89, n2460, n88, n2738, n87, n2737, n86, n2735,
         n85, n2732, n84, n2730, n83, n2729, n82, n2728, n81, n2727, n80,
         n2726, n79, n2724, n78, n2722, n77, n2721, n76, n2719, n75, n2717,
         n74, n2716, n73, n2714, n72, n2712, n71, n2711, n70, n2710, n69,
         n2709, n68, n2708, n67, n2707, n66, n2506, n65, n2505, n64, n2503,
         n63, n2502, n62, n2501, n61, n2767, n2766, n2765, n2756, n2755, n2753,
         n2740, n2831, n60, n2830, n59, n2828, n58, n2827, n57, n2826, n56,
         n2824, n55, n2823, n54, n2822, n53, n2821, n52, n2820, n51, n2819,
         n50, n2818, n49, n2817, n48, n2816, n47, n2815, n46, n2813, n2812,
         n2810, n2809, n2808, n2805, n2804, n2803, n2463, n2462, n2461, n2459,
         n2571, n2574, n2577, n2570, n2565, n2567, n2889, n9, N4718, n4844,
         n4841, n2434, n4845, n2431, n4846, n2450, n4843, n2440, n4768, n2439,
         n4759, n2438, n4750, n2437, n4741, n2436, n4732, n2435, n4723, n2433,
         n4722, n2432, n4721, n2430, n4720, n2429, n4719, n2428, n4710, n2427,
         n4701, n2426, n4692, n2425, n4683, n2424, n4674, n2423, n4665, n2422,
         n4656, n2421, n4647, n2420, n4638, n2419, n4629, n2418, n4620, n2417,
         n4611, n2416, n4602, n2415, n4593, n2414, n4584, n2413, n4575, n2412,
         n4566, n2411, n4557, n2410, n4548, n2409, n4539, n2408, n4530, n2407,
         n4521, n2406, n4512, n2405, n4503, n2404, n4494, n2403, n4485, n2402,
         n4476, n2401, n4467, n2400, n4458, n2399, n4449, n2398, n4440, n2397,
         n4431, n2448, n2447, n2446, n2445, n2444, n2443, n2442, n2441, n2524,
         n2530, n2674, n2672, n2671, n2670, n2669, n2668, n2667, n2666, n2665,
         n2664, n2662, n2661, n2660, n2657, n2656, n2655, n2654, n2653, n2652,
         n2651, n2650, n2649, n2648, n2647, n2646, n2645, n2644, n2534, n2533,
         n2532, n2531, n2673, n2663, n2659, n2658, n2643, n2474, n2516, n2802,
         n2801, n2799, n2798, n2796, n2795, n2793, n2791, n2790, n2789, n2788,
         n2787, n2786, n2785, n2784, n2781, n2779, n2778, n2777, n2776, n2774,
         n2773, n2772, n2771, n2478, n2477, n2476, n2475, n2473, n2548, n2547,
         n2546, n2545, n2520, n2519, n2518, n2517, n2515, n2800, n2797, n2794,
         n2792, n2783, n2782, n2780, n2775, n2544, n2858,
         \requesterAddressbuffer[3][0] , n2857, \requesterAddressbuffer[3][1] ,
         n2856, \requesterAddressbuffer[3][2] , n2855,
         \requesterAddressbuffer[3][3] , n2853, \requesterAddressbuffer[3][5] ,
         n2854, \requesterAddressbuffer[3][4] , n2875,
         \requesterAddressbuffer[6][1] , n2874, \requesterAddressbuffer[6][2] ,
         n2873, \requesterAddressbuffer[6][3] , n2872,
         \requesterAddressbuffer[6][4] , n2871, \requesterAddressbuffer[6][5] ,
         n2876, \requesterAddressbuffer[6][0] , n2870, n2869, n2868, n2867,
         n2866, n2865, n2576, n2860, n2859, n2864, n2863, n2862, n2861, n2846,
         n2845, n2844, n2843, n2842, n2841, n2528, n2527, n2526, n2525, n2523,
         n2522, n2883, n2884, n8, n2529, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2521, n2885, n6257,
         n2888, n5327, n2887, n5323, n2886, n5326, n2769, n2770, n2490, n2487,
         n2488, n2489, n2741, n2742, n2744, n2745, n2747, n2749, n2750, n2751,
         n2752, n2757, n2758, n2759, n2761, n2762, n2763, n2743, n2760, n2764,
         n2512, n2513, n2514, n2575, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n781, n782, n783, n784, n785, n788, n790, n791, n794, n797, n798,
         n801, n802, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n909, n910, n911, n912, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n926, n928, n929, n930, n932,
         n933, n934, n935, n936, n938, n940, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n972, n973, n974, n981, n982, n983, n984, n985, n998,
         n1031, n1086, n1132, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
         n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2449, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n1, n2, n3, n4, n5, n6, n7, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n780, n786, n787, n789, n792, n793, n795, n796, n799,
         n800, n803, n804, n805, n907, n908, n913, n914, n915, n925, n927,
         n931, n937, n939, n941, n971, n975, n976, n977, n978, n979, n980,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1133, n1134, n1155, n1199, n1215, n1246, n1662, n1794,
         n1846, n1919, n1988, n2098, n2158, n2955, n2956, n2964, n2965, n2966,
         n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n3058,
         n3059, n3060, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573;

  DFFNSRX2TS \dataoutbuffer_reg[0][0]  ( .D(n2834), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n698) );
  DFFNSRX2TS \dataoutbuffer_reg[0][1]  ( .D(n2833), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n699) );
  DFFNSRX2TS \dataoutbuffer_reg[0][2]  ( .D(n2832), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n700) );
  DFFNSRX2TS \dataoutbuffer_reg[0][5]  ( .D(n2829), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n701) );
  DFFNSRX2TS \dataoutbuffer_reg[0][9]  ( .D(n2825), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n702) );
  DFFNSRX2TS \dataoutbuffer_reg[0][20]  ( .D(n2814), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n703) );
  DFFNSRX2TS \dataoutbuffer_reg[0][23]  ( .D(n2811), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n704) );
  DFFNSRX2TS \dataoutbuffer_reg[0][27]  ( .D(n2807), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n705) );
  DFFNSRX2TS \dataoutbuffer_reg[0][28]  ( .D(n2806), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n706) );
  DFFNSRX2TS \dataoutbuffer_reg[0][21]  ( .D(n2813), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n753) );
  DFFNSRX2TS \dataoutbuffer_reg[0][22]  ( .D(n2812), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n754) );
  DFFNSRX2TS \dataoutbuffer_reg[0][24]  ( .D(n2810), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n755) );
  DFFNSRX2TS \dataoutbuffer_reg[0][25]  ( .D(n2809), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n756) );
  DFFNSRX2TS \dataoutbuffer_reg[0][26]  ( .D(n2808), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n757) );
  DFFNSRX2TS \dataoutbuffer_reg[0][29]  ( .D(n2805), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n758) );
  DFFNSRX2TS \dataoutbuffer_reg[0][30]  ( .D(n2804), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n759) );
  DFFNSRX2TS \dataoutbuffer_reg[0][31]  ( .D(n2803), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n760) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][1]  ( .D(n2463), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n761) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][2]  ( .D(n2462), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n762) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][3]  ( .D(n2461), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n763) );
  DFFNSRX2TS \destinationAddressbuffer_reg[0][5]  ( .D(n2459), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n764) );
  DFFNSRX2TS \dataoutbuffer_reg[3][7]  ( .D(n2731), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n692), .QN(n4654) );
  DFFNSRX2TS empty_reg_reg ( .D(n2885), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        n6257), .QN(n459) );
  DFFNSRX2TS \read_reg_reg[0]  ( .D(n2889), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n9), .QN(n458) );
  DFFNSRX2TS \read_reg_reg[2]  ( .D(n2884), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n8), .QN(n466) );
  DFFNSRX2TS \read_reg_reg[1]  ( .D(n2883), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n1), .QN(n4) );
  DFFNSRX2TS \write_reg_reg[0]  ( .D(n2888), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n3), .QN(n5327) );
  DFFNSRX2TS \write_reg_reg[2]  ( .D(n2886), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n493), .QN(n5326) );
  DFFNSRX2TS writeOut_reg ( .D(n679), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        writeOut), .QN(n4841) );
  DFFNSRX2TS \requesterAddressOut_reg[0]  ( .D(n2434), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[0]), .QN(n4845) );
  DFFNSRX2TS \requesterAddressOut_reg[3]  ( .D(n2431), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[3]), .QN(n4846) );
  DFFNSRX2TS readOut_reg ( .D(n2450), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        readOut), .QN(n4843) );
  DFFNSRX2TS \destinationAddressOut_reg[0]  ( .D(n2440), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[0]), .QN(n4768) );
  DFFNSRX2TS \destinationAddressOut_reg[1]  ( .D(n2439), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[1]), .QN(n4759) );
  DFFNSRX2TS \destinationAddressOut_reg[2]  ( .D(n2438), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[2]), .QN(n4750) );
  DFFNSRX2TS \destinationAddressOut_reg[3]  ( .D(n2437), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[3]), .QN(n4741) );
  DFFNSRX2TS \destinationAddressOut_reg[4]  ( .D(n2436), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[4]), .QN(n4732) );
  DFFNSRX2TS \destinationAddressOut_reg[5]  ( .D(n2435), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[5]), .QN(n4723) );
  DFFNSRX2TS \requesterAddressOut_reg[1]  ( .D(n2433), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[1]), .QN(n4722) );
  DFFNSRX2TS \requesterAddressOut_reg[2]  ( .D(n2432), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[2]), .QN(n4721) );
  DFFNSRX2TS \requesterAddressOut_reg[4]  ( .D(n2430), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[4]), .QN(n4720) );
  DFFNSRX2TS \requesterAddressOut_reg[5]  ( .D(n2429), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(requesterAddressOut[5]), .QN(n4719) );
  DFFNSRX2TS \dataOut_reg[0]  ( .D(n2428), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[0]), .QN(n4710) );
  DFFNSRX2TS \dataOut_reg[1]  ( .D(n2427), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[1]), .QN(n4701) );
  DFFNSRX2TS \dataOut_reg[2]  ( .D(n2426), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[2]), .QN(n4692) );
  DFFNSRX2TS \dataOut_reg[3]  ( .D(n2425), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[3]), .QN(n4683) );
  DFFNSRX2TS \dataOut_reg[4]  ( .D(n2424), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[4]), .QN(n4674) );
  DFFNSRX2TS \dataOut_reg[5]  ( .D(n2423), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[5]), .QN(n4665) );
  DFFNSRX2TS \dataOut_reg[6]  ( .D(n2422), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[6]), .QN(n4656) );
  DFFNSRX2TS \dataOut_reg[7]  ( .D(n2421), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[7]), .QN(n4647) );
  DFFNSRX2TS \dataOut_reg[8]  ( .D(n2420), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[8]), .QN(n4638) );
  DFFNSRX2TS \dataOut_reg[9]  ( .D(n2419), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[9]), .QN(n4629) );
  DFFNSRX2TS \dataOut_reg[10]  ( .D(n2418), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[10]), .QN(n4620) );
  DFFNSRX2TS \dataOut_reg[11]  ( .D(n2417), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[11]), .QN(n4611) );
  DFFNSRX2TS \dataOut_reg[12]  ( .D(n2416), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[12]), .QN(n4602) );
  DFFNSRX2TS \dataOut_reg[13]  ( .D(n2415), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[13]), .QN(n4593) );
  DFFNSRX2TS \dataOut_reg[14]  ( .D(n2414), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[14]), .QN(n4584) );
  DFFNSRX2TS \dataOut_reg[15]  ( .D(n2413), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[15]), .QN(n4575) );
  DFFNSRX2TS \dataOut_reg[16]  ( .D(n2412), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[16]), .QN(n4566) );
  DFFNSRX2TS \dataOut_reg[17]  ( .D(n2411), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[17]), .QN(n4557) );
  DFFNSRX2TS \dataOut_reg[18]  ( .D(n2410), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[18]), .QN(n4548) );
  DFFNSRX2TS \dataOut_reg[19]  ( .D(n2409), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[19]), .QN(n4539) );
  DFFNSRX2TS \dataOut_reg[20]  ( .D(n2408), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[20]), .QN(n4530) );
  DFFNSRX2TS \dataOut_reg[21]  ( .D(n2407), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[21]), .QN(n4521) );
  DFFNSRX2TS \dataOut_reg[22]  ( .D(n2406), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[22]), .QN(n4512) );
  DFFNSRX2TS \dataOut_reg[23]  ( .D(n2405), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[23]), .QN(n4503) );
  DFFNSRX2TS \dataOut_reg[24]  ( .D(n2404), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[24]), .QN(n4494) );
  DFFNSRX2TS \dataOut_reg[25]  ( .D(n2403), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[25]), .QN(n4485) );
  DFFNSRX2TS \dataOut_reg[26]  ( .D(n2402), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[26]), .QN(n4476) );
  DFFNSRX2TS \dataOut_reg[27]  ( .D(n2401), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[27]), .QN(n4467) );
  DFFNSRX2TS \dataOut_reg[28]  ( .D(n2400), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[28]), .QN(n4458) );
  DFFNSRX2TS \dataOut_reg[29]  ( .D(n2399), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[29]), .QN(n4449) );
  DFFNSRX2TS \dataOut_reg[30]  ( .D(n2398), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[30]), .QN(n4440) );
  DFFNSRX2TS \dataOut_reg[31]  ( .D(n2397), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(dataOut[31]), .QN(n4431) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][4]  ( .D(n2558), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n666) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][4]  ( .D(n2530), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n807) );
  DFFNSRXLTS \dataoutbuffer_reg[7][0]  ( .D(n2610), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n609) );
  DFFNSRXLTS \dataoutbuffer_reg[7][1]  ( .D(n2609), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n610) );
  DFFNSRXLTS \dataoutbuffer_reg[7][2]  ( .D(n2608), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n611) );
  DFFNSRXLTS \dataoutbuffer_reg[7][3]  ( .D(n2607), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n612) );
  DFFNSRXLTS \dataoutbuffer_reg[7][4]  ( .D(n2606), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n613) );
  DFFNSRXLTS \dataoutbuffer_reg[7][5]  ( .D(n2605), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n614) );
  DFFNSRXLTS \dataoutbuffer_reg[7][6]  ( .D(n2604), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n615) );
  DFFNSRXLTS \dataoutbuffer_reg[7][7]  ( .D(n2603), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n616) );
  DFFNSRXLTS \dataoutbuffer_reg[7][8]  ( .D(n2602), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n617) );
  DFFNSRXLTS \dataoutbuffer_reg[7][9]  ( .D(n2601), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n618) );
  DFFNSRXLTS \dataoutbuffer_reg[7][10]  ( .D(n2600), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n619) );
  DFFNSRXLTS \dataoutbuffer_reg[7][11]  ( .D(n2599), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n620) );
  DFFNSRXLTS \dataoutbuffer_reg[7][12]  ( .D(n2598), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n621) );
  DFFNSRXLTS \dataoutbuffer_reg[7][13]  ( .D(n2597), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n622) );
  DFFNSRXLTS \dataoutbuffer_reg[7][14]  ( .D(n2596), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n623) );
  DFFNSRXLTS \dataoutbuffer_reg[7][15]  ( .D(n2595), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n624) );
  DFFNSRXLTS \dataoutbuffer_reg[7][16]  ( .D(n2594), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n625) );
  DFFNSRXLTS \dataoutbuffer_reg[7][17]  ( .D(n2593), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n626) );
  DFFNSRXLTS \dataoutbuffer_reg[7][18]  ( .D(n2592), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n627) );
  DFFNSRXLTS \dataoutbuffer_reg[7][19]  ( .D(n2591), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n628) );
  DFFNSRXLTS \dataoutbuffer_reg[7][20]  ( .D(n2590), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n629) );
  DFFNSRXLTS \dataoutbuffer_reg[7][21]  ( .D(n2589), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n630) );
  DFFNSRXLTS \dataoutbuffer_reg[7][22]  ( .D(n2588), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n631) );
  DFFNSRXLTS \dataoutbuffer_reg[7][23]  ( .D(n2587), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n632) );
  DFFNSRXLTS \dataoutbuffer_reg[7][24]  ( .D(n2586), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n633) );
  DFFNSRXLTS \dataoutbuffer_reg[7][25]  ( .D(n2585), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n634) );
  DFFNSRXLTS \dataoutbuffer_reg[7][26]  ( .D(n2584), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n635) );
  DFFNSRXLTS \dataoutbuffer_reg[7][27]  ( .D(n2583), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n636) );
  DFFNSRXLTS \dataoutbuffer_reg[7][28]  ( .D(n2582), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n637) );
  DFFNSRXLTS \dataoutbuffer_reg[7][29]  ( .D(n2581), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n638) );
  DFFNSRXLTS \dataoutbuffer_reg[7][30]  ( .D(n2580), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n639) );
  DFFNSRXLTS \dataoutbuffer_reg[7][31]  ( .D(n2579), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n640) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][1]  ( .D(n2561), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n641) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][2]  ( .D(n2560), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n642) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][3]  ( .D(n2559), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n643) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][5]  ( .D(n2557), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n644) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][0]  ( .D(n2562), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n665) );
  DFFNSRXLTS \requesterAddressbuffer_reg[7][0]  ( .D(n2882), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n684) );
  DFFNSRXLTS \requesterAddressbuffer_reg[7][1]  ( .D(n2881), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n685) );
  DFFNSRXLTS \requesterAddressbuffer_reg[7][3]  ( .D(n2879), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n686) );
  DFFNSRXLTS \requesterAddressbuffer_reg[7][2]  ( .D(n2880), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n687) );
  DFFNSRXLTS \requesterAddressbuffer_reg[7][4]  ( .D(n2878), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n688) );
  DFFNSRXLTS \requesterAddressbuffer_reg[7][5]  ( .D(n2877), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n689) );
  DFFNSRXLTS \requesterAddressbuffer_reg[5][0]  ( .D(n2870), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n888) );
  DFFNSRXLTS \requesterAddressbuffer_reg[5][1]  ( .D(n2869), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n889) );
  DFFNSRXLTS \requesterAddressbuffer_reg[5][2]  ( .D(n2868), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n890) );
  DFFNSRXLTS \requesterAddressbuffer_reg[5][3]  ( .D(n2867), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n891) );
  DFFNSRXLTS \requesterAddressbuffer_reg[5][4]  ( .D(n2866), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n892) );
  DFFNSRXLTS \requesterAddressbuffer_reg[5][5]  ( .D(n2865), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n893) );
  DFFNSRXLTS \readOutbuffer_reg[4]  ( .D(n2567), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n769) );
  DFFNSRXLTS \requesterAddressbuffer_reg[2][2]  ( .D(n2850), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][2] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[2][3]  ( .D(n2849), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][3] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[2][5]  ( .D(n2847), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][5] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[2][0]  ( .D(n2852), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][0] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[2][1]  ( .D(n2851), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][1] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[2][4]  ( .D(n2848), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[2][4] ) );
  DFFNSRXLTS \dataoutbuffer_reg[1][0]  ( .D(n2802), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3092), .QN(n845) );
  DFFNSRXLTS \dataoutbuffer_reg[1][1]  ( .D(n2801), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3091), .QN(n846) );
  DFFNSRXLTS \dataoutbuffer_reg[1][3]  ( .D(n2799), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3089), .QN(n847) );
  DFFNSRXLTS \dataoutbuffer_reg[1][4]  ( .D(n2798), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3088), .QN(n848) );
  DFFNSRXLTS \dataoutbuffer_reg[1][6]  ( .D(n2796), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3086), .QN(n849) );
  DFFNSRXLTS \dataoutbuffer_reg[1][7]  ( .D(n2795), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3085), .QN(n850) );
  DFFNSRXLTS \dataoutbuffer_reg[1][9]  ( .D(n2793), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3083), .QN(n851) );
  DFFNSRXLTS \dataoutbuffer_reg[1][11]  ( .D(n2791), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3081), .QN(n852) );
  DFFNSRXLTS \dataoutbuffer_reg[1][12]  ( .D(n2790), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3080), .QN(n853) );
  DFFNSRXLTS \dataoutbuffer_reg[1][13]  ( .D(n2789), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3079), .QN(n854) );
  DFFNSRXLTS \dataoutbuffer_reg[1][14]  ( .D(n2788), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3078), .QN(n855) );
  DFFNSRXLTS \dataoutbuffer_reg[1][15]  ( .D(n2787), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3077), .QN(n856) );
  DFFNSRXLTS \dataoutbuffer_reg[1][16]  ( .D(n2786), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3076), .QN(n857) );
  DFFNSRXLTS \dataoutbuffer_reg[1][17]  ( .D(n2785), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3075), .QN(n858) );
  DFFNSRXLTS \dataoutbuffer_reg[1][18]  ( .D(n2784), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3074), .QN(n859) );
  DFFNSRXLTS \dataoutbuffer_reg[1][21]  ( .D(n2781), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3071), .QN(n860) );
  DFFNSRXLTS \dataoutbuffer_reg[1][23]  ( .D(n2779), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3069), .QN(n861) );
  DFFNSRXLTS \dataoutbuffer_reg[1][24]  ( .D(n2778), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3068), .QN(n862) );
  DFFNSRXLTS \dataoutbuffer_reg[1][25]  ( .D(n2777), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3067), .QN(n863) );
  DFFNSRXLTS \dataoutbuffer_reg[1][26]  ( .D(n2776), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3066), .QN(n864) );
  DFFNSRXLTS \dataoutbuffer_reg[1][28]  ( .D(n2774), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3064), .QN(n865) );
  DFFNSRXLTS \dataoutbuffer_reg[1][29]  ( .D(n2773), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3063), .QN(n866) );
  DFFNSRXLTS \dataoutbuffer_reg[1][30]  ( .D(n2772), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3062), .QN(n867) );
  DFFNSRXLTS \dataoutbuffer_reg[1][31]  ( .D(n2771), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3061), .QN(n868) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][0]  ( .D(n2478), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3098), .QN(n869) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][1]  ( .D(n2477), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3097), .QN(n870) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][2]  ( .D(n2476), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3096), .QN(n871) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][3]  ( .D(n2475), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3095), .QN(n872) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][5]  ( .D(n2473), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3093), .QN(n873) );
  DFFNSRXLTS \dataoutbuffer_reg[1][2]  ( .D(n2800), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3090), .QN(n874) );
  DFFNSRXLTS \dataoutbuffer_reg[1][5]  ( .D(n2797), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3087), .QN(n875) );
  DFFNSRXLTS \dataoutbuffer_reg[1][8]  ( .D(n2794), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3084), .QN(n876) );
  DFFNSRXLTS \dataoutbuffer_reg[1][10]  ( .D(n2792), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3082), .QN(n877) );
  DFFNSRXLTS \dataoutbuffer_reg[1][19]  ( .D(n2783), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3073), .QN(n878) );
  DFFNSRXLTS \dataoutbuffer_reg[1][20]  ( .D(n2782), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3072), .QN(n879) );
  DFFNSRXLTS \dataoutbuffer_reg[1][22]  ( .D(n2780), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3070), .QN(n880) );
  DFFNSRXLTS \dataoutbuffer_reg[1][27]  ( .D(n2775), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3065), .QN(n881) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][0]  ( .D(n2846), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2963), .QN(n895) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][1]  ( .D(n2845), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2961), .QN(n896) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][2]  ( .D(n2844), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2960), .QN(n897) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][3]  ( .D(n2843), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2962), .QN(n898) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][4]  ( .D(n2842), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2959), .QN(n899) );
  DFFNSRXLTS \requesterAddressbuffer_reg[1][5]  ( .D(n2841), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2958), .QN(n900) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][4]  ( .D(n2474), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3094), .QN(n844) );
  DFFNSRXLTS \readOutbuffer_reg[0]  ( .D(n2563), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n683) );
  DFFNSRXLTS \writeOutbuffer_reg[2]  ( .D(n2573), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n691) );
  DFFNSRXLTS \writeOutbuffer_reg[4]  ( .D(n2575), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n970) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][5]  ( .D(n2543), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3047) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][0]  ( .D(n2548), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3057) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][1]  ( .D(n2547), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3055) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][2]  ( .D(n2546), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3053) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][3]  ( .D(n2545), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3051) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][4]  ( .D(n2544), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3049) );
  DFFNSRXLTS \requesterAddressbuffer_reg[6][1]  ( .D(n2875), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][1] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[6][2]  ( .D(n2874), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][2] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[6][3]  ( .D(n2873), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][3] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[6][4]  ( .D(n2872), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][4] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[6][5]  ( .D(n2871), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][5] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[6][0]  ( .D(n2876), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[6][0] ) );
  DFFNSRXLTS \dataoutbuffer_reg[6][4]  ( .D(n2638), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3037), .QN(n606) );
  DFFNSRXLTS \dataoutbuffer_reg[6][18]  ( .D(n2624), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3009), .QN(n607) );
  DFFNSRXLTS \dataoutbuffer_reg[6][25]  ( .D(n2617), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2995), .QN(n608) );
  DFFNSRXLTS \dataoutbuffer_reg[6][0]  ( .D(n2642), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3045), .QN(n645) );
  DFFNSRXLTS \dataoutbuffer_reg[6][2]  ( .D(n2640), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3041), .QN(n646) );
  DFFNSRXLTS \dataoutbuffer_reg[6][3]  ( .D(n2639), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3039), .QN(n647) );
  DFFNSRXLTS \dataoutbuffer_reg[6][5]  ( .D(n2637), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3035), .QN(n648) );
  DFFNSRXLTS \dataoutbuffer_reg[6][7]  ( .D(n2635), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3031), .QN(n649) );
  DFFNSRXLTS \dataoutbuffer_reg[6][8]  ( .D(n2634), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3029), .QN(n650) );
  DFFNSRXLTS \dataoutbuffer_reg[6][9]  ( .D(n2633), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3027), .QN(n651) );
  DFFNSRXLTS \dataoutbuffer_reg[6][11]  ( .D(n2631), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3023), .QN(n652) );
  DFFNSRXLTS \dataoutbuffer_reg[6][14]  ( .D(n2628), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3017), .QN(n653) );
  DFFNSRXLTS \dataoutbuffer_reg[6][15]  ( .D(n2627), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3015), .QN(n654) );
  DFFNSRXLTS \dataoutbuffer_reg[6][16]  ( .D(n2626), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3013), .QN(n655) );
  DFFNSRXLTS \dataoutbuffer_reg[6][17]  ( .D(n2625), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3011), .QN(n656) );
  DFFNSRXLTS \dataoutbuffer_reg[6][19]  ( .D(n2623), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3007), .QN(n657) );
  DFFNSRXLTS \dataoutbuffer_reg[6][22]  ( .D(n2620), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3001), .QN(n658) );
  DFFNSRXLTS \dataoutbuffer_reg[6][24]  ( .D(n2618), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2997), .QN(n659) );
  DFFNSRXLTS \dataoutbuffer_reg[6][26]  ( .D(n2616), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2993), .QN(n660) );
  DFFNSRXLTS \dataoutbuffer_reg[6][27]  ( .D(n2615), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2991), .QN(n661) );
  DFFNSRXLTS \dataoutbuffer_reg[6][28]  ( .D(n2614), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2989), .QN(n662) );
  DFFNSRXLTS \dataoutbuffer_reg[6][30]  ( .D(n2612), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2985), .QN(n663) );
  DFFNSRXLTS \dataoutbuffer_reg[6][31]  ( .D(n2611), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2983), .QN(n664) );
  DFFNSRXLTS \dataoutbuffer_reg[6][1]  ( .D(n2641), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3043), .QN(n667) );
  DFFNSRXLTS \dataoutbuffer_reg[6][6]  ( .D(n2636), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3033), .QN(n668) );
  DFFNSRXLTS \dataoutbuffer_reg[6][10]  ( .D(n2632), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3025), .QN(n669) );
  DFFNSRXLTS \dataoutbuffer_reg[6][12]  ( .D(n2630), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3021), .QN(n670) );
  DFFNSRXLTS \dataoutbuffer_reg[6][13]  ( .D(n2629), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3019), .QN(n671) );
  DFFNSRXLTS \dataoutbuffer_reg[6][20]  ( .D(n2622), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3005), .QN(n672) );
  DFFNSRXLTS \dataoutbuffer_reg[6][21]  ( .D(n2621), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3003), .QN(n673) );
  DFFNSRXLTS \dataoutbuffer_reg[6][23]  ( .D(n2619), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2999), .QN(n674) );
  DFFNSRXLTS \dataoutbuffer_reg[6][29]  ( .D(n2613), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2987), .QN(n675) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][13]  ( .D(n2479), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3240), .QN(n565) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][13]  ( .D(n2507), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3186), .QN(n582) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][13]  ( .D(n2465), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3178), .QN(n597) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][6]  ( .D(n2486), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3233), .QN(n552) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][8]  ( .D(n2484), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3235), .QN(n553) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][10]  ( .D(n2482), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3237), .QN(n554) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][12]  ( .D(n2480), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3239), .QN(n555) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][7]  ( .D(n2485), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3234), .QN(n559) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][9]  ( .D(n2483), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3236), .QN(n560) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][11]  ( .D(n2481), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3238), .QN(n561) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][9]  ( .D(n2511), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3190), .QN(n581) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][10]  ( .D(n2510), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3189), .QN(n603) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][11]  ( .D(n2509), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3188), .QN(n604) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][12]  ( .D(n2508), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3187), .QN(n605) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][8]  ( .D(n2512), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3191), .QN(n967) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][7]  ( .D(n2513), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3192), .QN(n968) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][6]  ( .D(n2514), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3193), .QN(n969) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][1]  ( .D(n2491), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n718) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][0]  ( .D(n2492), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n717) );
  DFFNSRXLTS \dataoutbuffer_reg[2][31]  ( .D(n2739), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n697) );
  DFFNSRXLTS \dataoutbuffer_reg[2][30]  ( .D(n2740), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n752) );
  DFFNSRXLTS \dataoutbuffer_reg[2][29]  ( .D(n2741), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n949) );
  DFFNSRXLTS \dataoutbuffer_reg[2][28]  ( .D(n2742), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n950) );
  DFFNSRXLTS \dataoutbuffer_reg[2][27]  ( .D(n2743), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n964) );
  DFFNSRXLTS \dataoutbuffer_reg[2][26]  ( .D(n2744), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n951) );
  DFFNSRXLTS \dataoutbuffer_reg[2][25]  ( .D(n2745), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n952) );
  DFFNSRXLTS \dataoutbuffer_reg[2][24]  ( .D(n2746), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n696) );
  DFFNSRXLTS \dataoutbuffer_reg[2][23]  ( .D(n2747), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n953) );
  DFFNSRXLTS \dataoutbuffer_reg[2][22]  ( .D(n2748), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n695) );
  DFFNSRXLTS \dataoutbuffer_reg[2][21]  ( .D(n2749), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n954) );
  DFFNSRXLTS \dataoutbuffer_reg[2][20]  ( .D(n2750), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n955) );
  DFFNSRXLTS \dataoutbuffer_reg[2][19]  ( .D(n2751), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n956) );
  DFFNSRXLTS \dataoutbuffer_reg[2][18]  ( .D(n2752), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n957) );
  DFFNSRXLTS \dataoutbuffer_reg[2][17]  ( .D(n2753), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n751) );
  DFFNSRXLTS \dataoutbuffer_reg[2][16]  ( .D(n2754), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n694) );
  DFFNSRXLTS \dataoutbuffer_reg[2][15]  ( .D(n2755), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n750) );
  DFFNSRXLTS \dataoutbuffer_reg[2][14]  ( .D(n2756), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n749) );
  DFFNSRXLTS \dataoutbuffer_reg[2][13]  ( .D(n2757), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n958) );
  DFFNSRXLTS \dataoutbuffer_reg[2][12]  ( .D(n2758), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n959) );
  DFFNSRXLTS \dataoutbuffer_reg[2][11]  ( .D(n2759), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n960) );
  DFFNSRXLTS \dataoutbuffer_reg[2][10]  ( .D(n2760), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n965) );
  DFFNSRXLTS \dataoutbuffer_reg[2][9]  ( .D(n2761), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n961) );
  DFFNSRXLTS \dataoutbuffer_reg[2][8]  ( .D(n2762), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n962) );
  DFFNSRXLTS \dataoutbuffer_reg[2][7]  ( .D(n2763), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n963) );
  DFFNSRXLTS \dataoutbuffer_reg[2][6]  ( .D(n2764), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n966) );
  DFFNSRXLTS \dataoutbuffer_reg[2][5]  ( .D(n2765), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n748) );
  DFFNSRXLTS \dataoutbuffer_reg[2][4]  ( .D(n2766), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n747) );
  DFFNSRXLTS \dataoutbuffer_reg[2][3]  ( .D(n2767), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n746) );
  DFFNSRXLTS \dataoutbuffer_reg[2][2]  ( .D(n2768), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n693) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][5]  ( .D(n2487), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n946) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][4]  ( .D(n2488), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n947) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][3]  ( .D(n2489), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n948) );
  DFFNSRXLTS \destinationAddressbuffer_reg[2][2]  ( .D(n2490), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n945) );
  DFFNSRXLTS \dataoutbuffer_reg[2][1]  ( .D(n2769), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n943) );
  DFFNSRXLTS \dataoutbuffer_reg[2][0]  ( .D(n2770), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n944) );
  DFFNSRXLTS \write_reg_reg[1]  ( .D(n2887), .CKN(clk), .SN(1'b1), .RN(1'b1), 
        .Q(n469), .QN(n5323) );
  DFFNSRXLTS \requesterAddressbuffer_reg[0][3]  ( .D(n2837), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][3] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[0][2]  ( .D(n2838), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][2] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[0][0]  ( .D(n2840), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][0] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[0][1]  ( .D(n2839), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][1] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[0][5]  ( .D(n2835), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][5] ) );
  DFFNSRXLTS \requesterAddressbuffer_reg[0][4]  ( .D(n2836), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[0][4] ) );
  DFFNSRXLTS \destinationAddressOut_reg[7]  ( .D(n2447), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[7]) );
  DFFNSRXLTS \destinationAddressOut_reg[6]  ( .D(n2448), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[6]) );
  DFFNSRXLTS \destinationAddressOut_reg[13]  ( .D(n2441), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[13]) );
  DFFNSRXLTS \destinationAddressOut_reg[12]  ( .D(n2442), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[12]) );
  DFFNSRXLTS \destinationAddressOut_reg[11]  ( .D(n2443), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[11]) );
  DFFNSRXLTS \destinationAddressOut_reg[10]  ( .D(n2444), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[10]) );
  DFFNSRXLTS \destinationAddressOut_reg[9]  ( .D(n2445), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[9]) );
  DFFNSRXLTS \destinationAddressOut_reg[8]  ( .D(n2446), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(destinationAddressOut[8]) );
  DFFNSRXLTS \readOutbuffer_reg[7]  ( .D(n2570), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(readOutbuffer_7) );
  DFFNSRXLTS \readOutbuffer_reg[5]  ( .D(n2568), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n681) );
  DFFNSRXLTS \readOutbuffer_reg[6]  ( .D(n2569), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n677) );
  DFFNSRXLTS \readOutbuffer_reg[3]  ( .D(n2566), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n676) );
  DFFNSRXLTS \readOutbuffer_reg[1]  ( .D(n2564), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n682) );
  DFFNSRXLTS \readOutbuffer_reg[2]  ( .D(n2565), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(\readOutbuffer[2] ), .QN(n768) );
  DFFNSRXLTS full_reg_reg ( .D(N4718), .CKN(clk), .SN(1'b1), .RN(1'b1), .Q(
        n4844), .QN(n781) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][13]  ( .D(n2535), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3210), .QN(n580) );
  DFFNSRXLTS \writeOutbuffer_reg[5]  ( .D(n2576), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3177), .QN(n894) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][13]  ( .D(n2521), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3194), .QN(n910) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][12]  ( .D(n2522), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3196), .QN(n906) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][11]  ( .D(n2523), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3198), .QN(n905) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][10]  ( .D(n2524), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3200), .QN(n806) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][9]  ( .D(n2525), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3201), .QN(n904) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][8]  ( .D(n2526), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3203), .QN(n903) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][7]  ( .D(n2527), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3205), .QN(n902) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][6]  ( .D(n2528), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3207), .QN(n901) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][5]  ( .D(n2529), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n909) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][3]  ( .D(n2531), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n838) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][2]  ( .D(n2532), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n837) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][1]  ( .D(n2533), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n836) );
  DFFNSRXLTS \destinationAddressbuffer_reg[5][0]  ( .D(n2534), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .QN(n835) );
  DFFNSRXLTS \dataoutbuffer_reg[5][31]  ( .D(n2643), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n843) );
  DFFNSRXLTS \dataoutbuffer_reg[5][30]  ( .D(n2644), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n834) );
  DFFNSRXLTS \dataoutbuffer_reg[5][29]  ( .D(n2645), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n833) );
  DFFNSRXLTS \dataoutbuffer_reg[5][28]  ( .D(n2646), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n832) );
  DFFNSRXLTS \dataoutbuffer_reg[5][27]  ( .D(n2647), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n831) );
  DFFNSRXLTS \dataoutbuffer_reg[5][26]  ( .D(n2648), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n830) );
  DFFNSRXLTS \dataoutbuffer_reg[5][25]  ( .D(n2649), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n829) );
  DFFNSRXLTS \dataoutbuffer_reg[5][24]  ( .D(n2650), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n828) );
  DFFNSRXLTS \dataoutbuffer_reg[5][23]  ( .D(n2651), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n827) );
  DFFNSRXLTS \dataoutbuffer_reg[5][22]  ( .D(n2652), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n826) );
  DFFNSRXLTS \dataoutbuffer_reg[5][21]  ( .D(n2653), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n825) );
  DFFNSRXLTS \dataoutbuffer_reg[5][20]  ( .D(n2654), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n824) );
  DFFNSRXLTS \dataoutbuffer_reg[5][19]  ( .D(n2655), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n823) );
  DFFNSRXLTS \dataoutbuffer_reg[5][18]  ( .D(n2656), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n822) );
  DFFNSRXLTS \dataoutbuffer_reg[5][17]  ( .D(n2657), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n821) );
  DFFNSRXLTS \dataoutbuffer_reg[5][16]  ( .D(n2658), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n842) );
  DFFNSRXLTS \dataoutbuffer_reg[5][15]  ( .D(n2659), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n841) );
  DFFNSRXLTS \dataoutbuffer_reg[5][14]  ( .D(n2660), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n820) );
  DFFNSRXLTS \dataoutbuffer_reg[5][13]  ( .D(n2661), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n819) );
  DFFNSRXLTS \dataoutbuffer_reg[5][12]  ( .D(n2662), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n818) );
  DFFNSRXLTS \dataoutbuffer_reg[5][11]  ( .D(n2663), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n840) );
  DFFNSRXLTS \dataoutbuffer_reg[5][10]  ( .D(n2664), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .QN(n817) );
  DFFNSRXLTS \dataoutbuffer_reg[5][9]  ( .D(n2665), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n816) );
  DFFNSRXLTS \dataoutbuffer_reg[5][8]  ( .D(n2666), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n815) );
  DFFNSRXLTS \dataoutbuffer_reg[5][7]  ( .D(n2667), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n814) );
  DFFNSRXLTS \dataoutbuffer_reg[5][6]  ( .D(n2668), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n813) );
  DFFNSRXLTS \dataoutbuffer_reg[5][5]  ( .D(n2669), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n812) );
  DFFNSRXLTS \dataoutbuffer_reg[5][4]  ( .D(n2670), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n811) );
  DFFNSRXLTS \dataoutbuffer_reg[5][3]  ( .D(n2671), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n810) );
  DFFNSRXLTS \dataoutbuffer_reg[5][2]  ( .D(n2672), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n809) );
  DFFNSRXLTS \dataoutbuffer_reg[5][1]  ( .D(n2673), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n839) );
  DFFNSRXLTS \dataoutbuffer_reg[5][0]  ( .D(n2674), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n808) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][5]  ( .D(n2853), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][5] ), .QN(n886) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][4]  ( .D(n2854), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][4] ), .QN(n887) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][3]  ( .D(n2855), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][3] ), .QN(n885) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][2]  ( .D(n2856), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][2] ), .QN(n884) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][1]  ( .D(n2857), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][1] ), .QN(n883) );
  DFFNSRXLTS \requesterAddressbuffer_reg[3][0]  ( .D(n2858), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(\requesterAddressbuffer[3][0] ), .QN(n882) );
  DFFNSRXLTS \dataoutbuffer_reg[3][1]  ( .D(n2737), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n86), .QN(n720) );
  DFFNSRXLTS \dataoutbuffer_reg[3][0]  ( .D(n2738), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n87), .QN(n719) );
  DFFNSRXLTS \requesterAddressbuffer_reg[4][3]  ( .D(n2861), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2980) );
  DFFNSRXLTS \requesterAddressbuffer_reg[4][2]  ( .D(n2862), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2978) );
  DFFNSRXLTS \requesterAddressbuffer_reg[4][1]  ( .D(n2863), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2979) );
  DFFNSRXLTS \requesterAddressbuffer_reg[4][0]  ( .D(n2864), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2981) );
  DFFNSRXLTS \requesterAddressbuffer_reg[4][5]  ( .D(n2859), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2976) );
  DFFNSRXLTS \requesterAddressbuffer_reg[4][4]  ( .D(n2860), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n2977) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][13]  ( .D(n2451), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3232), .QN(n564) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][5]  ( .D(n2501), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n61), .QN(n745) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][4]  ( .D(n2502), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n62), .QN(n744) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][3]  ( .D(n2503), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n63), .QN(n743) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][2]  ( .D(n2504), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n90), .QN(n716) );
  DFFNSRXLTS \writeOutbuffer_reg[7]  ( .D(n2578), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3176), .QN(n678) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][13]  ( .D(n2549), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3195), .QN(n589) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][12]  ( .D(n2550), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3197), .QN(n588) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][11]  ( .D(n2551), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3199), .QN(n587) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][10]  ( .D(n2552), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n567), .QN(n586) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][9]  ( .D(n2553), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3202), .QN(n598) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][8]  ( .D(n2554), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3204), .QN(n585) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][7]  ( .D(n2555), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3206), .QN(n584) );
  DFFNSRXLTS \destinationAddressbuffer_reg[7][6]  ( .D(n2556), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3208), .QN(n583) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][12]  ( .D(n2466), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3179), .QN(n596) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][11]  ( .D(n2467), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3180), .QN(n595) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][10]  ( .D(n2468), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3181), .QN(n594) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][9]  ( .D(n2469), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3182), .QN(n593) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][1]  ( .D(n2505), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n64), .QN(n742) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][0]  ( .D(n2506), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n65), .QN(n741) );
  DFFNSRXLTS \dataoutbuffer_reg[3][31]  ( .D(n2707), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n66), .QN(n740) );
  DFFNSRXLTS \dataoutbuffer_reg[3][30]  ( .D(n2708), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n67), .QN(n739) );
  DFFNSRXLTS \dataoutbuffer_reg[3][29]  ( .D(n2709), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n68), .QN(n738) );
  DFFNSRXLTS \dataoutbuffer_reg[3][28]  ( .D(n2710), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n69), .QN(n737) );
  DFFNSRXLTS \dataoutbuffer_reg[3][27]  ( .D(n2711), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n70), .QN(n736) );
  DFFNSRXLTS \dataoutbuffer_reg[3][26]  ( .D(n2712), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n71), .QN(n735) );
  DFFNSRXLTS \dataoutbuffer_reg[3][25]  ( .D(n2713), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n91), .QN(n715) );
  DFFNSRXLTS \dataoutbuffer_reg[3][24]  ( .D(n2714), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n72), .QN(n734) );
  DFFNSRXLTS \dataoutbuffer_reg[3][23]  ( .D(n2715), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n92), .QN(n714) );
  DFFNSRXLTS \dataoutbuffer_reg[3][22]  ( .D(n2716), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n73), .QN(n733) );
  DFFNSRXLTS \dataoutbuffer_reg[3][21]  ( .D(n2717), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n74), .QN(n732) );
  DFFNSRXLTS \dataoutbuffer_reg[3][20]  ( .D(n2718), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n93), .QN(n713) );
  DFFNSRXLTS \dataoutbuffer_reg[3][19]  ( .D(n2719), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n75), .QN(n731) );
  DFFNSRXLTS \dataoutbuffer_reg[3][18]  ( .D(n2720), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n94), .QN(n712) );
  DFFNSRXLTS \dataoutbuffer_reg[3][17]  ( .D(n2721), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n76), .QN(n730) );
  DFFNSRXLTS \dataoutbuffer_reg[3][16]  ( .D(n2722), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n77), .QN(n729) );
  DFFNSRXLTS \dataoutbuffer_reg[3][15]  ( .D(n2723), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n95), .QN(n711) );
  DFFNSRXLTS \dataoutbuffer_reg[3][14]  ( .D(n2724), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n78), .QN(n728) );
  DFFNSRXLTS \dataoutbuffer_reg[3][13]  ( .D(n2725), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n96), .QN(n710) );
  DFFNSRXLTS \dataoutbuffer_reg[3][12]  ( .D(n2726), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n79), .QN(n727) );
  DFFNSRXLTS \dataoutbuffer_reg[3][11]  ( .D(n2727), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n80), .QN(n726) );
  DFFNSRXLTS \dataoutbuffer_reg[3][10]  ( .D(n2728), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n81), .QN(n725) );
  DFFNSRXLTS \dataoutbuffer_reg[3][9]  ( .D(n2729), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n82), .QN(n724) );
  DFFNSRXLTS \dataoutbuffer_reg[3][8]  ( .D(n2730), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n83), .QN(n723) );
  DFFNSRXLTS \dataoutbuffer_reg[3][6]  ( .D(n2732), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n84), .QN(n722) );
  DFFNSRXLTS \dataoutbuffer_reg[3][5]  ( .D(n2733), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n97), .QN(n709) );
  DFFNSRXLTS \dataoutbuffer_reg[3][4]  ( .D(n2734), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n98), .QN(n708) );
  DFFNSRXLTS \dataoutbuffer_reg[3][3]  ( .D(n2735), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n85), .QN(n721) );
  DFFNSRXLTS \dataoutbuffer_reg[3][2]  ( .D(n2736), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n99), .QN(n707) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][1]  ( .D(n2519), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3054) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][0]  ( .D(n2520), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3056) );
  DFFNSRXLTS \dataoutbuffer_reg[4][31]  ( .D(n2675), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2982) );
  DFFNSRXLTS \dataoutbuffer_reg[4][30]  ( .D(n2676), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2984) );
  DFFNSRXLTS \dataoutbuffer_reg[4][29]  ( .D(n2677), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2986) );
  DFFNSRXLTS \dataoutbuffer_reg[4][28]  ( .D(n2678), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2988) );
  DFFNSRXLTS \dataoutbuffer_reg[4][27]  ( .D(n2679), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2990) );
  DFFNSRXLTS \dataoutbuffer_reg[4][26]  ( .D(n2680), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2992) );
  DFFNSRXLTS \dataoutbuffer_reg[4][25]  ( .D(n2681), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2994) );
  DFFNSRXLTS \dataoutbuffer_reg[4][24]  ( .D(n2682), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2996) );
  DFFNSRXLTS \dataoutbuffer_reg[4][23]  ( .D(n2683), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n2998) );
  DFFNSRXLTS \dataoutbuffer_reg[4][22]  ( .D(n2684), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3000) );
  DFFNSRXLTS \dataoutbuffer_reg[4][21]  ( .D(n2685), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3002) );
  DFFNSRXLTS \dataoutbuffer_reg[4][20]  ( .D(n2686), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3004) );
  DFFNSRXLTS \dataoutbuffer_reg[4][19]  ( .D(n2687), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3006) );
  DFFNSRXLTS \dataoutbuffer_reg[4][18]  ( .D(n2688), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3008) );
  DFFNSRXLTS \dataoutbuffer_reg[4][17]  ( .D(n2689), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3010) );
  DFFNSRXLTS \dataoutbuffer_reg[4][16]  ( .D(n2690), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3012) );
  DFFNSRXLTS \dataoutbuffer_reg[4][15]  ( .D(n2691), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3014) );
  DFFNSRXLTS \dataoutbuffer_reg[4][14]  ( .D(n2692), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3016) );
  DFFNSRXLTS \dataoutbuffer_reg[4][13]  ( .D(n2693), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3018) );
  DFFNSRXLTS \dataoutbuffer_reg[4][12]  ( .D(n2694), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3020) );
  DFFNSRXLTS \dataoutbuffer_reg[4][11]  ( .D(n2695), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3022) );
  DFFNSRXLTS \dataoutbuffer_reg[4][10]  ( .D(n2696), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n3024) );
  DFFNSRXLTS \dataoutbuffer_reg[4][9]  ( .D(n2697), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3026) );
  DFFNSRXLTS \dataoutbuffer_reg[4][8]  ( .D(n2698), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3028) );
  DFFNSRXLTS \dataoutbuffer_reg[4][7]  ( .D(n2699), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3030) );
  DFFNSRXLTS \dataoutbuffer_reg[4][6]  ( .D(n2700), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3032) );
  DFFNSRXLTS \dataoutbuffer_reg[4][5]  ( .D(n2701), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3034) );
  DFFNSRXLTS \dataoutbuffer_reg[4][4]  ( .D(n2702), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3036) );
  DFFNSRXLTS \dataoutbuffer_reg[4][3]  ( .D(n2703), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3038) );
  DFFNSRXLTS \dataoutbuffer_reg[4][2]  ( .D(n2704), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3040) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][5]  ( .D(n2515), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3046) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][4]  ( .D(n2516), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3048) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][3]  ( .D(n2517), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3050) );
  DFFNSRXLTS \destinationAddressbuffer_reg[4][2]  ( .D(n2518), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3052) );
  DFFNSRXLTS \dataoutbuffer_reg[4][1]  ( .D(n2705), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3042) );
  DFFNSRXLTS \dataoutbuffer_reg[4][0]  ( .D(n2706), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n3044) );
  DFFNSRXLTS \writeOutbuffer_reg[1]  ( .D(n2572), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n690) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][8]  ( .D(n2470), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3183), .QN(n592) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][7]  ( .D(n2471), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3184), .QN(n591) );
  DFFNSRXLTS \destinationAddressbuffer_reg[1][6]  ( .D(n2472), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3185), .QN(n590) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][12]  ( .D(n2452), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3231), .QN(n568) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][11]  ( .D(n2453), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3230), .QN(n558) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][10]  ( .D(n2454), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3229), .QN(n563) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][9]  ( .D(n2455), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3228), .QN(n557) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][13]  ( .D(n2493), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3209), .QN(n571) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][12]  ( .D(n2494), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3211), .QN(n574) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][11]  ( .D(n2495), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3213), .QN(n576) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][10]  ( .D(n2496), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3215), .QN(n570) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][9]  ( .D(n2497), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3217), .QN(n573) );
  DFFNSRXLTS \writeOutbuffer_reg[0]  ( .D(n2571), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n765) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][8]  ( .D(n2456), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3227), .QN(n566) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][7]  ( .D(n2457), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3226), .QN(n556) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][6]  ( .D(n2458), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3225), .QN(n562) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][11]  ( .D(n2537), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3214), .QN(n579) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][9]  ( .D(n2539), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3218), .QN(n600) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][7]  ( .D(n2541), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3222), .QN(n577) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][6]  ( .D(n2542), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3224), .QN(n599) );
  DFFNSRXLTS \writeOutbuffer_reg[6]  ( .D(n2577), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n767) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][12]  ( .D(n2536), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3212), .QN(n602) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][10]  ( .D(n2538), .CKN(clk), 
        .SN(1'b1), .RN(1'b1), .Q(n3216), .QN(n601) );
  DFFNSRXLTS \destinationAddressbuffer_reg[6][8]  ( .D(n2540), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3220), .QN(n578) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][0]  ( .D(n2464), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n89) );
  DFFNSRXLTS \dataoutbuffer_reg[0][19]  ( .D(n2815), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n46) );
  DFFNSRXLTS \dataoutbuffer_reg[0][18]  ( .D(n2816), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n47) );
  DFFNSRXLTS \dataoutbuffer_reg[0][17]  ( .D(n2817), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n48) );
  DFFNSRXLTS \dataoutbuffer_reg[0][16]  ( .D(n2818), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n49) );
  DFFNSRXLTS \dataoutbuffer_reg[0][15]  ( .D(n2819), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n50) );
  DFFNSRXLTS \dataoutbuffer_reg[0][14]  ( .D(n2820), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n51) );
  DFFNSRXLTS \dataoutbuffer_reg[0][13]  ( .D(n2821), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n52) );
  DFFNSRXLTS \dataoutbuffer_reg[0][12]  ( .D(n2822), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n53) );
  DFFNSRXLTS \dataoutbuffer_reg[0][11]  ( .D(n2823), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n54) );
  DFFNSRXLTS \dataoutbuffer_reg[0][10]  ( .D(n2824), .CKN(clk), .SN(1'b1), 
        .RN(1'b1), .Q(n55) );
  DFFNSRXLTS \dataoutbuffer_reg[0][8]  ( .D(n2826), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n56) );
  DFFNSRXLTS \dataoutbuffer_reg[0][7]  ( .D(n2827), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n57) );
  DFFNSRXLTS \dataoutbuffer_reg[0][6]  ( .D(n2828), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n58) );
  DFFNSRXLTS \dataoutbuffer_reg[0][4]  ( .D(n2830), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n59) );
  DFFNSRXLTS \dataoutbuffer_reg[0][3]  ( .D(n2831), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .Q(n60) );
  DFFNSRXLTS \destinationAddressbuffer_reg[0][4]  ( .D(n2460), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n88) );
  DFFNSRXLTS \writeOutbuffer_reg[3]  ( .D(n2574), .CKN(clk), .SN(1'b1), .RN(
        1'b1), .QN(n766) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][8]  ( .D(n2498), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3219), .QN(n572) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][7]  ( .D(n2499), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3221), .QN(n569) );
  DFFNSRXLTS \destinationAddressbuffer_reg[3][6]  ( .D(n2500), .CKN(clk), .SN(
        1'b1), .RN(1'b1), .Q(n3223), .QN(n575) );
  NOR2BXLTS U2 ( .AN(n1822), .B(n1823), .Y(n1169) );
  INVX1TS U3 ( .A(n1823), .Y(n802) );
  NAND3X4TS U4 ( .A(n109), .B(n156), .C(n935), .Y(n1816) );
  INVX2TS U5 ( .A(n2064), .Y(n109) );
  XOR2X4TS U6 ( .A(n2057), .B(n5326), .Y(n1942) );
  OAI32X2TS U7 ( .A0(n2058), .A1(n986), .A2(n973), .B0(n157), .B1(n2059), .Y(
        n2057) );
  CLKBUFX2TS U8 ( .A(n3429), .Y(n3428) );
  NOR2BX1TS U9 ( .AN(n1893), .B(n1851), .Y(n1820) );
  NOR3X2TS U10 ( .A(n1820), .B(n1822), .C(n923), .Y(n1821) );
  CLKBUFX2TS U11 ( .A(n3138), .Y(n3136) );
  AOI2BB1X1TS U12 ( .A0N(n935), .A1N(n1963), .B0(n1866), .Y(n1864) );
  CLKINVX2TS U13 ( .A(n1800), .Y(n790) );
  AND3X2TS U14 ( .A(n1842), .B(n1843), .C(n1839), .Y(n1218) );
  NAND3X1TS U15 ( .A(n1895), .B(n1894), .C(n1942), .Y(n1843) );
  NAND2X1TS U16 ( .A(n2065), .B(n488), .Y(n2064) );
  AOI2BB1X1TS U17 ( .A0N(n2925), .A1N(n927), .B0(n2957), .Y(n2059) );
  AOI21X1TS U18 ( .A0(n916), .A1(n940), .B0(n3818), .Y(n1847) );
  CLKBUFX2TS U19 ( .A(n1219), .Y(n3418) );
  XOR2X1TS U20 ( .A(n2060), .B(n2061), .Y(n2011) );
  CLKBUFX2TS U21 ( .A(n1169), .Y(n3648) );
  NAND2X1TS U22 ( .A(n1816), .B(n2063), .Y(n1964) );
  OAI21X1TS U23 ( .A0(n1986), .A1(n103), .B0(n1977), .Y(n1800) );
  OA21XLTS U24 ( .A0(n1987), .A1(n1964), .B0(n1844), .Y(n1986) );
  CLKBUFX2TS U25 ( .A(n1151), .Y(n3730) );
  AND2X2TS U26 ( .A(n2011), .B(selectBit_WEST), .Y(n1941) );
  CLKBUFX2TS U27 ( .A(n3745), .Y(n3744) );
  CLKBUFX2TS U28 ( .A(n3616), .Y(n3613) );
  CLKBUFX2TS U29 ( .A(n1249), .Y(n3312) );
  AOI21X1TS U30 ( .A0(n916), .A1(n938), .B0(n797), .Y(n1831) );
  CLKBUFX2TS U31 ( .A(n3534), .Y(n3528) );
  CLKBUFX2TS U32 ( .A(n3582), .Y(n3576) );
  CLKBUFX2TS U33 ( .A(n3874), .Y(n3873) );
  CLKBUFX2TS U34 ( .A(n3773), .Y(n3769) );
  CLKBUFX2TS U35 ( .A(n3314), .Y(n3311) );
  CLKBUFX2TS U36 ( .A(n3673), .Y(n3672) );
  CLKBUFX2TS U37 ( .A(n3884), .Y(n3883) );
  CLKBUFX2TS U38 ( .A(n3551), .Y(n3544) );
  OAI221XLTS U39 ( .A0(n942), .A1(n929), .B0(n1851), .B1(n2010), .C0(n1853), 
        .Y(n1852) );
  NAND2X1TS U40 ( .A(n1834), .B(n1831), .Y(n1796) );
  CLKBUFX2TS U41 ( .A(n3547), .Y(n3537) );
  CLKBUFX2TS U42 ( .A(n3547), .Y(n3538) );
  AOI222XLTS U43 ( .A0(n4247), .A1(n3639), .B0(n4022), .B1(n3614), .C0(n3985), 
        .C1(n3771), .Y(n1916) );
  OAI221XLTS U44 ( .A0(n1802), .A1(n144), .B0(n162), .B1(n561), .C0(n2007), 
        .Y(n2481) );
  OAI221XLTS U45 ( .A0(n183), .A1(n146), .B0(n161), .B1(n560), .C0(n2005), .Y(
        n2483) );
  OAI221XLTS U46 ( .A0(n182), .A1(n137), .B0(n162), .B1(n559), .C0(n2003), .Y(
        n2485) );
  OAI221XLTS U47 ( .A0(n183), .A1(n148), .B0(n161), .B1(n555), .C0(n2008), .Y(
        n2480) );
  OAI221XLTS U48 ( .A0(n183), .A1(n160), .B0(n161), .B1(n691), .C0(n1804), .Y(
        n2573) );
  INVX2TS U49 ( .A(n115), .Y(n116) );
  NOR2BXLTS U50 ( .AN(n117), .B(n1989), .Y(n1827) );
  CLKINVX2TS U51 ( .A(n1860), .Y(n125) );
  INVX2TS U52 ( .A(n1892), .Y(n103) );
  AND2X2TS U53 ( .A(n986), .B(n1892), .Y(n2) );
  CLKBUFX2TS U54 ( .A(n801), .Y(n3774) );
  INVX2TS U55 ( .A(n1808), .Y(n163) );
  OAI22X1TS U56 ( .A0(n1864), .A1(n803), .B0(n105), .B1(n120), .Y(n1808) );
  NAND2X1TS U57 ( .A(n934), .B(n5323), .Y(n1860) );
  AND3X2TS U58 ( .A(n1824), .B(n126), .C(n1829), .Y(n5) );
  XNOR2X1TS U59 ( .A(n107), .B(n979), .Y(n6) );
  INVX2TS U60 ( .A(n1894), .Y(n926) );
  OAI22X1TS U61 ( .A0(n919), .A1(n103), .B0(n106), .B1(n1987), .Y(n1803) );
  AND2X2TS U62 ( .A(n2066), .B(n120), .Y(n7) );
  INVX1TS U63 ( .A(n1802), .Y(n181) );
  NAND2X1TS U64 ( .A(n919), .B(n1847), .Y(n1802) );
  CLKINVX2TS U65 ( .A(n181), .Y(n182) );
  CLKINVX2TS U66 ( .A(n174), .Y(n175) );
  AND2X2TS U67 ( .A(n6257), .B(n4572), .Y(n10) );
  AND2X2TS U68 ( .A(n459), .B(n4572), .Y(n11) );
  OR2X2TS U69 ( .A(n1143), .B(n8), .Y(n12) );
  INVXLTS U70 ( .A(readRequesterAddress[0]), .Y(n13) );
  INVXLTS U71 ( .A(n13), .Y(n14) );
  INVXLTS U72 ( .A(n13), .Y(n15) );
  INVXLTS U73 ( .A(n13), .Y(n16) );
  INVXLTS U74 ( .A(n13), .Y(n17) );
  INVXLTS U75 ( .A(readRequesterAddress[1]), .Y(n18) );
  INVXLTS U76 ( .A(n18), .Y(n19) );
  INVXLTS U77 ( .A(n18), .Y(n20) );
  INVXLTS U78 ( .A(n18), .Y(n21) );
  INVXLTS U79 ( .A(n18), .Y(n22) );
  INVXLTS U80 ( .A(readRequesterAddress[2]), .Y(n23) );
  INVXLTS U81 ( .A(n23), .Y(n24) );
  INVXLTS U82 ( .A(n23), .Y(n25) );
  INVXLTS U83 ( .A(n23), .Y(n26) );
  INVXLTS U84 ( .A(n23), .Y(n27) );
  INVXLTS U85 ( .A(readRequesterAddress[3]), .Y(n28) );
  INVXLTS U86 ( .A(n28), .Y(n29) );
  INVXLTS U87 ( .A(n28), .Y(n30) );
  INVXLTS U88 ( .A(n28), .Y(n31) );
  INVXLTS U89 ( .A(n28), .Y(n32) );
  INVXLTS U90 ( .A(readRequesterAddress[4]), .Y(n33) );
  INVXLTS U91 ( .A(n33), .Y(n34) );
  INVXLTS U92 ( .A(n33), .Y(n35) );
  INVXLTS U93 ( .A(n33), .Y(n36) );
  INVXLTS U94 ( .A(n33), .Y(n37) );
  INVXLTS U95 ( .A(readRequesterAddress[5]), .Y(n38) );
  INVXLTS U96 ( .A(n38), .Y(n39) );
  INVXLTS U97 ( .A(n38), .Y(n40) );
  INVXLTS U98 ( .A(n38), .Y(n41) );
  INVXLTS U99 ( .A(n38), .Y(n42) );
  INVXLTS U100 ( .A(n5327), .Y(n43) );
  INVXLTS U101 ( .A(n1), .Y(n44) );
  CLKBUFX2TS U102 ( .A(n1861), .Y(n45) );
  NAND2X1TS U103 ( .A(n1864), .B(n1861), .Y(n1807) );
  AOI21X1TS U104 ( .A0(n916), .A1(n119), .B0(n785), .Y(n1861) );
  CLKBUFX2TS U105 ( .A(n1839), .Y(n100) );
  NAND2X1TS U106 ( .A(n1839), .B(n935), .Y(n1799) );
  AOI21X1TS U107 ( .A0(n936), .A1(n940), .B0(n3861), .Y(n1839) );
  INVXLTS U108 ( .A(n7), .Y(n101) );
  INVXLTS U109 ( .A(n7), .Y(n102) );
  INVXLTS U110 ( .A(n103), .Y(n104) );
  INVXLTS U111 ( .A(n2), .Y(n105) );
  INVXLTS U112 ( .A(n2), .Y(n106) );
  CLKBUFX2TS U113 ( .A(n2034), .Y(n107) );
  INVXLTS U114 ( .A(n2055), .Y(n108) );
  INVXLTS U115 ( .A(n983), .Y(n110) );
  INVXLTS U116 ( .A(n110), .Y(n111) );
  INVXLTS U117 ( .A(n454), .Y(n112) );
  INVXLTS U118 ( .A(n1837), .Y(n113) );
  INVXLTS U119 ( .A(n113), .Y(n114) );
  INVX2TS U120 ( .A(n1942), .Y(n115) );
  INVXLTS U121 ( .A(n6), .Y(n117) );
  INVXLTS U122 ( .A(n6), .Y(n118) );
  INVXLTS U123 ( .A(n2025), .Y(n119) );
  INVXLTS U124 ( .A(n119), .Y(n120) );
  INVXLTS U125 ( .A(n112), .Y(n121) );
  INVXLTS U126 ( .A(n4), .Y(n122) );
  INVXLTS U127 ( .A(n466), .Y(n123) );
  INVXLTS U128 ( .A(n123), .Y(n124) );
  INVX2TS U129 ( .A(n125), .Y(n126) );
  INVXLTS U130 ( .A(n458), .Y(n127) );
  INVXLTS U131 ( .A(n127), .Y(n128) );
  INVXLTS U132 ( .A(n127), .Y(n129) );
  INVXLTS U133 ( .A(n11), .Y(n130) );
  INVXLTS U134 ( .A(n11), .Y(n131) );
  INVXLTS U135 ( .A(n777), .Y(n132) );
  INVXLTS U136 ( .A(n132), .Y(n133) );
  INVXLTS U137 ( .A(n132), .Y(n134) );
  INVXLTS U138 ( .A(n981), .Y(n135) );
  INVXLTS U139 ( .A(n135), .Y(n136) );
  INVXLTS U140 ( .A(n135), .Y(n137) );
  INVXLTS U141 ( .A(n982), .Y(n138) );
  INVXLTS U142 ( .A(n138), .Y(n139) );
  INVXLTS U143 ( .A(n138), .Y(n140) );
  INVXLTS U144 ( .A(destinationAddressIn_NORTH[13]), .Y(n141) );
  INVXLTS U145 ( .A(destinationAddressIn_NORTH[13]), .Y(n142) );
  INVXLTS U146 ( .A(destinationAddressIn_NORTH[11]), .Y(n143) );
  INVXLTS U147 ( .A(destinationAddressIn_NORTH[11]), .Y(n144) );
  INVXLTS U148 ( .A(destinationAddressIn_NORTH[9]), .Y(n145) );
  INVXLTS U149 ( .A(destinationAddressIn_NORTH[9]), .Y(n146) );
  INVXLTS U150 ( .A(destinationAddressIn_NORTH[12]), .Y(n147) );
  INVXLTS U151 ( .A(destinationAddressIn_NORTH[12]), .Y(n148) );
  INVXLTS U152 ( .A(destinationAddressIn_NORTH[10]), .Y(n149) );
  INVXLTS U153 ( .A(destinationAddressIn_NORTH[10]), .Y(n150) );
  INVXLTS U154 ( .A(destinationAddressIn_NORTH[8]), .Y(n151) );
  INVXLTS U155 ( .A(destinationAddressIn_NORTH[8]), .Y(n152) );
  INVXLTS U156 ( .A(n10), .Y(n153) );
  INVXLTS U157 ( .A(n10), .Y(n154) );
  INVXLTS U158 ( .A(n10), .Y(n155) );
  INVXLTS U159 ( .A(n979), .Y(n156) );
  INVXLTS U160 ( .A(n156), .Y(n157) );
  INVXLTS U161 ( .A(n984), .Y(n158) );
  INVXLTS U162 ( .A(n158), .Y(n159) );
  INVXLTS U163 ( .A(n158), .Y(n160) );
  INVXLTS U164 ( .A(n3831), .Y(n161) );
  INVXLTS U165 ( .A(n3827), .Y(n162) );
  INVXLTS U166 ( .A(n163), .Y(n164) );
  INVXLTS U167 ( .A(n163), .Y(n165) );
  INVXLTS U168 ( .A(n5), .Y(n166) );
  INVXLTS U169 ( .A(n5), .Y(n167) );
  INVXLTS U170 ( .A(n5), .Y(n168) );
  INVXLTS U171 ( .A(n1805), .Y(n169) );
  INVXLTS U172 ( .A(n169), .Y(n170) );
  INVXLTS U173 ( .A(n169), .Y(n171) );
  INVXLTS U174 ( .A(n3873), .Y(n172) );
  INVXLTS U175 ( .A(n3874), .Y(n173) );
  INVX2TS U176 ( .A(n1796), .Y(n174) );
  INVXLTS U177 ( .A(n174), .Y(n176) );
  INVXLTS U178 ( .A(n788), .Y(n177) );
  INVXLTS U179 ( .A(n3889), .Y(n178) );
  INVXLTS U180 ( .A(n3943), .Y(n179) );
  INVXLTS U181 ( .A(n3943), .Y(n180) );
  INVXLTS U182 ( .A(n181), .Y(n183) );
  INVXLTS U183 ( .A(n12), .Y(n184) );
  INVXLTS U184 ( .A(n12), .Y(n185) );
  INVXLTS U185 ( .A(n12), .Y(n186) );
  INVXLTS U186 ( .A(n121), .Y(n187) );
  INVXLTS U187 ( .A(n197), .Y(n188) );
  INVXLTS U188 ( .A(n188), .Y(n189) );
  INVXLTS U189 ( .A(n188), .Y(n190) );
  INVXLTS U190 ( .A(n188), .Y(n191) );
  INVXLTS U191 ( .A(n199), .Y(n192) );
  INVXLTS U192 ( .A(n192), .Y(n193) );
  INVXLTS U193 ( .A(n192), .Y(n194) );
  INVXLTS U194 ( .A(n112), .Y(n195) );
  INVXLTS U195 ( .A(n121), .Y(n196) );
  INVXLTS U196 ( .A(n195), .Y(n197) );
  INVXLTS U197 ( .A(n121), .Y(n198) );
  INVXLTS U198 ( .A(n195), .Y(n199) );
  NOR2X1TS U453 ( .A(n1086), .B(n2011), .Y(n1895) );
  OAI22X1TS U454 ( .A0(n1834), .A1(n803), .B0(n105), .B1(n456), .Y(n454) );
  INVX2TS U455 ( .A(n1797), .Y(n797) );
  CLKBUFX2TS U456 ( .A(n1836), .Y(n455) );
  AO21X1TS U457 ( .A0(n1893), .A1(n113), .B0(n1836), .Y(n1838) );
  INVX2TS U458 ( .A(n938), .Y(n456) );
  OAI22X1TS U459 ( .A0(n1834), .A1(n800), .B0(n106), .B1(n456), .Y(n1797) );
  AOI2BB1X1TS U460 ( .A0N(n102), .A1N(n1963), .B0(n1838), .Y(n1834) );
  AND3XLTS U461 ( .A(n1844), .B(n1839), .C(n102), .Y(n1219) );
  INVX2TS U462 ( .A(readIn_SOUTH), .Y(n457) );
  CLKBUFX2TS U463 ( .A(n1831), .Y(n460) );
  CLKBUFX2TS U464 ( .A(n1855), .Y(n461) );
  OAI21X1TS U465 ( .A0(n924), .A1(n928), .B0(n104), .Y(n1891) );
  NOR2X1TS U466 ( .A(n2067), .B(n4844), .Y(n1892) );
  INVX2TS U467 ( .A(n1132), .Y(n462) );
  CLKBUFX2TS U468 ( .A(n1880), .Y(n463) );
  OA22X1TS U469 ( .A0(n1821), .A1(n800), .B0(n1880), .B1(n105), .Y(n975) );
  OAI21X1TS U470 ( .A0(n1880), .A1(n1890), .B0(n1891), .Y(n1148) );
  OAI21X1TS U471 ( .A0(n463), .A1(n1918), .B0(n3122), .Y(n1823) );
  INVX2TS U472 ( .A(n2082), .Y(n464) );
  INVX2TS U473 ( .A(n2082), .Y(n465) );
  CLKBUFX2TS U474 ( .A(n1824), .Y(n467) );
  AOI21X1TS U475 ( .A0(n936), .A1(n938), .B0(n3600), .Y(n1824) );
  CLKBUFX2TS U476 ( .A(n2924), .Y(n468) );
  XOR2X1TS U477 ( .A(n156), .B(n972), .Y(n2061) );
  CLKBUFX2TS U478 ( .A(n2084), .Y(n776) );
  INVX2TS U479 ( .A(n776), .Y(n470) );
  INVX2TS U480 ( .A(n776), .Y(n471) );
  CLKBUFX2TS U481 ( .A(n2099), .Y(n779) );
  INVX2TS U482 ( .A(n779), .Y(n472) );
  INVX2TS U483 ( .A(n779), .Y(n473) );
  INVX2TS U484 ( .A(n779), .Y(n474) );
  AND2X2TS U485 ( .A(n1821), .B(n802), .Y(n1792) );
  INVX2TS U486 ( .A(n1792), .Y(n475) );
  INVX2TS U487 ( .A(n1792), .Y(n476) );
  INVX2TS U488 ( .A(n1792), .Y(n477) );
  CLKBUFX2TS U489 ( .A(n131), .Y(n912) );
  INVX2TS U490 ( .A(n912), .Y(n478) );
  INVX2TS U491 ( .A(n912), .Y(n479) );
  INVX2TS U492 ( .A(n912), .Y(n480) );
  CLKBUFX2TS U493 ( .A(n1847), .Y(n481) );
  CLKBUFX2TS U494 ( .A(n3831), .Y(n3818) );
  CLKBUFX2TS U495 ( .A(n1817), .Y(n482) );
  OAI21X1TS U496 ( .A0(n1889), .A1(n463), .B0(n3744), .Y(n1817) );
  CLKBUFX2TS U497 ( .A(selectBit_EAST), .Y(n483) );
  OA21XLTS U498 ( .A0(n2957), .A1(n2925), .B0(n483), .Y(n937) );
  CLKBUFX2TS U499 ( .A(n1827), .Y(n484) );
  AOI21X1TS U500 ( .A0(n1893), .A1(n1827), .B0(n922), .Y(n1829) );
  AOI21X1TS U501 ( .A0(n1827), .A1(n932), .B0(n918), .Y(n1859) );
  INVX2TS U502 ( .A(n1086), .Y(n485) );
  INVX2TS U503 ( .A(n926), .Y(n486) );
  XNOR2X1TS U504 ( .A(n2062), .B(n980), .Y(n1894) );
  AO21X2TS U505 ( .A0(n927), .A1(n931), .B0(n937), .Y(n2062) );
  INVXLTS U506 ( .A(selectBit_SOUTH), .Y(n487) );
  INVX2TS U507 ( .A(n487), .Y(n488) );
  XNOR2X1TS U508 ( .A(n974), .B(selectBit_SOUTH), .Y(n931) );
  NOR2X1TS U509 ( .A(selectBit_NORTH), .B(selectBit_SOUTH), .Y(n2925) );
  CLKBUFX2TS U510 ( .A(n2085), .Y(n778) );
  INVX2TS U511 ( .A(n778), .Y(n489) );
  INVX2TS U512 ( .A(n778), .Y(n490) );
  CLKBUFX2TS U513 ( .A(n2083), .Y(n771) );
  INVX2TS U514 ( .A(n771), .Y(n491) );
  INVX2TS U515 ( .A(n771), .Y(n492) );
  INVX2TS U516 ( .A(n493), .Y(n494) );
  CLKBUFX2TS U517 ( .A(cacheDataOut[7]), .Y(n495) );
  CLKBUFX2TS U518 ( .A(cacheDataOut[7]), .Y(n496) );
  CLKBUFX2TS U519 ( .A(cacheDataOut[31]), .Y(n497) );
  CLKBUFX2TS U520 ( .A(cacheDataOut[31]), .Y(n498) );
  CLKBUFX2TS U521 ( .A(cacheDataOut[30]), .Y(n499) );
  CLKBUFX2TS U522 ( .A(cacheDataOut[30]), .Y(n500) );
  CLKBUFX2TS U523 ( .A(cacheDataOut[29]), .Y(n501) );
  CLKBUFX2TS U524 ( .A(cacheDataOut[29]), .Y(n502) );
  CLKBUFX2TS U525 ( .A(cacheDataOut[28]), .Y(n503) );
  CLKBUFX2TS U526 ( .A(cacheDataOut[28]), .Y(n504) );
  CLKBUFX2TS U527 ( .A(cacheDataOut[27]), .Y(n505) );
  CLKBUFX2TS U528 ( .A(cacheDataOut[27]), .Y(n506) );
  CLKBUFX2TS U529 ( .A(cacheDataOut[26]), .Y(n507) );
  CLKBUFX2TS U530 ( .A(cacheDataOut[26]), .Y(n508) );
  CLKBUFX2TS U531 ( .A(cacheDataOut[25]), .Y(n509) );
  CLKBUFX2TS U532 ( .A(cacheDataOut[25]), .Y(n510) );
  CLKBUFX2TS U533 ( .A(cacheDataOut[24]), .Y(n511) );
  CLKBUFX2TS U534 ( .A(cacheDataOut[24]), .Y(n512) );
  CLKBUFX2TS U535 ( .A(cacheDataOut[23]), .Y(n513) );
  CLKBUFX2TS U536 ( .A(cacheDataOut[23]), .Y(n514) );
  CLKBUFX2TS U537 ( .A(cacheDataOut[22]), .Y(n515) );
  CLKBUFX2TS U538 ( .A(cacheDataOut[22]), .Y(n516) );
  CLKBUFX2TS U539 ( .A(cacheDataOut[21]), .Y(n517) );
  CLKBUFX2TS U540 ( .A(cacheDataOut[21]), .Y(n518) );
  CLKBUFX2TS U541 ( .A(cacheDataOut[20]), .Y(n519) );
  CLKBUFX2TS U542 ( .A(cacheDataOut[20]), .Y(n520) );
  CLKBUFX2TS U543 ( .A(cacheDataOut[19]), .Y(n521) );
  CLKBUFX2TS U544 ( .A(cacheDataOut[19]), .Y(n522) );
  CLKBUFX2TS U545 ( .A(cacheDataOut[18]), .Y(n523) );
  CLKBUFX2TS U546 ( .A(cacheDataOut[18]), .Y(n524) );
  CLKBUFX2TS U547 ( .A(cacheDataOut[17]), .Y(n525) );
  CLKBUFX2TS U548 ( .A(cacheDataOut[17]), .Y(n526) );
  CLKBUFX2TS U549 ( .A(cacheDataOut[16]), .Y(n527) );
  CLKBUFX2TS U550 ( .A(cacheDataOut[16]), .Y(n528) );
  CLKBUFX2TS U551 ( .A(cacheDataOut[15]), .Y(n529) );
  CLKBUFX2TS U552 ( .A(cacheDataOut[15]), .Y(n530) );
  CLKBUFX2TS U553 ( .A(cacheDataOut[14]), .Y(n531) );
  CLKBUFX2TS U554 ( .A(cacheDataOut[14]), .Y(n532) );
  CLKBUFX2TS U555 ( .A(cacheDataOut[13]), .Y(n533) );
  CLKBUFX2TS U556 ( .A(cacheDataOut[13]), .Y(n534) );
  CLKBUFX2TS U557 ( .A(cacheDataOut[12]), .Y(n535) );
  CLKBUFX2TS U558 ( .A(cacheDataOut[12]), .Y(n536) );
  CLKBUFX2TS U559 ( .A(cacheDataOut[11]), .Y(n537) );
  CLKBUFX2TS U560 ( .A(cacheDataOut[11]), .Y(n538) );
  CLKBUFX2TS U561 ( .A(cacheDataOut[10]), .Y(n539) );
  CLKBUFX2TS U562 ( .A(cacheDataOut[10]), .Y(n540) );
  CLKBUFX2TS U563 ( .A(cacheDataOut[9]), .Y(n541) );
  CLKBUFX2TS U564 ( .A(cacheDataOut[9]), .Y(n542) );
  CLKBUFX2TS U565 ( .A(cacheDataOut[8]), .Y(n543) );
  CLKBUFX2TS U566 ( .A(cacheDataOut[8]), .Y(n544) );
  CLKBUFX2TS U567 ( .A(cacheDataOut[6]), .Y(n545) );
  CLKBUFX2TS U568 ( .A(cacheDataOut[6]), .Y(n546) );
  CLKBUFX2TS U569 ( .A(cacheDataOut[5]), .Y(n547) );
  CLKBUFX2TS U570 ( .A(cacheDataOut[5]), .Y(n548) );
  CLKBUFX2TS U571 ( .A(cacheDataOut[4]), .Y(n549) );
  CLKBUFX2TS U572 ( .A(cacheDataOut[4]), .Y(n550) );
  CLKBUFX2TS U573 ( .A(cacheDataOut[3]), .Y(n551) );
  CLKBUFX2TS U574 ( .A(cacheDataOut[3]), .Y(n780) );
  CLKBUFX2TS U575 ( .A(cacheDataOut[2]), .Y(n786) );
  CLKBUFX2TS U576 ( .A(cacheDataOut[2]), .Y(n787) );
  CLKBUFX2TS U577 ( .A(cacheDataOut[1]), .Y(n789) );
  CLKBUFX2TS U578 ( .A(cacheDataOut[1]), .Y(n792) );
  CLKBUFX2TS U579 ( .A(cacheDataOut[0]), .Y(n793) );
  CLKBUFX2TS U580 ( .A(cacheDataOut[0]), .Y(n795) );
  CLKBUFX2TS U581 ( .A(n1810), .Y(n796) );
  CLKBUFX2TS U582 ( .A(n1810), .Y(n799) );
  INVX2TS U583 ( .A(n1892), .Y(n800) );
  INVX2TS U584 ( .A(n104), .Y(n803) );
  OA22X1TS U585 ( .A0(n1859), .A1(n800), .B0(n1890), .B1(n2025), .Y(n976) );
  CLKBUFX2TS U586 ( .A(n2087), .Y(n804) );
  CLKBUFX2TS U587 ( .A(n2087), .Y(n805) );
  AND2XLTS U588 ( .A(n1820), .B(n802), .Y(n1166) );
  CLKINVX2TS U589 ( .A(n1166), .Y(n907) );
  INVXLTS U590 ( .A(n1166), .Y(n908) );
  INVXLTS U591 ( .A(n1166), .Y(n913) );
  INVXLTS U592 ( .A(n1166), .Y(n914) );
  NOR2X2TS U593 ( .A(n974), .B(n985), .Y(n2957) );
  CLKINVX2TS U594 ( .A(selectBit_SOUTH), .Y(n985) );
  INVX2TS U595 ( .A(selectBit_EAST), .Y(n927) );
  CLKINVX2TS U596 ( .A(selectBit_NORTH), .Y(n974) );
  CLKBUFX2TS U597 ( .A(n1154), .Y(n3681) );
  CLKBUFX2TS U598 ( .A(n974), .Y(n915) );
  INVX2TS U599 ( .A(n1808), .Y(n785) );
  NOR3BX1TS U600 ( .AN(n45), .B(n1866), .C(n108), .Y(n1810) );
  NOR2BXLTS U601 ( .AN(n1847), .B(n1853), .Y(n1235) );
  OAI21X1TS U602 ( .A0(n114), .A1(n2010), .B0(n2056), .Y(n1866) );
  NOR2XLTS U603 ( .A(selectBit_NORTH), .B(n488), .Y(n925) );
  INVXLTS U604 ( .A(n1977), .Y(n791) );
  AND3XLTS U605 ( .A(n1827), .B(n1828), .C(n1824), .Y(n1187) );
  NOR2BXLTS U606 ( .AN(n467), .B(n1828), .Y(n1188) );
  NOR2XLTS U607 ( .A(n108), .B(n117), .Y(n1854) );
  NAND3XLTS U608 ( .A(n926), .B(n1941), .C(n1942), .Y(n2056) );
  NOR2X1TS U609 ( .A(n929), .B(n494), .Y(n1822) );
  AOI222XLTS U610 ( .A0(n4023), .A1(n3533), .B0(n3986), .B1(n3535), .C0(n4248), 
        .C1(n3579), .Y(n1940) );
  INVXLTS U611 ( .A(n3449), .Y(n3444) );
  INVXLTS U612 ( .A(n3448), .Y(n3445) );
  INVXLTS U613 ( .A(n3447), .Y(n3446) );
  INVXLTS U614 ( .A(n3397), .Y(n3392) );
  INVXLTS U615 ( .A(n3514), .Y(n3509) );
  INVXLTS U616 ( .A(n3396), .Y(n3393) );
  INVXLTS U617 ( .A(n3513), .Y(n3510) );
  INVXLTS U618 ( .A(n3395), .Y(n3394) );
  INVXLTS U619 ( .A(n3512), .Y(n3511) );
  INVX1TS U620 ( .A(n1807), .Y(n783) );
  CLKBUFX2TS U621 ( .A(n3139), .Y(n3134) );
  CLKBUFX2TS U622 ( .A(n3139), .Y(n3133) );
  CLKBUFX2TS U623 ( .A(n3138), .Y(n3135) );
  CLKBUFX2TS U624 ( .A(n3599), .Y(n3596) );
  CLKBUFX2TS U625 ( .A(n3598), .Y(n3597) );
  NOR3BX1TS U626 ( .AN(n1861), .B(n114), .C(n917), .Y(n1267) );
  NOR3BX1TS U627 ( .AN(n1831), .B(n1838), .C(n930), .Y(n1202) );
  AND2XLTS U628 ( .A(n921), .B(n100), .Y(n939) );
  CLKBUFX2TS U629 ( .A(n3335), .Y(n3332) );
  CLKBUFX2TS U630 ( .A(n3335), .Y(n3333) );
  CLKBUFX2TS U631 ( .A(n3121), .Y(n3116) );
  NAND3XLTS U632 ( .A(n1855), .B(n126), .C(n1859), .Y(n1805) );
  OAI21XLTS U633 ( .A0(n972), .A1(n2954), .B0(n2933), .Y(n2941) );
  NAND2XLTS U634 ( .A(n972), .B(n2954), .Y(n2933) );
  NOR2BXLTS U635 ( .AN(n1824), .B(n1860), .Y(n1185) );
  NOR2BXLTS U636 ( .AN(n1855), .B(n1860), .Y(n1249) );
  NOR2BXLTS U637 ( .AN(n1855), .B(n1858), .Y(n1251) );
  NAND2XLTS U638 ( .A(n1842), .B(n1893), .Y(n1813) );
  NOR2XLTS U639 ( .A(n1917), .B(n1823), .Y(n1171) );
  NOR2XLTS U640 ( .A(n1813), .B(n1817), .Y(n1153) );
  NOR2BXLTS U641 ( .AN(n1861), .B(n2056), .Y(n1265) );
  AND3XLTS U642 ( .A(n484), .B(n1858), .C(n461), .Y(n1252) );
  AND2XLTS U643 ( .A(n1836), .B(n460), .Y(n941) );
  INVX1TS U644 ( .A(n1230), .Y(n3401) );
  NAND3BXLTS U645 ( .AN(n1851), .B(n481), .C(n1853), .Y(n1230) );
  CLKINVX2TS U646 ( .A(n1182), .Y(n3600) );
  OAI22XLTS U647 ( .A0(n1829), .A1(n803), .B0(n1890), .B1(n1932), .Y(n1182) );
  NOR2BXLTS U648 ( .AN(n1879), .B(n1932), .Y(n1186) );
  NOR2BXLTS U649 ( .AN(n1879), .B(n463), .Y(n1152) );
  NOR3BXLTS U650 ( .AN(n1941), .B(n486), .C(n116), .Y(n1836) );
  OAI31XLTS U651 ( .A0(n934), .A1(n107), .A2(n936), .B0(n104), .Y(n1890) );
  OA21XLTS U652 ( .A0(n2942), .A1(n2943), .B0(n2944), .Y(n2932) );
  NAND3XLTS U653 ( .A(n115), .B(n486), .C(n1941), .Y(n1828) );
  NAND2XLTS U654 ( .A(n4194), .B(n922), .Y(n1825) );
  AOI32XLTS U655 ( .A0(n1842), .A1(n1843), .A2(n4200), .B0(n1844), .B1(n1845), 
        .Y(n1841) );
  OAI21XLTS U656 ( .A0(n2924), .A1(n973), .B0(n2952), .Y(n2954) );
  NOR2X1TS U657 ( .A(n985), .B(n2065), .Y(n2055) );
  AOI21XLTS U658 ( .A0(n985), .A1(n2065), .B0(n2055), .Y(n1989) );
  NAND3XLTS U659 ( .A(n1941), .B(n486), .C(n116), .Y(n1858) );
  INVXLTS U660 ( .A(n2010), .Y(n932) );
  OAI32XLTS U661 ( .A0(n4203), .A1(n920), .A2(n1851), .B0(n1852), .B1(n983), 
        .Y(n1850) );
  NOR2XLTS U662 ( .A(n1918), .B(n103), .Y(n1908) );
  NOR2BXLTS U663 ( .AN(n1879), .B(n120), .Y(n1250) );
  AOI32XLTS U664 ( .A0(n461), .A1(n1856), .A2(n1857), .B0(n3332), .B1(n682), 
        .Y(n2564) );
  NAND2XLTS U665 ( .A(n4194), .B(n918), .Y(n1856) );
  AOI32XLTS U666 ( .A0(n484), .A1(n1858), .A2(n4200), .B0(n1859), .B1(n1830), 
        .Y(n1857) );
  NAND2XLTS U667 ( .A(n104), .B(n4572), .Y(n1136) );
  OAI22XLTS U668 ( .A0(n1860), .A1(n998), .B0(n125), .B1(n983), .Y(n1830) );
  AOI22XLTS U669 ( .A0(n1816), .A1(n983), .B0(n933), .B1(n998), .Y(n1815) );
  NAND2X1TS U670 ( .A(n469), .B(n942), .Y(n1880) );
  NAND2X1TS U671 ( .A(n5323), .B(n942), .Y(n1932) );
  NAND3X1TS U672 ( .A(n124), .B(n129), .C(n122), .Y(n2099) );
  OAI211XLTS U673 ( .A0(n4570), .A1(n3925), .B0(n1276), .C0(n1277), .Y(n2835)
         );
  OAI211XLTS U674 ( .A0(n4567), .A1(n3925), .B0(n1274), .C0(n1275), .Y(n2836)
         );
  OAI211XLTS U675 ( .A0(n4563), .A1(n3926), .B0(n1272), .C0(n1273), .Y(n2837)
         );
  OAI211XLTS U676 ( .A0(n4560), .A1(n3926), .B0(n1270), .C0(n1271), .Y(n2838)
         );
  OAI211XLTS U677 ( .A0(n4556), .A1(n3926), .B0(n1268), .C0(n1269), .Y(n2839)
         );
  OAI211XLTS U678 ( .A0(n4553), .A1(n3926), .B0(n1263), .C0(n1264), .Y(n2840)
         );
  OAI211XLTS U679 ( .A0(n3393), .A1(n4347), .B0(n1406), .C0(n1407), .Y(n2770)
         );
  AOI22XLTS U680 ( .A0(n793), .A1(n3359), .B0(n4249), .B1(n3337), .Y(n1406) );
  OAI211XLTS U681 ( .A0(n3393), .A1(n4350), .B0(n1408), .C0(n1409), .Y(n2769)
         );
  AOI22XLTS U682 ( .A0(n789), .A1(n3358), .B0(n4252), .B1(n3337), .Y(n1408) );
  OAI211XLTS U683 ( .A0(n3391), .A1(n4365), .B0(n1418), .C0(n1419), .Y(n2764)
         );
  AOI22XLTS U684 ( .A0(n545), .A1(n3358), .B0(n4267), .B1(n3339), .Y(n1418) );
  OAI211XLTS U685 ( .A0(n3390), .A1(n4377), .B0(n1426), .C0(n1427), .Y(n2760)
         );
  AOI22XLTS U686 ( .A0(n539), .A1(n3359), .B0(n4279), .B1(n3339), .Y(n1426) );
  OAI211XLTS U687 ( .A0(n3386), .A1(n4428), .B0(n1460), .C0(n1461), .Y(n2743)
         );
  AOI22XLTS U688 ( .A0(n505), .A1(n3357), .B0(n4330), .B1(n3344), .Y(n1460) );
  OAI211XLTS U689 ( .A0(n3391), .A1(n4368), .B0(n1420), .C0(n1421), .Y(n2763)
         );
  AOI22XLTS U690 ( .A0(n495), .A1(n3361), .B0(n4270), .B1(n3339), .Y(n1420) );
  OAI211XLTS U691 ( .A0(n3391), .A1(n4371), .B0(n1422), .C0(n1423), .Y(n2762)
         );
  AOI22XLTS U692 ( .A0(n543), .A1(n3361), .B0(n4273), .B1(n3339), .Y(n1422) );
  OAI211XLTS U693 ( .A0(n3391), .A1(n4374), .B0(n1424), .C0(n1425), .Y(n2761)
         );
  AOI22XLTS U694 ( .A0(n541), .A1(n3364), .B0(n4276), .B1(n3342), .Y(n1424) );
  OAI211XLTS U695 ( .A0(n3390), .A1(n4380), .B0(n1428), .C0(n1429), .Y(n2759)
         );
  AOI22XLTS U696 ( .A0(n537), .A1(n3361), .B0(n4282), .B1(n3340), .Y(n1428) );
  OAI211XLTS U697 ( .A0(n3390), .A1(n4383), .B0(n1430), .C0(n1431), .Y(n2758)
         );
  AOI22XLTS U698 ( .A0(n535), .A1(n3361), .B0(n4285), .B1(n3340), .Y(n1430) );
  OAI211XLTS U699 ( .A0(n3390), .A1(n4386), .B0(n1432), .C0(n1433), .Y(n2757)
         );
  AOI22XLTS U700 ( .A0(n533), .A1(n3364), .B0(n4288), .B1(n3340), .Y(n1432) );
  OAI211XLTS U701 ( .A0(n3388), .A1(n4401), .B0(n1442), .C0(n1443), .Y(n2752)
         );
  AOI22XLTS U702 ( .A0(n523), .A1(n3364), .B0(n4303), .B1(n3341), .Y(n1442) );
  OAI211XLTS U703 ( .A0(n3388), .A1(n4404), .B0(n1444), .C0(n1445), .Y(n2751)
         );
  AOI22XLTS U704 ( .A0(n521), .A1(n3366), .B0(n4306), .B1(n3342), .Y(n1444) );
  OAI211XLTS U705 ( .A0(n3388), .A1(n4407), .B0(n1446), .C0(n1447), .Y(n2750)
         );
  AOI22XLTS U706 ( .A0(n519), .A1(n3360), .B0(n4309), .B1(n3342), .Y(n1446) );
  OAI211XLTS U707 ( .A0(n3388), .A1(n4410), .B0(n1448), .C0(n1449), .Y(n2749)
         );
  AOI22XLTS U708 ( .A0(n517), .A1(n3360), .B0(n4312), .B1(n3342), .Y(n1448) );
  OAI211XLTS U709 ( .A0(n3387), .A1(n4416), .B0(n1452), .C0(n1453), .Y(n2747)
         );
  AOI22XLTS U710 ( .A0(n513), .A1(n3357), .B0(n4318), .B1(n3343), .Y(n1452) );
  OAI211XLTS U711 ( .A0(n3387), .A1(n4422), .B0(n1456), .C0(n1457), .Y(n2745)
         );
  AOI22XLTS U712 ( .A0(n509), .A1(n3356), .B0(n4324), .B1(n3343), .Y(n1456) );
  OAI211XLTS U713 ( .A0(n3386), .A1(n4425), .B0(n1458), .C0(n1459), .Y(n2744)
         );
  AOI22XLTS U714 ( .A0(n507), .A1(n3362), .B0(n4327), .B1(n3344), .Y(n1458) );
  OAI211XLTS U715 ( .A0(n3386), .A1(n4432), .B0(n1462), .C0(n1463), .Y(n2742)
         );
  AOI22XLTS U716 ( .A0(n503), .A1(n3356), .B0(n4333), .B1(n3344), .Y(n1462) );
  OAI211XLTS U717 ( .A0(n3386), .A1(n4435), .B0(n1464), .C0(n1465), .Y(n2741)
         );
  AOI22XLTS U718 ( .A0(n501), .A1(n3356), .B0(n4336), .B1(n3344), .Y(n1464) );
  OAI211XLTS U719 ( .A0(n3384), .A1(n3957), .B0(n1996), .C0(n1997), .Y(n2489)
         );
  AOI22XLTS U720 ( .A0(n3355), .A1(n31), .B0(n3997), .B1(n3347), .Y(n1996) );
  OAI211XLTS U721 ( .A0(n3384), .A1(n3960), .B0(n1998), .C0(n1999), .Y(n2488)
         );
  AOI22XLTS U722 ( .A0(n3355), .A1(n36), .B0(n4000), .B1(n3350), .Y(n1998) );
  OAI211XLTS U723 ( .A0(n3384), .A1(n3963), .B0(n2000), .C0(n2001), .Y(n2487)
         );
  AOI22XLTS U724 ( .A0(n3353), .A1(n41), .B0(n4003), .B1(n3351), .Y(n2000) );
  OAI211XLTS U725 ( .A0(n3384), .A1(n3954), .B0(n1994), .C0(n1995), .Y(n2490)
         );
  AOI22XLTS U726 ( .A0(n3355), .A1(n26), .B0(n3994), .B1(n3350), .Y(n1994) );
  OAI211XLTS U727 ( .A0(n3385), .A1(n4438), .B0(n1466), .C0(n1467), .Y(n2740)
         );
  AOI22XLTS U728 ( .A0(n499), .A1(n3356), .B0(n4339), .B1(n3345), .Y(n1466) );
  OAI211XLTS U729 ( .A0(n3389), .A1(n4398), .B0(n1440), .C0(n1441), .Y(n2753)
         );
  AOI22XLTS U730 ( .A0(n525), .A1(n3363), .B0(n4300), .B1(n3341), .Y(n1440) );
  OAI211XLTS U731 ( .A0(n3389), .A1(n4392), .B0(n1436), .C0(n1437), .Y(n2755)
         );
  AOI22XLTS U732 ( .A0(n529), .A1(n3362), .B0(n4294), .B1(n3341), .Y(n1436) );
  OAI211XLTS U733 ( .A0(n3389), .A1(n4389), .B0(n1434), .C0(n1435), .Y(n2756)
         );
  AOI22XLTS U734 ( .A0(n531), .A1(n3363), .B0(n4291), .B1(n3340), .Y(n1434) );
  OAI211XLTS U735 ( .A0(n3392), .A1(n4362), .B0(n1416), .C0(n1417), .Y(n2765)
         );
  AOI22XLTS U736 ( .A0(n547), .A1(n3366), .B0(n4264), .B1(n3338), .Y(n1416) );
  OAI211XLTS U737 ( .A0(n3392), .A1(n4359), .B0(n1414), .C0(n1415), .Y(n2766)
         );
  AOI22XLTS U738 ( .A0(n549), .A1(n3358), .B0(n4261), .B1(n3338), .Y(n1414) );
  OAI211XLTS U739 ( .A0(n3392), .A1(n4356), .B0(n1412), .C0(n1413), .Y(n2767)
         );
  AOI22XLTS U740 ( .A0(n551), .A1(n3359), .B0(n4258), .B1(n3338), .Y(n1412) );
  OAI211XLTS U741 ( .A0(n3385), .A1(n3951), .B0(n1992), .C0(n1993), .Y(n2491)
         );
  AOI22XLTS U742 ( .A0(n3354), .A1(n21), .B0(n3991), .B1(n3345), .Y(n1992) );
  OAI211XLTS U743 ( .A0(n3385), .A1(n3948), .B0(n1990), .C0(n1991), .Y(n2492)
         );
  AOI22XLTS U744 ( .A0(n3355), .A1(n16), .B0(n3988), .B1(n3345), .Y(n1990) );
  OAI211XLTS U745 ( .A0(n3385), .A1(n4442), .B0(n1468), .C0(n1469), .Y(n2739)
         );
  AOI22XLTS U746 ( .A0(n497), .A1(n3359), .B0(n4342), .B1(n3345), .Y(n1468) );
  OAI211XLTS U747 ( .A0(n3387), .A1(n4419), .B0(n1454), .C0(n1455), .Y(n2746)
         );
  AOI22XLTS U748 ( .A0(n511), .A1(n3357), .B0(n4321), .B1(n3343), .Y(n1454) );
  OAI211XLTS U749 ( .A0(n3387), .A1(n4413), .B0(n1450), .C0(n1451), .Y(n2748)
         );
  AOI22XLTS U750 ( .A0(n515), .A1(n3357), .B0(n4315), .B1(n3343), .Y(n1450) );
  OAI211XLTS U751 ( .A0(n3389), .A1(n4395), .B0(n1438), .C0(n1439), .Y(n2754)
         );
  AOI22XLTS U752 ( .A0(n527), .A1(n3365), .B0(n4297), .B1(n3341), .Y(n1438) );
  OAI211XLTS U753 ( .A0(n3392), .A1(n4353), .B0(n1410), .C0(n1411), .Y(n2768)
         );
  AOI22XLTS U754 ( .A0(n786), .A1(n3358), .B0(n4255), .B1(n3338), .Y(n1410) );
  OAI211XLTS U755 ( .A0(n4188), .A1(n3393), .B0(n1242), .C0(n1243), .Y(n2848)
         );
  AOI22XLTS U756 ( .A0(n3354), .A1(n37), .B0(n3336), .B1(n4036), .Y(n1242) );
  OAI211XLTS U757 ( .A0(n4191), .A1(n3393), .B0(n1244), .C0(n1245), .Y(n2847)
         );
  AOI22XLTS U758 ( .A0(n3354), .A1(n42), .B0(n3337), .B1(n4039), .Y(n1244) );
  OAI211XLTS U759 ( .A0(n4179), .A1(n3394), .B0(n1236), .C0(n1237), .Y(n2851)
         );
  AOI22XLTS U760 ( .A0(n3353), .A1(n22), .B0(n3336), .B1(n4027), .Y(n1236) );
  OAI211XLTS U761 ( .A0(n4176), .A1(n3394), .B0(n1231), .C0(n1232), .Y(n2852)
         );
  AOI22XLTS U762 ( .A0(n3354), .A1(n17), .B0(n3337), .B1(n4024), .Y(n1231) );
  OAI211XLTS U763 ( .A0(n4185), .A1(n3394), .B0(n1240), .C0(n1241), .Y(n2849)
         );
  AOI22XLTS U764 ( .A0(n3353), .A1(n32), .B0(n3336), .B1(n4033), .Y(n1240) );
  OAI211XLTS U765 ( .A0(n4182), .A1(n3394), .B0(n1238), .C0(n1239), .Y(n2850)
         );
  AOI22XLTS U766 ( .A0(n3353), .A1(n27), .B0(n3336), .B1(n4030), .Y(n1238) );
  OAI211XLTS U767 ( .A0(n3925), .A1(n4448), .B0(n1280), .C0(n1281), .Y(n2833)
         );
  OAI211XLTS U768 ( .A0(n3925), .A1(n4445), .B0(n1278), .C0(n1279), .Y(n2834)
         );
  OAI211XLTS U769 ( .A0(n3918), .A1(n4224), .B0(n2045), .C0(n2046), .Y(n2459)
         );
  OAI211XLTS U770 ( .A0(n3918), .A1(n4218), .B0(n2041), .C0(n2042), .Y(n2461)
         );
  OAI211XLTS U771 ( .A0(n3918), .A1(n4215), .B0(n2039), .C0(n2040), .Y(n2462)
         );
  OAI211XLTS U772 ( .A0(n3929), .A1(n4212), .B0(n2037), .C0(n2038), .Y(n2463)
         );
  OAI211XLTS U773 ( .A0(n3928), .A1(n4550), .B0(n1340), .C0(n1341), .Y(n2803)
         );
  OAI211XLTS U774 ( .A0(n3931), .A1(n4546), .B0(n1338), .C0(n1339), .Y(n2804)
         );
  OAI211XLTS U775 ( .A0(n3927), .A1(n4543), .B0(n1336), .C0(n1337), .Y(n2805)
         );
  OAI211XLTS U776 ( .A0(n3930), .A1(n4533), .B0(n1330), .C0(n1331), .Y(n2808)
         );
  OAI211XLTS U777 ( .A0(n3919), .A1(n4529), .B0(n1328), .C0(n1329), .Y(n2809)
         );
  OAI211XLTS U778 ( .A0(n3919), .A1(n4526), .B0(n1326), .C0(n1327), .Y(n2810)
         );
  OAI211XLTS U779 ( .A0(n3919), .A1(n4519), .B0(n1322), .C0(n1323), .Y(n2812)
         );
  OAI211XLTS U780 ( .A0(n3920), .A1(n4516), .B0(n1320), .C0(n1321), .Y(n2813)
         );
  OAI211XLTS U781 ( .A0(n3920), .A1(n4509), .B0(n1316), .C0(n1317), .Y(n2815)
         );
  OAI211XLTS U782 ( .A0(n3920), .A1(n4506), .B0(n1314), .C0(n1315), .Y(n2816)
         );
  OAI211XLTS U783 ( .A0(n3921), .A1(n4502), .B0(n1312), .C0(n1313), .Y(n2817)
         );
  OAI211XLTS U784 ( .A0(n3921), .A1(n4499), .B0(n1310), .C0(n1311), .Y(n2818)
         );
  OAI211XLTS U785 ( .A0(n3921), .A1(n4496), .B0(n1308), .C0(n1309), .Y(n2819)
         );
  OAI211XLTS U786 ( .A0(n3921), .A1(n4492), .B0(n1306), .C0(n1307), .Y(n2820)
         );
  OAI211XLTS U787 ( .A0(n3922), .A1(n4489), .B0(n1304), .C0(n1305), .Y(n2821)
         );
  OAI211XLTS U788 ( .A0(n3922), .A1(n4486), .B0(n1302), .C0(n1303), .Y(n2822)
         );
  OAI211XLTS U789 ( .A0(n3922), .A1(n4482), .B0(n1300), .C0(n1301), .Y(n2823)
         );
  OAI211XLTS U790 ( .A0(n3922), .A1(n4479), .B0(n1298), .C0(n1299), .Y(n2824)
         );
  OAI211XLTS U791 ( .A0(n3923), .A1(n4472), .B0(n1294), .C0(n1295), .Y(n2826)
         );
  OAI211XLTS U792 ( .A0(n3923), .A1(n4469), .B0(n1292), .C0(n1293), .Y(n2827)
         );
  OAI211XLTS U793 ( .A0(n3923), .A1(n4465), .B0(n1290), .C0(n1291), .Y(n2828)
         );
  OAI211XLTS U794 ( .A0(n3924), .A1(n4459), .B0(n1286), .C0(n1287), .Y(n2830)
         );
  OAI211XLTS U795 ( .A0(n3924), .A1(n4455), .B0(n1284), .C0(n1285), .Y(n2831)
         );
  OAI211XLTS U796 ( .A0(n3918), .A1(n4221), .B0(n2043), .C0(n2044), .Y(n2460)
         );
  OAI211XLTS U797 ( .A0(n784), .A1(n4209), .B0(n2035), .C0(n2036), .Y(n2464)
         );
  OAI211XLTS U798 ( .A0(n3929), .A1(n4540), .B0(n1334), .C0(n1335), .Y(n2806)
         );
  OAI211XLTS U799 ( .A0(n3928), .A1(n4536), .B0(n1332), .C0(n1333), .Y(n2807)
         );
  OAI211XLTS U800 ( .A0(n3919), .A1(n4523), .B0(n1324), .C0(n1325), .Y(n2811)
         );
  OAI211XLTS U801 ( .A0(n3920), .A1(n4513), .B0(n1318), .C0(n1319), .Y(n2814)
         );
  OAI211XLTS U802 ( .A0(n3923), .A1(n4475), .B0(n1296), .C0(n1297), .Y(n2825)
         );
  OAI211XLTS U803 ( .A0(n3924), .A1(n4462), .B0(n1288), .C0(n1289), .Y(n2829)
         );
  OAI211XLTS U804 ( .A0(n3924), .A1(n4452), .B0(n1282), .C0(n1283), .Y(n2832)
         );
  AOI22XLTS U805 ( .A0(n1818), .A1(n1819), .B0(n3136), .B1(n677), .Y(n2569) );
  AOI2BB2XLTS U806 ( .B0(n1811), .B1(n1812), .A0N(n3744), .A1N(readOutbuffer_7), .Y(n2570) );
  XOR2XLTS U807 ( .A(n1132), .B(selectBit_WEST), .Y(n2951) );
  NOR2BXLTS U808 ( .AN(n2952), .B(n2924), .Y(n2950) );
  NAND2XLTS U809 ( .A(n4194), .B(n455), .Y(n1832) );
  OAI211XLTS U810 ( .A0(n3584), .A1(n909), .B0(n1930), .C0(n1931), .Y(n2529)
         );
  OAI211XLTS U811 ( .A0(n3124), .A1(n664), .B0(n1725), .C0(n1726), .Y(n2611)
         );
  OAI211XLTS U812 ( .A0(n3124), .A1(n663), .B0(n1723), .C0(n1724), .Y(n2612)
         );
  OAI211XLTS U813 ( .A0(n3584), .A1(n891), .B0(n1193), .C0(n1194), .Y(n2867)
         );
  OAI211XLTS U814 ( .A0(n3584), .A1(n889), .B0(n1189), .C0(n1190), .Y(n2869)
         );
  OAI211XLTS U815 ( .A0(n3320), .A1(n873), .B0(n2023), .C0(n2024), .Y(n2473)
         );
  OAI211XLTS U816 ( .A0(n3320), .A1(n898), .B0(n1257), .C0(n1258), .Y(n2843)
         );
  OAI211XLTS U817 ( .A0(n3320), .A1(n896), .B0(n1253), .C0(n1254), .Y(n2845)
         );
  OAI211XLTS U818 ( .A0(n3510), .A1(n4251), .B0(n1534), .C0(n1535), .Y(n2706)
         );
  OAI211XLTS U819 ( .A0(n3510), .A1(n4254), .B0(n1536), .C0(n1537), .Y(n2705)
         );
  OAI211XLTS U820 ( .A0(n3445), .A1(n4254), .B0(n1472), .C0(n1473), .Y(n2737)
         );
  OAI211XLTS U821 ( .A0(n3445), .A1(n4251), .B0(n1470), .C0(n1471), .Y(n2738)
         );
  OAI211XLTS U822 ( .A0(n3509), .A1(n4257), .B0(n1538), .C0(n1539), .Y(n2704)
         );
  OAI211XLTS U823 ( .A0(n3509), .A1(n4260), .B0(n1540), .C0(n1541), .Y(n2703)
         );
  OAI211XLTS U824 ( .A0(n3509), .A1(n4263), .B0(n1542), .C0(n1543), .Y(n2702)
         );
  OAI211XLTS U825 ( .A0(n3509), .A1(n4266), .B0(n1544), .C0(n1545), .Y(n2701)
         );
  OAI211XLTS U826 ( .A0(n3508), .A1(n4269), .B0(n1546), .C0(n1547), .Y(n2700)
         );
  OAI211XLTS U827 ( .A0(n3508), .A1(n4272), .B0(n1548), .C0(n1549), .Y(n2699)
         );
  OAI211XLTS U828 ( .A0(n3508), .A1(n4275), .B0(n1550), .C0(n1551), .Y(n2698)
         );
  OAI211XLTS U829 ( .A0(n3508), .A1(n4278), .B0(n1552), .C0(n1553), .Y(n2697)
         );
  OAI211XLTS U830 ( .A0(n3507), .A1(n4281), .B0(n1554), .C0(n1555), .Y(n2696)
         );
  OAI211XLTS U831 ( .A0(n3507), .A1(n4284), .B0(n1556), .C0(n1557), .Y(n2695)
         );
  OAI211XLTS U832 ( .A0(n3507), .A1(n4287), .B0(n1558), .C0(n1559), .Y(n2694)
         );
  OAI211XLTS U833 ( .A0(n3507), .A1(n4290), .B0(n1560), .C0(n1561), .Y(n2693)
         );
  OAI211XLTS U834 ( .A0(n3506), .A1(n4293), .B0(n1562), .C0(n1563), .Y(n2692)
         );
  OAI211XLTS U835 ( .A0(n3506), .A1(n4296), .B0(n1564), .C0(n1565), .Y(n2691)
         );
  OAI211XLTS U836 ( .A0(n3506), .A1(n4299), .B0(n1566), .C0(n1567), .Y(n2690)
         );
  OAI211XLTS U837 ( .A0(n3506), .A1(n4302), .B0(n1568), .C0(n1569), .Y(n2689)
         );
  OAI211XLTS U838 ( .A0(n3505), .A1(n4305), .B0(n1570), .C0(n1571), .Y(n2688)
         );
  OAI211XLTS U839 ( .A0(n3505), .A1(n4308), .B0(n1572), .C0(n1573), .Y(n2687)
         );
  OAI211XLTS U840 ( .A0(n3505), .A1(n4311), .B0(n1574), .C0(n1575), .Y(n2686)
         );
  OAI211XLTS U841 ( .A0(n3505), .A1(n4314), .B0(n1576), .C0(n1577), .Y(n2685)
         );
  OAI211XLTS U842 ( .A0(n3504), .A1(n4317), .B0(n1578), .C0(n1579), .Y(n2684)
         );
  OAI211XLTS U843 ( .A0(n3504), .A1(n4320), .B0(n1580), .C0(n1581), .Y(n2683)
         );
  OAI211XLTS U844 ( .A0(n3504), .A1(n4323), .B0(n1582), .C0(n1583), .Y(n2682)
         );
  OAI211XLTS U845 ( .A0(n3504), .A1(n4326), .B0(n1584), .C0(n1585), .Y(n2681)
         );
  OAI211XLTS U846 ( .A0(n3503), .A1(n4329), .B0(n1586), .C0(n1587), .Y(n2680)
         );
  OAI211XLTS U847 ( .A0(n3503), .A1(n4332), .B0(n1588), .C0(n1589), .Y(n2679)
         );
  OAI211XLTS U848 ( .A0(n3503), .A1(n4335), .B0(n1590), .C0(n1591), .Y(n2678)
         );
  OAI211XLTS U849 ( .A0(n3503), .A1(n4338), .B0(n1592), .C0(n1593), .Y(n2677)
         );
  OAI211XLTS U850 ( .A0(n3502), .A1(n4341), .B0(n1594), .C0(n1595), .Y(n2676)
         );
  OAI211XLTS U851 ( .A0(n3502), .A1(n4344), .B0(n1596), .C0(n1597), .Y(n2675)
         );
  OAI211XLTS U852 ( .A0(n3501), .A1(n4005), .B0(n1953), .C0(n1954), .Y(n2515)
         );
  OAI211XLTS U853 ( .A0(n3501), .A1(n3999), .B0(n1949), .C0(n1950), .Y(n2517)
         );
  OAI211XLTS U854 ( .A0(n3501), .A1(n3996), .B0(n1947), .C0(n1948), .Y(n2518)
         );
  OAI211XLTS U855 ( .A0(n3502), .A1(n3993), .B0(n1945), .C0(n1946), .Y(n2519)
         );
  OAI211XLTS U856 ( .A0(n3502), .A1(n3990), .B0(n1943), .C0(n1944), .Y(n2520)
         );
  OAI211XLTS U857 ( .A0(n3501), .A1(n4002), .B0(n1951), .C0(n1952), .Y(n2516)
         );
  OAI211XLTS U858 ( .A0(n3437), .A1(n3993), .B0(n1967), .C0(n1968), .Y(n2505)
         );
  OAI211XLTS U859 ( .A0(n3437), .A1(n3990), .B0(n1965), .C0(n1966), .Y(n2506)
         );
  OAI211XLTS U860 ( .A0(n3437), .A1(n4344), .B0(n1532), .C0(n1533), .Y(n2707)
         );
  OAI211XLTS U861 ( .A0(n3437), .A1(n4341), .B0(n1530), .C0(n1531), .Y(n2708)
         );
  OAI211XLTS U862 ( .A0(n3438), .A1(n4338), .B0(n1528), .C0(n1529), .Y(n2709)
         );
  OAI211XLTS U863 ( .A0(n3438), .A1(n4335), .B0(n1526), .C0(n1527), .Y(n2710)
         );
  OAI211XLTS U864 ( .A0(n3438), .A1(n4332), .B0(n1524), .C0(n1525), .Y(n2711)
         );
  OAI211XLTS U865 ( .A0(n3438), .A1(n4329), .B0(n1522), .C0(n1523), .Y(n2712)
         );
  OAI211XLTS U866 ( .A0(n3439), .A1(n4323), .B0(n1518), .C0(n1519), .Y(n2714)
         );
  OAI211XLTS U867 ( .A0(n3439), .A1(n4317), .B0(n1514), .C0(n1515), .Y(n2716)
         );
  OAI211XLTS U868 ( .A0(n3440), .A1(n4314), .B0(n1512), .C0(n1513), .Y(n2717)
         );
  OAI211XLTS U869 ( .A0(n3440), .A1(n4308), .B0(n1508), .C0(n1509), .Y(n2719)
         );
  OAI211XLTS U870 ( .A0(n3441), .A1(n4302), .B0(n1504), .C0(n1505), .Y(n2721)
         );
  OAI211XLTS U871 ( .A0(n3441), .A1(n4299), .B0(n1502), .C0(n1503), .Y(n2722)
         );
  OAI211XLTS U872 ( .A0(n3441), .A1(n4293), .B0(n1498), .C0(n1499), .Y(n2724)
         );
  OAI211XLTS U873 ( .A0(n3442), .A1(n4287), .B0(n1494), .C0(n1495), .Y(n2726)
         );
  OAI211XLTS U874 ( .A0(n3442), .A1(n4284), .B0(n1492), .C0(n1493), .Y(n2727)
         );
  OAI211XLTS U875 ( .A0(n3442), .A1(n4281), .B0(n1490), .C0(n1491), .Y(n2728)
         );
  OAI211XLTS U876 ( .A0(n3443), .A1(n4278), .B0(n1488), .C0(n1489), .Y(n2729)
         );
  OAI211XLTS U877 ( .A0(n3443), .A1(n4275), .B0(n1486), .C0(n1487), .Y(n2730)
         );
  OAI211XLTS U878 ( .A0(n3443), .A1(n4269), .B0(n1482), .C0(n1483), .Y(n2732)
         );
  OAI211XLTS U879 ( .A0(n3444), .A1(n4260), .B0(n1476), .C0(n1477), .Y(n2735)
         );
  OAI211XLTS U880 ( .A0(n3439), .A1(n4326), .B0(n1520), .C0(n1521), .Y(n2713)
         );
  OAI211XLTS U881 ( .A0(n3439), .A1(n4320), .B0(n1516), .C0(n1517), .Y(n2715)
         );
  OAI211XLTS U882 ( .A0(n3440), .A1(n4311), .B0(n1510), .C0(n1511), .Y(n2718)
         );
  OAI211XLTS U883 ( .A0(n3440), .A1(n4305), .B0(n1506), .C0(n1507), .Y(n2720)
         );
  OAI211XLTS U884 ( .A0(n3441), .A1(n4296), .B0(n1500), .C0(n1501), .Y(n2723)
         );
  OAI211XLTS U885 ( .A0(n3442), .A1(n4290), .B0(n1496), .C0(n1497), .Y(n2725)
         );
  OAI211XLTS U886 ( .A0(n3444), .A1(n4266), .B0(n1480), .C0(n1481), .Y(n2733)
         );
  OAI211XLTS U887 ( .A0(n3444), .A1(n4263), .B0(n1478), .C0(n1479), .Y(n2734)
         );
  OAI211XLTS U888 ( .A0(n3444), .A1(n4257), .B0(n1474), .C0(n1475), .Y(n2736)
         );
  OAI211XLTS U889 ( .A0(n3443), .A1(n4272), .B0(n1484), .C0(n1485), .Y(n2731)
         );
  OAI211XLTS U890 ( .A0(n3436), .A1(n4005), .B0(n1975), .C0(n1976), .Y(n2501)
         );
  OAI211XLTS U891 ( .A0(n3436), .A1(n4002), .B0(n1973), .C0(n1974), .Y(n2502)
         );
  OAI211XLTS U892 ( .A0(n3436), .A1(n3999), .B0(n1971), .C0(n1972), .Y(n2503)
         );
  OAI211XLTS U893 ( .A0(n3436), .A1(n3996), .B0(n1969), .C0(n1970), .Y(n2504)
         );
  OAI211XLTS U894 ( .A0(n3593), .A1(n843), .B0(n1660), .C0(n1661), .Y(n2643)
         );
  OAI211XLTS U895 ( .A0(n3590), .A1(n842), .B0(n1630), .C0(n1631), .Y(n2658)
         );
  OAI211XLTS U896 ( .A0(n3589), .A1(n841), .B0(n1628), .C0(n1629), .Y(n2659)
         );
  OAI211XLTS U897 ( .A0(n3588), .A1(n840), .B0(n1620), .C0(n1621), .Y(n2663)
         );
  OAI211XLTS U898 ( .A0(n3586), .A1(n839), .B0(n1600), .C0(n1601), .Y(n2673)
         );
  OAI211XLTS U899 ( .A0(n3593), .A1(n834), .B0(n1658), .C0(n1659), .Y(n2644)
         );
  OAI211XLTS U900 ( .A0(n3593), .A1(n833), .B0(n1656), .C0(n1657), .Y(n2645)
         );
  OAI211XLTS U901 ( .A0(n3593), .A1(n832), .B0(n1654), .C0(n1655), .Y(n2646)
         );
  OAI211XLTS U902 ( .A0(n3592), .A1(n831), .B0(n1652), .C0(n1653), .Y(n2647)
         );
  OAI211XLTS U903 ( .A0(n3592), .A1(n830), .B0(n1650), .C0(n1651), .Y(n2648)
         );
  OAI211XLTS U904 ( .A0(n3592), .A1(n829), .B0(n1648), .C0(n1649), .Y(n2649)
         );
  OAI211XLTS U905 ( .A0(n3592), .A1(n828), .B0(n1646), .C0(n1647), .Y(n2650)
         );
  OAI211XLTS U906 ( .A0(n3591), .A1(n827), .B0(n1644), .C0(n1645), .Y(n2651)
         );
  OAI211XLTS U907 ( .A0(n3591), .A1(n826), .B0(n1642), .C0(n1643), .Y(n2652)
         );
  OAI211XLTS U908 ( .A0(n3591), .A1(n825), .B0(n1640), .C0(n1641), .Y(n2653)
         );
  OAI211XLTS U909 ( .A0(n3591), .A1(n824), .B0(n1638), .C0(n1639), .Y(n2654)
         );
  OAI211XLTS U910 ( .A0(n3590), .A1(n823), .B0(n1636), .C0(n1637), .Y(n2655)
         );
  OAI211XLTS U911 ( .A0(n3590), .A1(n822), .B0(n1634), .C0(n1635), .Y(n2656)
         );
  OAI211XLTS U912 ( .A0(n3590), .A1(n821), .B0(n1632), .C0(n1633), .Y(n2657)
         );
  OAI211XLTS U913 ( .A0(n3589), .A1(n820), .B0(n1626), .C0(n1627), .Y(n2660)
         );
  OAI211XLTS U914 ( .A0(n3589), .A1(n819), .B0(n1624), .C0(n1625), .Y(n2661)
         );
  OAI211XLTS U915 ( .A0(n3588), .A1(n818), .B0(n1622), .C0(n1623), .Y(n2662)
         );
  OAI211XLTS U916 ( .A0(n3588), .A1(n817), .B0(n1618), .C0(n1619), .Y(n2664)
         );
  OAI211XLTS U917 ( .A0(n3588), .A1(n816), .B0(n1616), .C0(n1617), .Y(n2665)
         );
  OAI211XLTS U918 ( .A0(n3587), .A1(n815), .B0(n1614), .C0(n1615), .Y(n2666)
         );
  OAI211XLTS U919 ( .A0(n3587), .A1(n814), .B0(n1612), .C0(n1613), .Y(n2667)
         );
  OAI211XLTS U920 ( .A0(n3587), .A1(n813), .B0(n1610), .C0(n1611), .Y(n2668)
         );
  OAI211XLTS U921 ( .A0(n3587), .A1(n812), .B0(n1608), .C0(n1609), .Y(n2669)
         );
  OAI211XLTS U922 ( .A0(n3586), .A1(n811), .B0(n1606), .C0(n1607), .Y(n2670)
         );
  OAI211XLTS U923 ( .A0(n3586), .A1(n810), .B0(n1604), .C0(n1605), .Y(n2671)
         );
  OAI211XLTS U924 ( .A0(n3586), .A1(n809), .B0(n1602), .C0(n1603), .Y(n2672)
         );
  OAI211XLTS U925 ( .A0(n3585), .A1(n808), .B0(n1598), .C0(n1599), .Y(n2674)
         );
  OAI211XLTS U926 ( .A0(n3594), .A1(n838), .B0(n1926), .C0(n1927), .Y(n2531)
         );
  OAI211XLTS U927 ( .A0(n3594), .A1(n837), .B0(n1924), .C0(n1925), .Y(n2532)
         );
  OAI211XLTS U928 ( .A0(n3594), .A1(n836), .B0(n1922), .C0(n1923), .Y(n2533)
         );
  OAI211XLTS U929 ( .A0(n3594), .A1(n835), .B0(n1920), .C0(n1921), .Y(n2534)
         );
  OAI211XLTS U930 ( .A0(n3125), .A1(n675), .B0(n1721), .C0(n1722), .Y(n2613)
         );
  OAI211XLTS U931 ( .A0(n3126), .A1(n674), .B0(n1709), .C0(n1710), .Y(n2619)
         );
  OAI211XLTS U932 ( .A0(n3127), .A1(n673), .B0(n1705), .C0(n1706), .Y(n2621)
         );
  OAI211XLTS U933 ( .A0(n3127), .A1(n672), .B0(n1703), .C0(n1704), .Y(n2622)
         );
  OAI211XLTS U934 ( .A0(n3129), .A1(n671), .B0(n1689), .C0(n1690), .Y(n2629)
         );
  OAI211XLTS U935 ( .A0(n3129), .A1(n670), .B0(n1687), .C0(n1688), .Y(n2630)
         );
  OAI211XLTS U936 ( .A0(n3129), .A1(n669), .B0(n1683), .C0(n1684), .Y(n2632)
         );
  OAI211XLTS U937 ( .A0(n3130), .A1(n668), .B0(n1675), .C0(n1676), .Y(n2636)
         );
  OAI211XLTS U938 ( .A0(n3125), .A1(n662), .B0(n1719), .C0(n1720), .Y(n2614)
         );
  OAI211XLTS U939 ( .A0(n3125), .A1(n661), .B0(n1717), .C0(n1718), .Y(n2615)
         );
  OAI211XLTS U940 ( .A0(n3125), .A1(n660), .B0(n1715), .C0(n1716), .Y(n2616)
         );
  OAI211XLTS U941 ( .A0(n3126), .A1(n659), .B0(n1711), .C0(n1712), .Y(n2618)
         );
  OAI211XLTS U942 ( .A0(n3126), .A1(n658), .B0(n1707), .C0(n1708), .Y(n2620)
         );
  OAI211XLTS U943 ( .A0(n3127), .A1(n657), .B0(n1701), .C0(n1702), .Y(n2623)
         );
  OAI211XLTS U944 ( .A0(n3128), .A1(n656), .B0(n1697), .C0(n1698), .Y(n2625)
         );
  OAI211XLTS U945 ( .A0(n3128), .A1(n655), .B0(n1695), .C0(n1696), .Y(n2626)
         );
  OAI211XLTS U946 ( .A0(n3128), .A1(n654), .B0(n1693), .C0(n1694), .Y(n2627)
         );
  OAI211XLTS U947 ( .A0(n3128), .A1(n653), .B0(n1691), .C0(n1692), .Y(n2628)
         );
  OAI211XLTS U948 ( .A0(n3129), .A1(n652), .B0(n1685), .C0(n1686), .Y(n2631)
         );
  OAI211XLTS U949 ( .A0(n3130), .A1(n651), .B0(n1681), .C0(n1682), .Y(n2633)
         );
  OAI211XLTS U950 ( .A0(n3130), .A1(n650), .B0(n1679), .C0(n1680), .Y(n2634)
         );
  OAI211XLTS U951 ( .A0(n3130), .A1(n649), .B0(n1677), .C0(n1678), .Y(n2635)
         );
  OAI211XLTS U952 ( .A0(n3131), .A1(n648), .B0(n1673), .C0(n1674), .Y(n2637)
         );
  OAI211XLTS U953 ( .A0(n3126), .A1(n608), .B0(n1713), .C0(n1714), .Y(n2617)
         );
  OAI211XLTS U954 ( .A0(n3127), .A1(n607), .B0(n1699), .C0(n1700), .Y(n2624)
         );
  OAI211XLTS U955 ( .A0(n3131), .A1(n606), .B0(n1671), .C0(n1672), .Y(n2638)
         );
  OAI211XLTS U956 ( .A0(n3131), .A1(n647), .B0(n1669), .C0(n1670), .Y(n2639)
         );
  OAI211XLTS U957 ( .A0(n3131), .A1(n646), .B0(n1667), .C0(n1668), .Y(n2640)
         );
  OAI211XLTS U958 ( .A0(n3585), .A1(n890), .B0(n1191), .C0(n1192), .Y(n2868)
         );
  OAI211XLTS U959 ( .A0(n3585), .A1(n893), .B0(n1197), .C0(n1198), .Y(n2865)
         );
  OAI211XLTS U960 ( .A0(n3585), .A1(n892), .B0(n1195), .C0(n1196), .Y(n2866)
         );
  OAI211XLTS U961 ( .A0(n3589), .A1(n888), .B0(n1183), .C0(n1184), .Y(n2870)
         );
  OAI211XLTS U962 ( .A0(n3328), .A1(n881), .B0(n1396), .C0(n1397), .Y(n2775)
         );
  OAI211XLTS U963 ( .A0(n3327), .A1(n880), .B0(n1386), .C0(n1387), .Y(n2780)
         );
  OAI211XLTS U964 ( .A0(n3327), .A1(n879), .B0(n1382), .C0(n1383), .Y(n2782)
         );
  OAI211XLTS U965 ( .A0(n3326), .A1(n878), .B0(n1380), .C0(n1381), .Y(n2783)
         );
  OAI211XLTS U966 ( .A0(n3324), .A1(n877), .B0(n1362), .C0(n1363), .Y(n2792)
         );
  OAI211XLTS U967 ( .A0(n3323), .A1(n876), .B0(n1358), .C0(n1359), .Y(n2794)
         );
  OAI211XLTS U968 ( .A0(n3323), .A1(n875), .B0(n1352), .C0(n1353), .Y(n2797)
         );
  OAI211XLTS U969 ( .A0(n3322), .A1(n874), .B0(n1346), .C0(n1347), .Y(n2800)
         );
  OAI211XLTS U970 ( .A0(n3329), .A1(n868), .B0(n1404), .C0(n1405), .Y(n2771)
         );
  OAI211XLTS U971 ( .A0(n3329), .A1(n867), .B0(n1402), .C0(n1403), .Y(n2772)
         );
  OAI211XLTS U972 ( .A0(n3329), .A1(n866), .B0(n1400), .C0(n1401), .Y(n2773)
         );
  OAI211XLTS U973 ( .A0(n3329), .A1(n865), .B0(n1398), .C0(n1399), .Y(n2774)
         );
  OAI211XLTS U974 ( .A0(n3328), .A1(n864), .B0(n1394), .C0(n1395), .Y(n2776)
         );
  OAI211XLTS U975 ( .A0(n3328), .A1(n863), .B0(n1392), .C0(n1393), .Y(n2777)
         );
  OAI211XLTS U976 ( .A0(n3328), .A1(n862), .B0(n1390), .C0(n1391), .Y(n2778)
         );
  OAI211XLTS U977 ( .A0(n3327), .A1(n861), .B0(n1388), .C0(n1389), .Y(n2779)
         );
  OAI211XLTS U978 ( .A0(n3327), .A1(n860), .B0(n1384), .C0(n1385), .Y(n2781)
         );
  OAI211XLTS U979 ( .A0(n3326), .A1(n859), .B0(n1378), .C0(n1379), .Y(n2784)
         );
  OAI211XLTS U980 ( .A0(n3326), .A1(n858), .B0(n1376), .C0(n1377), .Y(n2785)
         );
  OAI211XLTS U981 ( .A0(n3326), .A1(n857), .B0(n1374), .C0(n1375), .Y(n2786)
         );
  OAI211XLTS U982 ( .A0(n3325), .A1(n856), .B0(n1372), .C0(n1373), .Y(n2787)
         );
  OAI211XLTS U983 ( .A0(n3325), .A1(n855), .B0(n1370), .C0(n1371), .Y(n2788)
         );
  OAI211XLTS U984 ( .A0(n3325), .A1(n854), .B0(n1368), .C0(n1369), .Y(n2789)
         );
  OAI211XLTS U985 ( .A0(n3324), .A1(n853), .B0(n1366), .C0(n1367), .Y(n2790)
         );
  OAI211XLTS U986 ( .A0(n3324), .A1(n852), .B0(n1364), .C0(n1365), .Y(n2791)
         );
  OAI211XLTS U987 ( .A0(n3324), .A1(n851), .B0(n1360), .C0(n1361), .Y(n2793)
         );
  OAI211XLTS U988 ( .A0(n3323), .A1(n850), .B0(n1356), .C0(n1357), .Y(n2795)
         );
  OAI211XLTS U989 ( .A0(n3323), .A1(n849), .B0(n1354), .C0(n1355), .Y(n2796)
         );
  OAI211XLTS U990 ( .A0(n3322), .A1(n848), .B0(n1350), .C0(n1351), .Y(n2798)
         );
  OAI211XLTS U991 ( .A0(n3322), .A1(n847), .B0(n1348), .C0(n1349), .Y(n2799)
         );
  OAI211XLTS U992 ( .A0(n3322), .A1(n846), .B0(n1344), .C0(n1345), .Y(n2801)
         );
  OAI211XLTS U993 ( .A0(n3321), .A1(n845), .B0(n1342), .C0(n1343), .Y(n2802)
         );
  OAI211XLTS U994 ( .A0(n3321), .A1(n897), .B0(n1255), .C0(n1256), .Y(n2844)
         );
  OAI211XLTS U995 ( .A0(n3321), .A1(n900), .B0(n1261), .C0(n1262), .Y(n2841)
         );
  OAI211XLTS U996 ( .A0(n3321), .A1(n899), .B0(n1259), .C0(n1260), .Y(n2842)
         );
  OAI211XLTS U997 ( .A0(n3325), .A1(n895), .B0(n1247), .C0(n1248), .Y(n2846)
         );
  OAI211XLTS U998 ( .A0(n3330), .A1(n872), .B0(n2019), .C0(n2020), .Y(n2475)
         );
  OAI211XLTS U999 ( .A0(n3330), .A1(n871), .B0(n2017), .C0(n2018), .Y(n2476)
         );
  OAI211XLTS U1000 ( .A0(n3330), .A1(n870), .B0(n2015), .C0(n2016), .Y(n2477)
         );
  OAI211XLTS U1001 ( .A0(n3330), .A1(n869), .B0(n2013), .C0(n2014), .Y(n2478)
         );
  OAI211XLTS U1002 ( .A0(n3132), .A1(n667), .B0(n1665), .C0(n1666), .Y(n2641)
         );
  OAI211XLTS U1003 ( .A0(n3132), .A1(n645), .B0(n1663), .C0(n1664), .Y(n2642)
         );
  OAI211XLTS U1004 ( .A0(n4041), .A1(n3510), .B0(n1213), .C0(n1214), .Y(n2859)
         );
  OAI211XLTS U1005 ( .A0(n4038), .A1(n3510), .B0(n1211), .C0(n1212), .Y(n2860)
         );
  OAI211XLTS U1006 ( .A0(n4035), .A1(n3511), .B0(n1209), .C0(n1210), .Y(n2861)
         );
  OAI211XLTS U1007 ( .A0(n4032), .A1(n3511), .B0(n1207), .C0(n1208), .Y(n2862)
         );
  OAI211XLTS U1008 ( .A0(n4029), .A1(n3511), .B0(n1205), .C0(n1206), .Y(n2863)
         );
  OAI211XLTS U1009 ( .A0(n4026), .A1(n3511), .B0(n1200), .C0(n1201), .Y(n2864)
         );
  OAI211XLTS U1010 ( .A0(n4035), .A1(n3446), .B0(n1224), .C0(n1225), .Y(n2855)
         );
  OAI211XLTS U1011 ( .A0(n4032), .A1(n3446), .B0(n1222), .C0(n1223), .Y(n2856)
         );
  OAI211XLTS U1012 ( .A0(n4029), .A1(n3446), .B0(n1220), .C0(n1221), .Y(n2857)
         );
  OAI211XLTS U1013 ( .A0(n4026), .A1(n3446), .B0(n1216), .C0(n1217), .Y(n2858)
         );
  OAI211XLTS U1014 ( .A0(n4038), .A1(n3445), .B0(n1226), .C0(n1227), .Y(n2854)
         );
  OAI211XLTS U1015 ( .A0(n4041), .A1(n3445), .B0(n1228), .C0(n1229), .Y(n2853)
         );
  OAI211XLTS U1016 ( .A0(n3595), .A1(n807), .B0(n1928), .C0(n1929), .Y(n2530)
         );
  INVXLTS U1017 ( .A(n3599), .Y(n3595) );
  OAI211XLTS U1018 ( .A0(n3331), .A1(n844), .B0(n2021), .C0(n2022), .Y(n2474)
         );
  INVXLTS U1019 ( .A(n3334), .Y(n3331) );
  OAI211XLTS U1020 ( .A0(n3738), .A1(n686), .B0(n1160), .C0(n1161), .Y(n2879)
         );
  OAI211XLTS U1021 ( .A0(n3739), .A1(n685), .B0(n1156), .C0(n1157), .Y(n2881)
         );
  OAI211XLTS U1022 ( .A0(n3740), .A1(n644), .B0(n1877), .C0(n1878), .Y(n2557)
         );
  OAI211XLTS U1023 ( .A0(n3743), .A1(n689), .B0(n1164), .C0(n1165), .Y(n2877)
         );
  OAI211XLTS U1024 ( .A0(n3747), .A1(n688), .B0(n1162), .C0(n1163), .Y(n2878)
         );
  OAI211XLTS U1025 ( .A0(n3747), .A1(n687), .B0(n1158), .C0(n1159), .Y(n2880)
         );
  OAI211XLTS U1026 ( .A0(n3733), .A1(n684), .B0(n1149), .C0(n1150), .Y(n2882)
         );
  OAI211XLTS U1027 ( .A0(n3737), .A1(n640), .B0(n1789), .C0(n1790), .Y(n2579)
         );
  OAI211XLTS U1028 ( .A0(n3737), .A1(n639), .B0(n1787), .C0(n1788), .Y(n2580)
         );
  OAI211XLTS U1029 ( .A0(n3736), .A1(n638), .B0(n1785), .C0(n1786), .Y(n2581)
         );
  OAI211XLTS U1030 ( .A0(n3736), .A1(n637), .B0(n1783), .C0(n1784), .Y(n2582)
         );
  OAI211XLTS U1031 ( .A0(n3736), .A1(n636), .B0(n1781), .C0(n1782), .Y(n2583)
         );
  OAI211XLTS U1032 ( .A0(n3736), .A1(n635), .B0(n1779), .C0(n1780), .Y(n2584)
         );
  OAI211XLTS U1033 ( .A0(n3735), .A1(n634), .B0(n1777), .C0(n1778), .Y(n2585)
         );
  OAI211XLTS U1034 ( .A0(n3735), .A1(n633), .B0(n1775), .C0(n1776), .Y(n2586)
         );
  OAI211XLTS U1035 ( .A0(n3735), .A1(n632), .B0(n1773), .C0(n1774), .Y(n2587)
         );
  OAI211XLTS U1036 ( .A0(n3735), .A1(n631), .B0(n1771), .C0(n1772), .Y(n2588)
         );
  OAI211XLTS U1037 ( .A0(n3734), .A1(n630), .B0(n1769), .C0(n1770), .Y(n2589)
         );
  OAI211XLTS U1038 ( .A0(n3734), .A1(n629), .B0(n1767), .C0(n1768), .Y(n2590)
         );
  OAI211XLTS U1039 ( .A0(n3734), .A1(n628), .B0(n1765), .C0(n1766), .Y(n2591)
         );
  OAI211XLTS U1040 ( .A0(n3734), .A1(n627), .B0(n1763), .C0(n1764), .Y(n2592)
         );
  OAI211XLTS U1041 ( .A0(n3733), .A1(n626), .B0(n1761), .C0(n1762), .Y(n2593)
         );
  OAI211XLTS U1042 ( .A0(n3733), .A1(n625), .B0(n1759), .C0(n1760), .Y(n2594)
         );
  OAI211XLTS U1043 ( .A0(n3733), .A1(n624), .B0(n1757), .C0(n1758), .Y(n2595)
         );
  OAI211XLTS U1044 ( .A0(n3732), .A1(n623), .B0(n1755), .C0(n1756), .Y(n2596)
         );
  OAI211XLTS U1045 ( .A0(n3732), .A1(n622), .B0(n1753), .C0(n1754), .Y(n2597)
         );
  OAI211XLTS U1046 ( .A0(n3732), .A1(n621), .B0(n1751), .C0(n1752), .Y(n2598)
         );
  OAI211XLTS U1047 ( .A0(n3732), .A1(n620), .B0(n1749), .C0(n1750), .Y(n2599)
         );
  OAI211XLTS U1048 ( .A0(n3731), .A1(n619), .B0(n1747), .C0(n1748), .Y(n2600)
         );
  OAI211XLTS U1049 ( .A0(n3731), .A1(n618), .B0(n1745), .C0(n1746), .Y(n2601)
         );
  OAI211XLTS U1050 ( .A0(n3731), .A1(n617), .B0(n1743), .C0(n1744), .Y(n2602)
         );
  OAI211XLTS U1051 ( .A0(n3731), .A1(n616), .B0(n1741), .C0(n1742), .Y(n2603)
         );
  OAI211XLTS U1052 ( .A0(n3743), .A1(n615), .B0(n1739), .C0(n1740), .Y(n2604)
         );
  OAI211XLTS U1053 ( .A0(n3740), .A1(n614), .B0(n1737), .C0(n1738), .Y(n2605)
         );
  OAI211XLTS U1054 ( .A0(n3741), .A1(n613), .B0(n1735), .C0(n1736), .Y(n2606)
         );
  OAI211XLTS U1055 ( .A0(n3742), .A1(n612), .B0(n1733), .C0(n1734), .Y(n2607)
         );
  OAI211XLTS U1056 ( .A0(n3741), .A1(n611), .B0(n1731), .C0(n1732), .Y(n2608)
         );
  OAI211XLTS U1057 ( .A0(n3742), .A1(n610), .B0(n1729), .C0(n1730), .Y(n2609)
         );
  OAI211XLTS U1058 ( .A0(n3739), .A1(n609), .B0(n1727), .C0(n1728), .Y(n2610)
         );
  OAI211XLTS U1059 ( .A0(n3737), .A1(n665), .B0(n1867), .C0(n1868), .Y(n2562)
         );
  OAI211XLTS U1060 ( .A0(n3738), .A1(n643), .B0(n1873), .C0(n1874), .Y(n2559)
         );
  OAI211XLTS U1061 ( .A0(n3738), .A1(n642), .B0(n1871), .C0(n1872), .Y(n2560)
         );
  OAI211XLTS U1062 ( .A0(n3737), .A1(n641), .B0(n1869), .C0(n1870), .Y(n2561)
         );
  OAI211XLTS U1063 ( .A0(n3738), .A1(n666), .B0(n1875), .C0(n1876), .Y(n2558)
         );
  INVXLTS U1064 ( .A(selectBit_EAST), .Y(n1031) );
  AOI32XLTS U1065 ( .A0(n481), .A1(n1848), .A2(n1849), .B0(n3827), .B1(n768), 
        .Y(n2565) );
  NAND2XLTS U1066 ( .A(readIn_SOUTH), .B(n1854), .Y(n1848) );
  AOI32XLTS U1067 ( .A0(n45), .A1(n1862), .A2(n1863), .B0(n3912), .B1(n683), 
        .Y(n2563) );
  AOI21XLTS U1068 ( .A0(readIn_NORTH), .A1(n1864), .B0(n1865), .Y(n1863) );
  INVXLTS U1069 ( .A(selectBit_WEST), .Y(n1086) );
  NAND4XLTS U1070 ( .A(n488), .B(n468), .C(n1031), .D(n915), .Y(n2074) );
  NAND2XLTS U1071 ( .A(n485), .B(readReady), .Y(n2952) );
  NAND4XLTS U1072 ( .A(n462), .B(n925), .C(n1031), .D(n1086), .Y(n2077) );
  NAND4XLTS U1073 ( .A(n485), .B(n925), .C(n1132), .D(n1031), .Y(n2076) );
  NAND3XLTS U1074 ( .A(n925), .B(n468), .C(n483), .Y(n2075) );
  OAI32XLTS U1075 ( .A0(n4843), .A1(n2067), .A2(n2068), .B0(n2069), .B1(n2070), 
        .Y(n2450) );
  NAND4XLTS U1076 ( .A(selectBit_NORTH), .B(n468), .C(n1031), .D(n985), .Y(
        n2073) );
  CLKBUFX2TS U1077 ( .A(n5323), .Y(n979) );
  CLKBUFX2TS U1078 ( .A(n5327), .Y(n986) );
  NAND2X1TS U1079 ( .A(n5326), .B(n157), .Y(n2025) );
  NAND3X1TS U1080 ( .A(n124), .B(n128), .C(n4), .Y(n2084) );
  NAND3X1TS U1081 ( .A(n1), .B(n128), .C(n8), .Y(n2086) );
  NAND3X1TS U1082 ( .A(n44), .B(n129), .C(n8), .Y(n2085) );
  NAND3X1TS U1083 ( .A(n9), .B(n466), .C(n44), .Y(n2083) );
  CLKBUFX2TS U1084 ( .A(n3772), .Y(n3767) );
  CLKBUFX2TS U1085 ( .A(n3770), .Y(n3765) );
  CLKBUFX2TS U1086 ( .A(n3771), .Y(n3764) );
  CLKBUFX2TS U1087 ( .A(n3770), .Y(n3768) );
  CLKBUFX2TS U1088 ( .A(n3770), .Y(n3766) );
  CLKBUFX2TS U1089 ( .A(n3771), .Y(n3763) );
  CLKBUFX2TS U1090 ( .A(n3942), .Y(n3933) );
  CLKBUFX2TS U1091 ( .A(n3843), .Y(n3834) );
  CLKBUFX2TS U1092 ( .A(n3941), .Y(n3936) );
  CLKBUFX2TS U1093 ( .A(n3940), .Y(n3939) );
  CLKBUFX2TS U1094 ( .A(n3940), .Y(n3938) );
  CLKBUFX2TS U1095 ( .A(n3944), .Y(n3937) );
  CLKBUFX2TS U1096 ( .A(n3941), .Y(n3935) );
  CLKBUFX2TS U1097 ( .A(n3942), .Y(n3934) );
  CLKBUFX2TS U1098 ( .A(n3842), .Y(n3836) );
  CLKBUFX2TS U1099 ( .A(n3842), .Y(n3837) );
  CLKBUFX2TS U1100 ( .A(n3841), .Y(n3839) );
  CLKBUFX2TS U1101 ( .A(n3841), .Y(n3838) );
  CLKBUFX2TS U1102 ( .A(n3843), .Y(n3835) );
  CLKBUFX2TS U1103 ( .A(n3945), .Y(n3940) );
  CLKBUFX2TS U1104 ( .A(n3944), .Y(n3941) );
  CLKBUFX2TS U1105 ( .A(n3944), .Y(n3942) );
  CLKBUFX2TS U1106 ( .A(n3845), .Y(n3842) );
  CLKBUFX2TS U1107 ( .A(n3846), .Y(n3840) );
  CLKBUFX2TS U1108 ( .A(n3846), .Y(n3841) );
  CLKBUFX2TS U1109 ( .A(n3845), .Y(n3843) );
  CLKBUFX2TS U1110 ( .A(n3773), .Y(n3770) );
  CLKBUFX2TS U1111 ( .A(n3773), .Y(n3771) );
  CLKBUFX2TS U1112 ( .A(n3150), .Y(n3148) );
  CLKBUFX2TS U1113 ( .A(n3898), .Y(n3896) );
  CLKBUFX2TS U1114 ( .A(n3899), .Y(n3895) );
  CLKBUFX2TS U1115 ( .A(n3899), .Y(n3894) );
  CLKBUFX2TS U1116 ( .A(n3900), .Y(n3893) );
  CLKBUFX2TS U1117 ( .A(n3900), .Y(n3892) );
  CLKBUFX2TS U1118 ( .A(n3901), .Y(n3891) );
  CLKBUFX2TS U1119 ( .A(n3901), .Y(n3890) );
  CLKBUFX2TS U1120 ( .A(n3898), .Y(n3897) );
  CLKBUFX2TS U1121 ( .A(n3797), .Y(n3795) );
  CLKBUFX2TS U1122 ( .A(n3798), .Y(n3794) );
  CLKBUFX2TS U1123 ( .A(n3799), .Y(n3793) );
  CLKBUFX2TS U1124 ( .A(n3799), .Y(n3792) );
  CLKBUFX2TS U1125 ( .A(n3800), .Y(n3791) );
  CLKBUFX2TS U1126 ( .A(n3797), .Y(n3796) );
  CLKBUFX2TS U1127 ( .A(n3153), .Y(n3143) );
  CLKBUFX2TS U1128 ( .A(n3153), .Y(n3142) );
  CLKBUFX2TS U1129 ( .A(n3154), .Y(n3141) );
  CLKBUFX2TS U1130 ( .A(n3151), .Y(n3147) );
  CLKBUFX2TS U1131 ( .A(n3151), .Y(n3146) );
  CLKBUFX2TS U1132 ( .A(n3152), .Y(n3145) );
  CLKBUFX2TS U1133 ( .A(n3152), .Y(n3144) );
  CLKBUFX2TS U1134 ( .A(n3154), .Y(n3140) );
  CLKBUFX2TS U1135 ( .A(n3787), .Y(n3777) );
  CLKBUFX2TS U1136 ( .A(n3786), .Y(n3778) );
  CLKBUFX2TS U1137 ( .A(n3785), .Y(n3780) );
  CLKBUFX2TS U1138 ( .A(n3787), .Y(n3776) );
  CLKBUFX2TS U1139 ( .A(n3786), .Y(n3779) );
  CLKBUFX2TS U1140 ( .A(n3150), .Y(n3149) );
  CLKBUFX2TS U1141 ( .A(n3498), .Y(n3484) );
  CLKBUFX2TS U1142 ( .A(n3498), .Y(n3485) );
  CLKBUFX2TS U1143 ( .A(n3382), .Y(n3367) );
  CLKBUFX2TS U1144 ( .A(n3382), .Y(n3368) );
  CLKBUFX2TS U1145 ( .A(n3772), .Y(n3762) );
  CLKBUFX2TS U1146 ( .A(n3773), .Y(n3772) );
  CLKBUFX2TS U1147 ( .A(n3497), .Y(n3486) );
  CLKBUFX2TS U1148 ( .A(n3381), .Y(n3369) );
  CLKBUFX2TS U1149 ( .A(n3497), .Y(n3487) );
  CLKBUFX2TS U1150 ( .A(n3496), .Y(n3488) );
  CLKBUFX2TS U1151 ( .A(n3496), .Y(n3489) );
  CLKBUFX2TS U1152 ( .A(n3495), .Y(n3490) );
  CLKBUFX2TS U1153 ( .A(n3495), .Y(n3491) );
  CLKBUFX2TS U1154 ( .A(n3494), .Y(n3492) );
  CLKBUFX2TS U1155 ( .A(n3886), .Y(n3877) );
  CLKBUFX2TS U1156 ( .A(n3886), .Y(n3878) );
  CLKBUFX2TS U1157 ( .A(n3885), .Y(n3879) );
  CLKBUFX2TS U1158 ( .A(n3885), .Y(n3880) );
  CLKBUFX2TS U1159 ( .A(n3886), .Y(n3881) );
  CLKBUFX2TS U1160 ( .A(n3884), .Y(n3882) );
  CLKBUFX2TS U1161 ( .A(n3380), .Y(n3371) );
  CLKBUFX2TS U1162 ( .A(n3379), .Y(n3374) );
  CLKBUFX2TS U1163 ( .A(n3378), .Y(n3376) );
  CLKBUFX2TS U1164 ( .A(n3380), .Y(n3372) );
  CLKBUFX2TS U1165 ( .A(n3378), .Y(n3375) );
  CLKBUFX2TS U1166 ( .A(n3379), .Y(n3373) );
  CLKBUFX2TS U1167 ( .A(n3381), .Y(n3370) );
  CLKBUFX2TS U1168 ( .A(n3494), .Y(n3493) );
  CLKBUFX2TS U1169 ( .A(n3785), .Y(n3781) );
  CLKBUFX2TS U1170 ( .A(n3814), .Y(n3805) );
  CLKBUFX2TS U1171 ( .A(n3784), .Y(n3782) );
  CLKBUFX2TS U1172 ( .A(n3814), .Y(n3806) );
  CLKBUFX2TS U1173 ( .A(n3813), .Y(n3807) );
  CLKBUFX2TS U1174 ( .A(n3813), .Y(n3808) );
  CLKBUFX2TS U1175 ( .A(n3812), .Y(n3809) );
  CLKBUFX2TS U1176 ( .A(n3816), .Y(n3810) );
  CLKBUFX2TS U1177 ( .A(n3812), .Y(n3811) );
  CLKBUFX2TS U1178 ( .A(n3784), .Y(n3783) );
  CLKBUFX2TS U1179 ( .A(n3943), .Y(n3932) );
  CLKBUFX2TS U1180 ( .A(n3944), .Y(n3943) );
  CLKBUFX2TS U1181 ( .A(n3844), .Y(n3833) );
  CLKBUFX2TS U1182 ( .A(n3845), .Y(n3844) );
  CLKBUFX2TS U1183 ( .A(n3929), .Y(n3921) );
  CLKBUFX2TS U1184 ( .A(n3929), .Y(n3922) );
  CLKBUFX2TS U1185 ( .A(n3930), .Y(n3919) );
  CLKBUFX2TS U1186 ( .A(n784), .Y(n3920) );
  CLKBUFX2TS U1187 ( .A(n3928), .Y(n3923) );
  CLKBUFX2TS U1188 ( .A(n3928), .Y(n3924) );
  CLKBUFX2TS U1189 ( .A(n3927), .Y(n3925) );
  CLKBUFX2TS U1190 ( .A(n3927), .Y(n3926) );
  INVX2TS U1191 ( .A(n4571), .Y(n4572) );
  CLKBUFX2TS U1192 ( .A(n3858), .Y(n3847) );
  CLKBUFX2TS U1193 ( .A(n3858), .Y(n3848) );
  CLKBUFX2TS U1194 ( .A(n3855), .Y(n3854) );
  CLKBUFX2TS U1195 ( .A(n3857), .Y(n3849) );
  CLKBUFX2TS U1196 ( .A(n3856), .Y(n3851) );
  CLKBUFX2TS U1197 ( .A(n3857), .Y(n3850) );
  CLKBUFX2TS U1198 ( .A(n3855), .Y(n3853) );
  CLKBUFX2TS U1199 ( .A(n3856), .Y(n3852) );
  INVX2TS U1200 ( .A(n4571), .Y(n4573) );
  CLKBUFX2TS U1201 ( .A(n3452), .Y(n3447) );
  CLKBUFX2TS U1202 ( .A(n3452), .Y(n3448) );
  CLKBUFX2TS U1203 ( .A(n3452), .Y(n3449) );
  CLKBUFX2TS U1204 ( .A(n3816), .Y(n3813) );
  CLKBUFX2TS U1205 ( .A(n3499), .Y(n3496) );
  CLKBUFX2TS U1206 ( .A(n3817), .Y(n3812) );
  CLKBUFX2TS U1207 ( .A(n1202), .Y(n3495) );
  CLKBUFX2TS U1208 ( .A(n3816), .Y(n3814) );
  CLKBUFX2TS U1209 ( .A(n3499), .Y(n3497) );
  CLKBUFX2TS U1210 ( .A(n1202), .Y(n3494) );
  CLKBUFX2TS U1211 ( .A(n3888), .Y(n3886) );
  CLKBUFX2TS U1212 ( .A(n3888), .Y(n3885) );
  CLKBUFX2TS U1213 ( .A(n3889), .Y(n3884) );
  CLKBUFX2TS U1214 ( .A(n3903), .Y(n3899) );
  CLKBUFX2TS U1215 ( .A(n3903), .Y(n3900) );
  CLKBUFX2TS U1216 ( .A(n3902), .Y(n3901) );
  CLKBUFX2TS U1217 ( .A(n3903), .Y(n3898) );
  CLKBUFX2TS U1218 ( .A(n3802), .Y(n3798) );
  CLKBUFX2TS U1219 ( .A(n3802), .Y(n3799) );
  CLKBUFX2TS U1220 ( .A(n798), .Y(n3800) );
  CLKBUFX2TS U1221 ( .A(n3802), .Y(n3797) );
  CLKBUFX2TS U1222 ( .A(n3383), .Y(n3380) );
  CLKBUFX2TS U1223 ( .A(n3383), .Y(n3378) );
  CLKBUFX2TS U1224 ( .A(n1233), .Y(n3379) );
  CLKBUFX2TS U1225 ( .A(n3383), .Y(n3381) );
  CLKBUFX2TS U1226 ( .A(n1233), .Y(n3377) );
  CLKBUFX2TS U1227 ( .A(n3789), .Y(n3784) );
  CLKBUFX2TS U1228 ( .A(n3789), .Y(n3785) );
  CLKBUFX2TS U1229 ( .A(n3786), .Y(n3787) );
  CLKBUFX2TS U1230 ( .A(n3789), .Y(n3786) );
  CLKBUFX2TS U1231 ( .A(n3499), .Y(n3498) );
  CLKBUFX2TS U1232 ( .A(n3383), .Y(n3382) );
  CLKBUFX2TS U1233 ( .A(n3931), .Y(n3929) );
  CLKBUFX2TS U1234 ( .A(n3931), .Y(n3928) );
  CLKBUFX2TS U1235 ( .A(n3931), .Y(n3927) );
  CLKBUFX2TS U1236 ( .A(n1267), .Y(n3153) );
  CLKBUFX2TS U1237 ( .A(n3156), .Y(n3151) );
  CLKBUFX2TS U1238 ( .A(n3156), .Y(n3152) );
  CLKBUFX2TS U1239 ( .A(n1267), .Y(n3154) );
  CLKBUFX2TS U1240 ( .A(n3156), .Y(n3155) );
  CLKBUFX2TS U1241 ( .A(n783), .Y(n3945) );
  CLKBUFX2TS U1242 ( .A(n783), .Y(n3944) );
  CLKBUFX2TS U1243 ( .A(n181), .Y(n3846) );
  CLKBUFX2TS U1244 ( .A(n181), .Y(n3845) );
  CLKBUFX2TS U1245 ( .A(n801), .Y(n3773) );
  CLKBUFX2TS U1246 ( .A(n3267), .Y(n3253) );
  CLKBUFX2TS U1247 ( .A(n3532), .Y(n3518) );
  CLKBUFX2TS U1248 ( .A(n3433), .Y(n3419) );
  CLKBUFX2TS U1249 ( .A(n3156), .Y(n3150) );
  CLKBUFX2TS U1250 ( .A(n3267), .Y(n3254) );
  CLKBUFX2TS U1251 ( .A(n3532), .Y(n3519) );
  CLKBUFX2TS U1252 ( .A(n3433), .Y(n3420) );
  CLKBUFX2TS U1253 ( .A(n3264), .Y(n3260) );
  CLKBUFX2TS U1254 ( .A(n3264), .Y(n3259) );
  CLKBUFX2TS U1255 ( .A(n3265), .Y(n3258) );
  CLKBUFX2TS U1256 ( .A(n3265), .Y(n3257) );
  CLKBUFX2TS U1257 ( .A(n3268), .Y(n3256) );
  CLKBUFX2TS U1258 ( .A(n3266), .Y(n3255) );
  CLKBUFX2TS U1259 ( .A(n3263), .Y(n3261) );
  CLKBUFX2TS U1260 ( .A(n3531), .Y(n3527) );
  CLKBUFX2TS U1261 ( .A(n3531), .Y(n3526) );
  CLKBUFX2TS U1262 ( .A(n3529), .Y(n3525) );
  CLKBUFX2TS U1263 ( .A(n3530), .Y(n3523) );
  CLKBUFX2TS U1264 ( .A(n3530), .Y(n3522) );
  CLKBUFX2TS U1265 ( .A(n3529), .Y(n3524) );
  CLKBUFX2TS U1266 ( .A(n3531), .Y(n3521) );
  CLKBUFX2TS U1267 ( .A(n3531), .Y(n3520) );
  CLKBUFX2TS U1268 ( .A(n3430), .Y(n3426) );
  CLKBUFX2TS U1269 ( .A(n3430), .Y(n3425) );
  CLKBUFX2TS U1270 ( .A(n3429), .Y(n3427) );
  CLKBUFX2TS U1271 ( .A(n3431), .Y(n3424) );
  CLKBUFX2TS U1272 ( .A(n3431), .Y(n3423) );
  CLKBUFX2TS U1273 ( .A(n3432), .Y(n3421) );
  CLKBUFX2TS U1274 ( .A(n3432), .Y(n3422) );
  CLKBUFX2TS U1275 ( .A(n3679), .Y(n3666) );
  CLKBUFX2TS U1276 ( .A(n3677), .Y(n3671) );
  CLKBUFX2TS U1277 ( .A(n3677), .Y(n3670) );
  CLKBUFX2TS U1278 ( .A(n3678), .Y(n3669) );
  CLKBUFX2TS U1279 ( .A(n3678), .Y(n3668) );
  CLKBUFX2TS U1280 ( .A(n3679), .Y(n3667) );
  CLKBUFX2TS U1281 ( .A(n3467), .Y(n3453) );
  CLKBUFX2TS U1282 ( .A(n3615), .Y(n3601) );
  CLKBUFX2TS U1283 ( .A(n3351), .Y(n3336) );
  CLKBUFX2TS U1284 ( .A(n3801), .Y(n3790) );
  CLKBUFX2TS U1285 ( .A(n798), .Y(n3801) );
  CLKBUFX2TS U1286 ( .A(n3467), .Y(n3454) );
  CLKBUFX2TS U1287 ( .A(n3351), .Y(n3337) );
  CLKBUFX2TS U1288 ( .A(n3615), .Y(n3602) );
  CLKBUFX2TS U1289 ( .A(n3350), .Y(n3339) );
  CLKBUFX2TS U1290 ( .A(n3348), .Y(n3342) );
  CLKBUFX2TS U1291 ( .A(n3348), .Y(n3344) );
  CLKBUFX2TS U1292 ( .A(n3466), .Y(n3455) );
  CLKBUFX2TS U1293 ( .A(n3466), .Y(n3456) );
  CLKBUFX2TS U1294 ( .A(n3465), .Y(n3457) );
  CLKBUFX2TS U1295 ( .A(n3465), .Y(n3458) );
  CLKBUFX2TS U1296 ( .A(n3467), .Y(n3459) );
  CLKBUFX2TS U1297 ( .A(n3464), .Y(n3460) );
  CLKBUFX2TS U1298 ( .A(n3349), .Y(n3340) );
  CLKBUFX2TS U1299 ( .A(n3348), .Y(n3345) );
  CLKBUFX2TS U1300 ( .A(n3348), .Y(n3343) );
  CLKBUFX2TS U1301 ( .A(n3349), .Y(n3341) );
  CLKBUFX2TS U1302 ( .A(n3350), .Y(n3338) );
  CLKBUFX2TS U1303 ( .A(n3788), .Y(n3775) );
  CLKBUFX2TS U1304 ( .A(n3785), .Y(n3788) );
  INVX2TS U1305 ( .A(n3660), .Y(n3659) );
  INVX2TS U1306 ( .A(n3662), .Y(n3657) );
  INVX2TS U1307 ( .A(n3661), .Y(n3658) );
  CLKBUFX2TS U1308 ( .A(n3873), .Y(n3861) );
  CLKBUFX2TS U1309 ( .A(n3830), .Y(n3823) );
  CLKBUFX2TS U1310 ( .A(n3829), .Y(n3824) );
  CLKBUFX2TS U1311 ( .A(n3830), .Y(n3822) );
  CLKBUFX2TS U1312 ( .A(n3832), .Y(n3821) );
  CLKBUFX2TS U1313 ( .A(n3317), .Y(n3301) );
  CLKBUFX2TS U1314 ( .A(n3917), .Y(n3904) );
  CLKBUFX2TS U1315 ( .A(n3916), .Y(n3906) );
  CLKBUFX2TS U1316 ( .A(n3916), .Y(n3905) );
  CLKBUFX2TS U1317 ( .A(n3915), .Y(n3907) );
  CLKBUFX2TS U1318 ( .A(n3828), .Y(n3820) );
  CLKBUFX2TS U1319 ( .A(n3831), .Y(n3819) );
  CLKBUFX2TS U1320 ( .A(n3829), .Y(n3825) );
  CLKBUFX2TS U1321 ( .A(n3317), .Y(n3302) );
  CLKBUFX2TS U1322 ( .A(n3915), .Y(n3908) );
  CLKBUFX2TS U1323 ( .A(n3828), .Y(n3826) );
  CLKBUFX2TS U1324 ( .A(n3313), .Y(n3308) );
  CLKBUFX2TS U1325 ( .A(n3313), .Y(n3307) );
  CLKBUFX2TS U1326 ( .A(n3315), .Y(n3306) );
  CLKBUFX2TS U1327 ( .A(n3315), .Y(n3305) );
  CLKBUFX2TS U1328 ( .A(n3316), .Y(n3304) );
  CLKBUFX2TS U1329 ( .A(n3316), .Y(n3303) );
  CLKBUFX2TS U1330 ( .A(n3312), .Y(n3309) );
  CLKBUFX2TS U1331 ( .A(n3577), .Y(n3573) );
  CLKBUFX2TS U1332 ( .A(n3577), .Y(n3572) );
  CLKBUFX2TS U1333 ( .A(n3578), .Y(n3571) );
  CLKBUFX2TS U1334 ( .A(n3579), .Y(n3569) );
  CLKBUFX2TS U1335 ( .A(n3579), .Y(n3568) );
  CLKBUFX2TS U1336 ( .A(n3578), .Y(n3570) );
  CLKBUFX2TS U1337 ( .A(n3580), .Y(n3567) );
  CLKBUFX2TS U1338 ( .A(n3580), .Y(n3566) );
  CLKBUFX2TS U1339 ( .A(n3576), .Y(n3574) );
  CLKBUFX2TS U1340 ( .A(n3913), .Y(n3911) );
  CLKBUFX2TS U1341 ( .A(n3914), .Y(n3909) );
  CLKBUFX2TS U1342 ( .A(n3728), .Y(n3714) );
  CLKBUFX2TS U1343 ( .A(n3913), .Y(n3910) );
  CLKBUFX2TS U1344 ( .A(n3725), .Y(n3722) );
  CLKBUFX2TS U1345 ( .A(n3728), .Y(n3721) );
  CLKBUFX2TS U1346 ( .A(n3727), .Y(n3720) );
  CLKBUFX2TS U1347 ( .A(n3726), .Y(n3719) );
  CLKBUFX2TS U1348 ( .A(n3726), .Y(n3718) );
  CLKBUFX2TS U1349 ( .A(n3727), .Y(n3717) );
  CLKBUFX2TS U1350 ( .A(n3727), .Y(n3716) );
  CLKBUFX2TS U1351 ( .A(n3728), .Y(n3715) );
  CLKBUFX2TS U1352 ( .A(n3263), .Y(n3262) );
  CLKBUFX2TS U1353 ( .A(n3250), .Y(n3171) );
  CLKBUFX2TS U1354 ( .A(n3250), .Y(n3172) );
  CLKBUFX2TS U1355 ( .A(n3249), .Y(n3173) );
  CLKBUFX2TS U1356 ( .A(n3548), .Y(n3536) );
  CLKBUFX2TS U1357 ( .A(n3548), .Y(n3535) );
  CLKBUFX2TS U1358 ( .A(n3252), .Y(n3242) );
  CLKBUFX2TS U1359 ( .A(n3248), .Y(n3241) );
  CLKBUFX2TS U1360 ( .A(n3247), .Y(n3244) );
  CLKBUFX2TS U1361 ( .A(n3247), .Y(n3243) );
  CLKBUFX2TS U1362 ( .A(n3248), .Y(n3175) );
  CLKBUFX2TS U1363 ( .A(n3249), .Y(n3174) );
  CLKBUFX2TS U1364 ( .A(n3464), .Y(n3461) );
  CLKBUFX2TS U1365 ( .A(n3283), .Y(n3270) );
  CLKBUFX2TS U1366 ( .A(n3283), .Y(n3271) );
  CLKBUFX2TS U1367 ( .A(n3697), .Y(n3683) );
  CLKBUFX2TS U1368 ( .A(n3697), .Y(n3684) );
  CLKBUFX2TS U1369 ( .A(n3247), .Y(n3245) );
  CLKBUFX2TS U1370 ( .A(n3282), .Y(n3272) );
  CLKBUFX2TS U1371 ( .A(n3282), .Y(n3273) );
  CLKBUFX2TS U1372 ( .A(n3696), .Y(n3685) );
  CLKBUFX2TS U1373 ( .A(n3887), .Y(n3876) );
  CLKBUFX2TS U1374 ( .A(n3888), .Y(n3887) );
  CLKBUFX2TS U1375 ( .A(n3576), .Y(n3575) );
  CLKBUFX2TS U1376 ( .A(n3545), .Y(n3543) );
  CLKBUFX2TS U1377 ( .A(n3551), .Y(n3541) );
  CLKBUFX2TS U1378 ( .A(n3551), .Y(n3542) );
  CLKBUFX2TS U1379 ( .A(n3546), .Y(n3540) );
  CLKBUFX2TS U1380 ( .A(n3546), .Y(n3539) );
  CLKBUFX2TS U1381 ( .A(n3312), .Y(n3310) );
  CLKBUFX2TS U1382 ( .A(n3280), .Y(n3278) );
  CLKBUFX2TS U1383 ( .A(n3286), .Y(n3276) );
  CLKBUFX2TS U1384 ( .A(n3286), .Y(n3277) );
  CLKBUFX2TS U1385 ( .A(n3281), .Y(n3275) );
  CLKBUFX2TS U1386 ( .A(n3281), .Y(n3274) );
  CLKBUFX2TS U1387 ( .A(n3871), .Y(n3865) );
  CLKBUFX2TS U1388 ( .A(n3873), .Y(n3862) );
  CLKBUFX2TS U1389 ( .A(n3870), .Y(n3868) );
  CLKBUFX2TS U1390 ( .A(n3870), .Y(n3867) );
  CLKBUFX2TS U1391 ( .A(n3871), .Y(n3866) );
  CLKBUFX2TS U1392 ( .A(n3872), .Y(n3864) );
  CLKBUFX2TS U1393 ( .A(n3872), .Y(n3863) );
  CLKBUFX2TS U1394 ( .A(n3611), .Y(n3606) );
  CLKBUFX2TS U1395 ( .A(n3611), .Y(n3605) );
  CLKBUFX2TS U1396 ( .A(n3612), .Y(n3604) );
  CLKBUFX2TS U1397 ( .A(n3699), .Y(n3692) );
  CLKBUFX2TS U1398 ( .A(n3699), .Y(n3691) );
  CLKBUFX2TS U1399 ( .A(n3694), .Y(n3690) );
  CLKBUFX2TS U1400 ( .A(n3694), .Y(n3689) );
  CLKBUFX2TS U1401 ( .A(n3695), .Y(n3688) );
  CLKBUFX2TS U1402 ( .A(n3695), .Y(n3687) );
  CLKBUFX2TS U1403 ( .A(n3696), .Y(n3686) );
  CLKBUFX2TS U1404 ( .A(n3610), .Y(n3608) );
  CLKBUFX2TS U1405 ( .A(n3610), .Y(n3607) );
  CLKBUFX2TS U1406 ( .A(n3612), .Y(n3603) );
  CLKBUFX2TS U1407 ( .A(n3725), .Y(n3723) );
  CLKBUFX2TS U1408 ( .A(n3815), .Y(n3804) );
  CLKBUFX2TS U1409 ( .A(n3816), .Y(n3815) );
  CLKBUFX2TS U1410 ( .A(n3930), .Y(n3918) );
  CLKBUFX2TS U1411 ( .A(n784), .Y(n3930) );
  CLKBUFX2TS U1412 ( .A(n3828), .Y(n3827) );
  CLKBUFX2TS U1413 ( .A(n3914), .Y(n3912) );
  INVX2TS U1414 ( .A(n3136), .Y(n3122) );
  INVX2TS U1415 ( .A(n3450), .Y(n3437) );
  INVX2TS U1416 ( .A(n3450), .Y(n3438) );
  INVX2TS U1417 ( .A(n3450), .Y(n3436) );
  INVX2TS U1418 ( .A(n3451), .Y(n3439) );
  INVX2TS U1419 ( .A(n3451), .Y(n3440) );
  INVX2TS U1420 ( .A(n3450), .Y(n3441) );
  INVX2TS U1421 ( .A(n3451), .Y(n3442) );
  INVX2TS U1422 ( .A(n3451), .Y(n3443) );
  INVX2TS U1423 ( .A(n3135), .Y(n3124) );
  INVX2TS U1424 ( .A(n3135), .Y(n3125) );
  INVX2TS U1425 ( .A(n3134), .Y(n3128) );
  INVX2TS U1426 ( .A(n3134), .Y(n3129) );
  INVX2TS U1427 ( .A(n3133), .Y(n3130) );
  INVX2TS U1428 ( .A(n3135), .Y(n3126) );
  INVX2TS U1429 ( .A(n3134), .Y(n3127) );
  INVX2TS U1430 ( .A(n3133), .Y(n3131) );
  INVX2TS U1431 ( .A(n3597), .Y(n3592) );
  INVX2TS U1432 ( .A(n3598), .Y(n3591) );
  INVX2TS U1433 ( .A(n3598), .Y(n3590) );
  INVX2TS U1434 ( .A(n3597), .Y(n3584) );
  INVX2TS U1435 ( .A(n3596), .Y(n3589) );
  INVX2TS U1436 ( .A(n3596), .Y(n3588) );
  INVX2TS U1437 ( .A(n3596), .Y(n3587) );
  INVX2TS U1438 ( .A(n3597), .Y(n3586) );
  INVX2TS U1439 ( .A(n3597), .Y(n3585) );
  INVX2TS U1440 ( .A(n3136), .Y(n3123) );
  INVX2TS U1441 ( .A(n3133), .Y(n3132) );
  INVX2TS U1442 ( .A(n3596), .Y(n3583) );
  CLKBUFX2TS U1443 ( .A(reset), .Y(n4571) );
  CLKBUFX2TS U1444 ( .A(n3859), .Y(n3858) );
  CLKBUFX2TS U1445 ( .A(n3860), .Y(n3857) );
  CLKBUFX2TS U1446 ( .A(n3860), .Y(n3855) );
  CLKBUFX2TS U1447 ( .A(n3860), .Y(n3856) );
  CLKBUFX2TS U1448 ( .A(n3481), .Y(n3471) );
  CLKBUFX2TS U1449 ( .A(n3629), .Y(n3618) );
  CLKBUFX2TS U1450 ( .A(n3481), .Y(n3472) );
  CLKBUFX2TS U1451 ( .A(n3478), .Y(n3477) );
  CLKBUFX2TS U1452 ( .A(n3479), .Y(n3476) );
  CLKBUFX2TS U1453 ( .A(n3479), .Y(n3475) );
  CLKBUFX2TS U1454 ( .A(n3480), .Y(n3474) );
  CLKBUFX2TS U1455 ( .A(n3480), .Y(n3473) );
  CLKBUFX2TS U1456 ( .A(n3563), .Y(n3552) );
  CLKBUFX2TS U1457 ( .A(n3561), .Y(n3553) );
  CLKBUFX2TS U1458 ( .A(n3561), .Y(n3554) );
  CLKBUFX2TS U1459 ( .A(n3560), .Y(n3555) );
  CLKBUFX2TS U1460 ( .A(n3709), .Y(n3708) );
  CLKBUFX2TS U1461 ( .A(n3627), .Y(n3619) );
  CLKBUFX2TS U1462 ( .A(n3626), .Y(n3621) );
  CLKBUFX2TS U1463 ( .A(n3626), .Y(n3622) );
  CLKBUFX2TS U1464 ( .A(n3625), .Y(n3624) );
  CLKBUFX2TS U1465 ( .A(n3712), .Y(n3700) );
  CLKBUFX2TS U1466 ( .A(n3712), .Y(n3701) );
  CLKBUFX2TS U1467 ( .A(n3711), .Y(n3702) );
  CLKBUFX2TS U1468 ( .A(n3713), .Y(n3703) );
  CLKBUFX2TS U1469 ( .A(n3711), .Y(n3704) );
  CLKBUFX2TS U1470 ( .A(n3710), .Y(n3705) );
  CLKBUFX2TS U1471 ( .A(n3710), .Y(n3706) );
  CLKBUFX2TS U1472 ( .A(n3709), .Y(n3707) );
  CLKBUFX2TS U1473 ( .A(n3627), .Y(n3620) );
  CLKBUFX2TS U1474 ( .A(n3625), .Y(n3623) );
  CLKBUFX2TS U1475 ( .A(n3560), .Y(n3556) );
  CLKBUFX2TS U1476 ( .A(n3559), .Y(n3557) );
  CLKBUFX2TS U1477 ( .A(n3559), .Y(n3558) );
  CLKBUFX2TS U1478 ( .A(n1070), .Y(n1059) );
  CLKBUFX2TS U1479 ( .A(n1068), .Y(n1060) );
  CLKBUFX2TS U1480 ( .A(n1068), .Y(n1061) );
  CLKBUFX2TS U1481 ( .A(n1067), .Y(n1062) );
  CLKBUFX2TS U1482 ( .A(n1066), .Y(n1065) );
  CLKBUFX2TS U1483 ( .A(n1067), .Y(n1063) );
  CLKBUFX2TS U1484 ( .A(n1066), .Y(n1064) );
  CLKBUFX2TS U1485 ( .A(n1057), .Y(n1045) );
  CLKBUFX2TS U1486 ( .A(n2167), .Y(n1046) );
  CLKBUFX2TS U1487 ( .A(n1056), .Y(n1047) );
  CLKBUFX2TS U1488 ( .A(n1056), .Y(n1048) );
  CLKBUFX2TS U1489 ( .A(n1058), .Y(n1049) );
  CLKBUFX2TS U1490 ( .A(n1055), .Y(n1050) );
  CLKBUFX2TS U1491 ( .A(n1054), .Y(n1053) );
  CLKBUFX2TS U1492 ( .A(n1055), .Y(n1051) );
  CLKBUFX2TS U1493 ( .A(n1054), .Y(n1052) );
  CLKBUFX2TS U1494 ( .A(n1084), .Y(n1073) );
  CLKBUFX2TS U1495 ( .A(n1082), .Y(n1074) );
  CLKBUFX2TS U1496 ( .A(n1082), .Y(n1075) );
  CLKBUFX2TS U1497 ( .A(n1081), .Y(n1076) );
  CLKBUFX2TS U1498 ( .A(n1080), .Y(n1079) );
  CLKBUFX2TS U1499 ( .A(n1081), .Y(n1077) );
  CLKBUFX2TS U1500 ( .A(n1080), .Y(n1078) );
  CLKBUFX2TS U1501 ( .A(n3665), .Y(n3660) );
  CLKBUFX2TS U1502 ( .A(n3665), .Y(n3661) );
  CLKBUFX2TS U1503 ( .A(n3665), .Y(n3662) );
  CLKBUFX2TS U1504 ( .A(n3517), .Y(n3514) );
  CLKBUFX2TS U1505 ( .A(n3517), .Y(n3512) );
  CLKBUFX2TS U1506 ( .A(n3517), .Y(n3513) );
  CLKBUFX2TS U1507 ( .A(n3400), .Y(n3395) );
  CLKBUFX2TS U1508 ( .A(n3400), .Y(n3396) );
  CLKBUFX2TS U1509 ( .A(n3400), .Y(n3397) );
  CLKBUFX2TS U1510 ( .A(n3832), .Y(n3830) );
  CLKBUFX2TS U1511 ( .A(n3832), .Y(n3829) );
  CLKBUFX2TS U1512 ( .A(n3832), .Y(n3828) );
  CLKBUFX2TS U1513 ( .A(n1185), .Y(n3579) );
  CLKBUFX2TS U1514 ( .A(n1185), .Y(n3580) );
  CLKBUFX2TS U1515 ( .A(n3582), .Y(n3581) );
  CLKBUFX2TS U1516 ( .A(n3875), .Y(n3869) );
  CLKBUFX2TS U1517 ( .A(n3875), .Y(n3870) );
  CLKBUFX2TS U1518 ( .A(n3915), .Y(n3914) );
  CLKBUFX2TS U1519 ( .A(n3916), .Y(n3913) );
  CLKBUFX2TS U1520 ( .A(n3729), .Y(n3727) );
  CLKBUFX2TS U1521 ( .A(n3549), .Y(n3547) );
  CLKBUFX2TS U1522 ( .A(n3550), .Y(n3545) );
  CLKBUFX2TS U1523 ( .A(n3549), .Y(n3546) );
  CLKBUFX2TS U1524 ( .A(n3549), .Y(n3548) );
  CLKBUFX2TS U1525 ( .A(n3251), .Y(n3248) );
  CLKBUFX2TS U1526 ( .A(n3251), .Y(n3249) );
  CLKBUFX2TS U1527 ( .A(n3252), .Y(n3247) );
  CLKBUFX2TS U1528 ( .A(n3681), .Y(n3674) );
  CLKBUFX2TS U1529 ( .A(n3616), .Y(n3614) );
  CLKBUFX2TS U1530 ( .A(n3468), .Y(n3466) );
  CLKBUFX2TS U1531 ( .A(n3468), .Y(n3465) );
  CLKBUFX2TS U1532 ( .A(n3468), .Y(n3467) );
  CLKBUFX2TS U1533 ( .A(n1249), .Y(n3313) );
  CLKBUFX2TS U1534 ( .A(n3269), .Y(n3264) );
  CLKBUFX2TS U1535 ( .A(n3285), .Y(n3280) );
  CLKBUFX2TS U1536 ( .A(n1249), .Y(n3315) );
  CLKBUFX2TS U1537 ( .A(n3268), .Y(n3266) );
  CLKBUFX2TS U1538 ( .A(n1249), .Y(n3314) );
  CLKBUFX2TS U1539 ( .A(n3269), .Y(n3265) );
  CLKBUFX2TS U1540 ( .A(n3313), .Y(n3316) );
  CLKBUFX2TS U1541 ( .A(n3284), .Y(n3281) );
  CLKBUFX2TS U1542 ( .A(n3312), .Y(n3317) );
  CLKBUFX2TS U1543 ( .A(n3268), .Y(n3267) );
  CLKBUFX2TS U1544 ( .A(n1204), .Y(n3464) );
  CLKBUFX2TS U1545 ( .A(n3533), .Y(n3530) );
  CLKBUFX2TS U1546 ( .A(n3534), .Y(n3529) );
  CLKBUFX2TS U1547 ( .A(n3533), .Y(n3531) );
  CLKBUFX2TS U1548 ( .A(n3533), .Y(n3532) );
  CLKBUFX2TS U1549 ( .A(n3435), .Y(n3430) );
  CLKBUFX2TS U1550 ( .A(n3434), .Y(n3433) );
  CLKBUFX2TS U1551 ( .A(n3435), .Y(n3431) );
  CLKBUFX2TS U1552 ( .A(n1235), .Y(n3348) );
  CLKBUFX2TS U1553 ( .A(n3352), .Y(n3349) );
  CLKBUFX2TS U1554 ( .A(n3352), .Y(n3350) );
  CLKBUFX2TS U1555 ( .A(n3434), .Y(n3432) );
  CLKBUFX2TS U1556 ( .A(n3284), .Y(n3282) );
  CLKBUFX2TS U1557 ( .A(n3352), .Y(n3351) );
  CLKBUFX2TS U1558 ( .A(n3616), .Y(n3615) );
  CLKBUFX2TS U1559 ( .A(n3617), .Y(n3611) );
  CLKBUFX2TS U1560 ( .A(n3681), .Y(n3675) );
  CLKBUFX2TS U1561 ( .A(n3729), .Y(n3726) );
  CLKBUFX2TS U1562 ( .A(n3681), .Y(n3676) );
  CLKBUFX2TS U1563 ( .A(n3680), .Y(n3677) );
  CLKBUFX2TS U1564 ( .A(n1153), .Y(n3694) );
  CLKBUFX2TS U1565 ( .A(n3680), .Y(n3678) );
  CLKBUFX2TS U1566 ( .A(n3729), .Y(n3728) );
  CLKBUFX2TS U1567 ( .A(n3698), .Y(n3695) );
  CLKBUFX2TS U1568 ( .A(n3698), .Y(n3696) );
  CLKBUFX2TS U1569 ( .A(n3680), .Y(n3679) );
  CLKBUFX2TS U1570 ( .A(n3617), .Y(n3610) );
  CLKBUFX2TS U1571 ( .A(n3617), .Y(n3612) );
  CLKBUFX2TS U1572 ( .A(n3284), .Y(n3283) );
  CLKBUFX2TS U1573 ( .A(n3269), .Y(n3263) );
  CLKBUFX2TS U1574 ( .A(n3698), .Y(n3697) );
  CLKBUFX2TS U1575 ( .A(n3435), .Y(n3429) );
  CLKBUFX2TS U1576 ( .A(n3251), .Y(n3250) );
  CLKBUFX2TS U1577 ( .A(n1235), .Y(n3347) );
  CLKBUFX2TS U1578 ( .A(n1202), .Y(n3500) );
  CLKBUFX2TS U1579 ( .A(n3582), .Y(n3578) );
  CLKBUFX2TS U1580 ( .A(n3582), .Y(n3577) );
  CLKBUFX2TS U1581 ( .A(n3874), .Y(n3871) );
  CLKBUFX2TS U1582 ( .A(n3874), .Y(n3872) );
  CLKBUFX2TS U1583 ( .A(n3917), .Y(n3916) );
  CLKBUFX2TS U1584 ( .A(n794), .Y(n3831) );
  CLKBUFX2TS U1585 ( .A(n3917), .Y(n3915) );
  CLKBUFX2TS U1586 ( .A(n3730), .Y(n3725) );
  CLKBUFX2TS U1587 ( .A(n1202), .Y(n3499) );
  CLKBUFX2TS U1588 ( .A(n1233), .Y(n3383) );
  CLKBUFX2TS U1589 ( .A(n797), .Y(n3803) );
  CLKBUFX2TS U1590 ( .A(n784), .Y(n3931) );
  CLKBUFX2TS U1591 ( .A(n798), .Y(n3802) );
  CLKBUFX2TS U1592 ( .A(n788), .Y(n3889) );
  CLKBUFX2TS U1593 ( .A(n788), .Y(n3888) );
  CLKBUFX2TS U1594 ( .A(n174), .Y(n3817) );
  CLKBUFX2TS U1595 ( .A(n174), .Y(n3816) );
  CLKBUFX2TS U1596 ( .A(n169), .Y(n3902) );
  CLKBUFX2TS U1597 ( .A(n169), .Y(n3903) );
  CLKBUFX2TS U1598 ( .A(n1792), .Y(n3789) );
  CLKBUFX2TS U1599 ( .A(n1267), .Y(n3156) );
  CLKBUFX2TS U1600 ( .A(n3644), .Y(n3637) );
  CLKBUFX2TS U1601 ( .A(n3645), .Y(n3635) );
  CLKBUFX2TS U1602 ( .A(n3645), .Y(n3634) );
  CLKBUFX2TS U1603 ( .A(n3646), .Y(n3632) );
  CLKBUFX2TS U1604 ( .A(n3643), .Y(n3638) );
  CLKBUFX2TS U1605 ( .A(n3644), .Y(n3636) );
  CLKBUFX2TS U1606 ( .A(n3646), .Y(n3633) );
  CLKBUFX2TS U1607 ( .A(n3416), .Y(n3402) );
  CLKBUFX2TS U1608 ( .A(n3416), .Y(n3403) );
  CLKBUFX2TS U1609 ( .A(n3411), .Y(n3410) );
  CLKBUFX2TS U1610 ( .A(n3413), .Y(n3409) );
  CLKBUFX2TS U1611 ( .A(n3413), .Y(n3408) );
  CLKBUFX2TS U1612 ( .A(n3414), .Y(n3407) );
  CLKBUFX2TS U1613 ( .A(n3414), .Y(n3406) );
  CLKBUFX2TS U1614 ( .A(n3415), .Y(n3404) );
  CLKBUFX2TS U1615 ( .A(n3415), .Y(n3405) );
  INVX2TS U1616 ( .A(n3663), .Y(n3649) );
  CLKBUFX2TS U1617 ( .A(n3664), .Y(n3663) );
  INVX2TS U1618 ( .A(n971), .Y(n3650) );
  INVX2TS U1619 ( .A(n3664), .Y(n3651) );
  INVX2TS U1620 ( .A(n3664), .Y(n3652) );
  INVX2TS U1621 ( .A(n3664), .Y(n3653) );
  INVX2TS U1622 ( .A(n3665), .Y(n3654) );
  INVX2TS U1623 ( .A(n3663), .Y(n3655) );
  INVX2TS U1624 ( .A(n971), .Y(n3656) );
  INVX2TS U1625 ( .A(n907), .Y(n801) );
  CLKBUFX2TS U1626 ( .A(n939), .Y(n3450) );
  CLKBUFX2TS U1627 ( .A(n939), .Y(n3451) );
  CLKBUFX2TS U1628 ( .A(n939), .Y(n3452) );
  CLKBUFX2TS U1629 ( .A(n3642), .Y(n3639) );
  CLKBUFX2TS U1630 ( .A(n3642), .Y(n3640) );
  CLKBUFX2TS U1631 ( .A(n3463), .Y(n3462) );
  CLKBUFX2TS U1632 ( .A(n1235), .Y(n3346) );
  CLKBUFX2TS U1633 ( .A(n3250), .Y(n3246) );
  CLKBUFX2TS U1634 ( .A(n3286), .Y(n3279) );
  CLKBUFX2TS U1635 ( .A(n3616), .Y(n3609) );
  CLKBUFX2TS U1636 ( .A(n3699), .Y(n3693) );
  CLKBUFX2TS U1637 ( .A(n3729), .Y(n3724) );
  INVX2TS U1638 ( .A(n3399), .Y(n3391) );
  INVX2TS U1639 ( .A(n3399), .Y(n3390) );
  INVX2TS U1640 ( .A(n3398), .Y(n3388) );
  INVX2TS U1641 ( .A(n3398), .Y(n3386) );
  INVX2TS U1642 ( .A(n3399), .Y(n3384) );
  INVX2TS U1643 ( .A(n3516), .Y(n3508) );
  INVX2TS U1644 ( .A(n3516), .Y(n3507) );
  INVX2TS U1645 ( .A(n3515), .Y(n3506) );
  INVX2TS U1646 ( .A(n3516), .Y(n3505) );
  INVX2TS U1647 ( .A(n3515), .Y(n3504) );
  INVX2TS U1648 ( .A(n3516), .Y(n3503) );
  INVX2TS U1649 ( .A(n3515), .Y(n3502) );
  INVX2TS U1650 ( .A(n3515), .Y(n3501) );
  INVX2TS U1651 ( .A(n3398), .Y(n3385) );
  INVX2TS U1652 ( .A(n3398), .Y(n3387) );
  INVX2TS U1653 ( .A(n3399), .Y(n3389) );
  CLKBUFX2TS U1654 ( .A(n3139), .Y(n3137) );
  CLKBUFX2TS U1655 ( .A(n3740), .Y(n3736) );
  CLKBUFX2TS U1656 ( .A(n3740), .Y(n3735) );
  CLKBUFX2TS U1657 ( .A(n3741), .Y(n3734) );
  CLKBUFX2TS U1658 ( .A(n3741), .Y(n3733) );
  CLKBUFX2TS U1659 ( .A(n3742), .Y(n3732) );
  CLKBUFX2TS U1660 ( .A(n3742), .Y(n3731) );
  INVX2TS U1661 ( .A(n3599), .Y(n3594) );
  INVX2TS U1662 ( .A(n3598), .Y(n3593) );
  INVX2TS U1663 ( .A(n3332), .Y(n3328) );
  INVX2TS U1664 ( .A(n3332), .Y(n3327) );
  INVX2TS U1665 ( .A(n3332), .Y(n3326) );
  INVX2TS U1666 ( .A(n3335), .Y(n3320) );
  INVX2TS U1667 ( .A(n3333), .Y(n3325) );
  INVX2TS U1668 ( .A(n3333), .Y(n3324) );
  INVX2TS U1669 ( .A(n3333), .Y(n3323) );
  INVX2TS U1670 ( .A(n976), .Y(n3322) );
  INVX2TS U1671 ( .A(n976), .Y(n3321) );
  INVX2TS U1672 ( .A(n3334), .Y(n3318) );
  INVX2TS U1673 ( .A(n3334), .Y(n3319) );
  CLKBUFX2TS U1674 ( .A(n3483), .Y(n3479) );
  CLKBUFX2TS U1675 ( .A(n1203), .Y(n3478) );
  CLKBUFX2TS U1676 ( .A(n3483), .Y(n3480) );
  CLKBUFX2TS U1677 ( .A(n3630), .Y(n3629) );
  CLKBUFX2TS U1678 ( .A(n3483), .Y(n3481) );
  CLKBUFX2TS U1679 ( .A(n3564), .Y(n3563) );
  CLKBUFX2TS U1680 ( .A(n3565), .Y(n3561) );
  CLKBUFX2TS U1681 ( .A(n3565), .Y(n3560) );
  CLKBUFX2TS U1682 ( .A(n3564), .Y(n3562) );
  CLKBUFX2TS U1683 ( .A(n3565), .Y(n3559) );
  CLKBUFX2TS U1684 ( .A(n3631), .Y(n3626) );
  CLKBUFX2TS U1685 ( .A(n3713), .Y(n3712) );
  CLKBUFX2TS U1686 ( .A(n1152), .Y(n3711) );
  CLKBUFX2TS U1687 ( .A(n3713), .Y(n3710) );
  CLKBUFX2TS U1688 ( .A(n3713), .Y(n3709) );
  CLKBUFX2TS U1689 ( .A(n3630), .Y(n3628) );
  CLKBUFX2TS U1690 ( .A(n3631), .Y(n3627) );
  CLKBUFX2TS U1691 ( .A(n3631), .Y(n3625) );
  CLKBUFX2TS U1692 ( .A(n791), .Y(n3859) );
  CLKBUFX2TS U1693 ( .A(n791), .Y(n3860) );
  CLKBUFX2TS U1694 ( .A(n3167), .Y(n3159) );
  CLKBUFX2TS U1695 ( .A(n3363), .Y(n3355) );
  CLKBUFX2TS U1696 ( .A(n3167), .Y(n3158) );
  CLKBUFX2TS U1697 ( .A(n3363), .Y(n3354) );
  CLKBUFX2TS U1698 ( .A(n3362), .Y(n3356) );
  CLKBUFX2TS U1699 ( .A(n3166), .Y(n3160) );
  CLKBUFX2TS U1700 ( .A(n3166), .Y(n3161) );
  CLKBUFX2TS U1701 ( .A(n3170), .Y(n3162) );
  CLKBUFX2TS U1702 ( .A(n3165), .Y(n3163) );
  CLKBUFX2TS U1703 ( .A(n3165), .Y(n3164) );
  CLKBUFX2TS U1704 ( .A(n3360), .Y(n3359) );
  CLKBUFX2TS U1705 ( .A(n3362), .Y(n3357) );
  CLKBUFX2TS U1706 ( .A(n3360), .Y(n3358) );
  INVX2TS U1707 ( .A(n3116), .Y(n3105) );
  INVX2TS U1708 ( .A(n3116), .Y(n3106) );
  INVX2TS U1709 ( .A(n3120), .Y(n3115) );
  INVX2TS U1710 ( .A(n3120), .Y(n3114) );
  INVX2TS U1711 ( .A(n3116), .Y(n3113) );
  INVX2TS U1712 ( .A(n3121), .Y(n3112) );
  INVX2TS U1713 ( .A(n3120), .Y(n3111) );
  INVX2TS U1714 ( .A(n3119), .Y(n3109) );
  INVX2TS U1715 ( .A(n3119), .Y(n3108) );
  INVX2TS U1716 ( .A(n3120), .Y(n3110) );
  INVX2TS U1717 ( .A(n3116), .Y(n3107) );
  CLKBUFX2TS U1718 ( .A(n3482), .Y(n3470) );
  CLKBUFX2TS U1719 ( .A(n3483), .Y(n3482) );
  CLKBUFX2TS U1720 ( .A(n2158), .Y(n1919) );
  CLKBUFX2TS U1721 ( .A(n2965), .Y(n1155) );
  CLKBUFX2TS U1722 ( .A(n2965), .Y(n1199) );
  CLKBUFX2TS U1723 ( .A(n2964), .Y(n1215) );
  CLKBUFX2TS U1724 ( .A(n2964), .Y(n1246) );
  CLKBUFX2TS U1725 ( .A(n2158), .Y(n1846) );
  CLKBUFX2TS U1726 ( .A(n2955), .Y(n1662) );
  CLKBUFX2TS U1727 ( .A(n2955), .Y(n1794) );
  CLKBUFX2TS U1728 ( .A(n3299), .Y(n3287) );
  CLKBUFX2TS U1729 ( .A(n3298), .Y(n3289) );
  CLKBUFX2TS U1730 ( .A(n1250), .Y(n3288) );
  CLKBUFX2TS U1731 ( .A(n3297), .Y(n3291) );
  CLKBUFX2TS U1732 ( .A(n3297), .Y(n3292) );
  CLKBUFX2TS U1733 ( .A(n3298), .Y(n3290) );
  CLKBUFX2TS U1734 ( .A(n3102), .Y(n2969) );
  CLKBUFX2TS U1735 ( .A(n3102), .Y(n2968) );
  CLKBUFX2TS U1736 ( .A(n3297), .Y(n3293) );
  CLKBUFX2TS U1737 ( .A(n3296), .Y(n3294) );
  CLKBUFX2TS U1738 ( .A(n3296), .Y(n3295) );
  CLKBUFX2TS U1739 ( .A(n1130), .Y(n1119) );
  CLKBUFX2TS U1740 ( .A(n3100), .Y(n3058) );
  CLKBUFX2TS U1741 ( .A(n3099), .Y(n2975) );
  CLKBUFX2TS U1742 ( .A(n3100), .Y(n2973) );
  CLKBUFX2TS U1743 ( .A(n3099), .Y(n2974) );
  CLKBUFX2TS U1744 ( .A(n3101), .Y(n2970) );
  CLKBUFX2TS U1745 ( .A(n3100), .Y(n2972) );
  CLKBUFX2TS U1746 ( .A(n3101), .Y(n2971) );
  CLKBUFX2TS U1747 ( .A(n1129), .Y(n1124) );
  CLKBUFX2TS U1748 ( .A(n1128), .Y(n1123) );
  CLKBUFX2TS U1749 ( .A(n1128), .Y(n1122) );
  CLKBUFX2TS U1750 ( .A(n1130), .Y(n1120) );
  CLKBUFX2TS U1751 ( .A(n1129), .Y(n1121) );
  INVX2TS U1752 ( .A(n1113), .Y(n1112) );
  INVX2TS U1753 ( .A(n1114), .Y(n1111) );
  INVX2TS U1754 ( .A(n1115), .Y(n1110) );
  CLKBUFX2TS U1755 ( .A(n1071), .Y(n1070) );
  CLKBUFX2TS U1756 ( .A(n1058), .Y(n1056) );
  CLKBUFX2TS U1757 ( .A(n1071), .Y(n1069) );
  CLKBUFX2TS U1758 ( .A(n1072), .Y(n1068) );
  CLKBUFX2TS U1759 ( .A(n1058), .Y(n1055) );
  CLKBUFX2TS U1760 ( .A(n1072), .Y(n1067) );
  CLKBUFX2TS U1761 ( .A(n1058), .Y(n1054) );
  CLKBUFX2TS U1762 ( .A(n1072), .Y(n1066) );
  CLKBUFX2TS U1763 ( .A(n1085), .Y(n1084) );
  CLKBUFX2TS U1764 ( .A(n1085), .Y(n1083) );
  CLKBUFX2TS U1765 ( .A(n1087), .Y(n1082) );
  CLKBUFX2TS U1766 ( .A(n1087), .Y(n1081) );
  CLKBUFX2TS U1767 ( .A(n1087), .Y(n1080) );
  CLKBUFX2TS U1768 ( .A(n3760), .Y(n3748) );
  CLKBUFX2TS U1769 ( .A(n3760), .Y(n3749) );
  CLKBUFX2TS U1770 ( .A(n3759), .Y(n3750) );
  CLKBUFX2TS U1771 ( .A(n3758), .Y(n3751) );
  CLKBUFX2TS U1772 ( .A(n3758), .Y(n3752) );
  CLKBUFX2TS U1773 ( .A(n3756), .Y(n3755) );
  CLKBUFX2TS U1774 ( .A(n3757), .Y(n3753) );
  CLKBUFX2TS U1775 ( .A(n3757), .Y(n3754) );
  CLKBUFX2TS U1776 ( .A(n2167), .Y(n1057) );
  CLKBUFX2TS U1777 ( .A(n1042), .Y(n1030) );
  CLKBUFX2TS U1778 ( .A(n1040), .Y(n1032) );
  CLKBUFX2TS U1779 ( .A(n1040), .Y(n1033) );
  CLKBUFX2TS U1780 ( .A(n1039), .Y(n1034) );
  CLKBUFX2TS U1781 ( .A(n1038), .Y(n1037) );
  CLKBUFX2TS U1782 ( .A(n1039), .Y(n1035) );
  CLKBUFX2TS U1783 ( .A(n1038), .Y(n1036) );
  CLKBUFX2TS U1784 ( .A(n1000), .Y(n988) );
  CLKBUFX2TS U1785 ( .A(n997), .Y(n989) );
  CLKBUFX2TS U1786 ( .A(n999), .Y(n990) );
  CLKBUFX2TS U1787 ( .A(n1011), .Y(n1003) );
  CLKBUFX2TS U1788 ( .A(n999), .Y(n991) );
  CLKBUFX2TS U1789 ( .A(n1011), .Y(n1004) );
  CLKBUFX2TS U1790 ( .A(n997), .Y(n992) );
  CLKBUFX2TS U1791 ( .A(n1010), .Y(n1005) );
  CLKBUFX2TS U1792 ( .A(n996), .Y(n995) );
  CLKBUFX2TS U1793 ( .A(n1009), .Y(n1008) );
  CLKBUFX2TS U1794 ( .A(n997), .Y(n993) );
  CLKBUFX2TS U1795 ( .A(n1010), .Y(n1006) );
  CLKBUFX2TS U1796 ( .A(n996), .Y(n994) );
  CLKBUFX2TS U1797 ( .A(n1009), .Y(n1007) );
  CLKBUFX2TS U1798 ( .A(n1099), .Y(n1088) );
  CLKBUFX2TS U1799 ( .A(n1027), .Y(n1017) );
  CLKBUFX2TS U1800 ( .A(n1097), .Y(n1089) );
  CLKBUFX2TS U1801 ( .A(n1026), .Y(n1018) );
  CLKBUFX2TS U1802 ( .A(n1097), .Y(n1090) );
  CLKBUFX2TS U1803 ( .A(n1026), .Y(n1019) );
  CLKBUFX2TS U1804 ( .A(n1096), .Y(n1091) );
  CLKBUFX2TS U1805 ( .A(n1025), .Y(n1020) );
  CLKBUFX2TS U1806 ( .A(n1095), .Y(n1094) );
  CLKBUFX2TS U1807 ( .A(n1024), .Y(n1023) );
  CLKBUFX2TS U1808 ( .A(n1096), .Y(n1092) );
  CLKBUFX2TS U1809 ( .A(n1025), .Y(n1021) );
  CLKBUFX2TS U1810 ( .A(n1095), .Y(n1093) );
  CLKBUFX2TS U1811 ( .A(n1024), .Y(n1022) );
  NOR2BX1TS U1812 ( .AN(n1847), .B(n929), .Y(n1233) );
  INVX2TS U1813 ( .A(n166), .Y(n798) );
  INVX2TS U1814 ( .A(n1810), .Y(n784) );
  INVX2TS U1815 ( .A(n1799), .Y(n788) );
  CLKBUFX2TS U1816 ( .A(n1154), .Y(n3680) );
  CLKBUFX2TS U1817 ( .A(n1151), .Y(n3729) );
  CLKBUFX2TS U1818 ( .A(n790), .Y(n3875) );
  CLKBUFX2TS U1819 ( .A(n975), .Y(n3138) );
  CLKBUFX2TS U1820 ( .A(n3648), .Y(n3642) );
  CLKBUFX2TS U1821 ( .A(n3647), .Y(n3645) );
  CLKBUFX2TS U1822 ( .A(n3648), .Y(n3643) );
  CLKBUFX2TS U1823 ( .A(n3647), .Y(n3644) );
  CLKBUFX2TS U1824 ( .A(n3647), .Y(n3646) );
  CLKBUFX2TS U1825 ( .A(n1187), .Y(n3551) );
  CLKBUFX2TS U1826 ( .A(n3682), .Y(n3673) );
  CLKBUFX2TS U1827 ( .A(n1154), .Y(n3682) );
  CLKBUFX2TS U1828 ( .A(n3418), .Y(n3411) );
  CLKBUFX2TS U1829 ( .A(n3418), .Y(n3412) );
  CLKBUFX2TS U1830 ( .A(n3417), .Y(n3416) );
  CLKBUFX2TS U1831 ( .A(n3418), .Y(n3413) );
  CLKBUFX2TS U1832 ( .A(n1251), .Y(n3286) );
  CLKBUFX2TS U1833 ( .A(n3417), .Y(n3414) );
  CLKBUFX2TS U1834 ( .A(n3417), .Y(n3415) );
  CLKBUFX2TS U1835 ( .A(n1153), .Y(n3699) );
  CLKBUFX2TS U1836 ( .A(n3469), .Y(n3463) );
  CLKBUFX2TS U1837 ( .A(n1204), .Y(n3469) );
  INVX2TS U1838 ( .A(n1814), .Y(n924) );
  CLKBUFX2TS U1839 ( .A(n1188), .Y(n3534) );
  CLKBUFX2TS U1840 ( .A(n1188), .Y(n3533) );
  CLKBUFX2TS U1841 ( .A(n1171), .Y(n3616) );
  CLKBUFX2TS U1842 ( .A(n1171), .Y(n3617) );
  CLKBUFX2TS U1843 ( .A(n1153), .Y(n3698) );
  CLKBUFX2TS U1844 ( .A(n1204), .Y(n3468) );
  CLKBUFX2TS U1845 ( .A(n1265), .Y(n3252) );
  CLKBUFX2TS U1846 ( .A(n1265), .Y(n3251) );
  CLKBUFX2TS U1847 ( .A(n1251), .Y(n3285) );
  CLKBUFX2TS U1848 ( .A(n1251), .Y(n3284) );
  CLKBUFX2TS U1849 ( .A(n1235), .Y(n3352) );
  CLKBUFX2TS U1850 ( .A(n1187), .Y(n3550) );
  CLKBUFX2TS U1851 ( .A(n1187), .Y(n3549) );
  CLKBUFX2TS U1852 ( .A(n1252), .Y(n3268) );
  CLKBUFX2TS U1853 ( .A(n1218), .Y(n3434) );
  CLKBUFX2TS U1854 ( .A(n1252), .Y(n3269) );
  CLKBUFX2TS U1855 ( .A(n1218), .Y(n3435) );
  CLKBUFX2TS U1856 ( .A(n1185), .Y(n3582) );
  INVX2TS U1857 ( .A(n1917), .Y(n923) );
  CLKBUFX2TS U1858 ( .A(n785), .Y(n3917) );
  CLKBUFX2TS U1859 ( .A(n790), .Y(n3874) );
  CLKBUFX2TS U1860 ( .A(n971), .Y(n3664) );
  CLKBUFX2TS U1861 ( .A(n941), .Y(n3516) );
  CLKBUFX2TS U1862 ( .A(n941), .Y(n3515) );
  CLKBUFX2TS U1863 ( .A(n3401), .Y(n3398) );
  CLKBUFX2TS U1864 ( .A(n3401), .Y(n3399) );
  INVX2TS U1865 ( .A(n1813), .Y(n928) );
  CLKBUFX2TS U1866 ( .A(n971), .Y(n3665) );
  CLKBUFX2TS U1867 ( .A(n941), .Y(n3517) );
  CLKBUFX2TS U1868 ( .A(n3401), .Y(n3400) );
  CLKBUFX2TS U1869 ( .A(n3642), .Y(n3641) );
  CLKBUFX2TS U1870 ( .A(n3335), .Y(n3334) );
  CLKBUFX2TS U1871 ( .A(n3600), .Y(n3599) );
  CLKBUFX2TS U1872 ( .A(n3600), .Y(n3598) );
  CLKBUFX2TS U1873 ( .A(n975), .Y(n3139) );
  CLKBUFX2TS U1874 ( .A(n3746), .Y(n3740) );
  CLKBUFX2TS U1875 ( .A(n3746), .Y(n3741) );
  CLKBUFX2TS U1876 ( .A(n3746), .Y(n3742) );
  CLKBUFX2TS U1877 ( .A(n3745), .Y(n3743) );
  INVX2TS U1878 ( .A(n1854), .Y(n929) );
  CLKBUFX2TS U1879 ( .A(n3739), .Y(n3737) );
  CLKBUFX2TS U1880 ( .A(n3739), .Y(n3738) );
  INVX2TS U1881 ( .A(n3333), .Y(n3330) );
  INVX2TS U1882 ( .A(n3334), .Y(n3329) );
  CLKBUFX2TS U1883 ( .A(n1117), .Y(n1113) );
  CLKBUFX2TS U1884 ( .A(n1117), .Y(n1114) );
  CLKBUFX2TS U1885 ( .A(n1117), .Y(n1115) );
  CLKBUFX2TS U1886 ( .A(n3300), .Y(n3297) );
  CLKBUFX2TS U1887 ( .A(n3300), .Y(n3298) );
  CLKBUFX2TS U1888 ( .A(n3300), .Y(n3296) );
  CLKBUFX2TS U1889 ( .A(n3103), .Y(n3102) );
  CLKBUFX2TS U1890 ( .A(n2090), .Y(n2965) );
  CLKBUFX2TS U1891 ( .A(n2090), .Y(n2964) );
  CLKBUFX2TS U1892 ( .A(n1133), .Y(n1128) );
  CLKBUFX2TS U1893 ( .A(n2966), .Y(n2956) );
  CLKBUFX2TS U1894 ( .A(n3103), .Y(n3099) );
  CLKBUFX2TS U1895 ( .A(n1133), .Y(n1130) );
  CLKBUFX2TS U1896 ( .A(n2966), .Y(n2158) );
  CLKBUFX2TS U1897 ( .A(n3103), .Y(n3100) );
  CLKBUFX2TS U1898 ( .A(n1133), .Y(n1129) );
  CLKBUFX2TS U1899 ( .A(n2966), .Y(n2955) );
  CLKBUFX2TS U1900 ( .A(n3103), .Y(n3101) );
  CLKBUFX2TS U1901 ( .A(n3366), .Y(n3361) );
  CLKBUFX2TS U1902 ( .A(n3169), .Y(n3166) );
  CLKBUFX2TS U1903 ( .A(n3170), .Y(n3165) );
  CLKBUFX2TS U1904 ( .A(n3365), .Y(n3362) );
  CLKBUFX2TS U1905 ( .A(n3366), .Y(n3360) );
  CLKBUFX2TS U1906 ( .A(n3169), .Y(n3167) );
  CLKBUFX2TS U1907 ( .A(n3365), .Y(n3363) );
  CLKBUFX2TS U1908 ( .A(n1203), .Y(n3483) );
  CLKBUFX2TS U1909 ( .A(n1186), .Y(n3564) );
  CLKBUFX2TS U1910 ( .A(n1186), .Y(n3565) );
  CLKBUFX2TS U1911 ( .A(n1152), .Y(n3713) );
  CLKBUFX2TS U1912 ( .A(n1170), .Y(n3630) );
  CLKBUFX2TS U1913 ( .A(n1170), .Y(n3631) );
  CLKBUFX2TS U1914 ( .A(n3168), .Y(n3157) );
  CLKBUFX2TS U1915 ( .A(n3169), .Y(n3168) );
  CLKBUFX2TS U1916 ( .A(n3364), .Y(n3353) );
  CLKBUFX2TS U1917 ( .A(n3365), .Y(n3364) );
  CLKBUFX2TS U1918 ( .A(n3119), .Y(n3117) );
  CLKBUFX2TS U1919 ( .A(n3119), .Y(n3118) );
  CLKBUFX2TS U1920 ( .A(n1250), .Y(n3299) );
  INVX2TS U1921 ( .A(n1816), .Y(n933) );
  CLKBUFX2TS U1922 ( .A(n2098), .Y(n1988) );
  CLKBUFX2TS U1923 ( .A(n4225), .Y(n4227) );
  CLKBUFX2TS U1924 ( .A(n4228), .Y(n4230) );
  CLKBUFX2TS U1925 ( .A(n3060), .Y(n3059) );
  CLKBUFX2TS U1926 ( .A(n1131), .Y(n1118) );
  CLKBUFX2TS U1927 ( .A(n1133), .Y(n1131) );
  CLKBUFX2TS U1928 ( .A(n1127), .Y(n1126) );
  CLKBUFX2TS U1929 ( .A(n1127), .Y(n1125) );
  INVX2TS U1930 ( .A(n1115), .Y(n1102) );
  INVX2TS U1931 ( .A(n977), .Y(n1103) );
  INVX2TS U1932 ( .A(n1117), .Y(n1104) );
  INVX2TS U1933 ( .A(n1116), .Y(n1105) );
  INVX2TS U1934 ( .A(n1116), .Y(n1106) );
  INVX2TS U1935 ( .A(n977), .Y(n1107) );
  INVX2TS U1936 ( .A(n1116), .Y(n1108) );
  INVX2TS U1937 ( .A(n1116), .Y(n1109) );
  CLKBUFX2TS U1938 ( .A(n3761), .Y(n3760) );
  CLKBUFX2TS U1939 ( .A(n1146), .Y(n3759) );
  CLKBUFX2TS U1940 ( .A(n3761), .Y(n3758) );
  CLKBUFX2TS U1941 ( .A(n3761), .Y(n3756) );
  CLKBUFX2TS U1942 ( .A(n3761), .Y(n3757) );
  CLKBUFX2TS U1943 ( .A(n1100), .Y(n1099) );
  CLKBUFX2TS U1944 ( .A(n1014), .Y(n1012) );
  CLKBUFX2TS U1945 ( .A(n1043), .Y(n1042) );
  CLKBUFX2TS U1946 ( .A(n1100), .Y(n1098) );
  CLKBUFX2TS U1947 ( .A(n2169), .Y(n1027) );
  CLKBUFX2TS U1948 ( .A(n1043), .Y(n1041) );
  CLKBUFX2TS U1949 ( .A(n1001), .Y(n999) );
  CLKBUFX2TS U1950 ( .A(n1101), .Y(n1097) );
  CLKBUFX2TS U1951 ( .A(n1015), .Y(n1011) );
  CLKBUFX2TS U1952 ( .A(n1029), .Y(n1026) );
  CLKBUFX2TS U1953 ( .A(n1044), .Y(n1040) );
  CLKBUFX2TS U1954 ( .A(n1001), .Y(n997) );
  CLKBUFX2TS U1955 ( .A(n1101), .Y(n1096) );
  CLKBUFX2TS U1956 ( .A(n1015), .Y(n1010) );
  CLKBUFX2TS U1957 ( .A(n1029), .Y(n1025) );
  CLKBUFX2TS U1958 ( .A(n1044), .Y(n1039) );
  CLKBUFX2TS U1959 ( .A(n1001), .Y(n996) );
  CLKBUFX2TS U1960 ( .A(n1101), .Y(n1095) );
  CLKBUFX2TS U1961 ( .A(n1015), .Y(n1009) );
  CLKBUFX2TS U1962 ( .A(n1029), .Y(n1024) );
  CLKBUFX2TS U1963 ( .A(n1044), .Y(n1038) );
  CLKBUFX2TS U1964 ( .A(n2164), .Y(n1085) );
  CLKBUFX2TS U1965 ( .A(n2164), .Y(n1087) );
  CLKBUFX2TS U1966 ( .A(n2166), .Y(n1071) );
  CLKBUFX2TS U1967 ( .A(n2167), .Y(n1058) );
  CLKBUFX2TS U1968 ( .A(n2166), .Y(n1072) );
  CLKBUFX2TS U1969 ( .A(n4228), .Y(n4229) );
  CLKBUFX2TS U1970 ( .A(n4225), .Y(n4226) );
  CLKBUFX2TS U1971 ( .A(n1000), .Y(n987) );
  CLKBUFX2TS U1972 ( .A(n2172), .Y(n1000) );
  CLKBUFX2TS U1973 ( .A(n1013), .Y(n1002) );
  CLKBUFX2TS U1974 ( .A(n1014), .Y(n1013) );
  CLKBUFX2TS U1975 ( .A(n1028), .Y(n1016) );
  CLKBUFX2TS U1976 ( .A(n2169), .Y(n1028) );
  INVX2TS U1977 ( .A(n4202), .Y(n4200) );
  NOR2X1TS U1978 ( .A(n1816), .B(n1817), .Y(n1151) );
  NOR3BX1TS U1979 ( .AN(n1831), .B(n114), .C(n1836), .Y(n1204) );
  AOI21X1TS U1980 ( .A0(n936), .A1(n119), .B0(n976), .Y(n1855) );
  XNOR2X1TS U1981 ( .A(n2940), .B(n2935), .Y(n1138) );
  XOR2X1TS U1982 ( .A(n469), .B(n2934), .Y(n2940) );
  OAI211X1TS U1983 ( .A0(n109), .A1(n118), .B0(n126), .C0(n1989), .Y(n1837) );
  NAND3X1TS U1984 ( .A(n115), .B(n486), .C(n1895), .Y(n1814) );
  OAI21X1TS U1985 ( .A0(n125), .A1(n2012), .B0(n1989), .Y(n1851) );
  NOR2X1TS U1986 ( .A(n109), .B(n117), .Y(n2012) );
  OR4X2TS U1987 ( .A(n482), .B(n928), .C(n924), .D(n933), .Y(n971) );
  NOR2X1TS U1988 ( .A(n118), .B(n1989), .Y(n1842) );
  NOR2X1TS U1989 ( .A(n2941), .B(n2932), .Y(n2934) );
  NAND3X1TS U1990 ( .A(n1895), .B(n115), .C(n926), .Y(n1917) );
  INVX2TS U1991 ( .A(n1852), .Y(n919) );
  INVX2TS U1992 ( .A(n1828), .Y(n922) );
  INVX2TS U1993 ( .A(n1803), .Y(n794) );
  INVX2TS U1994 ( .A(n1858), .Y(n918) );
  CLKBUFX2TS U1995 ( .A(n1169), .Y(n3647) );
  AO21X1TS U1996 ( .A0(n2934), .A1(n2935), .B0(n469), .Y(n2936) );
  INVX2TS U1997 ( .A(n2059), .Y(n972) );
  CLKBUFX2TS U1998 ( .A(n1219), .Y(n3417) );
  CLKBUFX2TS U1999 ( .A(n1148), .Y(n3745) );
  NAND2X1TS U2000 ( .A(n940), .B(n1879), .Y(n1977) );
  INVX2TS U2001 ( .A(n2055), .Y(n930) );
  INVX2TS U2002 ( .A(n2056), .Y(n917) );
  CLKBUFX2TS U2003 ( .A(n1148), .Y(n3746) );
  NAND2X1TS U2004 ( .A(n2055), .B(n118), .Y(n1963) );
  CLKBUFX2TS U2005 ( .A(n976), .Y(n3335) );
  CLKBUFX2TS U2006 ( .A(n3747), .Y(n3739) );
  CLKBUFX2TS U2007 ( .A(n1148), .Y(n3747) );
  NOR2BX1TS U2008 ( .AN(n1908), .B(n463), .Y(n1170) );
  NOR2BX1TS U2009 ( .AN(n1908), .B(n1932), .Y(n1203) );
  CLKBUFX2TS U2010 ( .A(n3121), .Y(n3120) );
  CLKBUFX2TS U2011 ( .A(n3121), .Y(n3119) );
  CLKBUFX2TS U2012 ( .A(destinationAddressIn_SOUTH[7]), .Y(n4228) );
  CLKBUFX2TS U2013 ( .A(destinationAddressIn_SOUTH[6]), .Y(n4225) );
  INVX2TS U2014 ( .A(n1853), .Y(n920) );
  CLKBUFX2TS U2015 ( .A(n1250), .Y(n3300) );
  CLKBUFX2TS U2016 ( .A(n1266), .Y(n3170) );
  CLKBUFX2TS U2017 ( .A(n1234), .Y(n3366) );
  CLKBUFX2TS U2018 ( .A(n1266), .Y(n3169) );
  CLKBUFX2TS U2019 ( .A(n1234), .Y(n3365) );
  CLKBUFX2TS U2020 ( .A(n2103), .Y(n1133) );
  CLKBUFX2TS U2021 ( .A(n2090), .Y(n2966) );
  CLKBUFX2TS U2022 ( .A(n2089), .Y(n3103) );
  CLKBUFX2TS U2023 ( .A(n1134), .Y(n1127) );
  CLKBUFX2TS U2024 ( .A(n2103), .Y(n1134) );
  CLKBUFX2TS U2025 ( .A(n2967), .Y(n2098) );
  CLKBUFX2TS U2026 ( .A(n2090), .Y(n2967) );
  CLKBUFX2TS U2027 ( .A(n3104), .Y(n3060) );
  CLKBUFX2TS U2028 ( .A(n2089), .Y(n3104) );
  CLKBUFX2TS U2029 ( .A(n977), .Y(n1116) );
  CLKBUFX2TS U2030 ( .A(n977), .Y(n1117) );
  NOR2X1TS U2031 ( .A(n2099), .B(n130), .Y(n2164) );
  NAND2X1TS U2032 ( .A(n800), .B(n4572), .Y(n1137) );
  CLKBUFX2TS U2033 ( .A(n4203), .Y(n4202) );
  NAND2X1TS U2034 ( .A(n804), .B(n478), .Y(n2167) );
  NAND2X1TS U2035 ( .A(n464), .B(n478), .Y(n2166) );
  INVX2TS U2036 ( .A(n4196), .Y(n4194) );
  INVX2TS U2037 ( .A(n1136), .Y(n782) );
  CLKBUFX2TS U2038 ( .A(n1146), .Y(n3761) );
  CLKBUFX2TS U2039 ( .A(n2163), .Y(n1100) );
  CLKBUFX2TS U2040 ( .A(n2170), .Y(n1014) );
  CLKBUFX2TS U2041 ( .A(n2168), .Y(n1043) );
  CLKBUFX2TS U2042 ( .A(n2163), .Y(n1101) );
  CLKBUFX2TS U2043 ( .A(n2170), .Y(n1015) );
  CLKBUFX2TS U2044 ( .A(n2169), .Y(n1029) );
  CLKBUFX2TS U2045 ( .A(n2168), .Y(n1044) );
  CLKBUFX2TS U2046 ( .A(n2172), .Y(n1001) );
  CLKBUFX2TS U2047 ( .A(n4171), .Y(n4172) );
  CLKBUFX2TS U2048 ( .A(n4168), .Y(n4169) );
  CLKBUFX2TS U2049 ( .A(n4165), .Y(n4166) );
  CLKBUFX2TS U2050 ( .A(n4162), .Y(n4163) );
  CLKBUFX2TS U2051 ( .A(n4159), .Y(n4160) );
  CLKBUFX2TS U2052 ( .A(n4156), .Y(n4157) );
  CLKBUFX2TS U2053 ( .A(n4150), .Y(n4151) );
  CLKBUFX2TS U2054 ( .A(n4147), .Y(n4148) );
  CLKBUFX2TS U2055 ( .A(n4144), .Y(n4145) );
  CLKBUFX2TS U2056 ( .A(n4141), .Y(n4142) );
  CLKBUFX2TS U2057 ( .A(n4138), .Y(n4139) );
  CLKBUFX2TS U2058 ( .A(n4135), .Y(n4136) );
  CLKBUFX2TS U2059 ( .A(n4129), .Y(n4130) );
  CLKBUFX2TS U2060 ( .A(n4126), .Y(n4127) );
  CLKBUFX2TS U2061 ( .A(n4123), .Y(n4124) );
  CLKBUFX2TS U2062 ( .A(n4120), .Y(n4121) );
  CLKBUFX2TS U2063 ( .A(n4117), .Y(n4118) );
  CLKBUFX2TS U2064 ( .A(n4114), .Y(n4115) );
  CLKBUFX2TS U2065 ( .A(n4111), .Y(n4112) );
  CLKBUFX2TS U2066 ( .A(n4108), .Y(n4109) );
  CLKBUFX2TS U2067 ( .A(n4105), .Y(n4106) );
  CLKBUFX2TS U2068 ( .A(n4102), .Y(n4103) );
  CLKBUFX2TS U2069 ( .A(n4099), .Y(n4100) );
  CLKBUFX2TS U2070 ( .A(n4096), .Y(n4097) );
  CLKBUFX2TS U2071 ( .A(n4093), .Y(n4094) );
  CLKBUFX2TS U2072 ( .A(n4087), .Y(n4088) );
  CLKBUFX2TS U2073 ( .A(n4084), .Y(n4085) );
  CLKBUFX2TS U2074 ( .A(n4081), .Y(n4082) );
  CLKBUFX2TS U2075 ( .A(n4078), .Y(n4079) );
  CLKBUFX2TS U2076 ( .A(n4153), .Y(n4154) );
  CLKBUFX2TS U2077 ( .A(n4132), .Y(n4133) );
  CLKBUFX2TS U2078 ( .A(n4090), .Y(n4091) );
  INVX2TS U2079 ( .A(n3963), .Y(n3961) );
  INVX2TS U2080 ( .A(n3957), .Y(n3955) );
  INVX2TS U2081 ( .A(n3951), .Y(n3949) );
  INVX2TS U2082 ( .A(n4442), .Y(n4439) );
  INVX2TS U2083 ( .A(n4438), .Y(n4436) );
  INVX2TS U2084 ( .A(n4435), .Y(n4433) );
  INVX2TS U2085 ( .A(n4425), .Y(n4423) );
  INVX2TS U2086 ( .A(n4419), .Y(n4417) );
  INVX2TS U2087 ( .A(n4413), .Y(n4411) );
  INVX2TS U2088 ( .A(n4410), .Y(n4408) );
  INVX2TS U2089 ( .A(n4404), .Y(n4402) );
  INVX2TS U2090 ( .A(n4398), .Y(n4396) );
  INVX2TS U2091 ( .A(n4395), .Y(n4393) );
  INVX2TS U2092 ( .A(n4389), .Y(n4387) );
  INVX2TS U2093 ( .A(n4383), .Y(n4381) );
  INVX2TS U2094 ( .A(n4380), .Y(n4378) );
  INVX2TS U2095 ( .A(n4377), .Y(n4375) );
  INVX2TS U2096 ( .A(n4371), .Y(n4369) );
  INVX2TS U2097 ( .A(n4365), .Y(n4363) );
  INVX2TS U2098 ( .A(n4356), .Y(n4354) );
  INVX2TS U2099 ( .A(n3960), .Y(n3958) );
  INVX2TS U2100 ( .A(n3948), .Y(n3946) );
  INVX2TS U2101 ( .A(n3954), .Y(n3952) );
  INVX2TS U2102 ( .A(n4422), .Y(n4420) );
  INVX2TS U2103 ( .A(n4401), .Y(n4399) );
  INVX2TS U2104 ( .A(n4392), .Y(n4390) );
  INVX2TS U2105 ( .A(n4386), .Y(n4384) );
  INVX2TS U2106 ( .A(n4359), .Y(n4357) );
  INVX2TS U2107 ( .A(n4432), .Y(n4429) );
  INVX2TS U2108 ( .A(n4428), .Y(n4426) );
  INVX2TS U2109 ( .A(n4416), .Y(n4414) );
  INVX2TS U2110 ( .A(n4407), .Y(n4405) );
  INVX2TS U2111 ( .A(n4374), .Y(n4372) );
  INVX2TS U2112 ( .A(n4362), .Y(n4360) );
  INVX2TS U2113 ( .A(n4353), .Y(n4351) );
  INVX2TS U2114 ( .A(n4350), .Y(n4348) );
  INVX2TS U2115 ( .A(n4347), .Y(n4345) );
  INVX2TS U2116 ( .A(n4368), .Y(n4366) );
  INVX2TS U2117 ( .A(n4002), .Y(n4000) );
  INVX2TS U2118 ( .A(n3990), .Y(n3988) );
  INVX2TS U2119 ( .A(n4005), .Y(n4003) );
  INVX2TS U2120 ( .A(n3999), .Y(n3997) );
  INVX2TS U2121 ( .A(n3996), .Y(n3994) );
  INVX2TS U2122 ( .A(n3993), .Y(n3991) );
  INVX2TS U2123 ( .A(n4038), .Y(n4036) );
  INVX2TS U2124 ( .A(n4029), .Y(n4027) );
  INVX2TS U2125 ( .A(n4026), .Y(n4024) );
  INVX2TS U2126 ( .A(n4041), .Y(n4039) );
  INVX2TS U2127 ( .A(n4035), .Y(n4033) );
  INVX2TS U2128 ( .A(n4032), .Y(n4030) );
  CLKBUFX2TS U2129 ( .A(n4054), .Y(n4055) );
  CLKBUFX2TS U2130 ( .A(n4042), .Y(n4043) );
  CLKBUFX2TS U2131 ( .A(n4057), .Y(n4058) );
  CLKBUFX2TS U2132 ( .A(n4051), .Y(n4052) );
  CLKBUFX2TS U2133 ( .A(n4048), .Y(n4049) );
  CLKBUFX2TS U2134 ( .A(n4045), .Y(n4046) );
  INVX2TS U2135 ( .A(n4191), .Y(n4189) );
  INVX2TS U2136 ( .A(n4185), .Y(n4183) );
  INVX2TS U2137 ( .A(n4188), .Y(n4186) );
  INVX2TS U2138 ( .A(n4182), .Y(n4180) );
  INVX2TS U2139 ( .A(n4179), .Y(n4177) );
  INVX2TS U2140 ( .A(n4176), .Y(n4174) );
  CLKBUFX2TS U2141 ( .A(n4075), .Y(n4076) );
  CLKBUFX2TS U2142 ( .A(n4072), .Y(n4073) );
  CLKBUFX2TS U2143 ( .A(n4066), .Y(n4067) );
  CLKBUFX2TS U2144 ( .A(n4069), .Y(n4070) );
  CLKBUFX2TS U2145 ( .A(n4063), .Y(n4064) );
  CLKBUFX2TS U2146 ( .A(n4060), .Y(n4061) );
  INVX2TS U2147 ( .A(n4344), .Y(n4342) );
  INVX2TS U2148 ( .A(n4341), .Y(n4339) );
  INVX2TS U2149 ( .A(n4338), .Y(n4336) );
  INVX2TS U2150 ( .A(n4335), .Y(n4333) );
  INVX2TS U2151 ( .A(n4332), .Y(n4330) );
  INVX2TS U2152 ( .A(n4329), .Y(n4327) );
  INVX2TS U2153 ( .A(n4326), .Y(n4324) );
  INVX2TS U2154 ( .A(n4323), .Y(n4321) );
  INVX2TS U2155 ( .A(n4320), .Y(n4318) );
  INVX2TS U2156 ( .A(n4317), .Y(n4315) );
  INVX2TS U2157 ( .A(n4314), .Y(n4312) );
  INVX2TS U2158 ( .A(n4311), .Y(n4309) );
  INVX2TS U2159 ( .A(n4308), .Y(n4306) );
  INVX2TS U2160 ( .A(n4305), .Y(n4303) );
  INVX2TS U2161 ( .A(n4302), .Y(n4300) );
  INVX2TS U2162 ( .A(n4299), .Y(n4297) );
  INVX2TS U2163 ( .A(n4296), .Y(n4294) );
  INVX2TS U2164 ( .A(n4293), .Y(n4291) );
  INVX2TS U2165 ( .A(n4290), .Y(n4288) );
  INVX2TS U2166 ( .A(n4287), .Y(n4285) );
  INVX2TS U2167 ( .A(n4284), .Y(n4282) );
  INVX2TS U2168 ( .A(n4281), .Y(n4279) );
  INVX2TS U2169 ( .A(n4278), .Y(n4276) );
  INVX2TS U2170 ( .A(n4275), .Y(n4273) );
  INVX2TS U2171 ( .A(n4272), .Y(n4270) );
  INVX2TS U2172 ( .A(n4269), .Y(n4267) );
  INVX2TS U2173 ( .A(n4266), .Y(n4264) );
  INVX2TS U2174 ( .A(n4263), .Y(n4261) );
  INVX2TS U2175 ( .A(n4260), .Y(n4258) );
  INVX2TS U2176 ( .A(n4257), .Y(n4255) );
  INVX2TS U2177 ( .A(n4254), .Y(n4252) );
  INVX2TS U2178 ( .A(n4251), .Y(n4249) );
  INVX2TS U2179 ( .A(n4543), .Y(n4541) );
  INVX2TS U2180 ( .A(n4523), .Y(n4520) );
  INVX2TS U2181 ( .A(n4516), .Y(n4514) );
  INVX2TS U2182 ( .A(n4513), .Y(n4510) );
  INVX2TS U2183 ( .A(n4489), .Y(n4487) );
  INVX2TS U2184 ( .A(n4486), .Y(n4483) );
  INVX2TS U2185 ( .A(n4479), .Y(n4477) );
  INVX2TS U2186 ( .A(n4465), .Y(n4463) );
  INVX2TS U2187 ( .A(n4448), .Y(n4446) );
  INVX2TS U2188 ( .A(n4550), .Y(n4547) );
  INVX2TS U2189 ( .A(n4546), .Y(n4544) );
  INVX2TS U2190 ( .A(n4540), .Y(n4537) );
  INVX2TS U2191 ( .A(n4536), .Y(n4534) );
  INVX2TS U2192 ( .A(n4533), .Y(n4531) );
  INVX2TS U2193 ( .A(n4526), .Y(n4524) );
  INVX2TS U2194 ( .A(n4519), .Y(n4517) );
  INVX2TS U2195 ( .A(n4509), .Y(n4507) );
  INVX2TS U2196 ( .A(n4502), .Y(n4500) );
  INVX2TS U2197 ( .A(n4499), .Y(n4497) );
  INVX2TS U2198 ( .A(n4496), .Y(n4493) );
  INVX2TS U2199 ( .A(n4492), .Y(n4490) );
  INVX2TS U2200 ( .A(n4482), .Y(n4480) );
  INVX2TS U2201 ( .A(n4475), .Y(n4473) );
  INVX2TS U2202 ( .A(n4472), .Y(n4470) );
  INVX2TS U2203 ( .A(n4469), .Y(n4466) );
  INVX2TS U2204 ( .A(n4462), .Y(n4460) );
  INVX2TS U2205 ( .A(n4455), .Y(n4453) );
  INVX2TS U2206 ( .A(n4452), .Y(n4450) );
  INVX2TS U2207 ( .A(n4445), .Y(n4443) );
  INVX2TS U2208 ( .A(n4529), .Y(n4527) );
  INVX2TS U2209 ( .A(n4506), .Y(n4504) );
  INVX2TS U2210 ( .A(n4459), .Y(n4456) );
  CLKBUFX2TS U2211 ( .A(n4192), .Y(n4193) );
  CLKBUFX2TS U2212 ( .A(n4020), .Y(n4021) );
  CLKBUFX2TS U2213 ( .A(n4012), .Y(n4013) );
  CLKBUFX2TS U2214 ( .A(n4022), .Y(n4023) );
  CLKBUFX2TS U2215 ( .A(destinationAddressIn_WEST[10]), .Y(n4016) );
  CLKBUFX2TS U2216 ( .A(n4006), .Y(n4007) );
  CLKBUFX2TS U2217 ( .A(n4018), .Y(n4019) );
  CLKBUFX2TS U2218 ( .A(destinationAddressIn_WEST[9]), .Y(n4014) );
  CLKBUFX2TS U2219 ( .A(n4009), .Y(n4010) );
  CLKBUFX2TS U2220 ( .A(n4246), .Y(n4247) );
  CLKBUFX2TS U2221 ( .A(n4240), .Y(n4241) );
  CLKBUFX2TS U2222 ( .A(n4234), .Y(n4235) );
  CLKBUFX2TS U2223 ( .A(n4243), .Y(n4244) );
  CLKBUFX2TS U2224 ( .A(n4237), .Y(n4238) );
  CLKBUFX2TS U2225 ( .A(n4231), .Y(n4232) );
  CLKBUFX2TS U2226 ( .A(n4204), .Y(n4205) );
  CLKBUFX2TS U2227 ( .A(n4204), .Y(n4206) );
  CLKBUFX2TS U2228 ( .A(n4243), .Y(n4245) );
  CLKBUFX2TS U2229 ( .A(n4231), .Y(n4233) );
  CLKBUFX2TS U2230 ( .A(n4246), .Y(n4248) );
  CLKBUFX2TS U2231 ( .A(n4237), .Y(n4239) );
  CLKBUFX2TS U2232 ( .A(n4240), .Y(n4242) );
  CLKBUFX2TS U2233 ( .A(n4234), .Y(n4236) );
  CLKBUFX2TS U2234 ( .A(n4057), .Y(n4059) );
  CLKBUFX2TS U2235 ( .A(n4051), .Y(n4053) );
  CLKBUFX2TS U2236 ( .A(n4168), .Y(n4170) );
  CLKBUFX2TS U2237 ( .A(n4165), .Y(n4167) );
  CLKBUFX2TS U2238 ( .A(n4156), .Y(n4158) );
  CLKBUFX2TS U2239 ( .A(n4141), .Y(n4143) );
  CLKBUFX2TS U2240 ( .A(n4135), .Y(n4137) );
  CLKBUFX2TS U2241 ( .A(n4129), .Y(n4131) );
  CLKBUFX2TS U2242 ( .A(n4120), .Y(n4122) );
  CLKBUFX2TS U2243 ( .A(n4114), .Y(n4116) );
  CLKBUFX2TS U2244 ( .A(n4111), .Y(n4113) );
  CLKBUFX2TS U2245 ( .A(n4108), .Y(n4110) );
  CLKBUFX2TS U2246 ( .A(n4102), .Y(n4104) );
  CLKBUFX2TS U2247 ( .A(n4096), .Y(n4098) );
  CLKBUFX2TS U2248 ( .A(n4087), .Y(n4089) );
  CLKBUFX2TS U2249 ( .A(n4054), .Y(n4056) );
  CLKBUFX2TS U2250 ( .A(n4045), .Y(n4047) );
  CLKBUFX2TS U2251 ( .A(n4042), .Y(n4044) );
  CLKBUFX2TS U2252 ( .A(n4048), .Y(n4050) );
  CLKBUFX2TS U2253 ( .A(n4153), .Y(n4155) );
  CLKBUFX2TS U2254 ( .A(n4132), .Y(n4134) );
  CLKBUFX2TS U2255 ( .A(n4123), .Y(n4125) );
  CLKBUFX2TS U2256 ( .A(n4117), .Y(n4119) );
  CLKBUFX2TS U2257 ( .A(n4090), .Y(n4092) );
  CLKBUFX2TS U2258 ( .A(n4162), .Y(n4164) );
  CLKBUFX2TS U2259 ( .A(n4159), .Y(n4161) );
  CLKBUFX2TS U2260 ( .A(n4147), .Y(n4149) );
  CLKBUFX2TS U2261 ( .A(n4138), .Y(n4140) );
  CLKBUFX2TS U2262 ( .A(n4105), .Y(n4107) );
  CLKBUFX2TS U2263 ( .A(n4093), .Y(n4095) );
  CLKBUFX2TS U2264 ( .A(n4081), .Y(n4083) );
  CLKBUFX2TS U2265 ( .A(n4078), .Y(n4080) );
  CLKBUFX2TS U2266 ( .A(n4171), .Y(n4173) );
  CLKBUFX2TS U2267 ( .A(n4150), .Y(n4152) );
  CLKBUFX2TS U2268 ( .A(n4144), .Y(n4146) );
  CLKBUFX2TS U2269 ( .A(n4126), .Y(n4128) );
  CLKBUFX2TS U2270 ( .A(n4084), .Y(n4086) );
  CLKBUFX2TS U2271 ( .A(n4099), .Y(n4101) );
  CLKBUFX2TS U2272 ( .A(destinationAddressIn_WEST[9]), .Y(n4015) );
  CLKBUFX2TS U2273 ( .A(n4009), .Y(n4011) );
  CLKBUFX2TS U2274 ( .A(destinationAddressIn_WEST[10]), .Y(n4017) );
  CLKBUFX2TS U2275 ( .A(n4006), .Y(n4008) );
  CLKBUFX2TS U2276 ( .A(n4072), .Y(n4074) );
  CLKBUFX2TS U2277 ( .A(n4063), .Y(n4065) );
  CLKBUFX2TS U2278 ( .A(n4060), .Y(n4062) );
  CLKBUFX2TS U2279 ( .A(n4075), .Y(n4077) );
  CLKBUFX2TS U2280 ( .A(n4069), .Y(n4071) );
  CLKBUFX2TS U2281 ( .A(n4066), .Y(n4068) );
  INVX2TS U2282 ( .A(n4221), .Y(n4219) );
  INVX2TS U2283 ( .A(n4209), .Y(n4207) );
  INVX2TS U2284 ( .A(n4224), .Y(n4222) );
  INVX2TS U2285 ( .A(n4218), .Y(n4216) );
  INVX2TS U2286 ( .A(n4215), .Y(n4213) );
  INVX2TS U2287 ( .A(n4212), .Y(n4210) );
  INVX2TS U2288 ( .A(n4570), .Y(n4568) );
  INVX2TS U2289 ( .A(n4567), .Y(n4564) );
  INVX2TS U2290 ( .A(n4560), .Y(n4558) );
  INVX2TS U2291 ( .A(n4563), .Y(n4561) );
  INVX2TS U2292 ( .A(n4556), .Y(n4554) );
  INVX2TS U2293 ( .A(n4553), .Y(n4551) );
  INVX2TS U2294 ( .A(n4196), .Y(n4195) );
  INVX2TS U2295 ( .A(n4550), .Y(n4549) );
  INVX2TS U2296 ( .A(n4546), .Y(n4545) );
  INVX2TS U2297 ( .A(n4543), .Y(n4542) );
  INVX2TS U2298 ( .A(n4540), .Y(n4538) );
  INVX2TS U2299 ( .A(n4536), .Y(n4535) );
  INVX2TS U2300 ( .A(n4533), .Y(n4532) );
  INVX2TS U2301 ( .A(n4529), .Y(n4528) );
  INVX2TS U2302 ( .A(n4526), .Y(n4525) );
  INVX2TS U2303 ( .A(n4523), .Y(n4522) );
  INVX2TS U2304 ( .A(n4519), .Y(n4518) );
  INVX2TS U2305 ( .A(n4516), .Y(n4515) );
  INVX2TS U2306 ( .A(n4513), .Y(n4511) );
  INVX2TS U2307 ( .A(n4509), .Y(n4508) );
  INVX2TS U2308 ( .A(n4506), .Y(n4505) );
  INVX2TS U2309 ( .A(n4502), .Y(n4501) );
  INVX2TS U2310 ( .A(n4499), .Y(n4498) );
  INVX2TS U2311 ( .A(n4496), .Y(n4495) );
  INVX2TS U2312 ( .A(n4492), .Y(n4491) );
  INVX2TS U2313 ( .A(n4489), .Y(n4488) );
  INVX2TS U2314 ( .A(n4486), .Y(n4484) );
  INVX2TS U2315 ( .A(n4482), .Y(n4481) );
  INVX2TS U2316 ( .A(n4479), .Y(n4478) );
  INVX2TS U2317 ( .A(n4475), .Y(n4474) );
  INVX2TS U2318 ( .A(n4472), .Y(n4471) );
  INVX2TS U2319 ( .A(n4469), .Y(n4468) );
  INVX2TS U2320 ( .A(n4465), .Y(n4464) );
  INVX2TS U2321 ( .A(n4462), .Y(n4461) );
  INVX2TS U2322 ( .A(n4459), .Y(n4457) );
  INVX2TS U2323 ( .A(n4455), .Y(n4454) );
  INVX2TS U2324 ( .A(n4452), .Y(n4451) );
  INVX2TS U2325 ( .A(n4448), .Y(n4447) );
  INVX2TS U2326 ( .A(n4445), .Y(n4444) );
  INVX2TS U2327 ( .A(n4199), .Y(n4197) );
  INVX2TS U2328 ( .A(n3987), .Y(n3985) );
  INVX2TS U2329 ( .A(n3981), .Y(n3979) );
  INVX2TS U2330 ( .A(n3975), .Y(n3973) );
  INVX2TS U2331 ( .A(n3969), .Y(n3967) );
  INVX2TS U2332 ( .A(n3984), .Y(n3982) );
  INVX2TS U2333 ( .A(n3978), .Y(n3976) );
  INVX2TS U2334 ( .A(n3972), .Y(n3970) );
  INVX2TS U2335 ( .A(n3966), .Y(n3964) );
  INVX2TS U2336 ( .A(n4442), .Y(n4441) );
  INVX2TS U2337 ( .A(n4438), .Y(n4437) );
  INVX2TS U2338 ( .A(n4435), .Y(n4434) );
  INVX2TS U2339 ( .A(n4432), .Y(n4430) );
  INVX2TS U2340 ( .A(n4428), .Y(n4427) );
  INVX2TS U2341 ( .A(n4425), .Y(n4424) );
  INVX2TS U2342 ( .A(n4419), .Y(n4418) );
  INVX2TS U2343 ( .A(n4416), .Y(n4415) );
  INVX2TS U2344 ( .A(n4413), .Y(n4412) );
  INVX2TS U2345 ( .A(n4410), .Y(n4409) );
  INVX2TS U2346 ( .A(n4407), .Y(n4406) );
  INVX2TS U2347 ( .A(n4404), .Y(n4403) );
  INVX2TS U2348 ( .A(n4398), .Y(n4397) );
  INVX2TS U2349 ( .A(n4395), .Y(n4394) );
  INVX2TS U2350 ( .A(n4392), .Y(n4391) );
  INVX2TS U2351 ( .A(n4389), .Y(n4388) );
  INVX2TS U2352 ( .A(n4386), .Y(n4385) );
  INVX2TS U2353 ( .A(n4383), .Y(n4382) );
  INVX2TS U2354 ( .A(n4380), .Y(n4379) );
  INVX2TS U2355 ( .A(n4377), .Y(n4376) );
  INVX2TS U2356 ( .A(n4374), .Y(n4373) );
  INVX2TS U2357 ( .A(n4371), .Y(n4370) );
  INVX2TS U2358 ( .A(n4368), .Y(n4367) );
  INVX2TS U2359 ( .A(n4365), .Y(n4364) );
  INVX2TS U2360 ( .A(n4362), .Y(n4361) );
  INVX2TS U2361 ( .A(n4356), .Y(n4355) );
  INVX2TS U2362 ( .A(n4353), .Y(n4352) );
  INVX2TS U2363 ( .A(n4350), .Y(n4349) );
  INVX2TS U2364 ( .A(n4347), .Y(n4346) );
  INVX2TS U2365 ( .A(n4422), .Y(n4421) );
  INVX2TS U2366 ( .A(n4401), .Y(n4400) );
  INVX2TS U2367 ( .A(n4359), .Y(n4358) );
  INVX2TS U2368 ( .A(n4567), .Y(n4565) );
  INVX2TS U2369 ( .A(n4556), .Y(n4555) );
  INVX2TS U2370 ( .A(n4553), .Y(n4552) );
  INVX2TS U2371 ( .A(n4570), .Y(n4569) );
  INVX2TS U2372 ( .A(n4563), .Y(n4562) );
  INVX2TS U2373 ( .A(n4560), .Y(n4559) );
  INVX2TS U2374 ( .A(n4221), .Y(n4220) );
  INVX2TS U2375 ( .A(n4218), .Y(n4217) );
  INVX2TS U2376 ( .A(n4215), .Y(n4214) );
  INVX2TS U2377 ( .A(n4212), .Y(n4211) );
  INVX2TS U2378 ( .A(n4209), .Y(n4208) );
  INVX2TS U2379 ( .A(n4224), .Y(n4223) );
  INVX2TS U2380 ( .A(n4199), .Y(n4198) );
  INVX2TS U2381 ( .A(n3981), .Y(n3980) );
  INVX2TS U2382 ( .A(n3966), .Y(n3965) );
  INVX2TS U2383 ( .A(n3984), .Y(n3983) );
  INVX2TS U2384 ( .A(n3975), .Y(n3974) );
  INVX2TS U2385 ( .A(n3972), .Y(n3971) );
  INVX2TS U2386 ( .A(n3987), .Y(n3986) );
  INVX2TS U2387 ( .A(n3978), .Y(n3977) );
  INVX2TS U2388 ( .A(n3969), .Y(n3968) );
  INVX2TS U2389 ( .A(n4041), .Y(n4040) );
  INVX2TS U2390 ( .A(n4035), .Y(n4034) );
  INVX2TS U2391 ( .A(n4038), .Y(n4037) );
  INVX2TS U2392 ( .A(n4032), .Y(n4031) );
  INVX2TS U2393 ( .A(n4029), .Y(n4028) );
  INVX2TS U2394 ( .A(n4026), .Y(n4025) );
  INVX2TS U2395 ( .A(n4005), .Y(n4004) );
  INVX2TS U2396 ( .A(n3999), .Y(n3998) );
  INVX2TS U2397 ( .A(n3996), .Y(n3995) );
  INVX2TS U2398 ( .A(n3993), .Y(n3992) );
  INVX2TS U2399 ( .A(n4002), .Y(n4001) );
  INVX2TS U2400 ( .A(n3990), .Y(n3989) );
  INVX2TS U2401 ( .A(n4338), .Y(n4337) );
  INVX2TS U2402 ( .A(n4320), .Y(n4319) );
  INVX2TS U2403 ( .A(n4314), .Y(n4313) );
  INVX2TS U2404 ( .A(n4311), .Y(n4310) );
  INVX2TS U2405 ( .A(n4290), .Y(n4289) );
  INVX2TS U2406 ( .A(n4287), .Y(n4286) );
  INVX2TS U2407 ( .A(n4281), .Y(n4280) );
  INVX2TS U2408 ( .A(n4269), .Y(n4268) );
  INVX2TS U2409 ( .A(n4254), .Y(n4253) );
  INVX2TS U2410 ( .A(n4344), .Y(n4343) );
  INVX2TS U2411 ( .A(n4341), .Y(n4340) );
  INVX2TS U2412 ( .A(n4335), .Y(n4334) );
  INVX2TS U2413 ( .A(n4332), .Y(n4331) );
  INVX2TS U2414 ( .A(n4329), .Y(n4328) );
  INVX2TS U2415 ( .A(n4323), .Y(n4322) );
  INVX2TS U2416 ( .A(n4317), .Y(n4316) );
  INVX2TS U2417 ( .A(n4308), .Y(n4307) );
  INVX2TS U2418 ( .A(n4302), .Y(n4301) );
  INVX2TS U2419 ( .A(n4299), .Y(n4298) );
  INVX2TS U2420 ( .A(n4296), .Y(n4295) );
  INVX2TS U2421 ( .A(n4293), .Y(n4292) );
  INVX2TS U2422 ( .A(n4284), .Y(n4283) );
  INVX2TS U2423 ( .A(n4278), .Y(n4277) );
  INVX2TS U2424 ( .A(n4275), .Y(n4274) );
  INVX2TS U2425 ( .A(n4272), .Y(n4271) );
  INVX2TS U2426 ( .A(n4266), .Y(n4265) );
  INVX2TS U2427 ( .A(n4260), .Y(n4259) );
  INVX2TS U2428 ( .A(n4257), .Y(n4256) );
  INVX2TS U2429 ( .A(n4251), .Y(n4250) );
  INVX2TS U2430 ( .A(n4326), .Y(n4325) );
  INVX2TS U2431 ( .A(n4305), .Y(n4304) );
  INVX2TS U2432 ( .A(n4263), .Y(n4262) );
  INVX2TS U2433 ( .A(n3960), .Y(n3959) );
  INVX2TS U2434 ( .A(n3948), .Y(n3947) );
  INVX2TS U2435 ( .A(n3963), .Y(n3962) );
  INVX2TS U2436 ( .A(n3957), .Y(n3956) );
  INVX2TS U2437 ( .A(n3954), .Y(n3953) );
  INVX2TS U2438 ( .A(n3951), .Y(n3950) );
  INVX2TS U2439 ( .A(n4191), .Y(n4190) );
  INVX2TS U2440 ( .A(n4188), .Y(n4187) );
  INVX2TS U2441 ( .A(n4182), .Y(n4181) );
  INVX2TS U2442 ( .A(n4185), .Y(n4184) );
  INVX2TS U2443 ( .A(n4179), .Y(n4178) );
  INVX2TS U2444 ( .A(n4176), .Y(n4175) );
  INVX2TS U2445 ( .A(n2948), .Y(n774) );
  INVX2TS U2446 ( .A(n2945), .Y(n773) );
  INVX2TS U2447 ( .A(n1932), .Y(n938) );
  INVX2TS U2448 ( .A(n1141), .Y(n775) );
  AOI21X1TS U2449 ( .A0(n915), .A1(n980), .B0(n2034), .Y(n2065) );
  AOI222XLTS U2450 ( .A0(n4193), .A1(n3449), .B0(n4198), .B1(n3428), .C0(n4206), .C1(n3411), .Y(n1801) );
  AOI222XLTS U2451 ( .A0(n4205), .A1(n3486), .B0(n4198), .B1(n3461), .C0(
        writeIn_WEST), .C1(n3514), .Y(n1798) );
  AOI222XLTS U2452 ( .A0(n4193), .A1(n3173), .B0(n4197), .B1(n3149), .C0(n4206), .C1(n796), .Y(n1809) );
  NOR3X1TS U2453 ( .A(n2938), .B(n986), .C(n2932), .Y(n2935) );
  NAND3X1TS U2454 ( .A(n926), .B(n1895), .C(n1942), .Y(n1853) );
  XNOR2X1TS U2455 ( .A(n43), .B(n2937), .Y(n1135) );
  NOR2X1TS U2456 ( .A(n2932), .B(n2938), .Y(n2937) );
  OAI21X1TS U2457 ( .A0(n979), .A1(n2064), .B0(n102), .Y(n2063) );
  NOR2X1TS U2458 ( .A(n974), .B(n986), .Y(n2034) );
  NOR2X1TS U2459 ( .A(n1964), .B(n927), .Y(n1893) );
  NAND2X1TS U2460 ( .A(n2062), .B(n43), .Y(n2060) );
  INVX2TS U2461 ( .A(n2064), .Y(n934) );
  AND3X2TS U2462 ( .A(n2924), .B(n927), .C(n925), .Y(n2067) );
  XOR2X1TS U2463 ( .A(n1138), .B(n1), .Y(n2939) );
  INVX2TS U2464 ( .A(n101), .Y(n935) );
  XOR2X1TS U2465 ( .A(n1139), .B(n466), .Y(n2928) );
  OAI22X1TS U2466 ( .A0(n773), .A1(n2941), .B0(n2946), .B1(n2933), .Y(n2943)
         );
  AOI32X1TS U2467 ( .A0(n2945), .A1(n1144), .A2(n775), .B0(n2946), .B1(n2933), 
        .Y(n2944) );
  AOI211XLTS U2468 ( .A0(n773), .A1(n2941), .B0(n1141), .C0(n2938), .Y(n2942)
         );
  OAI221XLTS U2469 ( .A0(n171), .A1(n984), .B0(n3320), .B1(n690), .C0(n1806), 
        .Y(n2572) );
  AOI222XLTS U2470 ( .A0(n4197), .A1(n3262), .B0(n4192), .B1(n3272), .C0(n4206), .C1(n3310), .Y(n1806) );
  AOI222XLTS U2471 ( .A0(n4205), .A1(n3369), .B0(n4192), .B1(n3347), .C0(n4197), .C1(n3397), .Y(n1804) );
  OAI221XLTS U2472 ( .A0(n475), .A1(n160), .B0(n3124), .B1(n767), .C0(n1793), 
        .Y(n2577) );
  AOI222XLTS U2473 ( .A0(n4205), .A1(n3639), .B0(n4192), .B1(n3613), .C0(n4197), .C1(n3774), .Y(n1793) );
  OAI22X1TS U2474 ( .A0(n102), .A1(n111), .B0(n935), .B1(n998), .Y(n1845) );
  NOR2X1TS U2475 ( .A(n1889), .B(n803), .Y(n1879) );
  INVX2TS U2476 ( .A(n1889), .Y(n936) );
  NOR2BX1TS U2477 ( .AN(n1908), .B(n2025), .Y(n1266) );
  NOR2BX1TS U2478 ( .AN(n1908), .B(n1987), .Y(n1234) );
  NOR2X1TS U2479 ( .A(n2073), .B(n153), .Y(n2103) );
  NOR2X1TS U2480 ( .A(n2074), .B(n154), .Y(n2090) );
  NOR2X1TS U2481 ( .A(n2076), .B(n155), .Y(n2089) );
  INVX2TS U2482 ( .A(n2088), .Y(n679) );
  AOI221X1TS U2483 ( .A0(writeIn_WEST), .A1(n3104), .B0(writeIn_SOUTH), .B1(
        n2967), .C0(n2091), .Y(n2088) );
  INVX2TS U2484 ( .A(writeIn_EAST), .Y(n4199) );
  INVX2TS U2485 ( .A(n2068), .Y(n3121) );
  NAND4BX1TS U2486 ( .AN(n153), .B(n2923), .C(n2075), .D(n2073), .Y(n2068) );
  AND3X2TS U2487 ( .A(n2076), .B(n2074), .C(n2077), .Y(n2923) );
  INVX2TS U2488 ( .A(n1918), .Y(n916) );
  OR2X2TS U2489 ( .A(n2075), .B(n155), .Y(n977) );
  OAI221XLTS U2490 ( .A0(n4203), .A1(n2075), .B0(n4196), .B1(n2076), .C0(n2077), .Y(n2071) );
  OAI22X1TS U2491 ( .A0(n843), .A1(n1071), .B0(n640), .B1(n1057), .Y(n2921) );
  OAI22X1TS U2492 ( .A0(n834), .A1(n1072), .B0(n639), .B1(n1057), .Y(n2915) );
  OAI22X1TS U2493 ( .A0(n833), .A1(n1071), .B0(n638), .B1(n1057), .Y(n2909) );
  OAI22X1TS U2494 ( .A0(n832), .A1(n2166), .B0(n637), .B1(n1056), .Y(n2903) );
  OAI22X1TS U2495 ( .A0(n831), .A1(n1059), .B0(n636), .B1(n1045), .Y(n2897) );
  OAI22X1TS U2496 ( .A0(n830), .A1(n1059), .B0(n635), .B1(n1045), .Y(n2891) );
  OAI22X1TS U2497 ( .A0(n829), .A1(n1059), .B0(n634), .B1(n1045), .Y(n2393) );
  OAI22X1TS U2498 ( .A0(n828), .A1(n1059), .B0(n633), .B1(n1045), .Y(n2387) );
  OAI22X1TS U2499 ( .A0(n827), .A1(n1070), .B0(n632), .B1(n1046), .Y(n2381) );
  OAI22X1TS U2500 ( .A0(n826), .A1(n1067), .B0(n631), .B1(n1046), .Y(n2375) );
  OAI22X1TS U2501 ( .A0(n825), .A1(n1066), .B0(n630), .B1(n1046), .Y(n2369) );
  OAI22X1TS U2502 ( .A0(n824), .A1(n1068), .B0(n629), .B1(n1046), .Y(n2363) );
  OAI22X1TS U2503 ( .A0(n823), .A1(n1069), .B0(n628), .B1(n1047), .Y(n2357) );
  OAI22X1TS U2504 ( .A0(n822), .A1(n1069), .B0(n627), .B1(n1047), .Y(n2351) );
  OAI22X1TS U2505 ( .A0(n821), .A1(n1069), .B0(n626), .B1(n1047), .Y(n2345) );
  OAI22X1TS U2506 ( .A0(n842), .A1(n1070), .B0(n625), .B1(n1047), .Y(n2339) );
  OAI22X1TS U2507 ( .A0(n841), .A1(n1069), .B0(n624), .B1(n1048), .Y(n2333) );
  OAI22X1TS U2508 ( .A0(n820), .A1(n1067), .B0(n623), .B1(n1048), .Y(n2327) );
  OAI22X1TS U2509 ( .A0(n819), .A1(n1066), .B0(n622), .B1(n1048), .Y(n2321) );
  OAI22X1TS U2510 ( .A0(n818), .A1(n1068), .B0(n621), .B1(n1048), .Y(n2315) );
  OAI22X1TS U2511 ( .A0(n840), .A1(n1060), .B0(n620), .B1(n1056), .Y(n2309) );
  OAI22X1TS U2512 ( .A0(n817), .A1(n1060), .B0(n619), .B1(n1055), .Y(n2303) );
  OAI22X1TS U2513 ( .A0(n816), .A1(n1060), .B0(n618), .B1(n1055), .Y(n2297) );
  OAI22X1TS U2514 ( .A0(n815), .A1(n1060), .B0(n617), .B1(n1054), .Y(n2291) );
  OAI22X1TS U2515 ( .A0(n814), .A1(n1061), .B0(n616), .B1(n1049), .Y(n2285) );
  OAI22X1TS U2516 ( .A0(n813), .A1(n1061), .B0(n615), .B1(n1049), .Y(n2279) );
  OAI22X1TS U2517 ( .A0(n812), .A1(n1061), .B0(n614), .B1(n1049), .Y(n2273) );
  OAI22X1TS U2518 ( .A0(n811), .A1(n1061), .B0(n613), .B1(n1049), .Y(n2267) );
  OAI22X1TS U2519 ( .A0(n810), .A1(n1062), .B0(n612), .B1(n1050), .Y(n2261) );
  OAI22X1TS U2520 ( .A0(n809), .A1(n1062), .B0(n611), .B1(n1050), .Y(n2255) );
  OAI22X1TS U2521 ( .A0(n839), .A1(n1062), .B0(n610), .B1(n1050), .Y(n2249) );
  OAI22X1TS U2522 ( .A0(n808), .A1(n1062), .B0(n609), .B1(n1050), .Y(n2243) );
  OAI22X1TS U2523 ( .A0(n893), .A1(n1063), .B0(n689), .B1(n1051), .Y(n2237) );
  OAI22X1TS U2524 ( .A0(n892), .A1(n1063), .B0(n688), .B1(n1051), .Y(n2231) );
  OAI22X1TS U2525 ( .A0(n890), .A1(n1063), .B0(n687), .B1(n1051), .Y(n2219) );
  OAI22X1TS U2526 ( .A0(n889), .A1(n1064), .B0(n685), .B1(n1052), .Y(n2213) );
  OAI22X1TS U2527 ( .A0(n909), .A1(n1064), .B0(n644), .B1(n1052), .Y(n2201) );
  OAI22X1TS U2528 ( .A0(n807), .A1(n1064), .B0(n666), .B1(n1052), .Y(n2195) );
  OAI22X1TS U2529 ( .A0(n838), .A1(n1065), .B0(n643), .B1(n1053), .Y(n2189) );
  OAI22X1TS U2530 ( .A0(n837), .A1(n1065), .B0(n642), .B1(n1053), .Y(n2183) );
  OAI22X1TS U2531 ( .A0(n836), .A1(n1065), .B0(n641), .B1(n1053), .Y(n2177) );
  OAI22X1TS U2532 ( .A0(n835), .A1(n1065), .B0(n665), .B1(n1053), .Y(n2165) );
  OAI22X1TS U2533 ( .A0(n891), .A1(n1063), .B0(n686), .B1(n1051), .Y(n2225) );
  OAI22X1TS U2534 ( .A0(n888), .A1(n1064), .B0(n684), .B1(n1052), .Y(n2207) );
  OAI22X1TS U2535 ( .A0(n111), .A1(n2073), .B0(n457), .B1(n2074), .Y(n2072) );
  NOR2X1TS U2536 ( .A(n2085), .B(n130), .Y(n2170) );
  NOR2X1TS U2537 ( .A(n2083), .B(n131), .Y(n2163) );
  NOR2X1TS U2538 ( .A(n2084), .B(n131), .Y(n2168) );
  NOR2X1TS U2539 ( .A(n2086), .B(n130), .Y(n2169) );
  NOR2X1TS U2540 ( .A(n2077), .B(n154), .Y(n2172) );
  NAND2X1TS U2541 ( .A(n185), .B(n478), .Y(n1146) );
  OAI21X1TS U2542 ( .A0(n124), .A1(n1145), .B0(n3756), .Y(n2884) );
  INVX2TS U2543 ( .A(requesterAddressIn_WEST[4]), .Y(n4038) );
  INVX2TS U2544 ( .A(requesterAddressIn_WEST[5]), .Y(n4041) );
  INVX2TS U2545 ( .A(requesterAddressIn_WEST[3]), .Y(n4035) );
  INVX2TS U2546 ( .A(requesterAddressIn_WEST[2]), .Y(n4032) );
  INVX2TS U2547 ( .A(requesterAddressIn_WEST[1]), .Y(n4029) );
  INVX2TS U2548 ( .A(requesterAddressIn_WEST[0]), .Y(n4026) );
  INVX2TS U2549 ( .A(requesterAddressIn_EAST[4]), .Y(n4188) );
  INVX2TS U2550 ( .A(requesterAddressIn_EAST[1]), .Y(n4179) );
  INVX2TS U2551 ( .A(requesterAddressIn_EAST[0]), .Y(n4176) );
  INVX2TS U2552 ( .A(requesterAddressIn_EAST[5]), .Y(n4191) );
  INVX2TS U2553 ( .A(requesterAddressIn_EAST[3]), .Y(n4185) );
  INVX2TS U2554 ( .A(requesterAddressIn_EAST[2]), .Y(n4182) );
  INVX2TS U2555 ( .A(destinationAddressIn_WEST[5]), .Y(n4005) );
  INVX2TS U2556 ( .A(destinationAddressIn_WEST[4]), .Y(n4002) );
  INVX2TS U2557 ( .A(destinationAddressIn_WEST[3]), .Y(n3999) );
  INVX2TS U2558 ( .A(destinationAddressIn_WEST[1]), .Y(n3993) );
  INVX2TS U2559 ( .A(destinationAddressIn_WEST[0]), .Y(n3990) );
  INVX2TS U2560 ( .A(dataIn_WEST[31]), .Y(n4344) );
  INVX2TS U2561 ( .A(dataIn_WEST[30]), .Y(n4341) );
  INVX2TS U2562 ( .A(dataIn_WEST[29]), .Y(n4338) );
  INVX2TS U2563 ( .A(dataIn_WEST[28]), .Y(n4335) );
  INVX2TS U2564 ( .A(dataIn_WEST[27]), .Y(n4332) );
  INVX2TS U2565 ( .A(dataIn_WEST[26]), .Y(n4329) );
  INVX2TS U2566 ( .A(dataIn_WEST[24]), .Y(n4323) );
  INVX2TS U2567 ( .A(dataIn_WEST[22]), .Y(n4317) );
  INVX2TS U2568 ( .A(dataIn_WEST[21]), .Y(n4314) );
  INVX2TS U2569 ( .A(dataIn_WEST[19]), .Y(n4308) );
  INVX2TS U2570 ( .A(dataIn_WEST[17]), .Y(n4302) );
  INVX2TS U2571 ( .A(dataIn_WEST[16]), .Y(n4299) );
  INVX2TS U2572 ( .A(dataIn_WEST[14]), .Y(n4293) );
  INVX2TS U2573 ( .A(dataIn_WEST[12]), .Y(n4287) );
  INVX2TS U2574 ( .A(dataIn_WEST[11]), .Y(n4284) );
  INVX2TS U2575 ( .A(dataIn_WEST[10]), .Y(n4281) );
  INVX2TS U2576 ( .A(dataIn_WEST[9]), .Y(n4278) );
  INVX2TS U2577 ( .A(dataIn_WEST[8]), .Y(n4275) );
  INVX2TS U2578 ( .A(dataIn_WEST[6]), .Y(n4269) );
  INVX2TS U2579 ( .A(dataIn_WEST[3]), .Y(n4260) );
  INVX2TS U2580 ( .A(dataIn_WEST[1]), .Y(n4254) );
  INVX2TS U2581 ( .A(dataIn_WEST[0]), .Y(n4251) );
  INVX2TS U2582 ( .A(destinationAddressIn_WEST[2]), .Y(n3996) );
  INVX2TS U2583 ( .A(dataIn_WEST[25]), .Y(n4326) );
  INVX2TS U2584 ( .A(dataIn_WEST[23]), .Y(n4320) );
  INVX2TS U2585 ( .A(dataIn_WEST[20]), .Y(n4311) );
  INVX2TS U2586 ( .A(dataIn_WEST[18]), .Y(n4305) );
  INVX2TS U2587 ( .A(dataIn_WEST[15]), .Y(n4296) );
  INVX2TS U2588 ( .A(dataIn_WEST[13]), .Y(n4290) );
  INVX2TS U2589 ( .A(dataIn_WEST[5]), .Y(n4266) );
  INVX2TS U2590 ( .A(dataIn_WEST[4]), .Y(n4263) );
  INVX2TS U2591 ( .A(dataIn_WEST[2]), .Y(n4257) );
  INVX2TS U2592 ( .A(dataIn_WEST[7]), .Y(n4272) );
  INVX2TS U2593 ( .A(destinationAddressIn_EAST[4]), .Y(n3960) );
  INVX2TS U2594 ( .A(destinationAddressIn_EAST[3]), .Y(n3957) );
  INVX2TS U2595 ( .A(destinationAddressIn_EAST[2]), .Y(n3954) );
  INVX2TS U2596 ( .A(destinationAddressIn_EAST[1]), .Y(n3951) );
  INVX2TS U2597 ( .A(destinationAddressIn_EAST[0]), .Y(n3948) );
  INVX2TS U2598 ( .A(destinationAddressIn_EAST[5]), .Y(n3963) );
  INVX2TS U2599 ( .A(readIn_WEST), .Y(n4196) );
  INVX2TS U2600 ( .A(destinationAddressIn_EAST[13]), .Y(n3987) );
  INVX2TS U2601 ( .A(destinationAddressIn_EAST[11]), .Y(n3981) );
  INVX2TS U2602 ( .A(destinationAddressIn_EAST[9]), .Y(n3975) );
  INVX2TS U2603 ( .A(destinationAddressIn_EAST[7]), .Y(n3969) );
  INVX2TS U2604 ( .A(destinationAddressIn_EAST[12]), .Y(n3984) );
  INVX2TS U2605 ( .A(destinationAddressIn_EAST[10]), .Y(n3978) );
  INVX2TS U2606 ( .A(destinationAddressIn_EAST[8]), .Y(n3972) );
  INVX2TS U2607 ( .A(destinationAddressIn_EAST[6]), .Y(n3966) );
  INVX2TS U2608 ( .A(dataIn_EAST[31]), .Y(n4442) );
  INVX2TS U2609 ( .A(dataIn_EAST[30]), .Y(n4438) );
  INVX2TS U2610 ( .A(dataIn_EAST[29]), .Y(n4435) );
  INVX2TS U2611 ( .A(dataIn_EAST[28]), .Y(n4432) );
  INVX2TS U2612 ( .A(dataIn_EAST[27]), .Y(n4428) );
  INVX2TS U2613 ( .A(dataIn_EAST[26]), .Y(n4425) );
  INVX2TS U2614 ( .A(dataIn_EAST[24]), .Y(n4419) );
  INVX2TS U2615 ( .A(dataIn_EAST[23]), .Y(n4416) );
  INVX2TS U2616 ( .A(dataIn_EAST[22]), .Y(n4413) );
  INVX2TS U2617 ( .A(dataIn_EAST[21]), .Y(n4410) );
  INVX2TS U2618 ( .A(dataIn_EAST[20]), .Y(n4407) );
  INVX2TS U2619 ( .A(dataIn_EAST[19]), .Y(n4404) );
  INVX2TS U2620 ( .A(dataIn_EAST[17]), .Y(n4398) );
  INVX2TS U2621 ( .A(dataIn_EAST[16]), .Y(n4395) );
  INVX2TS U2622 ( .A(dataIn_EAST[15]), .Y(n4392) );
  INVX2TS U2623 ( .A(dataIn_EAST[14]), .Y(n4389) );
  INVX2TS U2624 ( .A(dataIn_EAST[13]), .Y(n4386) );
  INVX2TS U2625 ( .A(dataIn_EAST[12]), .Y(n4383) );
  INVX2TS U2626 ( .A(dataIn_EAST[11]), .Y(n4380) );
  INVX2TS U2627 ( .A(dataIn_EAST[10]), .Y(n4377) );
  INVX2TS U2628 ( .A(dataIn_EAST[9]), .Y(n4374) );
  INVX2TS U2629 ( .A(dataIn_EAST[8]), .Y(n4371) );
  INVX2TS U2630 ( .A(dataIn_EAST[7]), .Y(n4368) );
  INVX2TS U2631 ( .A(dataIn_EAST[6]), .Y(n4365) );
  INVX2TS U2632 ( .A(dataIn_EAST[5]), .Y(n4362) );
  INVX2TS U2633 ( .A(dataIn_EAST[3]), .Y(n4356) );
  INVX2TS U2634 ( .A(dataIn_EAST[2]), .Y(n4353) );
  INVX2TS U2635 ( .A(dataIn_EAST[1]), .Y(n4350) );
  INVX2TS U2636 ( .A(dataIn_EAST[0]), .Y(n4347) );
  INVX2TS U2637 ( .A(dataIn_EAST[25]), .Y(n4422) );
  INVX2TS U2638 ( .A(dataIn_EAST[18]), .Y(n4401) );
  INVX2TS U2639 ( .A(dataIn_EAST[4]), .Y(n4359) );
  INVX2TS U2640 ( .A(requesterAddressIn_SOUTH[4]), .Y(n4567) );
  INVX2TS U2641 ( .A(requesterAddressIn_SOUTH[1]), .Y(n4556) );
  INVX2TS U2642 ( .A(requesterAddressIn_SOUTH[0]), .Y(n4553) );
  INVX2TS U2643 ( .A(requesterAddressIn_SOUTH[5]), .Y(n4570) );
  INVX2TS U2644 ( .A(requesterAddressIn_SOUTH[3]), .Y(n4563) );
  INVX2TS U2645 ( .A(requesterAddressIn_SOUTH[2]), .Y(n4560) );
  INVX2TS U2646 ( .A(destinationAddressIn_SOUTH[4]), .Y(n4221) );
  INVX2TS U2647 ( .A(destinationAddressIn_SOUTH[0]), .Y(n4209) );
  INVX2TS U2648 ( .A(destinationAddressIn_SOUTH[5]), .Y(n4224) );
  INVX2TS U2649 ( .A(destinationAddressIn_SOUTH[3]), .Y(n4218) );
  INVX2TS U2650 ( .A(destinationAddressIn_SOUTH[2]), .Y(n4215) );
  INVX2TS U2651 ( .A(destinationAddressIn_SOUTH[1]), .Y(n4212) );
  INVX2TS U2652 ( .A(dataIn_SOUTH[31]), .Y(n4550) );
  INVX2TS U2653 ( .A(dataIn_SOUTH[30]), .Y(n4546) );
  INVX2TS U2654 ( .A(dataIn_SOUTH[29]), .Y(n4543) );
  INVX2TS U2655 ( .A(dataIn_SOUTH[28]), .Y(n4540) );
  INVX2TS U2656 ( .A(dataIn_SOUTH[27]), .Y(n4536) );
  INVX2TS U2657 ( .A(dataIn_SOUTH[26]), .Y(n4533) );
  INVX2TS U2658 ( .A(dataIn_SOUTH[24]), .Y(n4526) );
  INVX2TS U2659 ( .A(dataIn_SOUTH[23]), .Y(n4523) );
  INVX2TS U2660 ( .A(dataIn_SOUTH[22]), .Y(n4519) );
  INVX2TS U2661 ( .A(dataIn_SOUTH[21]), .Y(n4516) );
  INVX2TS U2662 ( .A(dataIn_SOUTH[20]), .Y(n4513) );
  INVX2TS U2663 ( .A(dataIn_SOUTH[19]), .Y(n4509) );
  INVX2TS U2664 ( .A(dataIn_SOUTH[17]), .Y(n4502) );
  INVX2TS U2665 ( .A(dataIn_SOUTH[16]), .Y(n4499) );
  INVX2TS U2666 ( .A(dataIn_SOUTH[15]), .Y(n4496) );
  INVX2TS U2667 ( .A(dataIn_SOUTH[14]), .Y(n4492) );
  INVX2TS U2668 ( .A(dataIn_SOUTH[13]), .Y(n4489) );
  INVX2TS U2669 ( .A(dataIn_SOUTH[12]), .Y(n4486) );
  INVX2TS U2670 ( .A(dataIn_SOUTH[11]), .Y(n4482) );
  INVX2TS U2671 ( .A(dataIn_SOUTH[10]), .Y(n4479) );
  INVX2TS U2672 ( .A(dataIn_SOUTH[9]), .Y(n4475) );
  INVX2TS U2673 ( .A(dataIn_SOUTH[8]), .Y(n4472) );
  INVX2TS U2674 ( .A(dataIn_SOUTH[7]), .Y(n4469) );
  INVX2TS U2675 ( .A(dataIn_SOUTH[6]), .Y(n4465) );
  INVX2TS U2676 ( .A(dataIn_SOUTH[5]), .Y(n4462) );
  INVX2TS U2677 ( .A(dataIn_SOUTH[3]), .Y(n4455) );
  INVX2TS U2678 ( .A(dataIn_SOUTH[2]), .Y(n4452) );
  INVX2TS U2679 ( .A(dataIn_SOUTH[1]), .Y(n4448) );
  INVX2TS U2680 ( .A(dataIn_SOUTH[0]), .Y(n4445) );
  INVX2TS U2681 ( .A(dataIn_SOUTH[25]), .Y(n4529) );
  INVX2TS U2682 ( .A(dataIn_SOUTH[18]), .Y(n4506) );
  INVX2TS U2683 ( .A(dataIn_SOUTH[4]), .Y(n4459) );
  CLKBUFX2TS U2684 ( .A(writeIn_WEST), .Y(n4192) );
  CLKBUFX2TS U2685 ( .A(writeIn_SOUTH), .Y(n4204) );
  CLKBUFX2TS U2686 ( .A(destinationAddressIn_SOUTH[13]), .Y(n4246) );
  CLKBUFX2TS U2687 ( .A(destinationAddressIn_SOUTH[11]), .Y(n4240) );
  CLKBUFX2TS U2688 ( .A(destinationAddressIn_SOUTH[9]), .Y(n4234) );
  CLKBUFX2TS U2689 ( .A(destinationAddressIn_SOUTH[12]), .Y(n4243) );
  CLKBUFX2TS U2690 ( .A(destinationAddressIn_SOUTH[10]), .Y(n4237) );
  CLKBUFX2TS U2691 ( .A(destinationAddressIn_SOUTH[8]), .Y(n4231) );
  CLKBUFX2TS U2692 ( .A(requesterAddressIn_NORTH[4]), .Y(n4072) );
  CLKBUFX2TS U2693 ( .A(requesterAddressIn_NORTH[1]), .Y(n4063) );
  CLKBUFX2TS U2694 ( .A(requesterAddressIn_NORTH[0]), .Y(n4060) );
  CLKBUFX2TS U2695 ( .A(requesterAddressIn_NORTH[5]), .Y(n4075) );
  CLKBUFX2TS U2696 ( .A(requesterAddressIn_NORTH[3]), .Y(n4069) );
  CLKBUFX2TS U2697 ( .A(requesterAddressIn_NORTH[2]), .Y(n4066) );
  CLKBUFX2TS U2698 ( .A(destinationAddressIn_NORTH[4]), .Y(n4054) );
  CLKBUFX2TS U2699 ( .A(destinationAddressIn_NORTH[0]), .Y(n4042) );
  CLKBUFX2TS U2700 ( .A(destinationAddressIn_NORTH[5]), .Y(n4057) );
  CLKBUFX2TS U2701 ( .A(destinationAddressIn_NORTH[3]), .Y(n4051) );
  CLKBUFX2TS U2702 ( .A(destinationAddressIn_NORTH[2]), .Y(n4048) );
  CLKBUFX2TS U2703 ( .A(destinationAddressIn_NORTH[1]), .Y(n4045) );
  CLKBUFX2TS U2704 ( .A(dataIn_NORTH[31]), .Y(n4171) );
  CLKBUFX2TS U2705 ( .A(dataIn_NORTH[30]), .Y(n4168) );
  CLKBUFX2TS U2706 ( .A(dataIn_NORTH[29]), .Y(n4165) );
  CLKBUFX2TS U2707 ( .A(dataIn_NORTH[28]), .Y(n4162) );
  CLKBUFX2TS U2708 ( .A(dataIn_NORTH[27]), .Y(n4159) );
  CLKBUFX2TS U2709 ( .A(dataIn_NORTH[26]), .Y(n4156) );
  CLKBUFX2TS U2710 ( .A(dataIn_NORTH[24]), .Y(n4150) );
  CLKBUFX2TS U2711 ( .A(dataIn_NORTH[23]), .Y(n4147) );
  CLKBUFX2TS U2712 ( .A(dataIn_NORTH[22]), .Y(n4144) );
  CLKBUFX2TS U2713 ( .A(dataIn_NORTH[21]), .Y(n4141) );
  CLKBUFX2TS U2714 ( .A(dataIn_NORTH[20]), .Y(n4138) );
  CLKBUFX2TS U2715 ( .A(dataIn_NORTH[19]), .Y(n4135) );
  CLKBUFX2TS U2716 ( .A(dataIn_NORTH[17]), .Y(n4129) );
  CLKBUFX2TS U2717 ( .A(dataIn_NORTH[16]), .Y(n4126) );
  CLKBUFX2TS U2718 ( .A(dataIn_NORTH[15]), .Y(n4123) );
  CLKBUFX2TS U2719 ( .A(dataIn_NORTH[14]), .Y(n4120) );
  CLKBUFX2TS U2720 ( .A(dataIn_NORTH[13]), .Y(n4117) );
  CLKBUFX2TS U2721 ( .A(dataIn_NORTH[12]), .Y(n4114) );
  CLKBUFX2TS U2722 ( .A(dataIn_NORTH[11]), .Y(n4111) );
  CLKBUFX2TS U2723 ( .A(dataIn_NORTH[10]), .Y(n4108) );
  CLKBUFX2TS U2724 ( .A(dataIn_NORTH[9]), .Y(n4105) );
  CLKBUFX2TS U2725 ( .A(dataIn_NORTH[7]), .Y(n4099) );
  CLKBUFX2TS U2726 ( .A(dataIn_NORTH[6]), .Y(n4096) );
  CLKBUFX2TS U2727 ( .A(dataIn_NORTH[5]), .Y(n4093) );
  CLKBUFX2TS U2728 ( .A(dataIn_NORTH[3]), .Y(n4087) );
  CLKBUFX2TS U2729 ( .A(dataIn_NORTH[2]), .Y(n4084) );
  CLKBUFX2TS U2730 ( .A(dataIn_NORTH[1]), .Y(n4081) );
  CLKBUFX2TS U2731 ( .A(dataIn_NORTH[0]), .Y(n4078) );
  CLKBUFX2TS U2732 ( .A(dataIn_NORTH[25]), .Y(n4153) );
  CLKBUFX2TS U2733 ( .A(dataIn_NORTH[18]), .Y(n4132) );
  CLKBUFX2TS U2734 ( .A(dataIn_NORTH[4]), .Y(n4090) );
  CLKBUFX2TS U2735 ( .A(destinationAddressIn_WEST[13]), .Y(n4022) );
  CLKBUFX2TS U2736 ( .A(destinationAddressIn_WEST[11]), .Y(n4018) );
  CLKBUFX2TS U2737 ( .A(destinationAddressIn_WEST[7]), .Y(n4009) );
  CLKBUFX2TS U2738 ( .A(destinationAddressIn_WEST[12]), .Y(n4020) );
  CLKBUFX2TS U2739 ( .A(destinationAddressIn_WEST[8]), .Y(n4012) );
  CLKBUFX2TS U2740 ( .A(destinationAddressIn_WEST[6]), .Y(n4006) );
  CLKBUFX2TS U2741 ( .A(dataIn_NORTH[8]), .Y(n4102) );
  NOR2X1TS U2742 ( .A(n782), .B(n1140), .Y(n2885) );
  AOI31X1TS U2743 ( .A0(n773), .A1(n1141), .A2(n1142), .B0(n131), .Y(n1140) );
  XNOR2X1TS U2744 ( .A(n1143), .B(n1144), .Y(n1142) );
  INVX2TS U2745 ( .A(readIn_EAST), .Y(n4203) );
  NAND2X1TS U2746 ( .A(n43), .B(n128), .Y(n2948) );
  XOR2X1TS U2747 ( .A(n942), .B(n124), .Y(n1144) );
  XOR2X1TS U2748 ( .A(n2953), .B(n774), .Y(n2945) );
  XOR2X1TS U2749 ( .A(n122), .B(n157), .Y(n2953) );
  OAI21X1TS U2750 ( .A0(n129), .A1(n3), .B0(n2948), .Y(n1141) );
  CLKBUFX2TS U2751 ( .A(n2087), .Y(n978) );
  NOR2X1TS U2752 ( .A(n1143), .B(n466), .Y(n2087) );
  INVX2TS U2753 ( .A(n1987), .Y(n940) );
  OAI22X1TS U2754 ( .A0(n691), .A1(n2099), .B0(n690), .B1(n2083), .Y(n2094) );
  OAI22X1TS U2755 ( .A0(n765), .A1(n2084), .B0(n970), .B1(n2085), .Y(n2097) );
  OAI22X1TS U2756 ( .A0(n772), .A1(n766), .B0(n767), .B1(n2086), .Y(n2096) );
  OAI22X1TS U2757 ( .A0(n772), .A1(n676), .B0(n2082), .B1(n681), .Y(n2081) );
  OAI22X1TS U2758 ( .A0(n2083), .A1(n682), .B0(n2084), .B1(n683), .Y(n2080) );
  INVX2TS U2759 ( .A(n2086), .Y(n777) );
  INVX2TS U2760 ( .A(n2082), .Y(n770) );
  INVX2TS U2761 ( .A(n184), .Y(n772) );
  NOR2X1TS U2762 ( .A(readReady), .B(selectBit_WEST), .Y(n2924) );
  AOI222XLTS U2763 ( .A0(n4019), .A1(n3447), .B0(n3980), .B1(n3430), .C0(n4242), .C1(n3412), .Y(n1983) );
  AOI222XLTS U2764 ( .A0(n4007), .A1(n3449), .B0(n3965), .B1(n3428), .C0(n4227), .C1(n3411), .Y(n1978) );
  AOI222XLTS U2765 ( .A0(n4021), .A1(n3447), .B0(n3983), .B1(n3431), .C0(n4245), .C1(n3412), .Y(n1984) );
  AOI222XLTS U2766 ( .A0(n4014), .A1(n3448), .B0(n3974), .B1(n3431), .C0(n4236), .C1(n3412), .Y(n1981) );
  AOI222XLTS U2767 ( .A0(n4013), .A1(n3448), .B0(n3971), .B1(n3428), .C0(n4233), .C1(n3411), .Y(n1980) );
  AOI222XLTS U2768 ( .A0(n4023), .A1(n3447), .B0(n3986), .B1(n3434), .C0(n4248), .C1(n3417), .Y(n1985) );
  AOI222XLTS U2769 ( .A0(n4016), .A1(n3448), .B0(n3977), .B1(n3430), .C0(n4239), .C1(n3412), .Y(n1982) );
  AOI222XLTS U2770 ( .A0(n4010), .A1(n3449), .B0(n3968), .B1(n3428), .C0(n4230), .C1(n3418), .Y(n1979) );
  AOI222XLTS U2771 ( .A0(n4226), .A1(n3485), .B0(n3965), .B1(n3461), .C0(n4008), .C1(n3514), .Y(n1955) );
  AOI222XLTS U2772 ( .A0(n4229), .A1(n3485), .B0(n3968), .B1(n3461), .C0(n4011), .C1(n3514), .Y(n1956) );
  AOI222XLTS U2773 ( .A0(n4232), .A1(n3485), .B0(n3971), .B1(n3461), .C0(
        destinationAddressIn_WEST[8]), .C1(n3513), .Y(n1957) );
  AOI222XLTS U2774 ( .A0(n4244), .A1(n3484), .B0(n3983), .B1(n3462), .C0(
        destinationAddressIn_WEST[12]), .C1(n3512), .Y(n1961) );
  AOI222XLTS U2775 ( .A0(n4241), .A1(n3484), .B0(n3980), .B1(n3462), .C0(
        destinationAddressIn_WEST[11]), .C1(n3512), .Y(n1960) );
  AOI222XLTS U2776 ( .A0(n4238), .A1(n3484), .B0(n3977), .B1(n3462), .C0(n4017), .C1(n3513), .Y(n1959) );
  AOI222XLTS U2777 ( .A0(n4247), .A1(n3484), .B0(n3986), .B1(n3468), .C0(
        destinationAddressIn_WEST[13]), .C1(n3512), .Y(n1962) );
  AOI222XLTS U2778 ( .A0(n4235), .A1(n3485), .B0(n3974), .B1(n3462), .C0(n4015), .C1(n3513), .Y(n1958) );
  AOI222XLTS U2779 ( .A0(n4021), .A1(n3171), .B0(n3982), .B1(n3151), .C0(n4245), .C1(n796), .Y(n2053) );
  AOI222XLTS U2780 ( .A0(n4013), .A1(n3172), .B0(n3970), .B1(n3149), .C0(n4233), .C1(n796), .Y(n2049) );
  AOI222XLTS U2781 ( .A0(n4023), .A1(n3171), .B0(n3985), .B1(n1267), .C0(n4248), .C1(n799), .Y(n2054) );
  AOI222XLTS U2782 ( .A0(n4016), .A1(n3171), .B0(n3976), .B1(n3152), .C0(n4239), .C1(n796), .Y(n2051) );
  AOI222XLTS U2783 ( .A0(n4007), .A1(n3172), .B0(n3964), .B1(n3149), .C0(n4227), .C1(n1810), .Y(n2047) );
  AOI222XLTS U2784 ( .A0(n4019), .A1(n3171), .B0(n3979), .B1(n3151), .C0(n4242), .C1(n799), .Y(n2052) );
  AOI222XLTS U2785 ( .A0(n4014), .A1(n3172), .B0(n3973), .B1(n3152), .C0(n4236), .C1(n799), .Y(n2050) );
  AOI222XLTS U2786 ( .A0(n4010), .A1(n3172), .B0(n3967), .B1(n3149), .C0(n4230), .C1(n799), .Y(n2048) );
  XNOR2X1TS U2787 ( .A(n2929), .B(n2930), .Y(n1139) );
  XOR2X1TS U2788 ( .A(n494), .B(n2931), .Y(n2930) );
  OAI21X1TS U2789 ( .A0(n2934), .A1(n2935), .B0(n2936), .Y(n2929) );
  NOR2X1TS U2790 ( .A(n2932), .B(n2933), .Y(n2931) );
  AOI22X1TS U2791 ( .A0(n3629), .A1(n34), .B0(n4000), .B1(n3615), .Y(n1904) );
  AOI222XLTS U2792 ( .A0(n3049), .A1(n3138), .B0(n4220), .B1(n3644), .C0(n4055), .C1(n3783), .Y(n1905) );
  AOI22X1TS U2793 ( .A0(n3626), .A1(n30), .B0(n3997), .B1(n3614), .Y(n1902) );
  AOI222XLTS U2794 ( .A0(n3051), .A1(n3138), .B0(n4217), .B1(n3646), .C0(n4052), .C1(n3783), .Y(n1903) );
  AOI22X1TS U2795 ( .A0(n3625), .A1(n26), .B0(n3994), .B1(n3602), .Y(n1900) );
  AOI222XLTS U2796 ( .A0(n3053), .A1(n975), .B0(n4214), .B1(n3644), .C0(n4049), 
        .C1(n3783), .Y(n1901) );
  AOI22X1TS U2797 ( .A0(n3618), .A1(n20), .B0(n3991), .B1(n3614), .Y(n1898) );
  AOI222XLTS U2798 ( .A0(n3055), .A1(n3139), .B0(n4211), .B1(n3646), .C0(n4046), .C1(n3782), .Y(n1899) );
  AOI22X1TS U2799 ( .A0(n3627), .A1(n14), .B0(n3988), .B1(n3617), .Y(n1896) );
  AOI222XLTS U2800 ( .A0(n3057), .A1(n3137), .B0(n4208), .B1(n3642), .C0(n4043), .C1(n3782), .Y(n1897) );
  AOI22X1TS U2801 ( .A0(n3629), .A1(n41), .B0(n4003), .B1(n3602), .Y(n1906) );
  AOI222XLTS U2802 ( .A0(n3047), .A1(n3135), .B0(n4223), .B1(n3648), .C0(n4058), .C1(n3783), .Y(n1907) );
  AOI22X1TS U2803 ( .A0(n3618), .A1(n17), .B0(n3601), .B1(n4024), .Y(n1167) );
  AOI222XLTS U2804 ( .A0(\requesterAddressbuffer[6][0] ), .A1(n3137), .B0(
        n3647), .B1(n4552), .C0(n3782), .C1(n4062), .Y(n1168) );
  AOI22X1TS U2805 ( .A0(n3618), .A1(n42), .B0(n3602), .B1(n4039), .Y(n1180) );
  AOI222XLTS U2806 ( .A0(\requesterAddressbuffer[6][5] ), .A1(n3137), .B0(
        n3645), .B1(n4569), .C0(n3782), .C1(n4077), .Y(n1181) );
  AOI22X1TS U2807 ( .A0(n3618), .A1(n37), .B0(n3601), .B1(n4036), .Y(n1178) );
  AOI222XLTS U2808 ( .A0(\requesterAddressbuffer[6][4] ), .A1(n3136), .B0(
        n3641), .B1(n4565), .C0(n3781), .C1(n4074), .Y(n1179) );
  AOI22X1TS U2809 ( .A0(n3629), .A1(n32), .B0(n3601), .B1(n4033), .Y(n1176) );
  AOI222XLTS U2810 ( .A0(\requesterAddressbuffer[6][3] ), .A1(n3137), .B0(
        n3641), .B1(n4562), .C0(n3781), .C1(n4071), .Y(n1177) );
  AOI22X1TS U2811 ( .A0(n3630), .A1(n27), .B0(n3601), .B1(n4030), .Y(n1174) );
  AOI222XLTS U2812 ( .A0(\requesterAddressbuffer[6][2] ), .A1(n3134), .B0(
        n3641), .B1(n4559), .C0(n3781), .C1(n4068), .Y(n1175) );
  AOI22X1TS U2813 ( .A0(n3631), .A1(n19), .B0(n3602), .B1(n4027), .Y(n1172) );
  AOI222XLTS U2814 ( .A0(\requesterAddressbuffer[6][1] ), .A1(n3133), .B0(
        n3641), .B1(n4555), .C0(n3781), .C1(n4065), .Y(n1173) );
  OAI2BB2XLTS U2815 ( .B0(n5326), .B1(n2034), .A0N(n1880), .A1N(n2034), .Y(
        n2066) );
  OAI22X1TS U2816 ( .A0(n1136), .A1(n1139), .B0(n494), .B1(n1137), .Y(n2886)
         );
  NAND2X1TS U2817 ( .A(selectBit_EAST), .B(n1964), .Y(n2010) );
  INVX2TS U2818 ( .A(readReady), .Y(n1132) );
  OAI32X1TS U2819 ( .A0(n2926), .A1(n2927), .A2(n2928), .B0(n155), .B1(n781), 
        .Y(N4718) );
  XOR2X1TS U2820 ( .A(n1135), .B(n128), .Y(n2927) );
  NAND2X1TS U2821 ( .A(n2939), .B(n782), .Y(n2926) );
  OAI221XLTS U2822 ( .A0(n1805), .A1(n147), .B0(n3318), .B1(n596), .C0(n2032), 
        .Y(n2466) );
  AOI222XLTS U2823 ( .A0(n3982), .A1(n3264), .B0(destinationAddressIn_WEST[12]), .B1(n3270), .C0(destinationAddressIn_SOUTH[12]), .C1(n3311), .Y(n2032) );
  OAI221XLTS U2824 ( .A0(n170), .A1(n143), .B0(n3318), .B1(n595), .C0(n2031), 
        .Y(n2467) );
  AOI222XLTS U2825 ( .A0(n3979), .A1(n3265), .B0(destinationAddressIn_WEST[11]), .B1(n3270), .C0(destinationAddressIn_SOUTH[11]), .C1(n3311), .Y(n2031) );
  OAI221XLTS U2826 ( .A0(n171), .A1(n149), .B0(n3318), .B1(n594), .C0(n2030), 
        .Y(n2468) );
  AOI222XLTS U2827 ( .A0(n3976), .A1(n3264), .B0(n4017), .B1(n3270), .C0(
        destinationAddressIn_SOUTH[10]), .C1(n3311), .Y(n2030) );
  OAI221XLTS U2828 ( .A0(n1805), .A1(n145), .B0(n3319), .B1(n593), .C0(n2029), 
        .Y(n2469) );
  AOI222XLTS U2829 ( .A0(n3973), .A1(n3265), .B0(n4015), .B1(n3271), .C0(
        destinationAddressIn_SOUTH[9]), .C1(n3311), .Y(n2029) );
  OAI221XLTS U2830 ( .A0(n170), .A1(n151), .B0(n3319), .B1(n592), .C0(n2028), 
        .Y(n2470) );
  AOI222XLTS U2831 ( .A0(n3970), .A1(n3262), .B0(destinationAddressIn_WEST[8]), 
        .B1(n3271), .C0(destinationAddressIn_SOUTH[8]), .C1(n3310), .Y(n2028)
         );
  OAI221XLTS U2832 ( .A0(n171), .A1(n136), .B0(n3319), .B1(n591), .C0(n2027), 
        .Y(n2471) );
  AOI222XLTS U2833 ( .A0(n3967), .A1(n3262), .B0(n4011), .B1(n3271), .C0(n4228), .C1(n3310), .Y(n2027) );
  OAI221XLTS U2834 ( .A0(n171), .A1(n139), .B0(n3319), .B1(n590), .C0(n2026), 
        .Y(n2472) );
  AOI222XLTS U2835 ( .A0(n3964), .A1(n3262), .B0(n4008), .B1(n3271), .C0(n4225), .C1(n3310), .Y(n2026) );
  OAI221XLTS U2836 ( .A0(n170), .A1(n141), .B0(n3318), .B1(n597), .C0(n2033), 
        .Y(n2465) );
  AOI222XLTS U2837 ( .A0(n3985), .A1(n3268), .B0(destinationAddressIn_WEST[13]), .B1(n3270), .C0(destinationAddressIn_SOUTH[13]), .C1(n3315), .Y(n2033) );
  OAI221XLTS U2838 ( .A0(n182), .A1(n142), .B0(n162), .B1(n565), .C0(n2009), 
        .Y(n2479) );
  AOI222XLTS U2839 ( .A0(n4247), .A1(n3367), .B0(n4022), .B1(n3352), .C0(n3985), .C1(n3395), .Y(n2009) );
  AOI222XLTS U2840 ( .A0(n4241), .A1(n3367), .B0(n4018), .B1(n3346), .C0(n3979), .C1(n3395), .Y(n2007) );
  AOI222XLTS U2841 ( .A0(n4235), .A1(n3368), .B0(n4015), .B1(n3346), .C0(n3973), .C1(n3396), .Y(n2005) );
  AOI222XLTS U2842 ( .A0(n4229), .A1(n3368), .B0(n4011), .B1(n3347), .C0(n3967), .C1(n3397), .Y(n2003) );
  AOI222XLTS U2843 ( .A0(n4244), .A1(n3367), .B0(n4020), .B1(n3346), .C0(n3982), .C1(n3395), .Y(n2008) );
  OAI221XLTS U2844 ( .A0(n183), .A1(n150), .B0(n1803), .B1(n554), .C0(n2006), 
        .Y(n2482) );
  AOI222XLTS U2845 ( .A0(n4238), .A1(n3367), .B0(n4017), .B1(n3346), .C0(n3976), .C1(n3396), .Y(n2006) );
  OAI221XLTS U2846 ( .A0(n1802), .A1(n152), .B0(n161), .B1(n553), .C0(n2004), 
        .Y(n2484) );
  AOI222XLTS U2847 ( .A0(n4232), .A1(n3368), .B0(n4012), .B1(n3347), .C0(n3970), .C1(n3396), .Y(n2004) );
  OAI221XLTS U2848 ( .A0(n1802), .A1(n140), .B0(n162), .B1(n552), .C0(n2002), 
        .Y(n2486) );
  AOI222XLTS U2849 ( .A0(n4226), .A1(n3368), .B0(n4008), .B1(n3349), .C0(n3964), .C1(n3397), .Y(n2002) );
  OAI221XLTS U2850 ( .A0(n167), .A1(n142), .B0(n3595), .B1(n910), .C0(n1940), 
        .Y(n2521) );
  OAI221XLTS U2851 ( .A0(n168), .A1(n148), .B0(n3595), .B1(n906), .C0(n1939), 
        .Y(n2522) );
  AOI222XLTS U2852 ( .A0(n4021), .A1(n3529), .B0(n3983), .B1(n3535), .C0(n4245), .C1(n3577), .Y(n1939) );
  OAI221XLTS U2853 ( .A0(n166), .A1(n144), .B0(n3595), .B1(n905), .C0(n1938), 
        .Y(n2523) );
  AOI222XLTS U2854 ( .A0(n4019), .A1(n3530), .B0(n3980), .B1(n3535), .C0(n4242), .C1(n3580), .Y(n1938) );
  OAI221XLTS U2855 ( .A0(n167), .A1(n146), .B0(n3583), .B1(n904), .C0(n1936), 
        .Y(n2525) );
  AOI222XLTS U2856 ( .A0(n4014), .A1(n3532), .B0(n3974), .B1(n3536), .C0(n4236), .C1(n3578), .Y(n1936) );
  OAI221XLTS U2857 ( .A0(n168), .A1(n151), .B0(n3583), .B1(n903), .C0(n1935), 
        .Y(n2526) );
  AOI222XLTS U2858 ( .A0(n4013), .A1(n3528), .B0(n3971), .B1(n3536), .C0(n4233), .C1(n3575), .Y(n1935) );
  OAI221XLTS U2859 ( .A0(n166), .A1(n137), .B0(n3583), .B1(n902), .C0(n1934), 
        .Y(n2527) );
  AOI222XLTS U2860 ( .A0(n4010), .A1(n3528), .B0(n3968), .B1(n3536), .C0(n4230), .C1(n3575), .Y(n1934) );
  OAI221XLTS U2861 ( .A0(n167), .A1(n139), .B0(n3583), .B1(n901), .C0(n1933), 
        .Y(n2528) );
  AOI222XLTS U2862 ( .A0(n4007), .A1(n3528), .B0(n3965), .B1(n3536), .C0(n4227), .C1(n3575), .Y(n1933) );
  OAI221XLTS U2863 ( .A0(n168), .A1(n149), .B0(n1182), .B1(n806), .C0(n1937), 
        .Y(n2524) );
  AOI222XLTS U2864 ( .A0(n4016), .A1(n3529), .B0(n3977), .B1(n3535), .C0(n4239), .C1(n3581), .Y(n1937) );
  OAI221XLTS U2865 ( .A0(n477), .A1(n150), .B0(n3123), .B1(n601), .C0(n1913), 
        .Y(n2538) );
  AOI222XLTS U2866 ( .A0(n4238), .A1(n3639), .B0(n4017), .B1(n3610), .C0(n3976), .C1(n3769), .Y(n1913) );
  OAI221XLTS U2867 ( .A0(n477), .A1(n145), .B0(n3123), .B1(n600), .C0(n1912), 
        .Y(n2539) );
  AOI222XLTS U2868 ( .A0(n4235), .A1(n3640), .B0(n4015), .B1(n3614), .C0(n3973), .C1(n3769), .Y(n1912) );
  OAI221XLTS U2869 ( .A0(n476), .A1(n152), .B0(n3123), .B1(n578), .C0(n1911), 
        .Y(n2540) );
  AOI222XLTS U2870 ( .A0(n4232), .A1(n3640), .B0(n4012), .B1(n3611), .C0(n3970), .C1(n3774), .Y(n1911) );
  OAI221XLTS U2871 ( .A0(n476), .A1(n136), .B0(n3123), .B1(n577), .C0(n1910), 
        .Y(n2541) );
  AOI222XLTS U2872 ( .A0(n4229), .A1(n3640), .B0(n4011), .B1(n3613), .C0(n3967), .C1(n3774), .Y(n1910) );
  OAI221XLTS U2873 ( .A0(n166), .A1(n159), .B0(n3584), .B1(n894), .C0(n1795), 
        .Y(n2576) );
  AOI222XLTS U2874 ( .A0(n4193), .A1(n3534), .B0(n4198), .B1(n3537), .C0(n4205), .C1(n3575), .Y(n1795) );
  OAI221XLTS U2875 ( .A0(n477), .A1(n140), .B0(n3124), .B1(n599), .C0(n1909), 
        .Y(n2542) );
  AOI222XLTS U2876 ( .A0(n4226), .A1(n3639), .B0(n4008), .B1(n3612), .C0(n3964), .C1(n3774), .Y(n1909) );
  OAI221XLTS U2877 ( .A0(n476), .A1(n147), .B0(n3122), .B1(n602), .C0(n1915), 
        .Y(n2536) );
  AOI222XLTS U2878 ( .A0(n4244), .A1(n3640), .B0(n4020), .B1(n3612), .C0(n3982), .C1(n3769), .Y(n1915) );
  OAI221XLTS U2879 ( .A0(n477), .A1(n142), .B0(n3122), .B1(n580), .C0(n1916), 
        .Y(n2535) );
  OAI221XLTS U2880 ( .A0(n476), .A1(n143), .B0(n3122), .B1(n579), .C0(n1914), 
        .Y(n2537) );
  AOI222XLTS U2881 ( .A0(n4241), .A1(n1169), .B0(n4018), .B1(n3611), .C0(n3979), .C1(n3769), .Y(n1914) );
  OAI221XLTS U2882 ( .A0(n3662), .A1(n160), .B0(n3743), .B1(n678), .C0(n1791), 
        .Y(n2578) );
  AOI222XLTS U2883 ( .A0(n4193), .A1(n3673), .B0(n4198), .B1(n3685), .C0(n4206), .C1(n3723), .Y(n1791) );
  OAI221XLTS U2884 ( .A0(n3661), .A1(n145), .B0(n3747), .B1(n598), .C0(n1884), 
        .Y(n2553) );
  AOI222XLTS U2885 ( .A0(n4014), .A1(n3672), .B0(n3974), .B1(n3684), .C0(n4236), .C1(n3724), .Y(n1884) );
  OAI221XLTS U2886 ( .A0(n3660), .A1(n143), .B0(n3745), .B1(n587), .C0(n1886), 
        .Y(n2551) );
  AOI222XLTS U2887 ( .A0(n4019), .A1(n3672), .B0(n3980), .B1(n3683), .C0(n4242), .C1(n3724), .Y(n1886) );
  OAI221XLTS U2888 ( .A0(n3661), .A1(n149), .B0(n1148), .B1(n586), .C0(n1885), 
        .Y(n2552) );
  AOI222XLTS U2889 ( .A0(n4016), .A1(n3672), .B0(n3977), .B1(n3683), .C0(n4239), .C1(n3724), .Y(n1885) );
  OAI221XLTS U2890 ( .A0(n3661), .A1(n151), .B0(n3745), .B1(n585), .C0(n1883), 
        .Y(n2554) );
  AOI222XLTS U2891 ( .A0(n4013), .A1(n3674), .B0(n3971), .B1(n3684), .C0(n4233), .C1(n3723), .Y(n1883) );
  OAI221XLTS U2892 ( .A0(n3662), .A1(n136), .B0(n3743), .B1(n584), .C0(n1882), 
        .Y(n2555) );
  AOI222XLTS U2893 ( .A0(n4010), .A1(n3674), .B0(n3968), .B1(n3684), .C0(n4230), .C1(n3723), .Y(n1882) );
  OAI221XLTS U2894 ( .A0(n3662), .A1(n139), .B0(n3746), .B1(n583), .C0(n1881), 
        .Y(n2556) );
  AOI222XLTS U2895 ( .A0(n4007), .A1(n3674), .B0(n3965), .B1(n3684), .C0(n4227), .C1(n3723), .Y(n1881) );
  OAI221XLTS U2896 ( .A0(n3660), .A1(n141), .B0(n3744), .B1(n589), .C0(n1888), 
        .Y(n2549) );
  AOI222XLTS U2897 ( .A0(n4023), .A1(n3680), .B0(n3986), .B1(n3683), .C0(n4248), .C1(n3726), .Y(n1888) );
  OAI221XLTS U2898 ( .A0(n3660), .A1(n148), .B0(n3744), .B1(n588), .C0(n1887), 
        .Y(n2550) );
  AOI222XLTS U2899 ( .A0(n4021), .A1(n3672), .B0(n3983), .B1(n3683), .C0(n4245), .C1(n3724), .Y(n1887) );
  AOI22X1TS U2900 ( .A0(n3254), .A1(n4189), .B0(n3901), .B1(n4076), .Y(n1261)
         );
  AOI222XLTS U2901 ( .A0(n3302), .A1(n4569), .B0(n3294), .B1(n39), .C0(n3273), 
        .C1(n4040), .Y(n1262) );
  AOI22X1TS U2902 ( .A0(n3253), .A1(n4186), .B0(n3898), .B1(n4073), .Y(n1259)
         );
  AOI222XLTS U2903 ( .A0(n3301), .A1(n4565), .B0(n3294), .B1(n34), .C0(n3273), 
        .C1(n4037), .Y(n1260) );
  AOI22X1TS U2904 ( .A0(n3253), .A1(n4183), .B0(n3901), .B1(n4070), .Y(n1257)
         );
  AOI222XLTS U2905 ( .A0(n3301), .A1(n4562), .B0(n3293), .B1(n29), .C0(n3272), 
        .C1(n4034), .Y(n1258) );
  AOI22X1TS U2906 ( .A0(n3253), .A1(n4180), .B0(n3902), .B1(n4067), .Y(n1255)
         );
  AOI222XLTS U2907 ( .A0(n3301), .A1(n4559), .B0(n3293), .B1(n24), .C0(n3272), 
        .C1(n4031), .Y(n1256) );
  AOI22X1TS U2908 ( .A0(n3253), .A1(n4177), .B0(n3903), .B1(n4064), .Y(n1253)
         );
  AOI222XLTS U2909 ( .A0(n3301), .A1(n4555), .B0(n3293), .B1(n19), .C0(n3272), 
        .C1(n4028), .Y(n1254) );
  AOI22X1TS U2910 ( .A0(n3254), .A1(n4174), .B0(n3902), .B1(n4061), .Y(n1247)
         );
  AOI222XLTS U2911 ( .A0(n3302), .A1(n4552), .B0(n3294), .B1(n14), .C0(n3273), 
        .C1(n4025), .Y(n1248) );
  AOI22X1TS U2912 ( .A0(n3519), .A1(n4039), .B0(n3799), .B1(n4076), .Y(n1197)
         );
  AOI222XLTS U2913 ( .A0(n3581), .A1(n4568), .B0(n3557), .B1(n40), .C0(n3538), 
        .C1(n4190), .Y(n1198) );
  AOI22X1TS U2914 ( .A0(n3518), .A1(n4036), .B0(n3797), .B1(n4073), .Y(n1195)
         );
  AOI222XLTS U2915 ( .A0(n3581), .A1(n4564), .B0(n3557), .B1(n35), .C0(n3538), 
        .C1(n4187), .Y(n1196) );
  AOI22X1TS U2916 ( .A0(n3518), .A1(n4033), .B0(n3790), .B1(n4070), .Y(n1193)
         );
  AOI222XLTS U2917 ( .A0(n3577), .A1(n4561), .B0(n3556), .B1(n30), .C0(n3537), 
        .C1(n4184), .Y(n1194) );
  AOI22X1TS U2918 ( .A0(n3518), .A1(n4030), .B0(n3790), .B1(n4067), .Y(n1191)
         );
  AOI222XLTS U2919 ( .A0(n3578), .A1(n4558), .B0(n3556), .B1(n25), .C0(n3537), 
        .C1(n4181), .Y(n1192) );
  AOI22X1TS U2920 ( .A0(n3518), .A1(n4027), .B0(n3790), .B1(n4064), .Y(n1189)
         );
  AOI222XLTS U2921 ( .A0(n3576), .A1(n4554), .B0(n3556), .B1(n20), .C0(n3537), 
        .C1(n4178), .Y(n1190) );
  AOI22X1TS U2922 ( .A0(n3519), .A1(n4024), .B0(n3790), .B1(n4061), .Y(n1183)
         );
  AOI222XLTS U2923 ( .A0(n3581), .A1(n4551), .B0(n3557), .B1(n15), .C0(n3538), 
        .C1(n4175), .Y(n1184) );
  AOI222XLTS U2924 ( .A0(n4219), .A1(n3309), .B0(n3295), .B1(n36), .C0(n4001), 
        .C1(n3286), .Y(n2022) );
  AOI22X1TS U2925 ( .A0(n3961), .A1(n3427), .B0(n4222), .B1(n3410), .Y(n1975)
         );
  AOI222XLTS U2926 ( .A0(n3855), .A1(n40), .B0(n4059), .B1(n3876), .C0(n61), 
        .C1(n3861), .Y(n1976) );
  AOI22X1TS U2927 ( .A0(n3958), .A1(n3427), .B0(n4219), .B1(n3410), .Y(n1973)
         );
  AOI222XLTS U2928 ( .A0(n3848), .A1(n35), .B0(n4056), .B1(n3876), .C0(n62), 
        .C1(n3871), .Y(n1974) );
  AOI22X1TS U2929 ( .A0(n3955), .A1(n3427), .B0(n4216), .B1(n3410), .Y(n1971)
         );
  AOI222XLTS U2930 ( .A0(n3848), .A1(n30), .B0(n4053), .B1(n3876), .C0(n63), 
        .C1(n3869), .Y(n1972) );
  AOI22X1TS U2931 ( .A0(n3949), .A1(n3426), .B0(n4210), .B1(n3414), .Y(n1967)
         );
  AOI222XLTS U2932 ( .A0(n3847), .A1(n20), .B0(n4047), .B1(n3877), .C0(n64), 
        .C1(n3870), .Y(n1968) );
  AOI22X1TS U2933 ( .A0(n3946), .A1(n3426), .B0(n4207), .B1(n3416), .Y(n1965)
         );
  AOI222XLTS U2934 ( .A0(n3848), .A1(n15), .B0(n4044), .B1(n3877), .C0(n65), 
        .C1(n790), .Y(n1966) );
  AOI22X1TS U2935 ( .A0(n3952), .A1(n3427), .B0(n4213), .B1(n3410), .Y(n1969)
         );
  AOI222XLTS U2936 ( .A0(n3848), .A1(n25), .B0(n4050), .B1(n3876), .C0(n90), 
        .C1(n790), .Y(n1970) );
  AOI22X1TS U2937 ( .A0(n3470), .A1(n30), .B0(n3453), .B1(n4183), .Y(n1209) );
  AOI222XLTS U2938 ( .A0(n2980), .A1(n189), .B0(n3500), .B1(n4562), .C0(n3804), 
        .C1(n4071), .Y(n1210) );
  AOI22X1TS U2939 ( .A0(n3470), .A1(n25), .B0(n3453), .B1(n4180), .Y(n1207) );
  AOI222XLTS U2940 ( .A0(n2978), .A1(n187), .B0(n3500), .B1(n4559), .C0(n3804), 
        .C1(n4068), .Y(n1208) );
  AOI22X1TS U2941 ( .A0(n3470), .A1(n20), .B0(n3453), .B1(n4177), .Y(n1205) );
  AOI222XLTS U2942 ( .A0(n2979), .A1(n190), .B0(n3500), .B1(n4555), .C0(n3804), 
        .C1(n4065), .Y(n1206) );
  AOI22X1TS U2943 ( .A0(n3471), .A1(n15), .B0(n3454), .B1(n4174), .Y(n1200) );
  AOI222XLTS U2944 ( .A0(n2981), .A1(n194), .B0(n3495), .B1(n4552), .C0(n3804), 
        .C1(n4062), .Y(n1201) );
  AOI22X1TS U2945 ( .A0(n3419), .A1(n4183), .B0(n3402), .B1(n4561), .Y(n1224)
         );
  AOI222XLTS U2946 ( .A0(n3858), .A1(n29), .B0(n3883), .B1(n4070), .C0(
        \requesterAddressbuffer[3][3] ), .C1(n3862), .Y(n1225) );
  AOI22X1TS U2947 ( .A0(n3419), .A1(n4180), .B0(n3402), .B1(n4558), .Y(n1222)
         );
  AOI222XLTS U2948 ( .A0(n3859), .A1(n24), .B0(n3883), .B1(n4067), .C0(
        \requesterAddressbuffer[3][2] ), .C1(n3861), .Y(n1223) );
  AOI22X1TS U2949 ( .A0(n3419), .A1(n4177), .B0(n3402), .B1(n4554), .Y(n1220)
         );
  AOI222XLTS U2950 ( .A0(n3859), .A1(n19), .B0(n3883), .B1(n4064), .C0(
        \requesterAddressbuffer[3][1] ), .C1(n3862), .Y(n1221) );
  AOI22X1TS U2951 ( .A0(n3420), .A1(n4174), .B0(n3403), .B1(n4551), .Y(n1216)
         );
  AOI222XLTS U2952 ( .A0(n3847), .A1(n14), .B0(n3883), .B1(n4061), .C0(
        \requesterAddressbuffer[3][0] ), .C1(n3866), .Y(n1217) );
  AOI222XLTS U2953 ( .A0(\requesterAddressbuffer[2][1] ), .A1(n3827), .B0(
        n3378), .B1(n4555), .C0(n3833), .C1(n4065), .Y(n1237) );
  AOI222XLTS U2954 ( .A0(\requesterAddressbuffer[2][0] ), .A1(n3825), .B0(
        n3382), .B1(n4552), .C0(n3833), .C1(n4062), .Y(n1232) );
  AOI222XLTS U2955 ( .A0(\requesterAddressbuffer[2][3] ), .A1(n3826), .B0(
        n3382), .B1(n4562), .C0(n3833), .C1(n4071), .Y(n1241) );
  AOI222XLTS U2956 ( .A0(\requesterAddressbuffer[2][2] ), .A1(n3826), .B0(
        n3379), .B1(n4559), .C0(n3833), .C1(n4068), .Y(n1239) );
  AOI22X1TS U2957 ( .A0(n3471), .A1(n40), .B0(n3454), .B1(n4189), .Y(n1213) );
  AOI222XLTS U2958 ( .A0(n2976), .A1(n193), .B0(n3493), .B1(n4569), .C0(n3805), 
        .C1(n4077), .Y(n1214) );
  AOI22X1TS U2959 ( .A0(n3471), .A1(n35), .B0(n3453), .B1(n4186), .Y(n1211) );
  AOI222XLTS U2960 ( .A0(n2977), .A1(n187), .B0(n3494), .B1(n4565), .C0(n3805), 
        .C1(n4074), .Y(n1212) );
  AOI22X1TS U2961 ( .A0(n3419), .A1(n4186), .B0(n3402), .B1(n4564), .Y(n1226)
         );
  AOI222XLTS U2962 ( .A0(n3847), .A1(n34), .B0(n3887), .B1(n4073), .C0(
        \requesterAddressbuffer[3][4] ), .C1(n3862), .Y(n1227) );
  AOI22X1TS U2963 ( .A0(n3420), .A1(n4189), .B0(n3403), .B1(n4568), .Y(n1228)
         );
  AOI222XLTS U2964 ( .A0(n3847), .A1(n39), .B0(n788), .B1(n4076), .C0(
        \requesterAddressbuffer[3][5] ), .C1(n3863), .Y(n1229) );
  AOI222XLTS U2965 ( .A0(\requesterAddressbuffer[2][4] ), .A1(n3826), .B0(
        n1233), .B1(n4565), .C0(n3834), .C1(n4074), .Y(n1243) );
  AOI222XLTS U2966 ( .A0(\requesterAddressbuffer[2][5] ), .A1(n3826), .B0(
        n3379), .B1(n4569), .C0(n3834), .C1(n4077), .Y(n1245) );
  AOI22X1TS U2967 ( .A0(n3158), .A1(n39), .B0(n3154), .B1(n4189), .Y(n1276) );
  AOI222XLTS U2968 ( .A0(\requesterAddressbuffer[0][5] ), .A1(n3912), .B0(
        n3245), .B1(n4040), .C0(n3933), .C1(n4077), .Y(n1277) );
  AOI22X1TS U2969 ( .A0(n3157), .A1(n29), .B0(n3155), .B1(n4183), .Y(n1272) );
  AOI222XLTS U2970 ( .A0(\requesterAddressbuffer[0][3] ), .A1(n3912), .B0(
        n3246), .B1(n4034), .C0(n3932), .C1(n4071), .Y(n1273) );
  AOI22X1TS U2971 ( .A0(n3158), .A1(n34), .B0(n3155), .B1(n4186), .Y(n1274) );
  AOI222XLTS U2972 ( .A0(\requesterAddressbuffer[0][4] ), .A1(n3916), .B0(
        n3250), .B1(n4037), .C0(n3933), .C1(n4074), .Y(n1275) );
  AOI22X1TS U2973 ( .A0(n3157), .A1(n24), .B0(n3155), .B1(n4180), .Y(n1270) );
  AOI222XLTS U2974 ( .A0(\requesterAddressbuffer[0][2] ), .A1(n3914), .B0(
        n3246), .B1(n4031), .C0(n3932), .C1(n4068), .Y(n1271) );
  AOI22X1TS U2975 ( .A0(n3157), .A1(n22), .B0(n3155), .B1(n4177), .Y(n1268) );
  AOI222XLTS U2976 ( .A0(\requesterAddressbuffer[0][1] ), .A1(n3908), .B0(
        n3246), .B1(n4028), .C0(n3932), .C1(n4065), .Y(n1269) );
  AOI22X1TS U2977 ( .A0(n3158), .A1(n14), .B0(n3154), .B1(n4174), .Y(n1263) );
  AOI222XLTS U2978 ( .A0(\requesterAddressbuffer[0][0] ), .A1(n3910), .B0(
        n3246), .B1(n4025), .C0(n3932), .C1(n4062), .Y(n1264) );
  AOI22X1TS U2979 ( .A0(n3157), .A1(n39), .B0(n3961), .B1(n3148), .Y(n2045) );
  AOI222XLTS U2980 ( .A0(n3917), .A1(n764), .B0(n4004), .B1(n3173), .C0(n4059), 
        .C1(n3939), .Y(n2046) );
  AOI22X1TS U2981 ( .A0(n3159), .A1(n29), .B0(n3955), .B1(n3148), .Y(n2041) );
  AOI222XLTS U2982 ( .A0(n3914), .A1(n763), .B0(n3998), .B1(n3245), .C0(n4053), 
        .C1(n3939), .Y(n2042) );
  AOI22X1TS U2983 ( .A0(n3159), .A1(n24), .B0(n3952), .B1(n3148), .Y(n2039) );
  AOI222XLTS U2984 ( .A0(n3913), .A1(n762), .B0(n3995), .B1(n3245), .C0(n4050), 
        .C1(n3939), .Y(n2040) );
  AOI22X1TS U2985 ( .A0(n3158), .A1(n19), .B0(n3949), .B1(n3147), .Y(n2037) );
  AOI222XLTS U2986 ( .A0(n3904), .A1(n761), .B0(n3992), .B1(n3244), .C0(n4047), 
        .C1(n3938), .Y(n2038) );
  AOI22X1TS U2987 ( .A0(n498), .A1(n3164), .B0(n4439), .B1(n3147), .Y(n1340)
         );
  AOI222XLTS U2988 ( .A0(n3904), .A1(n760), .B0(n4343), .B1(n3244), .C0(n4173), 
        .C1(n3938), .Y(n1341) );
  AOI22X1TS U2989 ( .A0(n500), .A1(n3160), .B0(n4436), .B1(n3147), .Y(n1338)
         );
  AOI222XLTS U2990 ( .A0(n3904), .A1(n759), .B0(n4340), .B1(n3244), .C0(n4170), 
        .C1(n3938), .Y(n1339) );
  AOI22X1TS U2991 ( .A0(n502), .A1(n3160), .B0(n4433), .B1(n3146), .Y(n1336)
         );
  AOI222XLTS U2992 ( .A0(n3905), .A1(n758), .B0(n4337), .B1(n3248), .C0(n4167), 
        .C1(n3941), .Y(n1337) );
  AOI22X1TS U2993 ( .A0(n508), .A1(n3168), .B0(n4423), .B1(n3146), .Y(n1330)
         );
  AOI222XLTS U2994 ( .A0(n3904), .A1(n757), .B0(n4328), .B1(n3251), .C0(n4158), 
        .C1(n3942), .Y(n1331) );
  AOI22X1TS U2995 ( .A0(n510), .A1(n3160), .B0(n4420), .B1(n3145), .Y(n1328)
         );
  AOI222XLTS U2996 ( .A0(n3906), .A1(n756), .B0(n4325), .B1(n3249), .C0(n4155), 
        .C1(n3945), .Y(n1329) );
  AOI22X1TS U2997 ( .A0(n512), .A1(n3161), .B0(n4417), .B1(n3145), .Y(n1326)
         );
  AOI222XLTS U2998 ( .A0(n3906), .A1(n755), .B0(n4322), .B1(n3252), .C0(n4152), 
        .C1(n783), .Y(n1327) );
  AOI22X1TS U2999 ( .A0(n516), .A1(n3161), .B0(n4411), .B1(n3145), .Y(n1322)
         );
  AOI222XLTS U3000 ( .A0(n3906), .A1(n754), .B0(n4316), .B1(n3252), .C0(n4146), 
        .C1(n3941), .Y(n1323) );
  AOI22X1TS U3001 ( .A0(n518), .A1(n3166), .B0(n4408), .B1(n3144), .Y(n1320)
         );
  AOI222XLTS U3002 ( .A0(n3907), .A1(n753), .B0(n4313), .B1(n3243), .C0(n4143), 
        .C1(n3937), .Y(n1321) );
  AOI22X1TS U3003 ( .A0(n522), .A1(n1266), .B0(n4402), .B1(n3144), .Y(n1316)
         );
  AOI222XLTS U3004 ( .A0(n46), .A1(n163), .B0(n4307), .B1(n3243), .C0(n4137), 
        .C1(n3937), .Y(n1317) );
  AOI22X1TS U3005 ( .A0(n524), .A1(n3169), .B0(n4399), .B1(n3143), .Y(n1314)
         );
  AOI222XLTS U3006 ( .A0(n47), .A1(n163), .B0(n4304), .B1(n3242), .C0(n4134), 
        .C1(n3937), .Y(n1315) );
  AOI22X1TS U3007 ( .A0(n526), .A1(n3165), .B0(n4396), .B1(n3143), .Y(n1312)
         );
  AOI222XLTS U3008 ( .A0(n48), .A1(n3913), .B0(n4301), .B1(n3242), .C0(n4131), 
        .C1(n3943), .Y(n1313) );
  AOI22X1TS U3009 ( .A0(n528), .A1(n3166), .B0(n4393), .B1(n3143), .Y(n1310)
         );
  AOI222XLTS U3010 ( .A0(n49), .A1(n3915), .B0(n4298), .B1(n3242), .C0(n4128), 
        .C1(n3945), .Y(n1311) );
  AOI22X1TS U3011 ( .A0(n530), .A1(n3168), .B0(n4390), .B1(n3143), .Y(n1308)
         );
  AOI222XLTS U3012 ( .A0(n50), .A1(n3911), .B0(n4295), .B1(n3242), .C0(n4125), 
        .C1(n783), .Y(n1309) );
  AOI22X1TS U3013 ( .A0(n532), .A1(n3170), .B0(n4387), .B1(n3142), .Y(n1306)
         );
  AOI222XLTS U3014 ( .A0(n51), .A1(n3911), .B0(n4292), .B1(n3241), .C0(n4122), 
        .C1(n3945), .Y(n1307) );
  AOI22X1TS U3015 ( .A0(n534), .A1(n3167), .B0(n4384), .B1(n3142), .Y(n1304)
         );
  AOI222XLTS U3016 ( .A0(n52), .A1(n3911), .B0(n4289), .B1(n3241), .C0(n4119), 
        .C1(n3936), .Y(n1305) );
  AOI22X1TS U3017 ( .A0(n536), .A1(n3167), .B0(n4381), .B1(n3142), .Y(n1302)
         );
  AOI222XLTS U3018 ( .A0(n53), .A1(n3911), .B0(n4286), .B1(n3241), .C0(n4116), 
        .C1(n3936), .Y(n1303) );
  AOI22X1TS U3019 ( .A0(n538), .A1(n3168), .B0(n4378), .B1(n3142), .Y(n1300)
         );
  AOI222XLTS U3020 ( .A0(n54), .A1(n3910), .B0(n4283), .B1(n3241), .C0(n4113), 
        .C1(n3936), .Y(n1301) );
  AOI22X1TS U3021 ( .A0(n540), .A1(n3164), .B0(n4375), .B1(n3141), .Y(n1298)
         );
  AOI222XLTS U3022 ( .A0(n55), .A1(n3910), .B0(n4280), .B1(n3175), .C0(n4110), 
        .C1(n3936), .Y(n1299) );
  AOI22X1TS U3023 ( .A0(n544), .A1(n3162), .B0(n4369), .B1(n3141), .Y(n1294)
         );
  AOI222XLTS U3024 ( .A0(n56), .A1(n3910), .B0(n4274), .B1(n3175), .C0(n4104), 
        .C1(n3935), .Y(n1295) );
  AOI22X1TS U3025 ( .A0(n496), .A1(n3162), .B0(n4366), .B1(n3141), .Y(n1292)
         );
  AOI222XLTS U3026 ( .A0(n57), .A1(n3909), .B0(n4271), .B1(n3175), .C0(n4101), 
        .C1(n3935), .Y(n1293) );
  AOI22X1TS U3027 ( .A0(n546), .A1(n3163), .B0(n4363), .B1(n3141), .Y(n1290)
         );
  AOI222XLTS U3028 ( .A0(n58), .A1(n3909), .B0(n4268), .B1(n3243), .C0(n4098), 
        .C1(n3935), .Y(n1291) );
  AOI22X1TS U3029 ( .A0(n550), .A1(n3163), .B0(n4357), .B1(n3140), .Y(n1286)
         );
  AOI222XLTS U3030 ( .A0(n59), .A1(n3909), .B0(n4262), .B1(n3174), .C0(n4092), 
        .C1(n3934), .Y(n1287) );
  AOI22X1TS U3031 ( .A0(n780), .A1(n3164), .B0(n4354), .B1(n3140), .Y(n1284)
         );
  AOI222XLTS U3032 ( .A0(n60), .A1(n3909), .B0(n4259), .B1(n3174), .C0(n4089), 
        .C1(n3934), .Y(n1285) );
  AOI22X1TS U3033 ( .A0(n3159), .A1(n35), .B0(n3958), .B1(n3148), .Y(n2043) );
  AOI222XLTS U3034 ( .A0(n88), .A1(n3908), .B0(n4001), .B1(n3245), .C0(n4056), 
        .C1(n3939), .Y(n2044) );
  AOI22X1TS U3035 ( .A0(n3159), .A1(n15), .B0(n3946), .B1(n3147), .Y(n2035) );
  AOI222XLTS U3036 ( .A0(n89), .A1(n3912), .B0(n3989), .B1(n3244), .C0(n4044), 
        .C1(n3938), .Y(n2036) );
  AOI22X1TS U3037 ( .A0(n504), .A1(n3160), .B0(n4429), .B1(n3146), .Y(n1334)
         );
  AOI222XLTS U3038 ( .A0(n3905), .A1(n706), .B0(n4334), .B1(n3249), .C0(n4164), 
        .C1(n3940), .Y(n1335) );
  AOI22X1TS U3039 ( .A0(n506), .A1(n3161), .B0(n4426), .B1(n3146), .Y(n1332)
         );
  AOI222XLTS U3040 ( .A0(n3905), .A1(n705), .B0(n4331), .B1(n3247), .C0(n4161), 
        .C1(n3940), .Y(n1333) );
  AOI22X1TS U3041 ( .A0(n514), .A1(n3161), .B0(n4414), .B1(n3145), .Y(n1324)
         );
  AOI222XLTS U3042 ( .A0(n3906), .A1(n704), .B0(n4319), .B1(n3248), .C0(n4149), 
        .C1(n3942), .Y(n1325) );
  AOI22X1TS U3043 ( .A0(n520), .A1(n3170), .B0(n4405), .B1(n3144), .Y(n1318)
         );
  AOI222XLTS U3044 ( .A0(n3905), .A1(n703), .B0(n4310), .B1(n3243), .C0(n4140), 
        .C1(n3937), .Y(n1319) );
  AOI22X1TS U3045 ( .A0(n542), .A1(n3162), .B0(n4372), .B1(n3144), .Y(n1296)
         );
  AOI222XLTS U3046 ( .A0(n3908), .A1(n702), .B0(n4277), .B1(n3175), .C0(n4107), 
        .C1(n3935), .Y(n1297) );
  AOI22X1TS U3047 ( .A0(n548), .A1(n3162), .B0(n4360), .B1(n3140), .Y(n1288)
         );
  AOI222XLTS U3048 ( .A0(n3908), .A1(n701), .B0(n4265), .B1(n3174), .C0(n4095), 
        .C1(n3934), .Y(n1289) );
  AOI22X1TS U3049 ( .A0(n787), .A1(n3163), .B0(n4351), .B1(n3140), .Y(n1282)
         );
  AOI222XLTS U3050 ( .A0(n3907), .A1(n700), .B0(n4256), .B1(n3174), .C0(n4086), 
        .C1(n3934), .Y(n1283) );
  AOI22X1TS U3051 ( .A0(n792), .A1(n3163), .B0(n4348), .B1(n3153), .Y(n1280)
         );
  AOI222XLTS U3052 ( .A0(n3907), .A1(n699), .B0(n4253), .B1(n3173), .C0(n4083), 
        .C1(n3933), .Y(n1281) );
  AOI22X1TS U3053 ( .A0(n795), .A1(n3164), .B0(n4345), .B1(n3153), .Y(n1278)
         );
  AOI222XLTS U3054 ( .A0(n3907), .A1(n698), .B0(n4250), .B1(n3173), .C0(n4080), 
        .C1(n3933), .Y(n1279) );
  AOI22X1TS U3055 ( .A0(n4039), .A1(n3667), .B0(n4076), .B1(n3658), .Y(n1164)
         );
  AOI222XLTS U3056 ( .A0(n4568), .A1(n3715), .B0(n41), .B1(n3707), .C0(n4190), 
        .C1(n3686), .Y(n1165) );
  AOI22X1TS U3057 ( .A0(n4036), .A1(n3666), .B0(n4073), .B1(n3658), .Y(n1162)
         );
  AOI222XLTS U3058 ( .A0(n4564), .A1(n3714), .B0(n36), .B1(n3707), .C0(n4187), 
        .C1(n3686), .Y(n1163) );
  AOI22X1TS U3059 ( .A0(n4030), .A1(n3666), .B0(n4067), .B1(n3659), .Y(n1158)
         );
  AOI222XLTS U3060 ( .A0(n4558), .A1(n3714), .B0(n26), .B1(n3708), .C0(n4181), 
        .C1(n3686), .Y(n1159) );
  AOI22X1TS U3061 ( .A0(n4033), .A1(n3666), .B0(n4070), .B1(n3659), .Y(n1160)
         );
  AOI222XLTS U3062 ( .A0(n4561), .A1(n3714), .B0(n31), .B1(n3708), .C0(n4184), 
        .C1(n3685), .Y(n1161) );
  AOI22X1TS U3063 ( .A0(n4027), .A1(n3666), .B0(n4064), .B1(n3659), .Y(n1156)
         );
  AOI222XLTS U3064 ( .A0(n4554), .A1(n3714), .B0(n21), .B1(n3708), .C0(n4178), 
        .C1(n3685), .Y(n1157) );
  AOI22X1TS U3065 ( .A0(n4024), .A1(n3676), .B0(n4061), .B1(n3659), .Y(n1149)
         );
  AOI222XLTS U3066 ( .A0(n4551), .A1(n3720), .B0(n16), .B1(n3708), .C0(n4175), 
        .C1(n3690), .Y(n1150) );
  AOI22X1TS U3067 ( .A0(n4000), .A1(n3681), .B0(n4055), .B1(n3649), .Y(n1875)
         );
  AOI222XLTS U3068 ( .A0(n4219), .A1(n3722), .B0(n37), .B1(n1152), .C0(n3959), 
        .C1(n3699), .Y(n1876) );
  AOI22X1TS U3069 ( .A0(n3988), .A1(n3675), .B0(n4043), .B1(n3650), .Y(n1867)
         );
  AOI222XLTS U3070 ( .A0(n4207), .A1(n3725), .B0(n17), .B1(n3700), .C0(n3947), 
        .C1(n3693), .Y(n1868) );
  AOI22X1TS U3071 ( .A0(n4003), .A1(n1154), .B0(n4058), .B1(n3649), .Y(n1877)
         );
  AOI222XLTS U3072 ( .A0(n4222), .A1(n3722), .B0(n42), .B1(n1152), .C0(n3962), 
        .C1(n3685), .Y(n1878) );
  AOI22X1TS U3073 ( .A0(n3997), .A1(n3682), .B0(n4052), .B1(n3649), .Y(n1873)
         );
  AOI222XLTS U3074 ( .A0(n4216), .A1(n3722), .B0(n32), .B1(n3709), .C0(n3956), 
        .C1(n3693), .Y(n1874) );
  AOI22X1TS U3075 ( .A0(n3994), .A1(n3674), .B0(n4049), .B1(n3649), .Y(n1871)
         );
  AOI222XLTS U3076 ( .A0(n4213), .A1(n3722), .B0(n27), .B1(n3711), .C0(n3953), 
        .C1(n3693), .Y(n1872) );
  AOI22X1TS U3077 ( .A0(n3991), .A1(n3678), .B0(n4046), .B1(n3650), .Y(n1869)
         );
  AOI222XLTS U3078 ( .A0(n4210), .A1(n3727), .B0(n22), .B1(n3700), .C0(n3950), 
        .C1(n3693), .Y(n1870) );
  AOI22X1TS U3079 ( .A0(n4342), .A1(n3682), .B0(n4172), .B1(n3650), .Y(n1789)
         );
  AOI222XLTS U3080 ( .A0(n4549), .A1(n3726), .B0(n497), .B1(n3700), .C0(n4441), 
        .C1(n1153), .Y(n1790) );
  AOI22X1TS U3081 ( .A0(n4339), .A1(n3682), .B0(n4169), .B1(n3650), .Y(n1787)
         );
  AOI222XLTS U3082 ( .A0(n4545), .A1(n1151), .B0(n499), .B1(n3700), .C0(n4437), 
        .C1(n3695), .Y(n1788) );
  AOI22X1TS U3083 ( .A0(n4336), .A1(n3679), .B0(n4166), .B1(n3651), .Y(n1785)
         );
  AOI222XLTS U3084 ( .A0(n4542), .A1(n1151), .B0(n501), .B1(n3701), .C0(n4434), 
        .C1(n3697), .Y(n1786) );
  AOI22X1TS U3085 ( .A0(n4333), .A1(n3679), .B0(n4163), .B1(n3651), .Y(n1783)
         );
  AOI222XLTS U3086 ( .A0(n4538), .A1(n3730), .B0(n503), .B1(n3701), .C0(n4430), 
        .C1(n3698), .Y(n1784) );
  AOI22X1TS U3087 ( .A0(n4330), .A1(n3675), .B0(n4160), .B1(n3651), .Y(n1781)
         );
  AOI222XLTS U3088 ( .A0(n4535), .A1(n3730), .B0(n505), .B1(n3701), .C0(n4427), 
        .C1(n3695), .Y(n1782) );
  AOI22X1TS U3089 ( .A0(n4327), .A1(n3677), .B0(n4157), .B1(n3651), .Y(n1779)
         );
  AOI222XLTS U3090 ( .A0(n4532), .A1(n3728), .B0(n507), .B1(n3701), .C0(n4424), 
        .C1(n3696), .Y(n1780) );
  AOI22X1TS U3091 ( .A0(n4324), .A1(n3676), .B0(n4154), .B1(n3652), .Y(n1777)
         );
  AOI222XLTS U3092 ( .A0(n4528), .A1(n3721), .B0(n509), .B1(n3702), .C0(n4421), 
        .C1(n3697), .Y(n1778) );
  AOI22X1TS U3093 ( .A0(n4321), .A1(n3676), .B0(n4151), .B1(n3652), .Y(n1775)
         );
  AOI222XLTS U3094 ( .A0(n4525), .A1(n3721), .B0(n511), .B1(n3702), .C0(n4418), 
        .C1(n3696), .Y(n1776) );
  AOI22X1TS U3095 ( .A0(n4318), .A1(n3677), .B0(n4148), .B1(n3652), .Y(n1773)
         );
  AOI222XLTS U3096 ( .A0(n4522), .A1(n3721), .B0(n513), .B1(n3702), .C0(n4415), 
        .C1(n3692), .Y(n1774) );
  AOI22X1TS U3097 ( .A0(n4315), .A1(n3678), .B0(n4145), .B1(n3652), .Y(n1771)
         );
  AOI222XLTS U3098 ( .A0(n4518), .A1(n3721), .B0(n515), .B1(n3702), .C0(n4412), 
        .C1(n3692), .Y(n1772) );
  AOI22X1TS U3099 ( .A0(n4312), .A1(n3675), .B0(n4142), .B1(n3653), .Y(n1769)
         );
  AOI222XLTS U3100 ( .A0(n4515), .A1(n3720), .B0(n517), .B1(n3711), .C0(n4409), 
        .C1(n3692), .Y(n1770) );
  AOI22X1TS U3101 ( .A0(n4309), .A1(n3676), .B0(n4139), .B1(n3653), .Y(n1767)
         );
  AOI222XLTS U3102 ( .A0(n4511), .A1(n3720), .B0(n519), .B1(n3712), .C0(n4406), 
        .C1(n3692), .Y(n1768) );
  AOI22X1TS U3103 ( .A0(n4306), .A1(n3675), .B0(n4136), .B1(n3653), .Y(n1765)
         );
  AOI222XLTS U3104 ( .A0(n4508), .A1(n3720), .B0(n521), .B1(n3710), .C0(n4403), 
        .C1(n3691), .Y(n1766) );
  AOI22X1TS U3105 ( .A0(n4303), .A1(n3671), .B0(n4133), .B1(n3653), .Y(n1763)
         );
  AOI222XLTS U3106 ( .A0(n4505), .A1(n3719), .B0(n523), .B1(n3712), .C0(n4400), 
        .C1(n3691), .Y(n1764) );
  AOI22X1TS U3107 ( .A0(n4300), .A1(n3671), .B0(n4130), .B1(n3654), .Y(n1761)
         );
  AOI222XLTS U3108 ( .A0(n4501), .A1(n3719), .B0(n525), .B1(n3703), .C0(n4397), 
        .C1(n3691), .Y(n1762) );
  AOI22X1TS U3109 ( .A0(n4297), .A1(n3671), .B0(n4127), .B1(n3654), .Y(n1759)
         );
  AOI222XLTS U3110 ( .A0(n4498), .A1(n3719), .B0(n527), .B1(n3703), .C0(n4394), 
        .C1(n3691), .Y(n1760) );
  AOI22X1TS U3111 ( .A0(n4294), .A1(n3671), .B0(n4124), .B1(n3654), .Y(n1757)
         );
  AOI222XLTS U3112 ( .A0(n4495), .A1(n3719), .B0(n529), .B1(n3703), .C0(n4391), 
        .C1(n3690), .Y(n1758) );
  AOI22X1TS U3113 ( .A0(n4291), .A1(n3670), .B0(n4121), .B1(n3654), .Y(n1755)
         );
  AOI222XLTS U3114 ( .A0(n4491), .A1(n3718), .B0(n531), .B1(n3703), .C0(n4388), 
        .C1(n3690), .Y(n1756) );
  AOI22X1TS U3115 ( .A0(n4288), .A1(n3670), .B0(n4118), .B1(n3655), .Y(n1753)
         );
  AOI222XLTS U3116 ( .A0(n4488), .A1(n3718), .B0(n533), .B1(n3704), .C0(n4385), 
        .C1(n3690), .Y(n1754) );
  AOI22X1TS U3117 ( .A0(n4285), .A1(n3670), .B0(n4115), .B1(n3655), .Y(n1751)
         );
  AOI222XLTS U3118 ( .A0(n4484), .A1(n3718), .B0(n535), .B1(n3704), .C0(n4382), 
        .C1(n3689), .Y(n1752) );
  AOI22X1TS U3119 ( .A0(n4282), .A1(n3670), .B0(n4112), .B1(n3655), .Y(n1749)
         );
  AOI222XLTS U3120 ( .A0(n4481), .A1(n3718), .B0(n537), .B1(n3704), .C0(n4379), 
        .C1(n3689), .Y(n1750) );
  AOI22X1TS U3121 ( .A0(n4279), .A1(n3669), .B0(n4109), .B1(n3655), .Y(n1747)
         );
  AOI222XLTS U3122 ( .A0(n4478), .A1(n3717), .B0(n539), .B1(n3704), .C0(n4376), 
        .C1(n3689), .Y(n1748) );
  AOI22X1TS U3123 ( .A0(n4276), .A1(n3669), .B0(n4106), .B1(n3656), .Y(n1745)
         );
  AOI222XLTS U3124 ( .A0(n4474), .A1(n3717), .B0(n541), .B1(n3705), .C0(n4373), 
        .C1(n3689), .Y(n1746) );
  AOI22X1TS U3125 ( .A0(n4273), .A1(n3669), .B0(n4103), .B1(n3656), .Y(n1743)
         );
  AOI222XLTS U3126 ( .A0(n4471), .A1(n3717), .B0(n543), .B1(n3705), .C0(n4370), 
        .C1(n3688), .Y(n1744) );
  AOI22X1TS U3127 ( .A0(n4270), .A1(n3669), .B0(n4100), .B1(n3656), .Y(n1741)
         );
  AOI222XLTS U3128 ( .A0(n4468), .A1(n3717), .B0(n495), .B1(n3705), .C0(n4367), 
        .C1(n3688), .Y(n1742) );
  AOI22X1TS U3129 ( .A0(n4267), .A1(n3668), .B0(n4097), .B1(n3656), .Y(n1739)
         );
  AOI222XLTS U3130 ( .A0(n4464), .A1(n3716), .B0(n545), .B1(n3705), .C0(n4364), 
        .C1(n3688), .Y(n1740) );
  AOI22X1TS U3131 ( .A0(n4264), .A1(n3668), .B0(n4094), .B1(n3657), .Y(n1737)
         );
  AOI222XLTS U3132 ( .A0(n4461), .A1(n3716), .B0(n547), .B1(n3706), .C0(n4361), 
        .C1(n3688), .Y(n1738) );
  AOI22X1TS U3133 ( .A0(n4261), .A1(n3668), .B0(n4091), .B1(n3657), .Y(n1735)
         );
  AOI222XLTS U3134 ( .A0(n4457), .A1(n3716), .B0(n549), .B1(n3706), .C0(n4358), 
        .C1(n3687), .Y(n1736) );
  AOI22X1TS U3135 ( .A0(n4258), .A1(n3668), .B0(n4088), .B1(n3657), .Y(n1733)
         );
  AOI222XLTS U3136 ( .A0(n4454), .A1(n3716), .B0(n551), .B1(n3706), .C0(n4355), 
        .C1(n3687), .Y(n1734) );
  AOI22X1TS U3137 ( .A0(n4255), .A1(n3667), .B0(n4085), .B1(n3657), .Y(n1731)
         );
  AOI222XLTS U3138 ( .A0(n4451), .A1(n3715), .B0(n786), .B1(n3706), .C0(n4352), 
        .C1(n3687), .Y(n1732) );
  AOI22X1TS U3139 ( .A0(n4252), .A1(n3667), .B0(n4082), .B1(n3658), .Y(n1729)
         );
  AOI222XLTS U3140 ( .A0(n4447), .A1(n3715), .B0(n789), .B1(n3707), .C0(n4349), 
        .C1(n3687), .Y(n1730) );
  AOI22X1TS U3141 ( .A0(n4249), .A1(n3667), .B0(n4079), .B1(n3658), .Y(n1727)
         );
  AOI222XLTS U3142 ( .A0(n4444), .A1(n3715), .B0(n793), .B1(n3707), .C0(n4346), 
        .C1(n3686), .Y(n1728) );
  AOI22X1TS U3143 ( .A0(n4003), .A1(n3528), .B0(n4058), .B1(n3796), .Y(n1930)
         );
  AOI222XLTS U3144 ( .A0(n4222), .A1(n3574), .B0(n3556), .B1(n41), .C0(n3962), 
        .C1(n3538), .Y(n1931) );
  AOI22X1TS U3145 ( .A0(n4342), .A1(n3527), .B0(n4172), .B1(n3795), .Y(n1660)
         );
  AOI222XLTS U3146 ( .A0(n4547), .A1(n3573), .B0(n498), .B1(n3552), .C0(n4441), 
        .C1(n3543), .Y(n1661) );
  AOI22X1TS U3147 ( .A0(n4297), .A1(n3523), .B0(n4127), .B1(n3792), .Y(n1630)
         );
  AOI222XLTS U3148 ( .A0(n4497), .A1(n3569), .B0(n528), .B1(n3559), .C0(n4394), 
        .C1(n3547), .Y(n1631) );
  AOI22X1TS U3149 ( .A0(n4294), .A1(n3523), .B0(n4124), .B1(n3792), .Y(n1628)
         );
  AOI222XLTS U3150 ( .A0(n4493), .A1(n3569), .B0(n530), .B1(n3562), .C0(n4391), 
        .C1(n3542), .Y(n1629) );
  AOI22X1TS U3151 ( .A0(n4282), .A1(n3522), .B0(n4112), .B1(n3801), .Y(n1620)
         );
  AOI222XLTS U3152 ( .A0(n4480), .A1(n3568), .B0(n538), .B1(n3554), .C0(n4379), 
        .C1(n3541), .Y(n1621) );
  AOI22X1TS U3153 ( .A0(n4252), .A1(n3519), .B0(n4082), .B1(n3800), .Y(n1600)
         );
  AOI222XLTS U3154 ( .A0(n4446), .A1(n3579), .B0(n792), .B1(n3555), .C0(n4349), 
        .C1(n3539), .Y(n1601) );
  AOI22X1TS U3155 ( .A0(n3997), .A1(n3532), .B0(n4052), .B1(n3796), .Y(n1926)
         );
  AOI222XLTS U3156 ( .A0(n4216), .A1(n3574), .B0(n3558), .B1(n31), .C0(n3956), 
        .C1(n3544), .Y(n1927) );
  AOI22X1TS U3157 ( .A0(n3994), .A1(n3530), .B0(n4049), .B1(n3796), .Y(n1924)
         );
  AOI222XLTS U3158 ( .A0(n4213), .A1(n3574), .B0(n3558), .B1(n26), .C0(n3953), 
        .C1(n3544), .Y(n1925) );
  AOI22X1TS U3159 ( .A0(n3991), .A1(n3527), .B0(n4046), .B1(n3795), .Y(n1922)
         );
  AOI222XLTS U3160 ( .A0(n4210), .A1(n3573), .B0(n3558), .B1(n21), .C0(n3950), 
        .C1(n3544), .Y(n1923) );
  AOI22X1TS U3161 ( .A0(n3988), .A1(n3527), .B0(n4043), .B1(n3795), .Y(n1920)
         );
  AOI222XLTS U3162 ( .A0(n4207), .A1(n3573), .B0(n3557), .B1(n16), .C0(n3947), 
        .C1(n3544), .Y(n1921) );
  AOI22X1TS U3163 ( .A0(n4339), .A1(n3527), .B0(n4169), .B1(n3795), .Y(n1658)
         );
  AOI222XLTS U3164 ( .A0(n4544), .A1(n3573), .B0(n500), .B1(n3559), .C0(n4437), 
        .C1(n3543), .Y(n1659) );
  AOI22X1TS U3165 ( .A0(n4336), .A1(n3526), .B0(n4166), .B1(n3794), .Y(n1656)
         );
  AOI222XLTS U3166 ( .A0(n4541), .A1(n3572), .B0(n502), .B1(n3552), .C0(n4434), 
        .C1(n3543), .Y(n1657) );
  AOI22X1TS U3167 ( .A0(n4333), .A1(n3526), .B0(n4163), .B1(n3794), .Y(n1654)
         );
  AOI222XLTS U3168 ( .A0(n4537), .A1(n3572), .B0(n504), .B1(n3564), .C0(n4430), 
        .C1(n3543), .Y(n1655) );
  AOI22X1TS U3169 ( .A0(n4330), .A1(n3526), .B0(n4160), .B1(n3794), .Y(n1652)
         );
  AOI222XLTS U3170 ( .A0(n4534), .A1(n3572), .B0(n506), .B1(n3564), .C0(n4427), 
        .C1(n3545), .Y(n1653) );
  AOI22X1TS U3171 ( .A0(n4327), .A1(n3526), .B0(n4157), .B1(n3794), .Y(n1650)
         );
  AOI222XLTS U3172 ( .A0(n4531), .A1(n3572), .B0(n508), .B1(n3563), .C0(n4424), 
        .C1(n3545), .Y(n1651) );
  AOI22X1TS U3173 ( .A0(n4324), .A1(n3525), .B0(n4154), .B1(n3798), .Y(n1648)
         );
  AOI222XLTS U3174 ( .A0(n4527), .A1(n3571), .B0(n510), .B1(n3563), .C0(n4421), 
        .C1(n3547), .Y(n1649) );
  AOI22X1TS U3175 ( .A0(n4321), .A1(n3525), .B0(n4151), .B1(n3798), .Y(n1646)
         );
  AOI222XLTS U3176 ( .A0(n4524), .A1(n3571), .B0(n512), .B1(n3552), .C0(n4418), 
        .C1(n3545), .Y(n1647) );
  AOI22X1TS U3177 ( .A0(n4318), .A1(n3525), .B0(n4148), .B1(n3799), .Y(n1644)
         );
  AOI222XLTS U3178 ( .A0(n4520), .A1(n3571), .B0(n514), .B1(n3562), .C0(n4415), 
        .C1(n3546), .Y(n1645) );
  AOI22X1TS U3179 ( .A0(n4315), .A1(n3525), .B0(n4145), .B1(n3797), .Y(n1642)
         );
  AOI222XLTS U3180 ( .A0(n4517), .A1(n3571), .B0(n516), .B1(n3562), .C0(n4412), 
        .C1(n3550), .Y(n1643) );
  AOI22X1TS U3181 ( .A0(n4312), .A1(n3524), .B0(n4142), .B1(n3793), .Y(n1640)
         );
  AOI222XLTS U3182 ( .A0(n4514), .A1(n3570), .B0(n518), .B1(n3552), .C0(n4409), 
        .C1(n3548), .Y(n1641) );
  AOI22X1TS U3183 ( .A0(n4309), .A1(n3524), .B0(n4139), .B1(n3793), .Y(n1638)
         );
  AOI222XLTS U3184 ( .A0(n4510), .A1(n3570), .B0(n520), .B1(n3563), .C0(n4406), 
        .C1(n3550), .Y(n1639) );
  AOI22X1TS U3185 ( .A0(n4306), .A1(n3524), .B0(n4136), .B1(n3793), .Y(n1636)
         );
  AOI222XLTS U3186 ( .A0(n4507), .A1(n3570), .B0(n522), .B1(n3561), .C0(n4403), 
        .C1(n3546), .Y(n1637) );
  AOI22X1TS U3187 ( .A0(n4303), .A1(n3523), .B0(n4133), .B1(n3793), .Y(n1634)
         );
  AOI222XLTS U3188 ( .A0(n4504), .A1(n3569), .B0(n524), .B1(n3561), .C0(n4400), 
        .C1(n3548), .Y(n1635) );
  AOI22X1TS U3189 ( .A0(n4300), .A1(n3523), .B0(n4130), .B1(n3792), .Y(n1632)
         );
  AOI222XLTS U3190 ( .A0(n4500), .A1(n3569), .B0(n526), .B1(n3560), .C0(n4397), 
        .C1(n3550), .Y(n1633) );
  AOI22X1TS U3191 ( .A0(n4291), .A1(n3522), .B0(n4121), .B1(n3792), .Y(n1626)
         );
  AOI222XLTS U3192 ( .A0(n4490), .A1(n3568), .B0(n532), .B1(n3560), .C0(n4388), 
        .C1(n3542), .Y(n1627) );
  AOI22X1TS U3193 ( .A0(n4288), .A1(n3522), .B0(n4118), .B1(n3800), .Y(n1624)
         );
  AOI222XLTS U3194 ( .A0(n4487), .A1(n3568), .B0(n534), .B1(n3553), .C0(n4385), 
        .C1(n3542), .Y(n1625) );
  AOI22X1TS U3195 ( .A0(n4285), .A1(n3522), .B0(n4115), .B1(n3801), .Y(n1622)
         );
  AOI222XLTS U3196 ( .A0(n4483), .A1(n3568), .B0(n536), .B1(n3562), .C0(n4382), 
        .C1(n3541), .Y(n1623) );
  AOI22X1TS U3197 ( .A0(n4279), .A1(n3521), .B0(n4109), .B1(n5), .Y(n1618) );
  AOI222XLTS U3198 ( .A0(n4477), .A1(n3567), .B0(n540), .B1(n3554), .C0(n4376), 
        .C1(n3541), .Y(n1619) );
  AOI22X1TS U3199 ( .A0(n4276), .A1(n3524), .B0(n4106), .B1(n3791), .Y(n1616)
         );
  AOI222XLTS U3200 ( .A0(n4473), .A1(n3570), .B0(n542), .B1(n3553), .C0(n4373), 
        .C1(n3541), .Y(n1617) );
  AOI22X1TS U3201 ( .A0(n4273), .A1(n3521), .B0(n4103), .B1(n3791), .Y(n1614)
         );
  AOI222XLTS U3202 ( .A0(n4470), .A1(n3567), .B0(n544), .B1(n3554), .C0(n4370), 
        .C1(n3540), .Y(n1615) );
  AOI22X1TS U3203 ( .A0(n4270), .A1(n3521), .B0(n4100), .B1(n3791), .Y(n1612)
         );
  AOI222XLTS U3204 ( .A0(n4466), .A1(n3567), .B0(n496), .B1(n3553), .C0(n4367), 
        .C1(n3540), .Y(n1613) );
  AOI22X1TS U3205 ( .A0(n4267), .A1(n3521), .B0(n4097), .B1(n3791), .Y(n1610)
         );
  AOI222XLTS U3206 ( .A0(n4463), .A1(n3567), .B0(n546), .B1(n3553), .C0(n4364), 
        .C1(n3542), .Y(n1611) );
  AOI22X1TS U3207 ( .A0(n4264), .A1(n3520), .B0(n4094), .B1(n3801), .Y(n1608)
         );
  AOI222XLTS U3208 ( .A0(n4460), .A1(n3566), .B0(n548), .B1(n3555), .C0(n4361), 
        .C1(n3540), .Y(n1609) );
  AOI22X1TS U3209 ( .A0(n4261), .A1(n3520), .B0(n4091), .B1(n3800), .Y(n1606)
         );
  AOI222XLTS U3210 ( .A0(n4456), .A1(n3566), .B0(n550), .B1(n3555), .C0(n4358), 
        .C1(n3540), .Y(n1607) );
  AOI22X1TS U3211 ( .A0(n4258), .A1(n3520), .B0(n4088), .B1(n798), .Y(n1604)
         );
  AOI222XLTS U3212 ( .A0(n4453), .A1(n3566), .B0(n780), .B1(n3554), .C0(n4355), 
        .C1(n3539), .Y(n1605) );
  AOI22X1TS U3213 ( .A0(n4255), .A1(n3520), .B0(n4085), .B1(n3802), .Y(n1602)
         );
  AOI222XLTS U3214 ( .A0(n4450), .A1(n3566), .B0(n787), .B1(n3555), .C0(n4352), 
        .C1(n3539), .Y(n1603) );
  AOI22X1TS U3215 ( .A0(n4249), .A1(n3519), .B0(n4079), .B1(n3798), .Y(n1598)
         );
  AOI222XLTS U3216 ( .A0(n4443), .A1(n3580), .B0(n795), .B1(n3565), .C0(n4346), 
        .C1(n3539), .Y(n1599) );
  AOI22X1TS U3217 ( .A0(n4426), .A1(n3259), .B0(n4160), .B1(n3895), .Y(n1396)
         );
  AOI222XLTS U3218 ( .A0(n4534), .A1(n3307), .B0(n506), .B1(n3299), .C0(n4331), 
        .C1(n3280), .Y(n1397) );
  AOI22X1TS U3219 ( .A0(n4411), .A1(n3258), .B0(n4145), .B1(n3894), .Y(n1386)
         );
  AOI222XLTS U3220 ( .A0(n4517), .A1(n3314), .B0(n516), .B1(n3289), .C0(n4316), 
        .C1(n3281), .Y(n1387) );
  AOI22X1TS U3221 ( .A0(n4405), .A1(n3257), .B0(n4139), .B1(n3893), .Y(n1382)
         );
  AOI222XLTS U3222 ( .A0(n4510), .A1(n3315), .B0(n520), .B1(n3289), .C0(n4310), 
        .C1(n3285), .Y(n1383) );
  AOI22X1TS U3223 ( .A0(n4402), .A1(n3257), .B0(n4136), .B1(n3893), .Y(n1380)
         );
  AOI222XLTS U3224 ( .A0(n4507), .A1(n3314), .B0(n522), .B1(n3290), .C0(n4307), 
        .C1(n3282), .Y(n1381) );
  AOI22X1TS U3225 ( .A0(n4375), .A1(n3256), .B0(n4109), .B1(n3891), .Y(n1362)
         );
  AOI222XLTS U3226 ( .A0(n4477), .A1(n3304), .B0(n540), .B1(n3291), .C0(n4280), 
        .C1(n3276), .Y(n1363) );
  AOI22X1TS U3227 ( .A0(n4369), .A1(n3256), .B0(n4103), .B1(n3890), .Y(n1358)
         );
  AOI222XLTS U3228 ( .A0(n4470), .A1(n3304), .B0(n544), .B1(n3291), .C0(n4274), 
        .C1(n3275), .Y(n1359) );
  AOI22X1TS U3229 ( .A0(n4360), .A1(n3255), .B0(n4094), .B1(n3902), .Y(n1352)
         );
  AOI222XLTS U3230 ( .A0(n4460), .A1(n3303), .B0(n548), .B1(n3292), .C0(n4265), 
        .C1(n3275), .Y(n1353) );
  AOI22X1TS U3231 ( .A0(n4351), .A1(n3255), .B0(n4085), .B1(n3898), .Y(n1346)
         );
  AOI222XLTS U3232 ( .A0(n4450), .A1(n3303), .B0(n787), .B1(n3292), .C0(n4256), 
        .C1(n3274), .Y(n1347) );
  AOI22X1TS U3233 ( .A0(n3961), .A1(n3261), .B0(n4058), .B1(n3897), .Y(n2023)
         );
  AOI222XLTS U3234 ( .A0(n4222), .A1(n3309), .B0(n3293), .B1(n42), .C0(n4004), 
        .C1(n3273), .Y(n2024) );
  AOI22X1TS U3235 ( .A0(n3955), .A1(n3261), .B0(n4052), .B1(n3897), .Y(n2019)
         );
  AOI222XLTS U3236 ( .A0(n4216), .A1(n3309), .B0(n3295), .B1(n32), .C0(n3998), 
        .C1(n3279), .Y(n2020) );
  AOI22X1TS U3237 ( .A0(n3952), .A1(n3261), .B0(n4049), .B1(n3897), .Y(n2017)
         );
  AOI222XLTS U3238 ( .A0(n4213), .A1(n3309), .B0(n3295), .B1(n27), .C0(n3995), 
        .C1(n3279), .Y(n2018) );
  AOI22X1TS U3239 ( .A0(n3949), .A1(n3260), .B0(n4046), .B1(n3896), .Y(n2015)
         );
  AOI222XLTS U3240 ( .A0(n4210), .A1(n3308), .B0(n3295), .B1(n22), .C0(n3992), 
        .C1(n3279), .Y(n2016) );
  AOI22X1TS U3241 ( .A0(n3946), .A1(n3260), .B0(n4043), .B1(n3896), .Y(n2013)
         );
  AOI222XLTS U3242 ( .A0(n4207), .A1(n3308), .B0(n3294), .B1(n17), .C0(n3989), 
        .C1(n3279), .Y(n2014) );
  AOI22X1TS U3243 ( .A0(n4439), .A1(n3260), .B0(n4172), .B1(n3896), .Y(n1404)
         );
  AOI222XLTS U3244 ( .A0(n4547), .A1(n3308), .B0(n498), .B1(n3287), .C0(n4343), 
        .C1(n3278), .Y(n1405) );
  AOI22X1TS U3245 ( .A0(n4436), .A1(n3260), .B0(n4169), .B1(n3896), .Y(n1402)
         );
  AOI222XLTS U3246 ( .A0(n4544), .A1(n3308), .B0(n500), .B1(n3299), .C0(n4340), 
        .C1(n3278), .Y(n1403) );
  AOI22X1TS U3247 ( .A0(n4433), .A1(n3259), .B0(n4166), .B1(n3895), .Y(n1400)
         );
  AOI222XLTS U3248 ( .A0(n4541), .A1(n3307), .B0(n502), .B1(n3287), .C0(n4337), 
        .C1(n3278), .Y(n1401) );
  AOI22X1TS U3249 ( .A0(n4429), .A1(n3259), .B0(n4163), .B1(n3895), .Y(n1398)
         );
  AOI222XLTS U3250 ( .A0(n4537), .A1(n3307), .B0(n504), .B1(n3299), .C0(n4334), 
        .C1(n3278), .Y(n1399) );
  AOI22X1TS U3251 ( .A0(n4423), .A1(n3259), .B0(n4157), .B1(n3895), .Y(n1394)
         );
  AOI222XLTS U3252 ( .A0(n4531), .A1(n3307), .B0(n508), .B1(n3288), .C0(n4328), 
        .C1(n3280), .Y(n1395) );
  AOI22X1TS U3253 ( .A0(n4420), .A1(n3258), .B0(n4154), .B1(n3894), .Y(n1392)
         );
  AOI222XLTS U3254 ( .A0(n4527), .A1(n3312), .B0(n510), .B1(n3288), .C0(n4325), 
        .C1(n3282), .Y(n1393) );
  AOI22X1TS U3255 ( .A0(n4417), .A1(n3258), .B0(n4151), .B1(n3894), .Y(n1390)
         );
  AOI222XLTS U3256 ( .A0(n4524), .A1(n3316), .B0(n512), .B1(n3287), .C0(n4322), 
        .C1(n3280), .Y(n1391) );
  AOI22X1TS U3257 ( .A0(n4414), .A1(n3258), .B0(n4148), .B1(n3894), .Y(n1388)
         );
  AOI222XLTS U3258 ( .A0(n4520), .A1(n3317), .B0(n514), .B1(n3289), .C0(n4319), 
        .C1(n3283), .Y(n1389) );
  AOI22X1TS U3259 ( .A0(n4408), .A1(n3257), .B0(n4142), .B1(n3893), .Y(n1384)
         );
  AOI222XLTS U3260 ( .A0(n4514), .A1(n3314), .B0(n518), .B1(n3287), .C0(n4313), 
        .C1(n3285), .Y(n1385) );
  AOI22X1TS U3261 ( .A0(n4399), .A1(n3266), .B0(n4133), .B1(n3893), .Y(n1378)
         );
  AOI222XLTS U3262 ( .A0(n4504), .A1(n3306), .B0(n524), .B1(n3288), .C0(n4304), 
        .C1(n3281), .Y(n1379) );
  AOI22X1TS U3263 ( .A0(n4396), .A1(n3269), .B0(n4130), .B1(n3892), .Y(n1376)
         );
  AOI222XLTS U3264 ( .A0(n4500), .A1(n3306), .B0(n526), .B1(n3290), .C0(n4301), 
        .C1(n3283), .Y(n1377) );
  AOI22X1TS U3265 ( .A0(n4393), .A1(n1252), .B0(n4127), .B1(n3892), .Y(n1374)
         );
  AOI222XLTS U3266 ( .A0(n4497), .A1(n3306), .B0(n528), .B1(n3296), .C0(n4298), 
        .C1(n3285), .Y(n1375) );
  AOI22X1TS U3267 ( .A0(n4390), .A1(n1252), .B0(n4124), .B1(n3892), .Y(n1372)
         );
  AOI222XLTS U3268 ( .A0(n4493), .A1(n3306), .B0(n530), .B1(n3289), .C0(n4295), 
        .C1(n3277), .Y(n1373) );
  AOI22X1TS U3269 ( .A0(n4387), .A1(n3266), .B0(n4121), .B1(n3892), .Y(n1370)
         );
  AOI222XLTS U3270 ( .A0(n4490), .A1(n3305), .B0(n532), .B1(n3288), .C0(n4292), 
        .C1(n3277), .Y(n1371) );
  AOI22X1TS U3271 ( .A0(n4384), .A1(n3267), .B0(n4118), .B1(n3891), .Y(n1368)
         );
  AOI222XLTS U3272 ( .A0(n4487), .A1(n3305), .B0(n534), .B1(n3297), .C0(n4289), 
        .C1(n3277), .Y(n1369) );
  AOI22X1TS U3273 ( .A0(n4381), .A1(n3266), .B0(n4115), .B1(n3891), .Y(n1366)
         );
  AOI222XLTS U3274 ( .A0(n4483), .A1(n3305), .B0(n536), .B1(n3290), .C0(n4286), 
        .C1(n3276), .Y(n1367) );
  AOI22X1TS U3275 ( .A0(n4378), .A1(n3267), .B0(n4112), .B1(n3891), .Y(n1364)
         );
  AOI222XLTS U3276 ( .A0(n4480), .A1(n3305), .B0(n538), .B1(n3291), .C0(n4283), 
        .C1(n3276), .Y(n1365) );
  AOI22X1TS U3277 ( .A0(n4372), .A1(n3257), .B0(n4106), .B1(n3890), .Y(n1360)
         );
  AOI222XLTS U3278 ( .A0(n4473), .A1(n3313), .B0(n542), .B1(n3296), .C0(n4277), 
        .C1(n3276), .Y(n1361) );
  AOI22X1TS U3279 ( .A0(n4366), .A1(n3256), .B0(n4100), .B1(n3890), .Y(n1356)
         );
  AOI222XLTS U3280 ( .A0(n4466), .A1(n3304), .B0(n496), .B1(n3300), .C0(n4271), 
        .C1(n3275), .Y(n1357) );
  AOI22X1TS U3281 ( .A0(n4363), .A1(n3256), .B0(n4097), .B1(n3890), .Y(n1354)
         );
  AOI222XLTS U3282 ( .A0(n4463), .A1(n3304), .B0(n546), .B1(n3298), .C0(n4268), 
        .C1(n3277), .Y(n1355) );
  AOI22X1TS U3283 ( .A0(n4357), .A1(n3255), .B0(n4091), .B1(n3899), .Y(n1350)
         );
  AOI222XLTS U3284 ( .A0(n4456), .A1(n3303), .B0(n550), .B1(n3292), .C0(n4262), 
        .C1(n3275), .Y(n1351) );
  AOI22X1TS U3285 ( .A0(n4354), .A1(n3255), .B0(n4088), .B1(n3900), .Y(n1348)
         );
  AOI222XLTS U3286 ( .A0(n4453), .A1(n3303), .B0(n780), .B1(n3291), .C0(n4259), 
        .C1(n3274), .Y(n1349) );
  AOI22X1TS U3287 ( .A0(n4348), .A1(n3254), .B0(n4082), .B1(n3899), .Y(n1344)
         );
  AOI222XLTS U3288 ( .A0(n4446), .A1(n3302), .B0(n792), .B1(n3292), .C0(n4253), 
        .C1(n3274), .Y(n1345) );
  AOI22X1TS U3289 ( .A0(n4345), .A1(n3254), .B0(n4079), .B1(n3900), .Y(n1342)
         );
  AOI222XLTS U3290 ( .A0(n4443), .A1(n3302), .B0(n795), .B1(n3290), .C0(n4250), 
        .C1(n3274), .Y(n1343) );
  AOI22X1TS U3291 ( .A0(n4541), .A1(n3643), .B0(n4166), .B1(n3775), .Y(n1721)
         );
  AOI222XLTS U3292 ( .A0(n4434), .A1(n3772), .B0(n501), .B1(n3630), .C0(n4337), 
        .C1(n3609), .Y(n1722) );
  AOI22X1TS U3293 ( .A0(n4520), .A1(n3637), .B0(n4148), .B1(n3777), .Y(n1709)
         );
  AOI222XLTS U3294 ( .A0(n4415), .A1(n3767), .B0(n513), .B1(n3628), .C0(n4319), 
        .C1(n3608), .Y(n1710) );
  AOI22X1TS U3295 ( .A0(n4514), .A1(n3637), .B0(n4142), .B1(n3777), .Y(n1705)
         );
  AOI222XLTS U3296 ( .A0(n4409), .A1(n3767), .B0(n517), .B1(n3619), .C0(n4313), 
        .C1(n3607), .Y(n1706) );
  AOI22X1TS U3297 ( .A0(n4510), .A1(n3637), .B0(n4139), .B1(n3788), .Y(n1703)
         );
  AOI222XLTS U3298 ( .A0(n4406), .A1(n3767), .B0(n519), .B1(n3619), .C0(n4310), 
        .C1(n3607), .Y(n1704) );
  AOI22X1TS U3299 ( .A0(n4487), .A1(n3635), .B0(n4118), .B1(n3787), .Y(n1689)
         );
  AOI222XLTS U3300 ( .A0(n4385), .A1(n3765), .B0(n533), .B1(n3620), .C0(n4289), 
        .C1(n3605), .Y(n1690) );
  AOI22X1TS U3301 ( .A0(n4483), .A1(n3635), .B0(n4115), .B1(n3779), .Y(n1687)
         );
  AOI222XLTS U3302 ( .A0(n4382), .A1(n3765), .B0(n535), .B1(n3621), .C0(n4286), 
        .C1(n3605), .Y(n1688) );
  AOI22X1TS U3303 ( .A0(n4477), .A1(n3634), .B0(n4109), .B1(n3778), .Y(n1683)
         );
  AOI222XLTS U3304 ( .A0(n4376), .A1(n3764), .B0(n539), .B1(n3624), .C0(n4280), 
        .C1(n3604), .Y(n1684) );
  AOI22X1TS U3305 ( .A0(n4463), .A1(n3633), .B0(n4097), .B1(n3780), .Y(n1675)
         );
  AOI222XLTS U3306 ( .A0(n4364), .A1(n3763), .B0(n545), .B1(n3623), .C0(n4268), 
        .C1(n3605), .Y(n1676) );
  AOI22X1TS U3307 ( .A0(n4547), .A1(n3643), .B0(n4172), .B1(n3775), .Y(n1725)
         );
  AOI222XLTS U3308 ( .A0(n4441), .A1(n3772), .B0(n497), .B1(n3624), .C0(n4343), 
        .C1(n3613), .Y(n1726) );
  AOI22X1TS U3309 ( .A0(n4544), .A1(n3643), .B0(n4169), .B1(n3776), .Y(n1723)
         );
  AOI222XLTS U3310 ( .A0(n4437), .A1(n3770), .B0(n499), .B1(n3628), .C0(n4340), 
        .C1(n3615), .Y(n1724) );
  AOI22X1TS U3311 ( .A0(n4537), .A1(n3645), .B0(n4163), .B1(n3775), .Y(n1719)
         );
  AOI222XLTS U3312 ( .A0(n4430), .A1(n3771), .B0(n503), .B1(n3628), .C0(n4334), 
        .C1(n3609), .Y(n1720) );
  AOI22X1TS U3313 ( .A0(n4534), .A1(n3638), .B0(n4160), .B1(n3786), .Y(n1717)
         );
  AOI222XLTS U3314 ( .A0(n4427), .A1(n3768), .B0(n505), .B1(n3628), .C0(n4331), 
        .C1(n3609), .Y(n1718) );
  AOI22X1TS U3315 ( .A0(n4531), .A1(n3638), .B0(n4157), .B1(n3788), .Y(n1715)
         );
  AOI222XLTS U3316 ( .A0(n4424), .A1(n3768), .B0(n507), .B1(n3621), .C0(n4328), 
        .C1(n3609), .Y(n1716) );
  AOI22X1TS U3317 ( .A0(n4524), .A1(n3638), .B0(n4151), .B1(n3777), .Y(n1711)
         );
  AOI222XLTS U3318 ( .A0(n4418), .A1(n3768), .B0(n511), .B1(n3627), .C0(n4322), 
        .C1(n3608), .Y(n1712) );
  AOI22X1TS U3319 ( .A0(n4517), .A1(n3637), .B0(n4145), .B1(n3776), .Y(n1707)
         );
  AOI222XLTS U3320 ( .A0(n4412), .A1(n3767), .B0(n515), .B1(n3625), .C0(n4316), 
        .C1(n3608), .Y(n1708) );
  AOI22X1TS U3321 ( .A0(n4507), .A1(n3636), .B0(n4136), .B1(n3787), .Y(n1701)
         );
  AOI222XLTS U3322 ( .A0(n4403), .A1(n3766), .B0(n521), .B1(n3619), .C0(n4307), 
        .C1(n3607), .Y(n1702) );
  AOI22X1TS U3323 ( .A0(n4500), .A1(n3636), .B0(n4130), .B1(n3775), .Y(n1697)
         );
  AOI222XLTS U3324 ( .A0(n4397), .A1(n3766), .B0(n525), .B1(n3619), .C0(n4301), 
        .C1(n3606), .Y(n1698) );
  AOI22X1TS U3325 ( .A0(n4497), .A1(n3636), .B0(n4127), .B1(n3777), .Y(n1695)
         );
  AOI222XLTS U3326 ( .A0(n4394), .A1(n3766), .B0(n527), .B1(n3620), .C0(n4298), 
        .C1(n3606), .Y(n1696) );
  AOI22X1TS U3327 ( .A0(n4493), .A1(n3635), .B0(n4124), .B1(n3788), .Y(n1693)
         );
  AOI222XLTS U3328 ( .A0(n4391), .A1(n3765), .B0(n529), .B1(n3621), .C0(n4295), 
        .C1(n3606), .Y(n1694) );
  AOI22X1TS U3329 ( .A0(n4490), .A1(n3635), .B0(n4121), .B1(n3778), .Y(n1691)
         );
  AOI222XLTS U3330 ( .A0(n4388), .A1(n3765), .B0(n531), .B1(n3620), .C0(n4292), 
        .C1(n3606), .Y(n1692) );
  AOI22X1TS U3331 ( .A0(n4480), .A1(n3634), .B0(n4112), .B1(n3779), .Y(n1685)
         );
  AOI222XLTS U3332 ( .A0(n4379), .A1(n3764), .B0(n537), .B1(n3621), .C0(n4283), 
        .C1(n3605), .Y(n1686) );
  AOI22X1TS U3333 ( .A0(n4473), .A1(n3634), .B0(n4106), .B1(n3779), .Y(n1681)
         );
  AOI222XLTS U3334 ( .A0(n4373), .A1(n3764), .B0(n541), .B1(n3622), .C0(n4277), 
        .C1(n3604), .Y(n1682) );
  AOI22X1TS U3335 ( .A0(n4470), .A1(n3634), .B0(n4103), .B1(n3778), .Y(n1679)
         );
  AOI222XLTS U3336 ( .A0(n4370), .A1(n3764), .B0(n543), .B1(n3622), .C0(n4274), 
        .C1(n3604), .Y(n1680) );
  AOI22X1TS U3337 ( .A0(n4466), .A1(n3633), .B0(n4100), .B1(n3778), .Y(n1677)
         );
  AOI222XLTS U3338 ( .A0(n4367), .A1(n3763), .B0(n495), .B1(n3622), .C0(n4271), 
        .C1(n3604), .Y(n1678) );
  AOI22X1TS U3339 ( .A0(n4460), .A1(n3633), .B0(n4094), .B1(n3780), .Y(n1673)
         );
  AOI222XLTS U3340 ( .A0(n4361), .A1(n3763), .B0(n547), .B1(n3622), .C0(n4265), 
        .C1(n3603), .Y(n1674) );
  AOI22X1TS U3341 ( .A0(n4453), .A1(n3632), .B0(n4088), .B1(n3780), .Y(n1669)
         );
  AOI222XLTS U3342 ( .A0(n4355), .A1(n3762), .B0(n551), .B1(n3624), .C0(n4259), 
        .C1(n3603), .Y(n1670) );
  AOI22X1TS U3343 ( .A0(n4450), .A1(n3632), .B0(n4085), .B1(n3780), .Y(n1667)
         );
  AOI222XLTS U3344 ( .A0(n4352), .A1(n3762), .B0(n786), .B1(n3623), .C0(n4256), 
        .C1(n3613), .Y(n1668) );
  AOI22X1TS U3345 ( .A0(n4527), .A1(n3638), .B0(n4154), .B1(n3776), .Y(n1713)
         );
  AOI222XLTS U3346 ( .A0(n4421), .A1(n3768), .B0(n509), .B1(n3626), .C0(n4325), 
        .C1(n3608), .Y(n1714) );
  AOI22X1TS U3347 ( .A0(n4504), .A1(n3636), .B0(n4133), .B1(n3785), .Y(n1699)
         );
  AOI222XLTS U3348 ( .A0(n4400), .A1(n3766), .B0(n523), .B1(n3620), .C0(n4304), 
        .C1(n3607), .Y(n1700) );
  AOI22X1TS U3349 ( .A0(n4456), .A1(n3633), .B0(n4091), .B1(n3779), .Y(n1671)
         );
  AOI222XLTS U3350 ( .A0(n4358), .A1(n3763), .B0(n549), .B1(n3623), .C0(n4262), 
        .C1(n3603), .Y(n1672) );
  AOI22X1TS U3351 ( .A0(n793), .A1(n3478), .B0(n4345), .B1(n3454), .Y(n1534)
         );
  AOI222XLTS U3352 ( .A0(n3044), .A1(n190), .B0(n4444), .B1(n3486), .C0(n4080), 
        .C1(n3805), .Y(n1535) );
  AOI22X1TS U3353 ( .A0(n789), .A1(n3481), .B0(n4348), .B1(n3454), .Y(n1536)
         );
  AOI222XLTS U3354 ( .A0(n3042), .A1(n187), .B0(n4447), .B1(n3486), .C0(n4083), 
        .C1(n3805), .Y(n1537) );
  AOI22X1TS U3355 ( .A0(n786), .A1(n3482), .B0(n4351), .B1(n3455), .Y(n1538)
         );
  AOI222XLTS U3356 ( .A0(n3040), .A1(n199), .B0(n4451), .B1(n3487), .C0(n4086), 
        .C1(n3806), .Y(n1539) );
  AOI22X1TS U3357 ( .A0(n551), .A1(n3480), .B0(n4354), .B1(n3455), .Y(n1540)
         );
  AOI222XLTS U3358 ( .A0(n3038), .A1(n194), .B0(n4454), .B1(n3487), .C0(n4089), 
        .C1(n3806), .Y(n1541) );
  AOI22X1TS U3359 ( .A0(n549), .A1(n3479), .B0(n4357), .B1(n3455), .Y(n1542)
         );
  AOI222XLTS U3360 ( .A0(n3036), .A1(n3803), .B0(n4457), .B1(n3487), .C0(n4092), .C1(n3806), .Y(n1543) );
  AOI22X1TS U3361 ( .A0(n547), .A1(n3477), .B0(n4360), .B1(n3455), .Y(n1544)
         );
  AOI222XLTS U3362 ( .A0(n3034), .A1(n191), .B0(n4461), .B1(n3487), .C0(n4095), 
        .C1(n3806), .Y(n1545) );
  AOI22X1TS U3363 ( .A0(n545), .A1(n3482), .B0(n4363), .B1(n3456), .Y(n1546)
         );
  AOI222XLTS U3364 ( .A0(n3032), .A1(n199), .B0(n4464), .B1(n3500), .C0(n4098), 
        .C1(n3807), .Y(n1547) );
  AOI22X1TS U3365 ( .A0(n495), .A1(n3477), .B0(n4366), .B1(n3456), .Y(n1548)
         );
  AOI222XLTS U3366 ( .A0(n3030), .A1(n196), .B0(n4468), .B1(n3488), .C0(n4101), 
        .C1(n3807), .Y(n1549) );
  AOI22X1TS U3367 ( .A0(n543), .A1(n3477), .B0(n4369), .B1(n3456), .Y(n1550)
         );
  AOI222XLTS U3368 ( .A0(n3028), .A1(n194), .B0(n4471), .B1(n3488), .C0(n4104), 
        .C1(n3807), .Y(n1551) );
  AOI22X1TS U3369 ( .A0(n541), .A1(n3477), .B0(n4372), .B1(n3464), .Y(n1552)
         );
  AOI222XLTS U3370 ( .A0(n3026), .A1(n191), .B0(n4474), .B1(n3488), .C0(n4107), 
        .C1(n3807), .Y(n1553) );
  AOI22X1TS U3371 ( .A0(n539), .A1(n3478), .B0(n4375), .B1(n3456), .Y(n1554)
         );
  AOI222XLTS U3372 ( .A0(n3024), .A1(n198), .B0(n4478), .B1(n3488), .C0(n4110), 
        .C1(n3808), .Y(n1555) );
  AOI22X1TS U3373 ( .A0(n537), .A1(n3478), .B0(n4378), .B1(n3457), .Y(n1556)
         );
  AOI222XLTS U3374 ( .A0(n3022), .A1(n187), .B0(n4481), .B1(n3489), .C0(n4113), 
        .C1(n3808), .Y(n1557) );
  AOI22X1TS U3375 ( .A0(n535), .A1(n3482), .B0(n4381), .B1(n3457), .Y(n1558)
         );
  AOI222XLTS U3376 ( .A0(n3020), .A1(n112), .B0(n4484), .B1(n3489), .C0(n4116), 
        .C1(n3808), .Y(n1559) );
  AOI22X1TS U3377 ( .A0(n533), .A1(n3476), .B0(n4384), .B1(n3457), .Y(n1560)
         );
  AOI222XLTS U3378 ( .A0(n3018), .A1(n196), .B0(n4488), .B1(n3489), .C0(n4119), 
        .C1(n3808), .Y(n1561) );
  AOI22X1TS U3379 ( .A0(n531), .A1(n3476), .B0(n4387), .B1(n3457), .Y(n1562)
         );
  AOI222XLTS U3380 ( .A0(n3016), .A1(n3803), .B0(n4491), .B1(n3489), .C0(n4122), .C1(n3809), .Y(n1563) );
  AOI22X1TS U3381 ( .A0(n529), .A1(n3479), .B0(n4390), .B1(n3458), .Y(n1564)
         );
  AOI222XLTS U3382 ( .A0(n3014), .A1(n191), .B0(n4495), .B1(n3495), .C0(n4125), 
        .C1(n3809), .Y(n1565) );
  AOI22X1TS U3383 ( .A0(n527), .A1(n3476), .B0(n4393), .B1(n3458), .Y(n1566)
         );
  AOI222XLTS U3384 ( .A0(n3012), .A1(n190), .B0(n4498), .B1(n3497), .C0(n4128), 
        .C1(n3809), .Y(n1567) );
  AOI22X1TS U3385 ( .A0(n525), .A1(n3475), .B0(n4396), .B1(n3458), .Y(n1568)
         );
  AOI222XLTS U3386 ( .A0(n3010), .A1(n196), .B0(n4501), .B1(n3497), .C0(n4131), 
        .C1(n3809), .Y(n1569) );
  AOI22X1TS U3387 ( .A0(n523), .A1(n3476), .B0(n4399), .B1(n3458), .Y(n1570)
         );
  AOI222XLTS U3388 ( .A0(n3008), .A1(n198), .B0(n4505), .B1(n3496), .C0(n4134), 
        .C1(n3812), .Y(n1571) );
  AOI22X1TS U3389 ( .A0(n521), .A1(n3475), .B0(n4402), .B1(n1204), .Y(n1572)
         );
  AOI222XLTS U3390 ( .A0(n3006), .A1(n196), .B0(n4508), .B1(n3494), .C0(n4137), 
        .C1(n3817), .Y(n1573) );
  AOI22X1TS U3391 ( .A0(n519), .A1(n3475), .B0(n4405), .B1(n3466), .Y(n1574)
         );
  AOI222XLTS U3392 ( .A0(n3004), .A1(n193), .B0(n4511), .B1(n3498), .C0(n4140), 
        .C1(n3813), .Y(n1575) );
  AOI22X1TS U3393 ( .A0(n517), .A1(n3475), .B0(n4408), .B1(n3465), .Y(n1576)
         );
  AOI222XLTS U3394 ( .A0(n3002), .A1(n189), .B0(n4515), .B1(n3498), .C0(n4143), 
        .C1(n3814), .Y(n1577) );
  AOI22X1TS U3395 ( .A0(n515), .A1(n3474), .B0(n4411), .B1(n3463), .Y(n1578)
         );
  AOI222XLTS U3396 ( .A0(n3000), .A1(n198), .B0(n4518), .B1(n3490), .C0(n4146), 
        .C1(n3813), .Y(n1579) );
  AOI22X1TS U3397 ( .A0(n513), .A1(n3474), .B0(n4414), .B1(n3466), .Y(n1580)
         );
  AOI222XLTS U3398 ( .A0(n2998), .A1(n194), .B0(n4522), .B1(n3490), .C0(n4149), 
        .C1(n3814), .Y(n1581) );
  AOI22X1TS U3399 ( .A0(n511), .A1(n3474), .B0(n4417), .B1(n3465), .Y(n1582)
         );
  AOI222XLTS U3400 ( .A0(n2996), .A1(n191), .B0(n4525), .B1(n3490), .C0(n4152), 
        .C1(n3812), .Y(n1583) );
  AOI22X1TS U3401 ( .A0(n509), .A1(n3473), .B0(n4420), .B1(n3467), .Y(n1584)
         );
  AOI222XLTS U3402 ( .A0(n2994), .A1(n197), .B0(n4528), .B1(n3490), .C0(n4155), 
        .C1(n3817), .Y(n1585) );
  AOI22X1TS U3403 ( .A0(n507), .A1(n3480), .B0(n4423), .B1(n3469), .Y(n1586)
         );
  AOI222XLTS U3404 ( .A0(n2992), .A1(n797), .B0(n4532), .B1(n3491), .C0(n4158), 
        .C1(n3815), .Y(n1587) );
  AOI22X1TS U3405 ( .A0(n505), .A1(n3474), .B0(n4426), .B1(n3469), .Y(n1588)
         );
  AOI222XLTS U3406 ( .A0(n2990), .A1(n197), .B0(n4535), .B1(n3491), .C0(n4161), 
        .C1(n3815), .Y(n1589) );
  AOI22X1TS U3407 ( .A0(n503), .A1(n3473), .B0(n4429), .B1(n3463), .Y(n1590)
         );
  AOI222XLTS U3408 ( .A0(n2988), .A1(n197), .B0(n4538), .B1(n3491), .C0(n4164), 
        .C1(n3815), .Y(n1591) );
  AOI22X1TS U3409 ( .A0(n501), .A1(n3473), .B0(n4433), .B1(n3469), .Y(n1592)
         );
  AOI222XLTS U3410 ( .A0(n2986), .A1(n3803), .B0(n4542), .B1(n3491), .C0(n4167), .C1(n3817), .Y(n1593) );
  AOI22X1TS U3411 ( .A0(n499), .A1(n3473), .B0(n4436), .B1(n3459), .Y(n1594)
         );
  AOI222XLTS U3412 ( .A0(n2984), .A1(n190), .B0(n4545), .B1(n3492), .C0(n4170), 
        .C1(n3810), .Y(n1595) );
  AOI22X1TS U3413 ( .A0(n497), .A1(n3481), .B0(n4439), .B1(n3459), .Y(n1596)
         );
  AOI222XLTS U3414 ( .A0(n2982), .A1(n199), .B0(n4549), .B1(n3492), .C0(n4173), 
        .C1(n3810), .Y(n1597) );
  AOI22X1TS U3415 ( .A0(n3470), .A1(n40), .B0(n3961), .B1(n3460), .Y(n1953) );
  AOI222XLTS U3416 ( .A0(n3046), .A1(n3803), .B0(n4223), .B1(n3486), .C0(n4059), .C1(n3811), .Y(n1954) );
  AOI22X1TS U3417 ( .A0(n3472), .A1(n31), .B0(n3955), .B1(n3460), .Y(n1949) );
  AOI222XLTS U3418 ( .A0(n3050), .A1(n193), .B0(n4217), .B1(n3493), .C0(n4053), 
        .C1(n3811), .Y(n1950) );
  AOI22X1TS U3419 ( .A0(n3472), .A1(n25), .B0(n3952), .B1(n3460), .Y(n1947) );
  AOI222XLTS U3420 ( .A0(n3052), .A1(n189), .B0(n4214), .B1(n3493), .C0(n4050), 
        .C1(n3811), .Y(n1948) );
  AOI22X1TS U3421 ( .A0(n3471), .A1(n21), .B0(n3949), .B1(n3459), .Y(n1945) );
  AOI222XLTS U3422 ( .A0(n3054), .A1(n193), .B0(n4211), .B1(n3492), .C0(n4047), 
        .C1(n3810), .Y(n1946) );
  AOI22X1TS U3423 ( .A0(n3472), .A1(n16), .B0(n3946), .B1(n3459), .Y(n1943) );
  AOI222XLTS U3424 ( .A0(n3056), .A1(n189), .B0(n4208), .B1(n3492), .C0(n4044), 
        .C1(n3810), .Y(n1944) );
  AOI22X1TS U3425 ( .A0(n3472), .A1(n36), .B0(n3958), .B1(n3460), .Y(n1951) );
  AOI222XLTS U3426 ( .A0(n3048), .A1(n198), .B0(n4220), .B1(n3493), .C0(n4056), 
        .C1(n3811), .Y(n1952) );
  AOI22X1TS U3427 ( .A0(n4439), .A1(n3426), .B0(n4547), .B1(n3415), .Y(n1532)
         );
  AOI222XLTS U3428 ( .A0(n498), .A1(n3854), .B0(n4173), .B1(n3877), .C0(n66), 
        .C1(n3870), .Y(n1533) );
  AOI22X1TS U3429 ( .A0(n4436), .A1(n3426), .B0(n4544), .B1(n3415), .Y(n1530)
         );
  AOI222XLTS U3430 ( .A0(n500), .A1(n3860), .B0(n4170), .B1(n3877), .C0(n67), 
        .C1(n3869), .Y(n1531) );
  AOI22X1TS U3431 ( .A0(n4433), .A1(n3425), .B0(n4541), .B1(n3413), .Y(n1528)
         );
  AOI222XLTS U3432 ( .A0(n502), .A1(n3859), .B0(n4167), .B1(n3878), .C0(n68), 
        .C1(n3871), .Y(n1529) );
  AOI22X1TS U3433 ( .A0(n4429), .A1(n3425), .B0(n4537), .B1(n3413), .Y(n1526)
         );
  AOI222XLTS U3434 ( .A0(n504), .A1(n791), .B0(n4164), .B1(n3878), .C0(n69), 
        .C1(n3872), .Y(n1527) );
  AOI22X1TS U3435 ( .A0(n4426), .A1(n3425), .B0(n4534), .B1(n3414), .Y(n1524)
         );
  AOI222XLTS U3436 ( .A0(n506), .A1(n3857), .B0(n4161), .B1(n3878), .C0(n70), 
        .C1(n3872), .Y(n1525) );
  AOI22X1TS U3437 ( .A0(n4423), .A1(n3425), .B0(n4531), .B1(n3416), .Y(n1522)
         );
  AOI222XLTS U3438 ( .A0(n508), .A1(n3851), .B0(n4158), .B1(n3878), .C0(n71), 
        .C1(n3875), .Y(n1523) );
  AOI22X1TS U3439 ( .A0(n4417), .A1(n3424), .B0(n4524), .B1(n3409), .Y(n1518)
         );
  AOI222XLTS U3440 ( .A0(n512), .A1(n3857), .B0(n4152), .B1(n3879), .C0(n72), 
        .C1(n3869), .Y(n1519) );
  AOI22X1TS U3441 ( .A0(n4411), .A1(n3424), .B0(n4517), .B1(n3409), .Y(n1514)
         );
  AOI222XLTS U3442 ( .A0(n516), .A1(n791), .B0(n4146), .B1(n3879), .C0(n73), 
        .C1(n3868), .Y(n1515) );
  AOI22X1TS U3443 ( .A0(n4408), .A1(n3423), .B0(n4514), .B1(n3408), .Y(n1512)
         );
  AOI222XLTS U3444 ( .A0(n518), .A1(n3849), .B0(n4143), .B1(n3880), .C0(n74), 
        .C1(n3868), .Y(n1513) );
  AOI22X1TS U3445 ( .A0(n4402), .A1(n3423), .B0(n4507), .B1(n3408), .Y(n1508)
         );
  AOI222XLTS U3446 ( .A0(n522), .A1(n3849), .B0(n4137), .B1(n3880), .C0(n75), 
        .C1(n3867), .Y(n1509) );
  AOI22X1TS U3447 ( .A0(n4396), .A1(n3434), .B0(n4500), .B1(n3407), .Y(n1504)
         );
  AOI222XLTS U3448 ( .A0(n526), .A1(n3849), .B0(n4131), .B1(n3885), .C0(n76), 
        .C1(n3867), .Y(n1505) );
  AOI22X1TS U3449 ( .A0(n4393), .A1(n3433), .B0(n4497), .B1(n3407), .Y(n1502)
         );
  AOI222XLTS U3450 ( .A0(n528), .A1(n3850), .B0(n4128), .B1(n3887), .C0(n77), 
        .C1(n3867), .Y(n1503) );
  AOI22X1TS U3451 ( .A0(n4387), .A1(n3435), .B0(n4490), .B1(n3406), .Y(n1498)
         );
  AOI222XLTS U3452 ( .A0(n532), .A1(n3850), .B0(n4122), .B1(n3885), .C0(n78), 
        .C1(n3866), .Y(n1499) );
  AOI22X1TS U3453 ( .A0(n4381), .A1(n1218), .B0(n4483), .B1(n3406), .Y(n1494)
         );
  AOI222XLTS U3454 ( .A0(n536), .A1(n3851), .B0(n4116), .B1(n3881), .C0(n79), 
        .C1(n3865), .Y(n1495) );
  AOI22X1TS U3455 ( .A0(n4378), .A1(n3433), .B0(n4480), .B1(n3406), .Y(n1492)
         );
  AOI222XLTS U3456 ( .A0(n538), .A1(n3851), .B0(n4113), .B1(n3881), .C0(n80), 
        .C1(n3865), .Y(n1493) );
  AOI22X1TS U3457 ( .A0(n4375), .A1(n3422), .B0(n4477), .B1(n3405), .Y(n1490)
         );
  AOI222XLTS U3458 ( .A0(n540), .A1(n3854), .B0(n4110), .B1(n3881), .C0(n81), 
        .C1(n3865), .Y(n1491) );
  AOI22X1TS U3459 ( .A0(n4372), .A1(n3423), .B0(n4473), .B1(n3408), .Y(n1488)
         );
  AOI222XLTS U3460 ( .A0(n542), .A1(n3852), .B0(n4107), .B1(n3884), .C0(n82), 
        .C1(n3865), .Y(n1489) );
  AOI22X1TS U3461 ( .A0(n4369), .A1(n3422), .B0(n4470), .B1(n3405), .Y(n1486)
         );
  AOI222XLTS U3462 ( .A0(n544), .A1(n3852), .B0(n4104), .B1(n3884), .C0(n83), 
        .C1(n3864), .Y(n1487) );
  AOI22X1TS U3463 ( .A0(n4363), .A1(n3422), .B0(n4463), .B1(n3405), .Y(n1482)
         );
  AOI222XLTS U3464 ( .A0(n546), .A1(n3853), .B0(n4098), .B1(n3888), .C0(n84), 
        .C1(n3864), .Y(n1483) );
  AOI22X1TS U3465 ( .A0(n4354), .A1(n3421), .B0(n4453), .B1(n3404), .Y(n1476)
         );
  AOI222XLTS U3466 ( .A0(n780), .A1(n3854), .B0(n4089), .B1(n3882), .C0(n85), 
        .C1(n3864), .Y(n1477) );
  AOI22X1TS U3467 ( .A0(n4348), .A1(n3420), .B0(n4446), .B1(n3403), .Y(n1472)
         );
  AOI222XLTS U3468 ( .A0(n792), .A1(n3853), .B0(n4083), .B1(n3889), .C0(n86), 
        .C1(n3863), .Y(n1473) );
  AOI22X1TS U3469 ( .A0(n4345), .A1(n3420), .B0(n4443), .B1(n3403), .Y(n1470)
         );
  AOI222XLTS U3470 ( .A0(n795), .A1(n3854), .B0(n4080), .B1(n3886), .C0(n87), 
        .C1(n3862), .Y(n1471) );
  AOI22X1TS U3471 ( .A0(n4420), .A1(n3424), .B0(n4527), .B1(n3409), .Y(n1520)
         );
  AOI222XLTS U3472 ( .A0(n510), .A1(n3858), .B0(n4155), .B1(n3879), .C0(n91), 
        .C1(n3875), .Y(n1521) );
  AOI22X1TS U3473 ( .A0(n4414), .A1(n3424), .B0(n4520), .B1(n3409), .Y(n1516)
         );
  AOI222XLTS U3474 ( .A0(n514), .A1(n3855), .B0(n4149), .B1(n3879), .C0(n92), 
        .C1(n3868), .Y(n1517) );
  AOI22X1TS U3475 ( .A0(n4405), .A1(n3423), .B0(n4510), .B1(n3408), .Y(n1510)
         );
  AOI222XLTS U3476 ( .A0(n520), .A1(n3849), .B0(n4140), .B1(n3880), .C0(n93), 
        .C1(n3868), .Y(n1511) );
  AOI22X1TS U3477 ( .A0(n4399), .A1(n3432), .B0(n4504), .B1(n3407), .Y(n1506)
         );
  AOI222XLTS U3478 ( .A0(n524), .A1(n3850), .B0(n4134), .B1(n3880), .C0(n94), 
        .C1(n3867), .Y(n1507) );
  AOI22X1TS U3479 ( .A0(n4390), .A1(n3432), .B0(n4493), .B1(n3407), .Y(n1500)
         );
  AOI222XLTS U3480 ( .A0(n530), .A1(n3851), .B0(n4125), .B1(n3887), .C0(n95), 
        .C1(n3866), .Y(n1501) );
  AOI22X1TS U3481 ( .A0(n4384), .A1(n1218), .B0(n4487), .B1(n3406), .Y(n1496)
         );
  AOI222XLTS U3482 ( .A0(n534), .A1(n3850), .B0(n4119), .B1(n3881), .C0(n96), 
        .C1(n3866), .Y(n1497) );
  AOI22X1TS U3483 ( .A0(n4360), .A1(n3421), .B0(n4460), .B1(n3404), .Y(n1480)
         );
  AOI222XLTS U3484 ( .A0(n548), .A1(n3852), .B0(n4095), .B1(n3882), .C0(n97), 
        .C1(n3864), .Y(n1481) );
  AOI22X1TS U3485 ( .A0(n4357), .A1(n3421), .B0(n4456), .B1(n3404), .Y(n1478)
         );
  AOI222XLTS U3486 ( .A0(n550), .A1(n3853), .B0(n4092), .B1(n3882), .C0(n98), 
        .C1(n3863), .Y(n1479) );
  AOI22X1TS U3487 ( .A0(n4351), .A1(n3421), .B0(n4450), .B1(n3404), .Y(n1474)
         );
  AOI222XLTS U3488 ( .A0(n787), .A1(n3853), .B0(n4086), .B1(n3882), .C0(n99), 
        .C1(n3863), .Y(n1475) );
  AOI22X1TS U3489 ( .A0(n4366), .A1(n3422), .B0(n4466), .B1(n3405), .Y(n1484)
         );
  AOI222XLTS U3490 ( .A0(n496), .A1(n3852), .B0(n4101), .B1(n3889), .C0(n3861), 
        .C1(n692), .Y(n1485) );
  AOI222XLTS U3491 ( .A0(n794), .A1(n966), .B0(n4464), .B1(n3374), .C0(n4098), 
        .C1(n3836), .Y(n1419) );
  AOI222XLTS U3492 ( .A0(n3827), .A1(n965), .B0(n4478), .B1(n3371), .C0(n4110), 
        .C1(n3837), .Y(n1427) );
  AOI222XLTS U3493 ( .A0(n3823), .A1(n964), .B0(n4535), .B1(n3376), .C0(n4161), 
        .C1(n3846), .Y(n1461) );
  AOI222XLTS U3494 ( .A0(n3829), .A1(n963), .B0(n4468), .B1(n3371), .C0(n4101), 
        .C1(n3836), .Y(n1421) );
  AOI222XLTS U3495 ( .A0(n3828), .A1(n962), .B0(n4471), .B1(n3371), .C0(n4104), 
        .C1(n3836), .Y(n1423) );
  AOI222XLTS U3496 ( .A0(n3829), .A1(n961), .B0(n4474), .B1(n3371), .C0(n4107), 
        .C1(n3836), .Y(n1425) );
  AOI222XLTS U3497 ( .A0(n794), .A1(n960), .B0(n4481), .B1(n3372), .C0(n4113), 
        .C1(n3837), .Y(n1429) );
  AOI222XLTS U3498 ( .A0(n3830), .A1(n959), .B0(n4484), .B1(n3372), .C0(n4116), 
        .C1(n3837), .Y(n1431) );
  AOI222XLTS U3499 ( .A0(n3830), .A1(n958), .B0(n4488), .B1(n3372), .C0(n4119), 
        .C1(n3837), .Y(n1433) );
  AOI222XLTS U3500 ( .A0(n3821), .A1(n957), .B0(n4505), .B1(n3373), .C0(n4134), 
        .C1(n3839), .Y(n1443) );
  AOI222XLTS U3501 ( .A0(n3821), .A1(n956), .B0(n4508), .B1(n3374), .C0(n4137), 
        .C1(n3839), .Y(n1445) );
  AOI222XLTS U3502 ( .A0(n3821), .A1(n955), .B0(n4511), .B1(n3374), .C0(n4140), 
        .C1(n3839), .Y(n1447) );
  AOI222XLTS U3503 ( .A0(n3822), .A1(n954), .B0(n4515), .B1(n3374), .C0(n4143), 
        .C1(n3839), .Y(n1449) );
  AOI222XLTS U3504 ( .A0(n3822), .A1(n953), .B0(n4522), .B1(n3375), .C0(n4149), 
        .C1(n3844), .Y(n1453) );
  AOI222XLTS U3505 ( .A0(n3823), .A1(n952), .B0(n4528), .B1(n3375), .C0(n4155), 
        .C1(n3844), .Y(n1457) );
  AOI222XLTS U3506 ( .A0(n3823), .A1(n951), .B0(n4532), .B1(n3376), .C0(n4158), 
        .C1(n3842), .Y(n1459) );
  AOI222XLTS U3507 ( .A0(n3823), .A1(n950), .B0(n4538), .B1(n3376), .C0(n4164), 
        .C1(n3843), .Y(n1463) );
  AOI222XLTS U3508 ( .A0(n3821), .A1(n949), .B0(n4542), .B1(n3376), .C0(n4167), 
        .C1(n3846), .Y(n1465) );
  AOI222XLTS U3509 ( .A0(n3825), .A1(n948), .B0(n4217), .B1(n3377), .C0(n4053), 
        .C1(n3840), .Y(n1997) );
  AOI222XLTS U3510 ( .A0(n3824), .A1(n947), .B0(n4220), .B1(n3377), .C0(n4056), 
        .C1(n3842), .Y(n1999) );
  AOI222XLTS U3511 ( .A0(n3818), .A1(n946), .B0(n4223), .B1(n3369), .C0(n4059), 
        .C1(n3841), .Y(n2001) );
  AOI222XLTS U3512 ( .A0(n3825), .A1(n945), .B0(n4214), .B1(n3377), .C0(n4050), 
        .C1(n3843), .Y(n1995) );
  AOI222XLTS U3513 ( .A0(n3818), .A1(n944), .B0(n4444), .B1(n3369), .C0(n4080), 
        .C1(n3834), .Y(n1407) );
  AOI222XLTS U3514 ( .A0(n3818), .A1(n943), .B0(n4447), .B1(n3369), .C0(n4083), 
        .C1(n3834), .Y(n1409) );
  AOI22X1TS U3515 ( .A0(n3958), .A1(n3261), .B0(n4055), .B1(n3897), .Y(n2021)
         );
  AOI22X1TS U3516 ( .A0(n4000), .A1(n3534), .B0(n4055), .B1(n3796), .Y(n1928)
         );
  AOI222XLTS U3517 ( .A0(n4219), .A1(n3574), .B0(n3558), .B1(n37), .C0(n3959), 
        .C1(n3551), .Y(n1929) );
  AOI222XLTS U3518 ( .A0(n3824), .A1(n752), .B0(n4545), .B1(n3377), .C0(n4170), 
        .C1(n3840), .Y(n1467) );
  AOI222XLTS U3519 ( .A0(n3820), .A1(n751), .B0(n4501), .B1(n3373), .C0(n4131), 
        .C1(n3838), .Y(n1441) );
  AOI222XLTS U3520 ( .A0(n3820), .A1(n750), .B0(n4495), .B1(n3373), .C0(n4125), 
        .C1(n3838), .Y(n1437) );
  AOI222XLTS U3521 ( .A0(n3820), .A1(n749), .B0(n4491), .B1(n3372), .C0(n4122), 
        .C1(n3838), .Y(n1435) );
  AOI222XLTS U3522 ( .A0(n3819), .A1(n748), .B0(n4461), .B1(n3370), .C0(n4095), 
        .C1(n3835), .Y(n1417) );
  AOI222XLTS U3523 ( .A0(n3819), .A1(n747), .B0(n4457), .B1(n3370), .C0(n4092), 
        .C1(n3835), .Y(n1415) );
  AOI222XLTS U3524 ( .A0(n3819), .A1(n746), .B0(n4454), .B1(n3370), .C0(n4089), 
        .C1(n3835), .Y(n1413) );
  AOI222XLTS U3525 ( .A0(n3825), .A1(n718), .B0(n4211), .B1(n3380), .C0(n4047), 
        .C1(n3840), .Y(n1993) );
  AOI222XLTS U3526 ( .A0(n3824), .A1(n717), .B0(n4208), .B1(n3381), .C0(n4044), 
        .C1(n3841), .Y(n1991) );
  AOI222XLTS U3527 ( .A0(n3824), .A1(n697), .B0(n4549), .B1(n3380), .C0(n4173), 
        .C1(n3840), .Y(n1469) );
  AOI222XLTS U3528 ( .A0(n3822), .A1(n696), .B0(n4525), .B1(n3375), .C0(n4152), 
        .C1(n3844), .Y(n1455) );
  AOI222XLTS U3529 ( .A0(n3822), .A1(n695), .B0(n4518), .B1(n3375), .C0(n4146), 
        .C1(n3845), .Y(n1451) );
  AOI222XLTS U3530 ( .A0(n3820), .A1(n694), .B0(n4498), .B1(n3373), .C0(n4128), 
        .C1(n3838), .Y(n1439) );
  AOI222XLTS U3531 ( .A0(n3819), .A1(n693), .B0(n4451), .B1(n3370), .C0(n4086), 
        .C1(n3835), .Y(n1411) );
  AOI22X1TS U3532 ( .A0(n4446), .A1(n3632), .B0(n4082), .B1(n3789), .Y(n1665)
         );
  AOI222XLTS U3533 ( .A0(n4349), .A1(n3762), .B0(n789), .B1(n3623), .C0(n4253), 
        .C1(n3610), .Y(n1666) );
  AOI22X1TS U3534 ( .A0(n4443), .A1(n3632), .B0(n4079), .B1(n3776), .Y(n1663)
         );
  AOI222XLTS U3535 ( .A0(n4346), .A1(n3762), .B0(n793), .B1(n3624), .C0(n4250), 
        .C1(n3603), .Y(n1664) );
  OAI33XLTS U3536 ( .A0(n4202), .A1(n455), .A2(n114), .B0(n998), .B1(n108), 
        .B2(n1838), .Y(n1835) );
  NAND2X1TS U3537 ( .A(readReady), .B(n3), .Y(n1889) );
  INVX2TS U3538 ( .A(n4202), .Y(n4201) );
  OAI22X1TS U3539 ( .A0(n1136), .A1(n1138), .B0(n5323), .B1(n1137), .Y(n2887)
         );
  OAI22X1TS U3540 ( .A0(n1135), .A1(n1136), .B0(n980), .B1(n1137), .Y(n2888)
         );
  CLKBUFX2TS U3541 ( .A(n5327), .Y(n980) );
  NAND2X1TS U3542 ( .A(n4194), .B(n917), .Y(n1862) );
  OAI33XLTS U3543 ( .A0(n4202), .A1(n917), .A2(n1837), .B0(n457), .B1(n930), 
        .B2(n1866), .Y(n1865) );
  AOI21X1TS U3544 ( .A0(n4195), .A1(n920), .B0(n1850), .Y(n1849) );
  NAND2X1TS U3545 ( .A(n462), .B(n980), .Y(n1918) );
  AOI221X1TS U3546 ( .A0(n1102), .A1(n4437), .B0(n1126), .B1(n4168), .C0(n2916), .Y(n2912) );
  OAI22X1TS U3547 ( .A0(n4440), .A1(n3115), .B0(n739), .B1(n3748), .Y(n2916)
         );
  AOI221X1TS U3548 ( .A0(n1102), .A1(n4434), .B0(n1126), .B1(n4165), .C0(n2910), .Y(n2906) );
  OAI22X1TS U3549 ( .A0(n4449), .A1(n3115), .B0(n738), .B1(n3748), .Y(n2910)
         );
  AOI221X1TS U3550 ( .A0(n1102), .A1(n4430), .B0(n1126), .B1(n4162), .C0(n2904), .Y(n2900) );
  OAI22X1TS U3551 ( .A0(n4458), .A1(n3115), .B0(n737), .B1(n3748), .Y(n2904)
         );
  AOI221X1TS U3552 ( .A0(n1103), .A1(n4427), .B0(n1125), .B1(n4159), .C0(n2898), .Y(n2894) );
  OAI22X1TS U3553 ( .A0(n4467), .A1(n3115), .B0(n736), .B1(n3749), .Y(n2898)
         );
  AOI221X1TS U3554 ( .A0(n1103), .A1(n4424), .B0(n1125), .B1(n4156), .C0(n2892), .Y(n2396) );
  OAI22X1TS U3555 ( .A0(n4476), .A1(n3114), .B0(n735), .B1(n3749), .Y(n2892)
         );
  AOI221X1TS U3556 ( .A0(n1103), .A1(n4421), .B0(n1125), .B1(n4153), .C0(n2394), .Y(n2390) );
  OAI22X1TS U3557 ( .A0(n4485), .A1(n3114), .B0(n715), .B1(n3749), .Y(n2394)
         );
  AOI221X1TS U3558 ( .A0(n1103), .A1(n4418), .B0(n1125), .B1(n4150), .C0(n2388), .Y(n2384) );
  OAI22X1TS U3559 ( .A0(n4494), .A1(n3114), .B0(n734), .B1(n3749), .Y(n2388)
         );
  AOI221X1TS U3560 ( .A0(n1104), .A1(n4415), .B0(n2103), .B1(n4147), .C0(n2382), .Y(n2378) );
  OAI22X1TS U3561 ( .A0(n4503), .A1(n3114), .B0(n714), .B1(n3750), .Y(n2382)
         );
  AOI221X1TS U3562 ( .A0(n1104), .A1(n4412), .B0(n1127), .B1(n4144), .C0(n2376), .Y(n2372) );
  OAI22X1TS U3563 ( .A0(n4512), .A1(n3113), .B0(n733), .B1(n3750), .Y(n2376)
         );
  AOI221X1TS U3564 ( .A0(n1104), .A1(n4409), .B0(n2103), .B1(n4141), .C0(n2370), .Y(n2366) );
  OAI22X1TS U3565 ( .A0(n4521), .A1(n3113), .B0(n732), .B1(n3750), .Y(n2370)
         );
  AOI221X1TS U3566 ( .A0(n1104), .A1(n4406), .B0(n1130), .B1(n4138), .C0(n2364), .Y(n2360) );
  OAI22X1TS U3567 ( .A0(n4530), .A1(n3113), .B0(n713), .B1(n3750), .Y(n2364)
         );
  AOI221X1TS U3568 ( .A0(n1105), .A1(n4403), .B0(n1128), .B1(n4135), .C0(n2358), .Y(n2354) );
  OAI22X1TS U3569 ( .A0(n4539), .A1(n3113), .B0(n731), .B1(n3759), .Y(n2358)
         );
  AOI221X1TS U3570 ( .A0(n1105), .A1(n4400), .B0(n1128), .B1(n4132), .C0(n2352), .Y(n2348) );
  OAI22X1TS U3571 ( .A0(n4548), .A1(n3112), .B0(n712), .B1(n3760), .Y(n2352)
         );
  AOI221X1TS U3572 ( .A0(n1105), .A1(n4397), .B0(n1129), .B1(n4129), .C0(n2346), .Y(n2342) );
  OAI22X1TS U3573 ( .A0(n4557), .A1(n3112), .B0(n730), .B1(n3758), .Y(n2346)
         );
  AOI221X1TS U3574 ( .A0(n1105), .A1(n4394), .B0(n1131), .B1(n4126), .C0(n2340), .Y(n2336) );
  OAI22X1TS U3575 ( .A0(n4566), .A1(n3112), .B0(n729), .B1(n1146), .Y(n2340)
         );
  AOI221X1TS U3576 ( .A0(n1106), .A1(n4391), .B0(n1127), .B1(n4123), .C0(n2334), .Y(n2330) );
  OAI22X1TS U3577 ( .A0(n4575), .A1(n3112), .B0(n711), .B1(n3757), .Y(n2334)
         );
  AOI221X1TS U3578 ( .A0(n1106), .A1(n4388), .B0(n1134), .B1(n4120), .C0(n2328), .Y(n2324) );
  OAI22X1TS U3579 ( .A0(n4584), .A1(n3111), .B0(n728), .B1(n3759), .Y(n2328)
         );
  AOI221X1TS U3580 ( .A0(n1106), .A1(n4385), .B0(n1134), .B1(n4117), .C0(n2322), .Y(n2318) );
  OAI22X1TS U3581 ( .A0(n4593), .A1(n3111), .B0(n710), .B1(n3760), .Y(n2322)
         );
  AOI221X1TS U3582 ( .A0(n1106), .A1(n4382), .B0(n1134), .B1(n4114), .C0(n2316), .Y(n2312) );
  OAI22X1TS U3583 ( .A0(n4602), .A1(n3111), .B0(n727), .B1(n3758), .Y(n2316)
         );
  AOI221X1TS U3584 ( .A0(n1107), .A1(n4379), .B0(n1124), .B1(n4111), .C0(n2310), .Y(n2306) );
  OAI22X1TS U3585 ( .A0(n4611), .A1(n3111), .B0(n726), .B1(n3756), .Y(n2310)
         );
  AOI221X1TS U3586 ( .A0(n1107), .A1(n4376), .B0(n1124), .B1(n4108), .C0(n2304), .Y(n2300) );
  OAI22X1TS U3587 ( .A0(n4620), .A1(n3110), .B0(n725), .B1(n3757), .Y(n2304)
         );
  AOI221X1TS U3588 ( .A0(n1107), .A1(n4373), .B0(n1124), .B1(n4105), .C0(n2298), .Y(n2294) );
  OAI22X1TS U3589 ( .A0(n4629), .A1(n3110), .B0(n724), .B1(n3759), .Y(n2298)
         );
  AOI221X1TS U3590 ( .A0(n1107), .A1(n4370), .B0(n1124), .B1(n4102), .C0(n2292), .Y(n2288) );
  OAI22X1TS U3591 ( .A0(n4638), .A1(n3110), .B0(n723), .B1(n3756), .Y(n2292)
         );
  AOI221X1TS U3592 ( .A0(n1108), .A1(n4364), .B0(n1123), .B1(n4096), .C0(n2280), .Y(n2276) );
  OAI22X1TS U3593 ( .A0(n4656), .A1(n3109), .B0(n722), .B1(n3751), .Y(n2280)
         );
  AOI221X1TS U3594 ( .A0(n1108), .A1(n4361), .B0(n1123), .B1(n4093), .C0(n2274), .Y(n2270) );
  OAI22X1TS U3595 ( .A0(n4665), .A1(n3109), .B0(n709), .B1(n3751), .Y(n2274)
         );
  AOI221X1TS U3596 ( .A0(n1108), .A1(n4358), .B0(n1123), .B1(n4090), .C0(n2268), .Y(n2264) );
  OAI22X1TS U3597 ( .A0(n4674), .A1(n3109), .B0(n708), .B1(n3751), .Y(n2268)
         );
  AOI221X1TS U3598 ( .A0(n1109), .A1(n4355), .B0(n1122), .B1(n4087), .C0(n2262), .Y(n2258) );
  OAI22X1TS U3599 ( .A0(n4683), .A1(n3108), .B0(n721), .B1(n3752), .Y(n2262)
         );
  AOI221X1TS U3600 ( .A0(n1109), .A1(n4352), .B0(n1122), .B1(n4084), .C0(n2256), .Y(n2252) );
  OAI22X1TS U3601 ( .A0(n4692), .A1(n3108), .B0(n707), .B1(n3752), .Y(n2256)
         );
  AOI221X1TS U3602 ( .A0(n1109), .A1(n4349), .B0(n1122), .B1(n4081), .C0(n2250), .Y(n2246) );
  OAI22X1TS U3603 ( .A0(n4701), .A1(n3108), .B0(n720), .B1(n3752), .Y(n2250)
         );
  AOI221X1TS U3604 ( .A0(n1109), .A1(n4346), .B0(n1122), .B1(n4078), .C0(n2244), .Y(n2240) );
  OAI22X1TS U3605 ( .A0(n4710), .A1(n3108), .B0(n719), .B1(n3752), .Y(n2244)
         );
  AOI221X1TS U3606 ( .A0(n1111), .A1(n3962), .B0(n1121), .B1(n4057), .C0(n2202), .Y(n2198) );
  OAI22X1TS U3607 ( .A0(n4723), .A1(n3107), .B0(n745), .B1(n3754), .Y(n2202)
         );
  AOI221X1TS U3608 ( .A0(n1111), .A1(n3959), .B0(n1121), .B1(n4054), .C0(n2196), .Y(n2192) );
  OAI22X1TS U3609 ( .A0(n4732), .A1(n3107), .B0(n744), .B1(n3754), .Y(n2196)
         );
  AOI221X1TS U3610 ( .A0(n1112), .A1(n3956), .B0(n1120), .B1(n4051), .C0(n2190), .Y(n2186) );
  OAI22X1TS U3611 ( .A0(n4741), .A1(n3110), .B0(n743), .B1(n3755), .Y(n2190)
         );
  AOI221X1TS U3612 ( .A0(n1112), .A1(n3953), .B0(n1120), .B1(n4048), .C0(n2184), .Y(n2180) );
  OAI22X1TS U3613 ( .A0(n4750), .A1(n3107), .B0(n716), .B1(n3755), .Y(n2184)
         );
  AOI221X1TS U3614 ( .A0(n1112), .A1(n3947), .B0(n1120), .B1(n4042), .C0(n2171), .Y(n2160) );
  OAI22X1TS U3615 ( .A0(n4768), .A1(n3107), .B0(n741), .B1(n3755), .Y(n2171)
         );
  AOI221X1TS U3616 ( .A0(n1108), .A1(n4367), .B0(n1123), .B1(n4099), .C0(n2286), .Y(n2282) );
  OAI22X1TS U3617 ( .A0(n4647), .A1(n3109), .B0(n4654), .B1(n3751), .Y(n2286)
         );
  INVX2TS U3618 ( .A(n2100), .Y(n911) );
  OAI221XLTS U3619 ( .A0(n4199), .A1(n2075), .B0(n159), .B1(n2073), .C0(n6257), 
        .Y(n2100) );
  AOI221X1TS U3620 ( .A0(n1102), .A1(n4441), .B0(n1126), .B1(n4171), .C0(n2922), .Y(n2918) );
  OAI22X1TS U3621 ( .A0(n4431), .A1(n3106), .B0(n740), .B1(n3748), .Y(n2922)
         );
  AOI221X1TS U3622 ( .A0(n1110), .A1(n4190), .B0(n1129), .B1(n4075), .C0(n2238), .Y(n2234) );
  OAI22X1TS U3623 ( .A0(n3106), .A1(n4719), .B0(n886), .B1(n3753), .Y(n2238)
         );
  AOI221X1TS U3624 ( .A0(n1110), .A1(n4187), .B0(n1131), .B1(n4072), .C0(n2232), .Y(n2228) );
  OAI22X1TS U3625 ( .A0(n3106), .A1(n4720), .B0(n887), .B1(n3753), .Y(n2232)
         );
  AOI221X1TS U3626 ( .A0(n1110), .A1(n4181), .B0(n1130), .B1(n4066), .C0(n2220), .Y(n2216) );
  OAI22X1TS U3627 ( .A0(n3105), .A1(n4721), .B0(n884), .B1(n3753), .Y(n2220)
         );
  AOI221X1TS U3628 ( .A0(n1111), .A1(n4178), .B0(n1121), .B1(n4063), .C0(n2214), .Y(n2210) );
  OAI22X1TS U3629 ( .A0(n3105), .A1(n4722), .B0(n883), .B1(n3754), .Y(n2214)
         );
  AOI221X1TS U3630 ( .A0(n1112), .A1(n3950), .B0(n1120), .B1(n4045), .C0(n2178), .Y(n2174) );
  OAI22X1TS U3631 ( .A0(n4759), .A1(n3106), .B0(n742), .B1(n3755), .Y(n2178)
         );
  AOI221X1TS U3632 ( .A0(n1110), .A1(n4184), .B0(n1131), .B1(n4069), .C0(n2226), .Y(n2222) );
  OAI22X1TS U3633 ( .A0(n3105), .A1(n4846), .B0(n885), .B1(n3753), .Y(n2226)
         );
  AOI221X1TS U3634 ( .A0(n1111), .A1(n4175), .B0(n1121), .B1(n4060), .C0(n2208), .Y(n2204) );
  OAI22X1TS U3635 ( .A0(n3105), .A1(n4845), .B0(n882), .B1(n3754), .Y(n2208)
         );
  NAND4X1TS U3636 ( .A(n2917), .B(n2918), .C(n2919), .D(n2920), .Y(n2397) );
  AOI222XLTS U3637 ( .A0(n1043), .A1(n760), .B0(n1016), .B1(n2983), .C0(n1002), 
        .C1(n2982), .Y(n2919) );
  AOI221X1TS U3638 ( .A0(n1099), .A1(n3061), .B0(n1085), .B1(n697), .C0(n2921), 
        .Y(n2920) );
  AOI222XLTS U3639 ( .A0(n2158), .A1(n4549), .B0(n2970), .B1(n4342), .C0(n987), 
        .C1(cacheDataOut[31]), .Y(n2917) );
  NAND4X1TS U3640 ( .A(n2911), .B(n2912), .C(n2913), .D(n2914), .Y(n2398) );
  AOI222XLTS U3641 ( .A0(n1043), .A1(n759), .B0(n1016), .B1(n2985), .C0(n1002), 
        .C1(n2984), .Y(n2913) );
  AOI221X1TS U3642 ( .A0(n1098), .A1(n3062), .B0(n1087), .B1(n752), .C0(n2915), 
        .Y(n2914) );
  AOI222XLTS U3643 ( .A0(n2956), .A1(n4545), .B0(n3059), .B1(n4339), .C0(n987), 
        .C1(cacheDataOut[30]), .Y(n2911) );
  NAND4X1TS U3644 ( .A(n2905), .B(n2906), .C(n2907), .D(n2908), .Y(n2399) );
  AOI222XLTS U3645 ( .A0(n1044), .A1(n758), .B0(n1016), .B1(n2987), .C0(n1002), 
        .C1(n2986), .Y(n2907) );
  AOI221X1TS U3646 ( .A0(n1100), .A1(n3063), .B0(n1085), .B1(n949), .C0(n2909), 
        .Y(n2908) );
  AOI222XLTS U3647 ( .A0(n2098), .A1(n4542), .B0(n3059), .B1(n4336), .C0(n987), 
        .C1(cacheDataOut[29]), .Y(n2905) );
  NAND4X1TS U3648 ( .A(n2899), .B(n2900), .C(n2901), .D(n2902), .Y(n2400) );
  AOI222XLTS U3649 ( .A0(n2168), .A1(n706), .B0(n1016), .B1(n2989), .C0(n1002), 
        .C1(n2988), .Y(n2901) );
  AOI221X1TS U3650 ( .A0(n1101), .A1(n3064), .B0(n2164), .B1(n950), .C0(n2903), 
        .Y(n2902) );
  AOI222XLTS U3651 ( .A0(n2966), .A1(n4538), .B0(n3059), .B1(n4333), .C0(n987), 
        .C1(cacheDataOut[28]), .Y(n2899) );
  NAND4X1TS U3652 ( .A(n2893), .B(n2894), .C(n2895), .D(n2896), .Y(n2401) );
  AOI222XLTS U3653 ( .A0(n1030), .A1(n705), .B0(n1029), .B1(n2991), .C0(n1012), 
        .C1(n2990), .Y(n2895) );
  AOI221X1TS U3654 ( .A0(n1088), .A1(n3065), .B0(n1073), .B1(n964), .C0(n2897), 
        .Y(n2896) );
  AOI222XLTS U3655 ( .A0(n2967), .A1(n4535), .B0(n3059), .B1(n4330), .C0(n999), 
        .C1(cacheDataOut[27]), .Y(n2893) );
  NAND4X1TS U3656 ( .A(n2395), .B(n2396), .C(n2449), .D(n2890), .Y(n2402) );
  AOI222XLTS U3657 ( .A0(n1030), .A1(n757), .B0(n1028), .B1(n2993), .C0(n1009), 
        .C1(n2992), .Y(n2449) );
  AOI221X1TS U3658 ( .A0(n1088), .A1(n3066), .B0(n1073), .B1(n951), .C0(n2891), 
        .Y(n2890) );
  AOI222XLTS U3659 ( .A0(n2967), .A1(n4532), .B0(n3100), .B1(n4327), .C0(n997), 
        .C1(cacheDataOut[26]), .Y(n2395) );
  NAND4X1TS U3660 ( .A(n2389), .B(n2390), .C(n2391), .D(n2392), .Y(n2403) );
  AOI222XLTS U3661 ( .A0(n1030), .A1(n756), .B0(n1027), .B1(n2995), .C0(n1014), 
        .C1(n2994), .Y(n2391) );
  AOI221X1TS U3662 ( .A0(n1088), .A1(n3067), .B0(n1073), .B1(n952), .C0(n2393), 
        .Y(n2392) );
  AOI222XLTS U3663 ( .A0(n2098), .A1(n4528), .B0(n3101), .B1(n4324), .C0(n1001), .C1(cacheDataOut[25]), .Y(n2389) );
  NAND4X1TS U3664 ( .A(n2383), .B(n2384), .C(n2385), .D(n2386), .Y(n2404) );
  AOI222XLTS U3665 ( .A0(n1030), .A1(n755), .B0(n1028), .B1(n2997), .C0(n1009), 
        .C1(n2996), .Y(n2385) );
  AOI221X1TS U3666 ( .A0(n1088), .A1(n3068), .B0(n1073), .B1(n696), .C0(n2387), 
        .Y(n2386) );
  AOI222XLTS U3667 ( .A0(n2098), .A1(n4525), .B0(n3102), .B1(n4321), .C0(n996), 
        .C1(cacheDataOut[24]), .Y(n2383) );
  NAND4X1TS U3668 ( .A(n2377), .B(n2378), .C(n2379), .D(n2380), .Y(n2405) );
  AOI222XLTS U3669 ( .A0(n1042), .A1(n704), .B0(n1017), .B1(n2999), .C0(n1012), 
        .C1(n2998), .Y(n2379) );
  AOI221X1TS U3670 ( .A0(n1099), .A1(n3069), .B0(n1084), .B1(n953), .C0(n2381), 
        .Y(n2380) );
  AOI222XLTS U3671 ( .A0(n1155), .A1(n4522), .B0(n3060), .B1(n4318), .C0(n996), 
        .C1(cacheDataOut[23]), .Y(n2377) );
  NAND4X1TS U3672 ( .A(n2371), .B(n2372), .C(n2373), .D(n2374), .Y(n2406) );
  AOI222XLTS U3673 ( .A0(n1040), .A1(n754), .B0(n1017), .B1(n3001), .C0(n1012), 
        .C1(n3000), .Y(n2373) );
  AOI221X1TS U3674 ( .A0(n1096), .A1(n3070), .B0(n1082), .B1(n695), .C0(n2375), 
        .Y(n2374) );
  AOI222XLTS U3675 ( .A0(n1155), .A1(n4518), .B0(n3104), .B1(n4315), .C0(n1000), .C1(cacheDataOut[22]), .Y(n2371) );
  NAND4X1TS U3676 ( .A(n2365), .B(n2366), .C(n2367), .D(n2368), .Y(n2407) );
  AOI222XLTS U3677 ( .A0(n1039), .A1(n753), .B0(n1017), .B1(n3003), .C0(n1011), 
        .C1(n3002), .Y(n2367) );
  AOI221X1TS U3678 ( .A0(n1095), .A1(n3071), .B0(n1081), .B1(n954), .C0(n2369), 
        .Y(n2368) );
  AOI222XLTS U3679 ( .A0(n1155), .A1(n4515), .B0(n3060), .B1(n4312), .C0(n999), 
        .C1(cacheDataOut[21]), .Y(n2365) );
  NAND4X1TS U3680 ( .A(n2359), .B(n2360), .C(n2361), .D(n2362), .Y(n2408) );
  AOI222XLTS U3681 ( .A0(n1038), .A1(n703), .B0(n1017), .B1(n3005), .C0(n1010), 
        .C1(n3004), .Y(n2361) );
  AOI221X1TS U3682 ( .A0(n1099), .A1(n3072), .B0(n1080), .B1(n955), .C0(n2363), 
        .Y(n2362) );
  AOI222XLTS U3683 ( .A0(n1155), .A1(n4511), .B0(n3104), .B1(n4309), .C0(n1000), .C1(cacheDataOut[20]), .Y(n2359) );
  NAND4X1TS U3684 ( .A(n2353), .B(n2354), .C(n2355), .D(n2356), .Y(n2409) );
  AOI222XLTS U3685 ( .A0(n1041), .A1(n46), .B0(n1027), .B1(n3007), .C0(n1014), 
        .C1(n3006), .Y(n2355) );
  AOI221X1TS U3686 ( .A0(n1098), .A1(n3073), .B0(n1083), .B1(n956), .C0(n2357), 
        .Y(n2356) );
  AOI222XLTS U3687 ( .A0(n1199), .A1(n4508), .B0(n3102), .B1(n4306), .C0(n988), 
        .C1(cacheDataOut[19]), .Y(n2353) );
  NAND4X1TS U3688 ( .A(n2347), .B(n2348), .C(n2349), .D(n2350), .Y(n2410) );
  AOI222XLTS U3689 ( .A0(n1041), .A1(n47), .B0(n1024), .B1(n3009), .C0(n1011), 
        .C1(n3008), .Y(n2349) );
  AOI221X1TS U3690 ( .A0(n1098), .A1(n3074), .B0(n1083), .B1(n957), .C0(n2351), 
        .Y(n2350) );
  AOI222XLTS U3691 ( .A0(n1199), .A1(n4505), .B0(n3058), .B1(n4303), .C0(n988), 
        .C1(cacheDataOut[18]), .Y(n2347) );
  NAND4X1TS U3692 ( .A(n2341), .B(n2342), .C(n2343), .D(n2344), .Y(n2411) );
  AOI222XLTS U3693 ( .A0(n1041), .A1(n48), .B0(n1024), .B1(n3011), .C0(n1015), 
        .C1(n3010), .Y(n2343) );
  AOI221X1TS U3694 ( .A0(n1100), .A1(n3075), .B0(n1083), .B1(n751), .C0(n2345), 
        .Y(n2344) );
  AOI222XLTS U3695 ( .A0(n1199), .A1(n4501), .B0(n3058), .B1(n4300), .C0(n988), 
        .C1(cacheDataOut[17]), .Y(n2341) );
  NAND4X1TS U3696 ( .A(n2335), .B(n2336), .C(n2337), .D(n2338), .Y(n2412) );
  AOI222XLTS U3697 ( .A0(n1042), .A1(n49), .B0(n1026), .B1(n3013), .C0(n1012), 
        .C1(n3012), .Y(n2337) );
  AOI221X1TS U3698 ( .A0(n1097), .A1(n3076), .B0(n1084), .B1(n694), .C0(n2339), 
        .Y(n2338) );
  AOI222XLTS U3699 ( .A0(n1199), .A1(n4498), .B0(n3058), .B1(n4297), .C0(n988), 
        .C1(cacheDataOut[16]), .Y(n2335) );
  NAND4X1TS U3700 ( .A(n2329), .B(n2330), .C(n2331), .D(n2332), .Y(n2413) );
  AOI222XLTS U3701 ( .A0(n1041), .A1(n50), .B0(n1027), .B1(n3015), .C0(n1010), 
        .C1(n3014), .Y(n2331) );
  AOI221X1TS U3702 ( .A0(n1098), .A1(n3077), .B0(n1083), .B1(n750), .C0(n2333), 
        .Y(n2332) );
  AOI222XLTS U3703 ( .A0(n1215), .A1(n4495), .B0(n3058), .B1(n4294), .C0(n989), 
        .C1(cacheDataOut[15]), .Y(n2329) );
  NAND4X1TS U3704 ( .A(n2323), .B(n2324), .C(n2325), .D(n2326), .Y(n2414) );
  AOI222XLTS U3705 ( .A0(n1040), .A1(n51), .B0(n1028), .B1(n3017), .C0(n1013), 
        .C1(n3016), .Y(n2325) );
  AOI221X1TS U3706 ( .A0(n1097), .A1(n3078), .B0(n1082), .B1(n749), .C0(n2327), 
        .Y(n2326) );
  AOI222XLTS U3707 ( .A0(n1215), .A1(n4491), .B0(n3099), .B1(n4291), .C0(n989), 
        .C1(cacheDataOut[14]), .Y(n2323) );
  NAND4X1TS U3708 ( .A(n2317), .B(n2318), .C(n2319), .D(n2320), .Y(n2415) );
  AOI222XLTS U3709 ( .A0(n1039), .A1(n52), .B0(n1026), .B1(n3019), .C0(n1013), 
        .C1(n3018), .Y(n2319) );
  AOI221X1TS U3710 ( .A0(n1096), .A1(n3079), .B0(n1081), .B1(n958), .C0(n2321), 
        .Y(n2320) );
  AOI222XLTS U3711 ( .A0(n1215), .A1(n4488), .B0(n3099), .B1(n4288), .C0(n989), 
        .C1(cacheDataOut[13]), .Y(n2317) );
  NAND4X1TS U3712 ( .A(n2311), .B(n2312), .C(n2313), .D(n2314), .Y(n2416) );
  AOI222XLTS U3713 ( .A0(n1038), .A1(n53), .B0(n1025), .B1(n3021), .C0(n1013), 
        .C1(n3020), .Y(n2313) );
  AOI221X1TS U3714 ( .A0(n1095), .A1(n3080), .B0(n1080), .B1(n959), .C0(n2315), 
        .Y(n2314) );
  AOI222XLTS U3715 ( .A0(n1215), .A1(n4484), .B0(n3101), .B1(n4285), .C0(n989), 
        .C1(cacheDataOut[12]), .Y(n2311) );
  NAND4X1TS U3716 ( .A(n2305), .B(n2306), .C(n2307), .D(n2308), .Y(n2417) );
  AOI222XLTS U3717 ( .A0(n1032), .A1(n54), .B0(n1018), .B1(n3023), .C0(n1003), 
        .C1(n3022), .Y(n2307) );
  AOI221X1TS U3718 ( .A0(n1089), .A1(n3081), .B0(n1074), .B1(n960), .C0(n2309), 
        .Y(n2308) );
  AOI222XLTS U3719 ( .A0(n1246), .A1(n4481), .B0(n3060), .B1(n4282), .C0(n990), 
        .C1(cacheDataOut[11]), .Y(n2305) );
  NAND4X1TS U3720 ( .A(n2299), .B(n2300), .C(n2301), .D(n2302), .Y(n2418) );
  AOI222XLTS U3721 ( .A0(n1032), .A1(n55), .B0(n1018), .B1(n3025), .C0(n1003), 
        .C1(n3024), .Y(n2301) );
  AOI221X1TS U3722 ( .A0(n1089), .A1(n3082), .B0(n1074), .B1(n965), .C0(n2303), 
        .Y(n2302) );
  AOI222XLTS U3723 ( .A0(n1246), .A1(n4478), .B0(n2975), .B1(n4279), .C0(n990), 
        .C1(cacheDataOut[10]), .Y(n2299) );
  NAND4X1TS U3724 ( .A(n2293), .B(n2294), .C(n2295), .D(n2296), .Y(n2419) );
  AOI222XLTS U3725 ( .A0(n1032), .A1(n702), .B0(n1018), .B1(n3027), .C0(n1003), 
        .C1(n3026), .Y(n2295) );
  AOI221X1TS U3726 ( .A0(n1089), .A1(n3083), .B0(n1074), .B1(n961), .C0(n2297), 
        .Y(n2296) );
  AOI222XLTS U3727 ( .A0(n1246), .A1(n4474), .B0(n2975), .B1(n4276), .C0(n990), 
        .C1(cacheDataOut[9]), .Y(n2293) );
  NAND4X1TS U3728 ( .A(n2287), .B(n2288), .C(n2289), .D(n2290), .Y(n2420) );
  AOI222XLTS U3729 ( .A0(n1032), .A1(n56), .B0(n1018), .B1(n3029), .C0(n1003), 
        .C1(n3028), .Y(n2289) );
  AOI221X1TS U3730 ( .A0(n1089), .A1(n3084), .B0(n1074), .B1(n962), .C0(n2291), 
        .Y(n2290) );
  AOI222XLTS U3731 ( .A0(n1246), .A1(n4471), .B0(n2975), .B1(n4273), .C0(n990), 
        .C1(cacheDataOut[8]), .Y(n2287) );
  NAND4X1TS U3732 ( .A(n2281), .B(n2282), .C(n2283), .D(n2284), .Y(n2421) );
  AOI222XLTS U3733 ( .A0(n1033), .A1(n57), .B0(n1019), .B1(n3031), .C0(n1004), 
        .C1(n3030), .Y(n2283) );
  AOI221X1TS U3734 ( .A0(n1090), .A1(n3085), .B0(n1075), .B1(n963), .C0(n2285), 
        .Y(n2284) );
  AOI222XLTS U3735 ( .A0(n2956), .A1(n4468), .B0(n2975), .B1(n4270), .C0(n991), 
        .C1(cacheDataOut[7]), .Y(n2281) );
  NAND4X1TS U3736 ( .A(n2275), .B(n2276), .C(n2277), .D(n2278), .Y(n2422) );
  AOI222XLTS U3737 ( .A0(n1033), .A1(n58), .B0(n1019), .B1(n3033), .C0(n1004), 
        .C1(n3032), .Y(n2277) );
  AOI221X1TS U3738 ( .A0(n1090), .A1(n3086), .B0(n1075), .B1(n966), .C0(n2279), 
        .Y(n2278) );
  AOI222XLTS U3739 ( .A0(n2956), .A1(n4464), .B0(n2974), .B1(n4267), .C0(n991), 
        .C1(cacheDataOut[6]), .Y(n2275) );
  NAND4X1TS U3740 ( .A(n2269), .B(n2270), .C(n2271), .D(n2272), .Y(n2423) );
  AOI222XLTS U3741 ( .A0(n1033), .A1(n701), .B0(n1019), .B1(n3035), .C0(n1004), 
        .C1(n3034), .Y(n2271) );
  AOI221X1TS U3742 ( .A0(n1090), .A1(n3087), .B0(n1075), .B1(n748), .C0(n2273), 
        .Y(n2272) );
  AOI222XLTS U3743 ( .A0(n2956), .A1(n4461), .B0(n2974), .B1(n4264), .C0(n991), 
        .C1(cacheDataOut[5]), .Y(n2269) );
  NAND4X1TS U3744 ( .A(n2263), .B(n2264), .C(n2265), .D(n2266), .Y(n2424) );
  AOI222XLTS U3745 ( .A0(n1033), .A1(n59), .B0(n1019), .B1(n3037), .C0(n1004), 
        .C1(n3036), .Y(n2265) );
  AOI221X1TS U3746 ( .A0(n1090), .A1(n3088), .B0(n1075), .B1(n747), .C0(n2267), 
        .Y(n2266) );
  AOI222XLTS U3747 ( .A0(n2955), .A1(n4457), .B0(n2974), .B1(n4261), .C0(n991), 
        .C1(cacheDataOut[4]), .Y(n2263) );
  NAND4X1TS U3748 ( .A(n2257), .B(n2258), .C(n2259), .D(n2260), .Y(n2425) );
  AOI222XLTS U3749 ( .A0(n1034), .A1(n60), .B0(n1020), .B1(n3039), .C0(n1005), 
        .C1(n3038), .Y(n2259) );
  AOI221X1TS U3750 ( .A0(n1091), .A1(n3089), .B0(n1076), .B1(n746), .C0(n2261), 
        .Y(n2260) );
  AOI222XLTS U3751 ( .A0(n2965), .A1(n4454), .B0(n2973), .B1(n4258), .C0(n992), 
        .C1(cacheDataOut[3]), .Y(n2257) );
  NAND4X1TS U3752 ( .A(n2251), .B(n2252), .C(n2253), .D(n2254), .Y(n2426) );
  AOI222XLTS U3753 ( .A0(n1034), .A1(n700), .B0(n1020), .B1(n3041), .C0(n1005), 
        .C1(n3040), .Y(n2253) );
  AOI221X1TS U3754 ( .A0(n1091), .A1(n3090), .B0(n1076), .B1(n693), .C0(n2255), 
        .Y(n2254) );
  AOI222XLTS U3755 ( .A0(n2964), .A1(n4451), .B0(n2973), .B1(n4255), .C0(n992), 
        .C1(cacheDataOut[2]), .Y(n2251) );
  NAND4X1TS U3756 ( .A(n2245), .B(n2246), .C(n2247), .D(n2248), .Y(n2427) );
  AOI222XLTS U3757 ( .A0(n1034), .A1(n699), .B0(n1020), .B1(n3043), .C0(n1005), 
        .C1(n3042), .Y(n2247) );
  AOI221X1TS U3758 ( .A0(n1091), .A1(n3091), .B0(n1076), .B1(n943), .C0(n2249), 
        .Y(n2248) );
  AOI222XLTS U3759 ( .A0(n2965), .A1(n4447), .B0(n2973), .B1(n4252), .C0(n992), 
        .C1(cacheDataOut[1]), .Y(n2245) );
  NAND4X1TS U3760 ( .A(n2239), .B(n2240), .C(n2241), .D(n2242), .Y(n2428) );
  AOI222XLTS U3761 ( .A0(n1034), .A1(n698), .B0(n1020), .B1(n3045), .C0(n1005), 
        .C1(n3044), .Y(n2241) );
  AOI221X1TS U3762 ( .A0(n1091), .A1(n3092), .B0(n1076), .B1(n944), .C0(n2243), 
        .Y(n2242) );
  AOI222XLTS U3763 ( .A0(n2964), .A1(n4444), .B0(n2973), .B1(n4249), .C0(n992), 
        .C1(cacheDataOut[0]), .Y(n2239) );
  NAND4X1TS U3764 ( .A(n2233), .B(n2234), .C(n2235), .D(n2236), .Y(n2429) );
  AOI222XLTS U3765 ( .A0(n1035), .A1(\requesterAddressbuffer[0][5] ), .B0(
        n1021), .B1(\requesterAddressbuffer[6][5] ), .C0(n1006), .C1(n2976), 
        .Y(n2235) );
  AOI221X1TS U3766 ( .A0(n1092), .A1(n2958), .B0(n1077), .B1(
        \requesterAddressbuffer[2][5] ), .C0(n2237), .Y(n2236) );
  AOI222XLTS U3767 ( .A0(n1662), .A1(n4568), .B0(n2972), .B1(n4040), .C0(n993), 
        .C1(readRequesterAddress[5]), .Y(n2233) );
  NAND4X1TS U3768 ( .A(n2227), .B(n2228), .C(n2229), .D(n2230), .Y(n2430) );
  AOI222XLTS U3769 ( .A0(n1035), .A1(\requesterAddressbuffer[0][4] ), .B0(
        n1021), .B1(\requesterAddressbuffer[6][4] ), .C0(n1006), .C1(n2977), 
        .Y(n2229) );
  AOI221X1TS U3770 ( .A0(n1092), .A1(n2959), .B0(n1077), .B1(
        \requesterAddressbuffer[2][4] ), .C0(n2231), .Y(n2230) );
  AOI222XLTS U3771 ( .A0(n1662), .A1(n4564), .B0(n2972), .B1(n4037), .C0(n993), 
        .C1(readRequesterAddress[4]), .Y(n2227) );
  NAND4X1TS U3772 ( .A(n2215), .B(n2216), .C(n2217), .D(n2218), .Y(n2432) );
  AOI222XLTS U3773 ( .A0(n1035), .A1(\requesterAddressbuffer[0][2] ), .B0(
        n1021), .B1(\requesterAddressbuffer[6][2] ), .C0(n1006), .C1(n2978), 
        .Y(n2217) );
  AOI221X1TS U3774 ( .A0(n1092), .A1(n2960), .B0(n1077), .B1(
        \requesterAddressbuffer[2][2] ), .C0(n2219), .Y(n2218) );
  AOI222XLTS U3775 ( .A0(n1662), .A1(n4558), .B0(n2972), .B1(n4031), .C0(n993), 
        .C1(readRequesterAddress[2]), .Y(n2215) );
  NAND4X1TS U3776 ( .A(n2209), .B(n2210), .C(n2211), .D(n2212), .Y(n2433) );
  AOI222XLTS U3777 ( .A0(n1036), .A1(\requesterAddressbuffer[0][1] ), .B0(
        n1022), .B1(\requesterAddressbuffer[6][1] ), .C0(n1007), .C1(n2979), 
        .Y(n2211) );
  AOI221X1TS U3778 ( .A0(n1093), .A1(n2961), .B0(n1078), .B1(
        \requesterAddressbuffer[2][1] ), .C0(n2213), .Y(n2212) );
  AOI222XLTS U3779 ( .A0(n1794), .A1(n4554), .B0(n2971), .B1(n4028), .C0(n994), 
        .C1(readRequesterAddress[1]), .Y(n2209) );
  NAND4X1TS U3780 ( .A(n2197), .B(n2198), .C(n2199), .D(n2200), .Y(n2435) );
  AOI222XLTS U3781 ( .A0(n1036), .A1(n764), .B0(n1022), .B1(n3047), .C0(n1007), 
        .C1(n3046), .Y(n2199) );
  AOI221X1TS U3782 ( .A0(n1093), .A1(n3093), .B0(n1078), .B1(n946), .C0(n2201), 
        .Y(n2200) );
  AOI222XLTS U3783 ( .A0(n1794), .A1(n4223), .B0(n2971), .B1(n4004), .C0(n994), 
        .C1(readRequesterAddress[5]), .Y(n2197) );
  NAND4X1TS U3784 ( .A(n2191), .B(n2192), .C(n2193), .D(n2194), .Y(n2436) );
  AOI222XLTS U3785 ( .A0(n1036), .A1(n88), .B0(n1022), .B1(n3049), .C0(n1007), 
        .C1(n3048), .Y(n2193) );
  AOI221X1TS U3786 ( .A0(n1093), .A1(n3094), .B0(n1078), .B1(n947), .C0(n2195), 
        .Y(n2194) );
  AOI222XLTS U3787 ( .A0(n1794), .A1(n4220), .B0(n2971), .B1(n4001), .C0(n994), 
        .C1(readRequesterAddress[4]), .Y(n2191) );
  NAND4X1TS U3788 ( .A(n2185), .B(n2186), .C(n2187), .D(n2188), .Y(n2437) );
  AOI222XLTS U3789 ( .A0(n1037), .A1(n763), .B0(n1023), .B1(n3051), .C0(n1008), 
        .C1(n3050), .Y(n2187) );
  AOI221X1TS U3790 ( .A0(n1094), .A1(n3095), .B0(n1079), .B1(n948), .C0(n2189), 
        .Y(n2188) );
  AOI222XLTS U3791 ( .A0(n1846), .A1(n4217), .B0(n2974), .B1(n3998), .C0(n995), 
        .C1(readRequesterAddress[3]), .Y(n2185) );
  NAND4X1TS U3792 ( .A(n2179), .B(n2180), .C(n2181), .D(n2182), .Y(n2438) );
  AOI222XLTS U3793 ( .A0(n1037), .A1(n762), .B0(n1023), .B1(n3053), .C0(n1008), 
        .C1(n3052), .Y(n2181) );
  AOI221X1TS U3794 ( .A0(n1094), .A1(n3096), .B0(n1079), .B1(n945), .C0(n2183), 
        .Y(n2182) );
  AOI222XLTS U3795 ( .A0(n1846), .A1(n4214), .B0(n2970), .B1(n3995), .C0(n995), 
        .C1(readRequesterAddress[2]), .Y(n2179) );
  NAND4X1TS U3796 ( .A(n2173), .B(n2174), .C(n2175), .D(n2176), .Y(n2439) );
  AOI222XLTS U3797 ( .A0(n1037), .A1(n761), .B0(n1023), .B1(n3055), .C0(n1008), 
        .C1(n3054), .Y(n2175) );
  AOI221X1TS U3798 ( .A0(n1094), .A1(n3097), .B0(n1079), .B1(n718), .C0(n2177), 
        .Y(n2176) );
  AOI222XLTS U3799 ( .A0(n1846), .A1(n4211), .B0(n2970), .B1(n3992), .C0(n995), 
        .C1(readRequesterAddress[1]), .Y(n2173) );
  NAND4X1TS U3800 ( .A(n2159), .B(n2160), .C(n2161), .D(n2162), .Y(n2440) );
  AOI222XLTS U3801 ( .A0(n1037), .A1(n89), .B0(n1023), .B1(n3057), .C0(n1008), 
        .C1(n3056), .Y(n2161) );
  AOI221X1TS U3802 ( .A0(n1094), .A1(n3098), .B0(n1079), .B1(n717), .C0(n2165), 
        .Y(n2162) );
  AOI222XLTS U3803 ( .A0(n1846), .A1(n4208), .B0(n2970), .B1(n3989), .C0(n995), 
        .C1(readRequesterAddress[0]), .Y(n2159) );
  NAND4X1TS U3804 ( .A(n2221), .B(n2222), .C(n2223), .D(n2224), .Y(n2431) );
  AOI222XLTS U3805 ( .A0(n1035), .A1(\requesterAddressbuffer[0][3] ), .B0(
        n1021), .B1(\requesterAddressbuffer[6][3] ), .C0(n1006), .C1(n2980), 
        .Y(n2223) );
  AOI221X1TS U3806 ( .A0(n1092), .A1(n2962), .B0(n1077), .B1(
        \requesterAddressbuffer[2][3] ), .C0(n2225), .Y(n2224) );
  AOI222XLTS U3807 ( .A0(n1662), .A1(n4561), .B0(n2972), .B1(n4034), .C0(n993), 
        .C1(readRequesterAddress[3]), .Y(n2221) );
  NAND4X1TS U3808 ( .A(n2203), .B(n2204), .C(n2205), .D(n2206), .Y(n2434) );
  AOI222XLTS U3809 ( .A0(n1036), .A1(\requesterAddressbuffer[0][0] ), .B0(
        n1022), .B1(\requesterAddressbuffer[6][0] ), .C0(n1007), .C1(n2981), 
        .Y(n2205) );
  AOI221X1TS U3810 ( .A0(n1093), .A1(n2963), .B0(n1078), .B1(
        \requesterAddressbuffer[2][0] ), .C0(n2207), .Y(n2206) );
  AOI222XLTS U3811 ( .A0(n1794), .A1(n4551), .B0(n2971), .B1(n4025), .C0(n994), 
        .C1(readRequesterAddress[0]), .Y(n2203) );
  OAI21X1TS U3812 ( .A0(n153), .A1(n911), .B0(n680), .Y(n2091) );
  INVX2TS U3813 ( .A(n2092), .Y(n680) );
  OAI33XLTS U3814 ( .A0(n4841), .A1(n2067), .A2(n2068), .B0(n2093), .B1(n4571), 
        .B2(n911), .Y(n2092) );
  NOR4XLTS U3815 ( .A(n2094), .B(n2095), .C(n2096), .D(n2097), .Y(n2093) );
  INVX2TS U3816 ( .A(writeIn_NORTH), .Y(n984) );
  NOR4BX1TS U3817 ( .AN(n2078), .B(n2079), .C(n2080), .D(n2081), .Y(n2069) );
  OAI31X1TS U3818 ( .A0(n2071), .A1(n459), .A2(n2072), .B0(n4573), .Y(n2070)
         );
  OAI22X1TS U3819 ( .A0(n2085), .A1(n769), .B0(n2086), .B1(n677), .Y(n2079) );
  OAI211X1TS U3820 ( .A0(n3987), .A1(n1113), .B0(n2151), .C0(n2152), .Y(n2441)
         );
  AOI22X1TS U3821 ( .A0(n478), .A1(n2153), .B0(n3117), .B1(
        destinationAddressOut[13]), .Y(n2151) );
  AOI222XLTS U3822 ( .A0(n1919), .A1(n4247), .B0(n1119), .B1(
        destinationAddressIn_NORTH[13]), .C0(n2969), .C1(n4022), .Y(n2152) );
  NAND4X1TS U3823 ( .A(n2154), .B(n2155), .C(n2156), .D(n2157), .Y(n2153) );
  OAI211X1TS U3824 ( .A0(n3984), .A1(n1113), .B0(n2144), .C0(n2145), .Y(n2442)
         );
  AOI22X1TS U3825 ( .A0(n480), .A1(n2146), .B0(n3117), .B1(
        destinationAddressOut[12]), .Y(n2144) );
  AOI222XLTS U3826 ( .A0(n1919), .A1(n4244), .B0(n1119), .B1(
        destinationAddressIn_NORTH[12]), .C0(n2969), .C1(n4020), .Y(n2145) );
  NAND4X1TS U3827 ( .A(n2147), .B(n2148), .C(n2149), .D(n2150), .Y(n2146) );
  OAI211X1TS U3828 ( .A0(n3981), .A1(n1113), .B0(n2137), .C0(n2138), .Y(n2443)
         );
  AOI22X1TS U3829 ( .A0(n479), .A1(n2139), .B0(n3117), .B1(
        destinationAddressOut[11]), .Y(n2137) );
  AOI222XLTS U3830 ( .A0(n1919), .A1(n4241), .B0(n1119), .B1(
        destinationAddressIn_NORTH[11]), .C0(n2969), .C1(n4018), .Y(n2138) );
  NAND4X1TS U3831 ( .A(n2140), .B(n2141), .C(n2142), .D(n2143), .Y(n2139) );
  OAI211X1TS U3832 ( .A0(n3978), .A1(n1114), .B0(n2130), .C0(n2131), .Y(n2444)
         );
  AOI22X1TS U3833 ( .A0(n480), .A1(n2132), .B0(n3117), .B1(
        destinationAddressOut[10]), .Y(n2130) );
  AOI222XLTS U3834 ( .A0(n1919), .A1(n4238), .B0(n1119), .B1(
        destinationAddressIn_NORTH[10]), .C0(n2968), .C1(
        destinationAddressIn_WEST[10]), .Y(n2131) );
  NAND4X1TS U3835 ( .A(n2133), .B(n2134), .C(n2135), .D(n2136), .Y(n2132) );
  OAI211X1TS U3836 ( .A0(n3975), .A1(n1114), .B0(n2123), .C0(n2124), .Y(n2445)
         );
  AOI22X1TS U3837 ( .A0(n479), .A1(n2125), .B0(n3118), .B1(
        destinationAddressOut[9]), .Y(n2123) );
  AOI222XLTS U3838 ( .A0(n1988), .A1(n4235), .B0(n1118), .B1(
        destinationAddressIn_NORTH[9]), .C0(n2969), .C1(
        destinationAddressIn_WEST[9]), .Y(n2124) );
  NAND4X1TS U3839 ( .A(n2126), .B(n2127), .C(n2128), .D(n2129), .Y(n2125) );
  OAI211X1TS U3840 ( .A0(n3972), .A1(n1114), .B0(n2116), .C0(n2117), .Y(n2446)
         );
  AOI22X1TS U3841 ( .A0(n480), .A1(n2118), .B0(n3118), .B1(
        destinationAddressOut[8]), .Y(n2116) );
  AOI222XLTS U3842 ( .A0(n1988), .A1(n4232), .B0(n1118), .B1(
        destinationAddressIn_NORTH[8]), .C0(n2968), .C1(n4012), .Y(n2117) );
  NAND4X1TS U3843 ( .A(n2119), .B(n2120), .C(n2121), .D(n2122), .Y(n2118) );
  OAI211X1TS U3844 ( .A0(n3969), .A1(n1115), .B0(n2109), .C0(n2110), .Y(n2447)
         );
  AOI22X1TS U3845 ( .A0(n479), .A1(n2111), .B0(n3118), .B1(
        destinationAddressOut[7]), .Y(n2109) );
  AOI222XLTS U3846 ( .A0(n1988), .A1(n4229), .B0(n1118), .B1(
        destinationAddressIn_NORTH[7]), .C0(n2968), .C1(n4009), .Y(n2110) );
  NAND4X1TS U3847 ( .A(n2112), .B(n2113), .C(n2114), .D(n2115), .Y(n2111) );
  OAI211X1TS U3848 ( .A0(n3966), .A1(n1115), .B0(n2101), .C0(n2102), .Y(n2448)
         );
  AOI22X1TS U3849 ( .A0(n480), .A1(n2104), .B0(n3118), .B1(
        destinationAddressOut[6]), .Y(n2101) );
  AOI222XLTS U3850 ( .A0(n1988), .A1(n4226), .B0(n1118), .B1(
        destinationAddressIn_NORTH[6]), .C0(n2968), .C1(n4006), .Y(n2102) );
  NAND4X1TS U3851 ( .A(n2105), .B(n2106), .C(n2107), .D(n2108), .Y(n2104) );
  INVX2TS U3852 ( .A(readIn_SOUTH), .Y(n998) );
  INVX2TS U3853 ( .A(readIn_NORTH), .Y(n983) );
  INVX2TS U3854 ( .A(destinationAddressIn_NORTH[7]), .Y(n981) );
  INVX2TS U3855 ( .A(destinationAddressIn_NORTH[6]), .Y(n982) );
  OAI21X1TS U3856 ( .A0(n6257), .A1(n1143), .B0(n4573), .Y(n1145) );
  NOR2X1TS U3857 ( .A(n1147), .B(n1145), .Y(n2883) );
  AOI21X1TS U3858 ( .A0(n9), .A1(n479), .B0(n122), .Y(n1147) );
  OAI22X1TS U3859 ( .A0(n154), .A1(n129), .B0(n127), .B1(n130), .Y(n2889) );
  INVX2TS U3860 ( .A(n5326), .Y(n942) );
  XNOR2X1TS U3861 ( .A(n2947), .B(n1144), .Y(n2946) );
  OAI22X1TS U3862 ( .A0(n1), .A1(n2948), .B0(n979), .B1(n2949), .Y(n2947) );
  NOR2X1TS U3863 ( .A(n774), .B(n44), .Y(n2949) );
  NAND2X1TS U3864 ( .A(n494), .B(n469), .Y(n1987) );
  NAND2X1TS U3865 ( .A(n9), .B(n122), .Y(n1143) );
  AO22X1TS U3866 ( .A0(n3177), .A1(n770), .B0(n3176), .B1(n978), .Y(n2095) );
  AOI22X1TS U3867 ( .A0(n489), .A1(n3186), .B0(n470), .B1(n3232), .Y(n2154) );
  AOI22X1TS U3868 ( .A0(n489), .A1(n3187), .B0(n470), .B1(n3231), .Y(n2147) );
  AOI22X1TS U3869 ( .A0(n489), .A1(n3188), .B0(n470), .B1(n3230), .Y(n2140) );
  AOI22X1TS U3870 ( .A0(n489), .A1(n3189), .B0(n470), .B1(n3229), .Y(n2133) );
  AOI22X1TS U3871 ( .A0(n490), .A1(n3190), .B0(n471), .B1(n3228), .Y(n2126) );
  AOI22X1TS U3872 ( .A0(n490), .A1(n3191), .B0(n471), .B1(n3227), .Y(n2119) );
  AOI22X1TS U3873 ( .A0(n490), .A1(n3192), .B0(n471), .B1(n3226), .Y(n2112) );
  AOI22X1TS U3874 ( .A0(n490), .A1(n3193), .B0(n471), .B1(n3225), .Y(n2105) );
  AOI22X1TS U3875 ( .A0(n491), .A1(n3178), .B0(n472), .B1(n3240), .Y(n2157) );
  AOI22X1TS U3876 ( .A0(n491), .A1(n3179), .B0(n472), .B1(n3239), .Y(n2150) );
  AOI22X1TS U3877 ( .A0(n491), .A1(n3180), .B0(n472), .B1(n3238), .Y(n2143) );
  AOI22X1TS U3878 ( .A0(n491), .A1(n3181), .B0(n473), .B1(n3237), .Y(n2136) );
  AOI22X1TS U3879 ( .A0(n492), .A1(n3182), .B0(n474), .B1(n3236), .Y(n2129) );
  AOI22X1TS U3880 ( .A0(n492), .A1(n3183), .B0(n473), .B1(n3235), .Y(n2122) );
  AOI22X1TS U3881 ( .A0(n492), .A1(n3184), .B0(n474), .B1(n3234), .Y(n2115) );
  AOI22X1TS U3882 ( .A0(n492), .A1(n3185), .B0(n474), .B1(n3233), .Y(n2108) );
  AOI22X1TS U3883 ( .A0(n133), .A1(n3210), .B0(n3209), .B1(n186), .Y(n2155) );
  AOI22X1TS U3884 ( .A0(n134), .A1(n3212), .B0(n3211), .B1(n184), .Y(n2148) );
  AOI22X1TS U3885 ( .A0(n134), .A1(n3214), .B0(n3213), .B1(n185), .Y(n2141) );
  AOI22X1TS U3886 ( .A0(n133), .A1(n3216), .B0(n3215), .B1(n186), .Y(n2134) );
  AOI22X1TS U3887 ( .A0(n133), .A1(n3218), .B0(n3217), .B1(n184), .Y(n2127) );
  AOI22X1TS U3888 ( .A0(n134), .A1(n3220), .B0(n3219), .B1(n185), .Y(n2120) );
  AOI22X1TS U3889 ( .A0(n133), .A1(n3222), .B0(n3221), .B1(n186), .Y(n2113) );
  AOI22X1TS U3890 ( .A0(n134), .A1(n3224), .B0(n3223), .B1(n184), .Y(n2106) );
  AOI22X1TS U3891 ( .A0(n978), .A1(n3195), .B0(n465), .B1(n3194), .Y(n2156) );
  AOI22X1TS U3892 ( .A0(n804), .A1(n3197), .B0(n770), .B1(n3196), .Y(n2149) );
  AOI22X1TS U3893 ( .A0(n805), .A1(n3199), .B0(n464), .B1(n3198), .Y(n2142) );
  AOI22X1TS U3894 ( .A0(n978), .A1(n567), .B0(n465), .B1(n3200), .Y(n2135) );
  AOI22X1TS U3895 ( .A0(n804), .A1(n3202), .B0(n770), .B1(n3201), .Y(n2128) );
  AOI22X1TS U3896 ( .A0(n805), .A1(n3204), .B0(n464), .B1(n3203), .Y(n2121) );
  AOI22X1TS U3897 ( .A0(n978), .A1(n3206), .B0(n465), .B1(n3205), .Y(n2114) );
  AOI22X1TS U3898 ( .A0(n804), .A1(n3208), .B0(n770), .B1(n3207), .Y(n2107) );
  NAND3X1TS U3899 ( .A(n4), .B(n9), .C(n8), .Y(n2082) );
  AOI221X1TS U3900 ( .A0(n473), .A1(\readOutbuffer[2] ), .B0(n805), .B1(
        readOutbuffer_7), .C0(n6257), .Y(n2078) );
  INVX2TS U3901 ( .A(n2062), .Y(n973) );
  NOR2X1TS U3902 ( .A(n156), .B(n972), .Y(n2058) );
  AOI21X1TS U3903 ( .A0(n1842), .A1(n932), .B0(n921), .Y(n1844) );
  NAND2X1TS U3904 ( .A(n4195), .B(n921), .Y(n1840) );
  INVX2TS U3905 ( .A(n1843), .Y(n921) );
  CLKBUFX2TS U3906 ( .A(n794), .Y(n3832) );
  AOI21XLTS U3907 ( .A0(n4195), .A1(n924), .B0(n482), .Y(n1811) );
  AOI32XLTS U3908 ( .A0(n1813), .A1(n1814), .A2(n1815), .B0(n4201), .B1(n928), 
        .Y(n1812) );
  NOR2X1TS U3909 ( .A(n1814), .B(n482), .Y(n1154) );
  AOI32XLTS U3910 ( .A0(n467), .A1(n1825), .A2(n1826), .B0(n3599), .B1(n681), 
        .Y(n2568) );
  AOI32XLTS U3911 ( .A0(n484), .A1(n1828), .A2(n4200), .B0(n1829), .B1(n1830), 
        .Y(n1826) );
  AOI21XLTS U3912 ( .A0(readIn_NORTH), .A1(n1834), .B0(n1835), .Y(n1833) );
  OAI221XLTS U3913 ( .A0(n176), .A1(n140), .B0(n1797), .B1(n969), .C0(n1955), 
        .Y(n2514) );
  OAI221XLTS U3914 ( .A0(n175), .A1(n137), .B0(n454), .B1(n968), .C0(n1956), 
        .Y(n2513) );
  OAI221XLTS U3915 ( .A0(n176), .A1(n152), .B0(n1797), .B1(n967), .C0(n1957), 
        .Y(n2512) );
  OAI221XLTS U3916 ( .A0(n1796), .A1(n146), .B0(n195), .B1(n581), .C0(n1958), 
        .Y(n2511) );
  OAI221XLTS U3917 ( .A0(n176), .A1(n150), .B0(n1797), .B1(n603), .C0(n1959), 
        .Y(n2510) );
  OAI221XLTS U3918 ( .A0(n1796), .A1(n144), .B0(n454), .B1(n604), .C0(n1960), 
        .Y(n2509) );
  OAI221XLTS U3919 ( .A0(n176), .A1(n147), .B0(n188), .B1(n605), .C0(n1961), 
        .Y(n2508) );
  OAI221XLTS U3920 ( .A0(n1796), .A1(n141), .B0(n192), .B1(n582), .C0(n1962), 
        .Y(n2507) );
  OAI221XLTS U3921 ( .A0(n175), .A1(n160), .B0(n454), .B1(n970), .C0(n1798), 
        .Y(n2575) );
  OAI221XLTS U3922 ( .A0(n179), .A1(n139), .B0(n165), .B1(n562), .C0(n2047), 
        .Y(n2458) );
  OAI221XLTS U3923 ( .A0(n180), .A1(n136), .B0(n164), .B1(n556), .C0(n2048), 
        .Y(n2457) );
  OAI221XLTS U3924 ( .A0(n179), .A1(n151), .B0(n165), .B1(n566), .C0(n2049), 
        .Y(n2456) );
  OAI221XLTS U3925 ( .A0(n180), .A1(n145), .B0(n164), .B1(n557), .C0(n2050), 
        .Y(n2455) );
  OAI221XLTS U3926 ( .A0(n179), .A1(n149), .B0(n165), .B1(n563), .C0(n2051), 
        .Y(n2454) );
  OAI221XLTS U3927 ( .A0(n180), .A1(n143), .B0(n164), .B1(n558), .C0(n2052), 
        .Y(n2453) );
  OAI221XLTS U3928 ( .A0(n179), .A1(n148), .B0(n165), .B1(n568), .C0(n2053), 
        .Y(n2452) );
  OAI221XLTS U3929 ( .A0(n180), .A1(n142), .B0(n164), .B1(n564), .C0(n2054), 
        .Y(n2451) );
  OAI221XLTS U3930 ( .A0(n1807), .A1(n159), .B0(n1808), .B1(n765), .C0(n1809), 
        .Y(n2571) );
  AOI21XLTS U3931 ( .A0(readIn_SOUTH), .A1(n1822), .B0(n1823), .Y(n1818) );
  OAI211XLTS U3932 ( .A0(n908), .A1(n3948), .B0(n1896), .C0(n1897), .Y(n2548)
         );
  OAI211XLTS U3933 ( .A0(n913), .A1(n3951), .B0(n1898), .C0(n1899), .Y(n2547)
         );
  OAI211XLTS U3934 ( .A0(n914), .A1(n3954), .B0(n1900), .C0(n1901), .Y(n2546)
         );
  OAI211XLTS U3935 ( .A0(n908), .A1(n3957), .B0(n1902), .C0(n1903), .Y(n2545)
         );
  OAI211XLTS U3936 ( .A0(n913), .A1(n3960), .B0(n1904), .C0(n1905), .Y(n2544)
         );
  OAI211XLTS U3937 ( .A0(n914), .A1(n3963), .B0(n1906), .C0(n1907), .Y(n2543)
         );
  OAI211XLTS U3938 ( .A0(n4176), .A1(n908), .B0(n1167), .C0(n1168), .Y(n2876)
         );
  OAI211XLTS U3939 ( .A0(n4179), .A1(n908), .B0(n1172), .C0(n1173), .Y(n2875)
         );
  OAI211XLTS U3940 ( .A0(n4182), .A1(n913), .B0(n1174), .C0(n1175), .Y(n2874)
         );
  OAI211XLTS U3941 ( .A0(n4185), .A1(n913), .B0(n1176), .C0(n1177), .Y(n2873)
         );
  OAI211XLTS U3942 ( .A0(n4188), .A1(n914), .B0(n1178), .C0(n1179), .Y(n2872)
         );
  OAI211XLTS U3943 ( .A0(n4191), .A1(n914), .B0(n1180), .C0(n1181), .Y(n2871)
         );
  AOI222XLTS U3944 ( .A0(n4200), .A1(n1820), .B0(readIn_NORTH), .B1(n1821), 
        .C0(n4195), .C1(n923), .Y(n1819) );
  AOI32XLTS U3945 ( .A0(n100), .A1(n1840), .A2(n1841), .B0(n3869), .B1(n676), 
        .Y(n2566) );
  OAI221XLTS U3946 ( .A0(n177), .A1(n140), .B0(n173), .B1(n575), .C0(n1978), 
        .Y(n2500) );
  OAI221XLTS U3947 ( .A0(n178), .A1(n137), .B0(n172), .B1(n569), .C0(n1979), 
        .Y(n2499) );
  OAI221XLTS U3948 ( .A0(n177), .A1(n152), .B0(n173), .B1(n572), .C0(n1980), 
        .Y(n2498) );
  OAI221XLTS U3949 ( .A0(n178), .A1(n146), .B0(n172), .B1(n573), .C0(n1981), 
        .Y(n2497) );
  OAI221XLTS U3950 ( .A0(n177), .A1(n150), .B0(n173), .B1(n570), .C0(n1982), 
        .Y(n2496) );
  OAI221XLTS U3951 ( .A0(n178), .A1(n144), .B0(n172), .B1(n576), .C0(n1983), 
        .Y(n2495) );
  OAI221XLTS U3952 ( .A0(n177), .A1(n147), .B0(n173), .B1(n574), .C0(n1984), 
        .Y(n2494) );
  OAI221XLTS U3953 ( .A0(n178), .A1(n141), .B0(n172), .B1(n571), .C0(n1985), 
        .Y(n2493) );
  OAI221XLTS U3954 ( .A0(n1799), .A1(n984), .B0(n1800), .B1(n766), .C0(n1801), 
        .Y(n2574) );
  AOI32XLTS U3955 ( .A0(n460), .A1(n1832), .A2(n1833), .B0(n112), .B1(n769), 
        .Y(n2567) );
  OA22XLTS U3956 ( .A0(n973), .A1(n2950), .B0(n2951), .B1(n2062), .Y(n2938) );
endmodule


module router ( clk, localRouterAddress, destinationAddressIn_NORTH, 
        requesterAddressIn_NORTH, readIn_NORTH, writeIn_NORTH, dataIn_NORTH, 
        destinationAddressOut_NORTH, requesterAddressOut_NORTH, readOut_NORTH, 
        writeOut_NORTH, dataOut_NORTH, destinationAddressIn_SOUTH, 
        requesterAddressIn_SOUTH, readIn_SOUTH, writeIn_SOUTH, dataIn_SOUTH, 
        destinationAddressOut_SOUTH, requesterAddressOut_SOUTH, readOut_SOUTH, 
        writeOut_SOUTH, dataOut_SOUTH, destinationAddressIn_EAST, 
        requesterAddressIn_EAST, readIn_EAST, writeIn_EAST, dataIn_EAST, 
        destinationAddressOut_EAST, requesterAddressOut_EAST, readOut_EAST, 
        writeOut_EAST, dataOut_EAST, destinationAddressIn_WEST, 
        requesterAddressIn_WEST, readIn_WEST, writeIn_WEST, dataIn_WEST, 
        destinationAddressOut_WEST, requesterAddressOut_WEST, readOut_WEST, 
        writeOut_WEST, dataOut_WEST, cacheDataIn_A, cacheAddressIn_A, 
        cacheDataOut_A, memWrite_A, portA_writtenTo, cacheDataIn_B, 
        cacheAddressIn_B, cacheDataOut_B, memWrite_B, portB_writtenTo, 
        reset_BAR );
  input [5:0] localRouterAddress;
  input [13:0] destinationAddressIn_NORTH;
  input [5:0] requesterAddressIn_NORTH;
  input [31:0] dataIn_NORTH;
  output [13:0] destinationAddressOut_NORTH;
  output [5:0] requesterAddressOut_NORTH;
  output [31:0] dataOut_NORTH;
  input [13:0] destinationAddressIn_SOUTH;
  input [5:0] requesterAddressIn_SOUTH;
  input [31:0] dataIn_SOUTH;
  output [13:0] destinationAddressOut_SOUTH;
  output [5:0] requesterAddressOut_SOUTH;
  output [31:0] dataOut_SOUTH;
  input [13:0] destinationAddressIn_EAST;
  input [5:0] requesterAddressIn_EAST;
  input [31:0] dataIn_EAST;
  output [13:0] destinationAddressOut_EAST;
  output [5:0] requesterAddressOut_EAST;
  output [31:0] dataOut_EAST;
  input [13:0] destinationAddressIn_WEST;
  input [5:0] requesterAddressIn_WEST;
  input [31:0] dataIn_WEST;
  output [13:0] destinationAddressOut_WEST;
  output [5:0] requesterAddressOut_WEST;
  output [31:0] dataOut_WEST;
  output [31:0] cacheDataIn_A;
  output [7:0] cacheAddressIn_A;
  input [31:0] cacheDataOut_A;
  output [31:0] cacheDataIn_B;
  output [7:0] cacheAddressIn_B;
  input [31:0] cacheDataOut_B;
  input clk, readIn_NORTH, writeIn_NORTH, readIn_SOUTH, writeIn_SOUTH,
         readIn_EAST, writeIn_EAST, readIn_WEST, writeIn_WEST, portA_writtenTo,
         portB_writtenTo, reset_BAR;
  output readOut_NORTH, writeOut_NORTH, readOut_SOUTH, writeOut_SOUTH,
         readOut_EAST, writeOut_EAST, readOut_WEST, writeOut_WEST, memWrite_A,
         memWrite_B;
  wire   reset, memRead_NORTH, memWrite_NORTH, memRead_SOUTH, memWrite_SOUTH,
         memRead_EAST, memWrite_EAST, memRead_WEST, memWrite_WEST,
         readReady_NORTH, readReady_SOUTH, readReady_EAST, readReady_WEST,
         writeInBuffer_SOUTH, readInBuffer_EAST, writeInBuffer_EAST,
         readInBuffer_WEST, writeInBuffer_WEST,
         destinationAddressInBuffer_NORTH_5,
         destinationAddressInBuffer_NORTH_4,
         destinationAddressInBuffer_NORTH_3,
         destinationAddressInBuffer_NORTH_2,
         destinationAddressInBuffer_NORTH_1,
         destinationAddressInBuffer_NORTH_0, n2, n1, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408;
  wire   [3:0] outputPortSelect_NORTH;
  wire   [3:0] outputPortSelect_SOUTH;
  wire   [3:0] outputPortSelect_EAST;
  wire   [3:0] outputPortSelect_WEST;
  wire   [5:0] cacheRequesterAddress_NORTH;
  wire   [31:0] cacheDataOut_NORTH;
  wire   [5:0] requesterAddressInBuffer_SOUTH;
  wire   [31:0] dataInBuffer_SOUTH;
  wire   [5:0] cacheRequesterAddress_SOUTH;
  wire   [31:0] cacheDataOut_SOUTH;
  wire   [31:0] dataInBuffer_EAST;
  wire   [5:0] cacheRequesterAddress_EAST;
  wire   [31:0] cacheDataOut_EAST;
  wire   [31:0] dataInBuffer_WEST;
  wire   [5:0] cacheRequesterAddress_WEST;
  wire   [31:0] cacheDataOut_WEST;
  wire   [13:0] destinationAddressInBuffer_SOUTH;
  wire   [5:0] requesterAddressInBuffer_EAST;
  wire   [31:0] dataInBuffer_NORTH;
  wire   [5:0] requesterAddressInBuffer_NORTH;
  wire   [5:0] requesterAddressInBuffer_WEST;
  wire   [13:0] destinationAddressInBuffer_WEST;
  wire   [13:0] destinationAddressInBuffer_EAST;
  assign reset = reset_BAR;

  incomingPortHandler_0 inNorth ( .clk(clk), .reset(n384), 
        .localRouterAddress({n17, n15, n13, localRouterAddress[2:0]}), 
        .destinationAddressIn({destinationAddressIn_NORTH[13:8], 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .requesterAddressIn({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .readIn(readIn_NORTH), .writeIn(
        writeIn_NORTH), .outputPortSelect(outputPortSelect_NORTH), .memRead(
        memRead_NORTH), .memWrite(memWrite_NORTH) );
  incomingPortHandler_3 inSouth ( .clk(clk), .reset(n382), 
        .localRouterAddress({n17, n15, n13, localRouterAddress[2:0]}), 
        .destinationAddressIn({destinationAddressIn_SOUTH[13:8], 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .requesterAddressIn({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .readIn(readIn_SOUTH), .writeIn(
        writeIn_SOUTH), .outputPortSelect(outputPortSelect_SOUTH), .memRead(
        memRead_SOUTH), .memWrite(memWrite_SOUTH) );
  incomingPortHandler_2 inEast ( .clk(clk), .reset(n383), .localRouterAddress(
        {n16, n14, n12, localRouterAddress[2:0]}), .destinationAddressIn({
        destinationAddressIn_EAST[13:8], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .requesterAddressIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .readIn(readIn_EAST), .writeIn(writeIn_EAST), .outputPortSelect(
        outputPortSelect_EAST), .memRead(memRead_EAST), .memWrite(
        memWrite_EAST) );
  incomingPortHandler_1 inWest ( .clk(clk), .reset(n385), .localRouterAddress(
        {n16, n14, n12, localRouterAddress[2:0]}), .destinationAddressIn({
        destinationAddressIn_WEST[13:8], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .requesterAddressIn({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .readIn(readIn_WEST), .writeIn(writeIn_WEST), .outputPortSelect(
        outputPortSelect_WEST), .memRead(memRead_WEST), .memWrite(
        memWrite_WEST) );
  cacheAccessArbiter cacheController ( .clk(clk), .reset(n385), 
        .cacheAddressIn_NORTH({n94, n91, n145, n144, n143, n142, n141, n140}), 
        .requesterAddressIn_NORTH({n151, n150, n149, n148, n147, n146}), 
        .memRead_NORTH(memRead_NORTH), .memWrite_NORTH(memWrite_NORTH), 
        .dataIn_NORTH({n183, n182, n181, n180, n179, n178, n177, n176, n175, 
        n174, n173, n172, n171, n170, n169, n168, n167, n166, n165, n164, n163, 
        n162, n161, n160, n159, n158, n157, n156, n155, n154, n153, n152}), 
        .readReady_NORTH(readReady_NORTH), .requesterAddressOut_NORTH(
        cacheRequesterAddress_NORTH), .cacheDataOut_NORTH(cacheDataOut_NORTH), 
        .cacheAddressIn_SOUTH({n202, n201, n200, n199, n197, n195, n194, n193}), .requesterAddressIn_SOUTH({n378, n376, n374, n372, n370, n368}), 
        .memRead_SOUTH(memRead_SOUTH), .memWrite_SOUTH(memWrite_SOUTH), 
        .dataIn_SOUTH({n367, n365, n363, n361, n359, n357, n356, n354, n352, 
        n351, n349, n347, n346, n344, n342, n340, n339, n337, n336, n334, n332, 
        n330, n328, n327, n325, n323, n321, n319, n318, n316, n314, n312}), 
        .readReady_SOUTH(readReady_SOUTH), .requesterAddressOut_SOUTH(
        cacheRequesterAddress_SOUTH), .cacheDataOut_SOUTH(cacheDataOut_SOUTH), 
        .cacheAddressIn_EAST(destinationAddressInBuffer_EAST[7:0]), 
        .requesterAddressIn_EAST(requesterAddressInBuffer_EAST), 
        .memRead_EAST(memRead_EAST), .memWrite_EAST(memWrite_EAST), 
        .dataIn_EAST({n310, n308, n306, n304, n302, n300, n298, n296, n294, 
        n292, n290, n288, n286, n284, n282, n280, n278, n276, n274, n272, n270, 
        n268, n266, n264, n262, n260, n258, n256, n254, n252, n250, n248}), 
        .readReady_EAST(readReady_EAST), .requesterAddressOut_EAST(
        cacheRequesterAddress_EAST), .cacheDataOut_EAST(cacheDataOut_EAST), 
        .cacheAddressIn_WEST(destinationAddressInBuffer_WEST[7:0]), 
        .requesterAddressIn_WEST({n138, n136, n134, n132, n130, n128}), 
        .memRead_WEST(memRead_WEST), .memWrite_WEST(memWrite_WEST), 
        .dataIn_WEST(dataInBuffer_WEST), .readReady_WEST(readReady_WEST), 
        .requesterAddressOut_WEST(cacheRequesterAddress_WEST), 
        .cacheDataOut_WEST(cacheDataOut_WEST), .cacheDataIn_A(cacheDataIn_A), 
        .cacheAddressIn_A(cacheAddressIn_A), .cacheDataOut_A(cacheDataOut_A), 
        .memWrite_A(memWrite_A), .cacheDataIn_B(cacheDataIn_B), 
        .cacheAddressIn_B(cacheAddressIn_B), .cacheDataOut_B(cacheDataOut_B), 
        .memWrite_B(memWrite_B) );
  outputPortArbiter_0 outNorth ( .clk(clk), .reset(n386), .selectBit_NORTH(
        outputPortSelect_NORTH[0]), .destinationAddressIn_NORTH({n83, n6, n75, 
        n71, n87, n79, n95, n92, destinationAddressInBuffer_NORTH_5, n144, 
        destinationAddressInBuffer_NORTH_3, n142, n141, 
        destinationAddressInBuffer_NORTH_0}), .requesterAddressIn_NORTH({
        requesterAddressInBuffer_NORTH[5], n150, n149, n148, n147, n146}), 
        .readIn_NORTH(n103), .writeIn_NORTH(n28), .dataIn_NORTH({
        dataInBuffer_NORTH[31], n182, n181, n180, dataInBuffer_NORTH[27], n178, 
        n177, n176, n175, n174, n173, n172, n171, n170, n169, n168, n167, n166, 
        n165, n164, n163, n162, dataInBuffer_NORTH[9], n160, n159, n158, 
        dataInBuffer_NORTH[5], n156, n155, n154, dataInBuffer_NORTH[1], n152}), 
        .selectBit_SOUTH(outputPortSelect_SOUTH[0]), 
        .destinationAddressIn_SOUTH({n213, n211, n209, n207, n205, n203, 
        destinationAddressInBuffer_SOUTH[7:6], n200, n198, n196, n195, n194, 
        n192}), .requesterAddressIn_SOUTH({n377, n375, n373, n371, n369, 
        requesterAddressInBuffer_SOUTH[0]}), .readIn_SOUTH(n99), 
        .writeIn_SOUTH(n191), .dataIn_SOUTH({n366, n364, n362, n360, n358, 
        dataInBuffer_SOUTH[26], n355, n353, dataInBuffer_SOUTH[23], n350, n348, 
        dataInBuffer_SOUTH[20], n345, n343, n341, dataInBuffer_SOUTH[16], n338, 
        dataInBuffer_SOUTH[14], n335, n333, n331, n329, dataInBuffer_SOUTH[9], 
        n326, n324, n322, n320, dataInBuffer_SOUTH[4], n317, n315, n313, n311}), .selectBit_EAST(outputPortSelect_EAST[0]), .destinationAddressIn_EAST({
        destinationAddressInBuffer_EAST[13:8], n111, n110, n109, n108, n107, 
        n106, n105, n104}), .requesterAddressIn_EAST({n189, n188, n187, n186, 
        n185, n184}), .readIn_EAST(readInBuffer_EAST), .writeIn_EAST(
        writeInBuffer_EAST), .dataIn_EAST({n309, n307, n305, n303, n301, n299, 
        n297, n295, n293, n291, n289, n287, n285, n283, n281, n279, n277, n275, 
        n273, n271, n269, n267, n265, n263, n261, n259, n257, n255, n253, n251, 
        n249, n247}), .selectBit_WEST(outputPortSelect_WEST[0]), 
        .destinationAddressIn_WEST({destinationAddressInBuffer_WEST[13:11], 
        n123, n121, n120, n119, n118, n117, n116, n115, n114, n113, n112}), 
        .requesterAddressIn_WEST({n139, n137, n135, n133, n131, n129}), 
        .readIn_WEST(readInBuffer_WEST), .dataIn_WEST({n246, n245, n244, n243, 
        n242, n241, n240, n239, n238, n237, n236, n235, n234, n233, n232, n231, 
        n230, n229, n228, n227, n226, n225, n224, n223, n222, n221, n220, n219, 
        n218, n217, n216, n215}), .readReady(readReady_NORTH), 
        .readRequesterAddress(cacheRequesterAddress_NORTH), .cacheDataOut(
        cacheDataOut_NORTH), .destinationAddressOut(
        destinationAddressOut_NORTH), .requesterAddressOut(
        requesterAddressOut_NORTH), .readOut(readOut_NORTH), .writeOut(
        writeOut_NORTH), .dataOut(dataOut_NORTH), .writeIn_WEST_BAR(n65) );
  outputPortArbiter_3 outSouth ( .clk(clk), .reset(n380), .selectBit_NORTH(
        outputPortSelect_NORTH[1]), .destinationAddressIn_NORTH({n7, n69, n8, 
        n9, n10, n11, n94, n91, n145, destinationAddressInBuffer_NORTH_4, n143, 
        destinationAddressInBuffer_NORTH_2, destinationAddressInBuffer_NORTH_1, 
        n140}), .requesterAddressIn_NORTH({n151, 
        requesterAddressInBuffer_NORTH[4:0]}), .readIn_NORTH(n102), 
        .writeIn_NORTH(n3), .dataIn_NORTH({n183, dataInBuffer_NORTH[30:28], 
        n179, dataInBuffer_NORTH[26:10], n161, dataInBuffer_NORTH[8:6], n157, 
        dataInBuffer_NORTH[4:2], n153, dataInBuffer_NORTH[0]}), 
        .selectBit_SOUTH(outputPortSelect_SOUTH[1]), 
        .destinationAddressIn_SOUTH({n213, n211, n209, n207, n205, n203, 
        destinationAddressInBuffer_SOUTH[7:5], n198, n196, 
        destinationAddressInBuffer_SOUTH[2:1], n192}), 
        .requesterAddressIn_SOUTH({n377, n375, n373, n371, n369, 
        requesterAddressInBuffer_SOUTH[0]}), .readIn_SOUTH(n98), 
        .writeIn_SOUTH(n191), .dataIn_SOUTH({n366, n364, n362, n360, n358, 
        dataInBuffer_SOUTH[26], n355, n353, dataInBuffer_SOUTH[23], n350, n348, 
        dataInBuffer_SOUTH[20], n345, n343, n341, dataInBuffer_SOUTH[16], n338, 
        dataInBuffer_SOUTH[14], n335, n333, n331, n329, dataInBuffer_SOUTH[9], 
        n326, n324, n322, n320, dataInBuffer_SOUTH[4], n317, n315, n313, n311}), .selectBit_EAST(outputPortSelect_EAST[1]), .destinationAddressIn_EAST({
        destinationAddressInBuffer_EAST[13:8], n111, n110, n109, n108, n107, 
        n106, n105, n104}), .requesterAddressIn_EAST({n189, n188, n187, n186, 
        n185, n184}), .readIn_EAST(readInBuffer_EAST), .writeIn_EAST(
        writeInBuffer_EAST), .dataIn_EAST({n309, n307, n305, n303, n301, n299, 
        n297, n295, n293, n291, n289, n287, n285, n283, n281, n279, n277, n275, 
        n273, n271, n269, n267, n265, n263, n261, n259, n257, n255, n253, n251, 
        n249, n247}), .selectBit_WEST(outputPortSelect_WEST[1]), 
        .destinationAddressIn_WEST({destinationAddressInBuffer_WEST[13:11], 
        n123, n121, n120, destinationAddressInBuffer_WEST[7:6], n117, n116, 
        n115, n114, n113, n112}), .requesterAddressIn_WEST({n139, n137, n135, 
        n133, n131, n129}), .readIn_WEST(readInBuffer_WEST), .dataIn_WEST({
        n246, n245, n244, n243, n242, n241, n240, n239, n238, n237, n236, n235, 
        n234, n233, n232, n231, n230, n229, n228, n227, n226, n225, n224, n223, 
        n222, n221, n220, n219, n218, n217, n216, n215}), .readReady(
        readReady_SOUTH), .readRequesterAddress(cacheRequesterAddress_SOUTH), 
        .cacheDataOut(cacheDataOut_SOUTH), .destinationAddressOut(
        destinationAddressOut_SOUTH), .requesterAddressOut(
        requesterAddressOut_SOUTH), .readOut(readOut_SOUTH), .writeOut(
        writeOut_SOUTH), .dataOut(dataOut_SOUTH), .writeIn_WEST_BAR(n65) );
  outputPortArbiter_2 outEast ( .clk(clk), .reset(n381), .selectBit_NORTH(
        outputPortSelect_NORTH[2]), .destinationAddressIn_NORTH({n85, n68, n77, 
        n73, n89, n81, n93, n90, n145, destinationAddressInBuffer_NORTH_4, 
        n143, destinationAddressInBuffer_NORTH_2, 
        destinationAddressInBuffer_NORTH_1, n140}), .requesterAddressIn_NORTH(
        {n151, requesterAddressInBuffer_NORTH[4:0]}), .readIn_NORTH(n18), 
        .writeIn_NORTH(n3), .dataIn_NORTH({n183, dataInBuffer_NORTH[30:28], 
        n179, dataInBuffer_NORTH[26:10], n161, dataInBuffer_NORTH[8:6], n157, 
        dataInBuffer_NORTH[4:2], n153, dataInBuffer_NORTH[0]}), 
        .selectBit_SOUTH(outputPortSelect_SOUTH[2]), 
        .destinationAddressIn_SOUTH({n214, n212, n210, n208, n206, n204, n202, 
        n201, destinationAddressInBuffer_SOUTH[5:0]}), 
        .requesterAddressIn_SOUTH({n378, n376, n374, n372, n370, n368}), 
        .readIn_SOUTH(n5), .writeIn_SOUTH(n190), .dataIn_SOUTH({n367, n365, 
        n363, n361, n359, n357, n356, n354, n352, n351, n349, n347, n346, n344, 
        n342, n340, n339, n337, n336, n334, n332, n330, n328, n327, n325, n323, 
        n321, n319, n318, n316, n314, n312}), .selectBit_EAST(
        outputPortSelect_EAST[2]), .destinationAddressIn_EAST({
        destinationAddressInBuffer_EAST[13:8], n111, n110, n109, n108, n107, 
        n106, n105, n104}), .requesterAddressIn_EAST({n189, n188, n187, n186, 
        n185, n184}), .readIn_EAST(readInBuffer_EAST), .writeIn_EAST(
        writeInBuffer_EAST), .dataIn_EAST({n309, n307, n305, n303, n301, n299, 
        n297, n295, n293, n291, n289, n287, n285, n283, n281, n279, n277, n275, 
        n273, n271, n269, n267, n265, n263, n261, n259, n257, n255, n253, n251, 
        n249, n247}), .selectBit_WEST(outputPortSelect_WEST[2]), 
        .destinationAddressIn_WEST({n127, n126, n125, n124, n122, n120, n119, 
        n118, n117, n116, n115, n114, n113, n112}), .requesterAddressIn_WEST({
        n139, n137, n135, n133, n131, n129}), .readIn_WEST(readInBuffer_WEST), 
        .writeIn_WEST(writeInBuffer_WEST), .dataIn_WEST({n246, n245, n244, 
        n243, n242, n241, n240, n239, n238, n237, n236, n235, n234, n233, n232, 
        n231, n230, n229, n228, n227, n226, n225, n224, n223, n222, n221, n220, 
        n219, n218, n217, n216, n215}), .readReady(readReady_EAST), 
        .readRequesterAddress(cacheRequesterAddress_EAST), .cacheDataOut(
        cacheDataOut_EAST), .destinationAddressOut(destinationAddressOut_EAST), 
        .requesterAddressOut(requesterAddressOut_EAST), .readOut(readOut_EAST), 
        .writeOut(writeOut_EAST), .dataOut(dataOut_EAST) );
  outputPortArbiter_1 outWest ( .clk(clk), .reset(n379), .selectBit_NORTH(
        outputPortSelect_NORTH[3]), .destinationAddressIn_NORTH({n84, n67, n76, 
        n72, n88, n80, n95, n92, n145, destinationAddressInBuffer_NORTH_4, 
        n143, destinationAddressInBuffer_NORTH_2, 
        destinationAddressInBuffer_NORTH_1, n140}), .requesterAddressIn_NORTH(
        {n151, requesterAddressInBuffer_NORTH[4:0]}), .readIn_NORTH(n101), 
        .writeIn_NORTH(n28), .dataIn_NORTH({n183, dataInBuffer_NORTH[30:28], 
        n179, dataInBuffer_NORTH[26:10], n161, dataInBuffer_NORTH[8:6], n157, 
        dataInBuffer_NORTH[4:2], n153, dataInBuffer_NORTH[0]}), 
        .selectBit_SOUTH(outputPortSelect_SOUTH[3]), 
        .destinationAddressIn_SOUTH({n214, n212, n210, n208, n206, n204, n202, 
        n201, n200, n199, n197, n195, n194, n193}), .requesterAddressIn_SOUTH(
        {n378, n376, n374, n372, n370, n368}), .readIn_SOUTH(n97), 
        .writeIn_SOUTH(n190), .dataIn_SOUTH({n367, n365, n363, n361, n359, 
        n357, n356, n354, n352, n351, n349, n347, n346, n344, n342, n340, n339, 
        n337, n336, n334, n332, n330, n328, n327, n325, n323, n321, n319, n318, 
        n316, n314, n312}), .selectBit_EAST(outputPortSelect_EAST[3]), 
        .destinationAddressIn_EAST({destinationAddressInBuffer_EAST[13:8], 
        n111, n110, n109, n108, n107, n106, n105, n104}), 
        .requesterAddressIn_EAST({n189, n188, n187, n186, n185, n184}), 
        .readIn_EAST(readInBuffer_EAST), .writeIn_EAST(writeInBuffer_EAST), 
        .dataIn_EAST({n309, n307, n305, n303, n301, n299, n297, n295, n293, 
        n291, n289, n287, n285, n283, n281, n279, n277, n275, n273, n271, n269, 
        n267, n265, n263, n261, n259, n257, n255, n253, n251, n249, n247}), 
        .selectBit_WEST(outputPortSelect_WEST[3]), .destinationAddressIn_WEST(
        {n127, n126, n125, n124, n122, destinationAddressInBuffer_WEST[8], 
        n119, n118, n117, n116, n115, n114, n113, n112}), 
        .requesterAddressIn_WEST({n139, n137, n135, n133, n131, n129}), 
        .readIn_WEST(readInBuffer_WEST), .writeIn_WEST(writeInBuffer_WEST), 
        .dataIn_WEST({n246, n245, n244, n243, n242, n241, n240, n239, n238, 
        n237, n236, n235, n234, n233, n232, n231, n230, n229, n228, n227, n226, 
        n225, n224, n223, n222, n221, n220, n219, n218, n217, n216, n215}), 
        .readReady(readReady_WEST), .readRequesterAddress(
        cacheRequesterAddress_WEST), .cacheDataOut(cacheDataOut_WEST), 
        .destinationAddressOut(destinationAddressOut_WEST), 
        .requesterAddressOut(requesterAddressOut_WEST), .readOut(readOut_WEST), 
        .writeOut(writeOut_WEST), .dataOut(dataOut_WEST) );
  DFFTRX2TS \dataInBuffer_EAST_reg[23]  ( .D(dataIn_EAST[23]), .RN(n395), .CK(
        clk), .Q(dataInBuffer_EAST[23]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[22]  ( .D(dataIn_EAST[22]), .RN(n395), .CK(
        clk), .Q(dataInBuffer_EAST[22]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[21]  ( .D(dataIn_EAST[21]), .RN(n395), .CK(
        clk), .Q(dataInBuffer_EAST[21]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[20]  ( .D(dataIn_EAST[20]), .RN(n395), .CK(
        clk), .Q(dataInBuffer_EAST[20]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[19]  ( .D(dataIn_EAST[19]), .RN(n396), .CK(
        clk), .Q(dataInBuffer_EAST[19]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[18]  ( .D(dataIn_EAST[18]), .RN(n396), .CK(
        clk), .Q(dataInBuffer_EAST[18]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[17]  ( .D(dataIn_EAST[17]), .RN(n396), .CK(
        clk), .Q(dataInBuffer_EAST[17]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[16]  ( .D(dataIn_EAST[16]), .RN(n396), .CK(
        clk), .Q(dataInBuffer_EAST[16]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[15]  ( .D(dataIn_EAST[15]), .RN(n397), .CK(
        clk), .Q(dataInBuffer_EAST[15]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[14]  ( .D(dataIn_EAST[14]), .RN(n397), .CK(
        clk), .Q(dataInBuffer_EAST[14]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[13]  ( .D(dataIn_EAST[13]), .RN(n397), .CK(
        clk), .Q(dataInBuffer_EAST[13]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[12]  ( .D(dataIn_EAST[12]), .RN(n397), .CK(
        clk), .Q(dataInBuffer_EAST[12]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[11]  ( .D(dataIn_EAST[11]), .RN(n398), .CK(
        clk), .Q(dataInBuffer_EAST[11]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[10]  ( .D(dataIn_EAST[10]), .RN(n398), .CK(
        clk), .Q(dataInBuffer_EAST[10]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[9]  ( .D(dataIn_EAST[9]), .RN(n398), .CK(
        clk), .Q(dataInBuffer_EAST[9]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[8]  ( .D(dataIn_EAST[8]), .RN(n398), .CK(
        clk), .Q(dataInBuffer_EAST[8]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[7]  ( .D(dataIn_EAST[7]), .RN(n399), .CK(
        clk), .Q(dataInBuffer_EAST[7]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[6]  ( .D(dataIn_EAST[6]), .RN(n399), .CK(
        clk), .Q(dataInBuffer_EAST[6]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[5]  ( .D(dataIn_EAST[5]), .RN(n399), .CK(
        clk), .Q(dataInBuffer_EAST[5]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[4]  ( .D(dataIn_EAST[4]), .RN(n399), .CK(
        clk), .Q(dataInBuffer_EAST[4]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[3]  ( .D(dataIn_EAST[3]), .RN(n400), .CK(
        clk), .Q(dataInBuffer_EAST[3]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[2]  ( .D(dataIn_EAST[2]), .RN(n400), .CK(
        clk), .Q(dataInBuffer_EAST[2]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[1]  ( .D(dataIn_EAST[1]), .RN(n400), .CK(
        clk), .Q(dataInBuffer_EAST[1]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[0]  ( .D(dataIn_EAST[0]), .RN(n400), .CK(
        clk), .Q(dataInBuffer_EAST[0]) );
  DFFTRX2TS writeInBuffer_WEST_reg ( .D(writeIn_WEST), .RN(n56), .CK(clk), .Q(
        writeInBuffer_WEST), .QN(n65) );
  DFFTRX2TS \requesterAddressInBuffer_WEST_reg[5]  ( .D(
        requesterAddressIn_WEST[5]), .RN(n55), .CK(clk), .Q(
        requesterAddressInBuffer_WEST[5]) );
  DFFTRX2TS \requesterAddressInBuffer_WEST_reg[4]  ( .D(
        requesterAddressIn_WEST[4]), .RN(n27), .CK(clk), .Q(
        requesterAddressInBuffer_WEST[4]) );
  DFFTRX2TS \requesterAddressInBuffer_WEST_reg[3]  ( .D(
        requesterAddressIn_WEST[3]), .RN(n388), .CK(clk), .Q(
        requesterAddressInBuffer_WEST[3]) );
  DFFTRX2TS \requesterAddressInBuffer_WEST_reg[2]  ( .D(
        requesterAddressIn_WEST[2]), .RN(n394), .CK(clk), .Q(
        requesterAddressInBuffer_WEST[2]) );
  DFFTRX2TS \requesterAddressInBuffer_WEST_reg[1]  ( .D(
        requesterAddressIn_WEST[1]), .RN(n46), .CK(clk), .Q(
        requesterAddressInBuffer_WEST[1]) );
  DFFTRX2TS \requesterAddressInBuffer_WEST_reg[0]  ( .D(
        requesterAddressIn_WEST[0]), .RN(n53), .CK(clk), .Q(
        requesterAddressInBuffer_WEST[0]) );
  DFFTRX2TS \requesterAddressInBuffer_NORTH_reg[3]  ( .D(
        requesterAddressIn_NORTH[3]), .RN(n50), .CK(clk), .Q(
        requesterAddressInBuffer_NORTH[3]) );
  DFFTRX2TS \requesterAddressInBuffer_NORTH_reg[0]  ( .D(
        requesterAddressIn_NORTH[0]), .RN(n57), .CK(clk), .Q(
        requesterAddressInBuffer_NORTH[0]) );
  DFFTRX2TS readInBuffer_WEST_reg ( .D(readIn_WEST), .RN(n35), .CK(clk), .Q(
        readInBuffer_WEST) );
  DFFTRX2TS \destinationAddressInBuffer_WEST_reg[13]  ( .D(
        destinationAddressIn_WEST[13]), .RN(n393), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[13]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[22]  ( .D(dataIn_WEST[22]), .RN(n52), .CK(
        clk), .Q(dataInBuffer_WEST[22]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[21]  ( .D(dataIn_WEST[21]), .RN(n47), .CK(
        clk), .Q(dataInBuffer_WEST[21]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[20]  ( .D(dataIn_WEST[20]), .RN(n45), .CK(
        clk), .Q(dataInBuffer_WEST[20]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[19]  ( .D(dataIn_WEST[19]), .RN(n23), .CK(
        clk), .Q(dataInBuffer_WEST[19]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[18]  ( .D(dataIn_WEST[18]), .RN(n49), .CK(
        clk), .Q(dataInBuffer_WEST[18]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[17]  ( .D(dataIn_WEST[17]), .RN(n39), .CK(
        clk), .Q(dataInBuffer_WEST[17]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[16]  ( .D(dataIn_WEST[16]), .RN(n41), .CK(
        clk), .Q(dataInBuffer_WEST[16]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[15]  ( .D(dataIn_WEST[15]), .RN(n387), .CK(
        clk), .Q(dataInBuffer_WEST[15]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[14]  ( .D(dataIn_WEST[14]), .RN(n390), .CK(
        clk), .Q(dataInBuffer_WEST[14]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[13]  ( .D(dataIn_WEST[13]), .RN(n408), .CK(
        clk), .Q(dataInBuffer_WEST[13]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[12]  ( .D(dataIn_WEST[12]), .RN(n26), .CK(
        clk), .Q(dataInBuffer_WEST[12]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[9]  ( .D(dataIn_WEST[9]), .RN(n33), .CK(clk), .Q(dataInBuffer_WEST[9]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[1]  ( .D(dataIn_WEST[1]), .RN(n30), .CK(clk), .Q(dataInBuffer_WEST[1]) );
  DFFTRX2TS writeInBuffer_SOUTH_reg ( .D(writeIn_SOUTH), .RN(n42), .CK(clk), 
        .Q(writeInBuffer_SOUTH) );
  DFFTRX2TS writeInBuffer_NORTH_reg ( .D(writeIn_NORTH), .RN(n401), .CK(clk), 
        .Q(n3), .QN(n4) );
  DFFTRX2TS writeInBuffer_EAST_reg ( .D(writeIn_EAST), .RN(n389), .CK(clk), 
        .Q(writeInBuffer_EAST) );
  DFFTRX2TS \requesterAddressInBuffer_SOUTH_reg[5]  ( .D(
        requesterAddressIn_SOUTH[5]), .RN(n22), .CK(clk), .Q(
        requesterAddressInBuffer_SOUTH[5]) );
  DFFTRX2TS \requesterAddressInBuffer_SOUTH_reg[4]  ( .D(
        requesterAddressIn_SOUTH[4]), .RN(n408), .CK(clk), .Q(
        requesterAddressInBuffer_SOUTH[4]) );
  DFFTRX2TS \requesterAddressInBuffer_SOUTH_reg[3]  ( .D(
        requesterAddressIn_SOUTH[3]), .RN(n64), .CK(clk), .Q(
        requesterAddressInBuffer_SOUTH[3]) );
  DFFTRX2TS \requesterAddressInBuffer_SOUTH_reg[2]  ( .D(
        requesterAddressIn_SOUTH[2]), .RN(n22), .CK(clk), .Q(
        requesterAddressInBuffer_SOUTH[2]) );
  DFFTRX2TS \requesterAddressInBuffer_SOUTH_reg[1]  ( .D(
        requesterAddressIn_SOUTH[1]), .RN(n21), .CK(clk), .Q(
        requesterAddressInBuffer_SOUTH[1]) );
  DFFTRX2TS \requesterAddressInBuffer_SOUTH_reg[0]  ( .D(
        requesterAddressIn_SOUTH[0]), .RN(n394), .CK(clk), .Q(
        requesterAddressInBuffer_SOUTH[0]) );
  DFFTRX2TS \requesterAddressInBuffer_NORTH_reg[5]  ( .D(
        requesterAddressIn_NORTH[5]), .RN(n54), .CK(clk), .Q(
        requesterAddressInBuffer_NORTH[5]) );
  DFFTRX2TS \requesterAddressInBuffer_NORTH_reg[4]  ( .D(
        requesterAddressIn_NORTH[4]), .RN(n47), .CK(clk), .Q(
        requesterAddressInBuffer_NORTH[4]) );
  DFFTRX2TS \requesterAddressInBuffer_NORTH_reg[2]  ( .D(
        requesterAddressIn_NORTH[2]), .RN(n45), .CK(clk), .Q(
        requesterAddressInBuffer_NORTH[2]) );
  DFFTRX2TS \requesterAddressInBuffer_NORTH_reg[1]  ( .D(
        requesterAddressIn_NORTH[1]), .RN(n20), .CK(clk), .Q(
        requesterAddressInBuffer_NORTH[1]) );
  DFFTRX2TS \requesterAddressInBuffer_EAST_reg[5]  ( .D(
        requesterAddressIn_EAST[5]), .RN(n43), .CK(clk), .Q(
        requesterAddressInBuffer_EAST[5]) );
  DFFTRX2TS \requesterAddressInBuffer_EAST_reg[4]  ( .D(
        requesterAddressIn_EAST[4]), .RN(n55), .CK(clk), .Q(
        requesterAddressInBuffer_EAST[4]) );
  DFFTRX2TS \requesterAddressInBuffer_EAST_reg[3]  ( .D(
        requesterAddressIn_EAST[3]), .RN(n393), .CK(clk), .Q(
        requesterAddressInBuffer_EAST[3]) );
  DFFTRX2TS \requesterAddressInBuffer_EAST_reg[2]  ( .D(
        requesterAddressIn_EAST[2]), .RN(n407), .CK(clk), .Q(
        requesterAddressInBuffer_EAST[2]) );
  DFFTRX2TS \requesterAddressInBuffer_EAST_reg[1]  ( .D(
        requesterAddressIn_EAST[1]), .RN(n36), .CK(clk), .Q(
        requesterAddressInBuffer_EAST[1]) );
  DFFTRX2TS \requesterAddressInBuffer_EAST_reg[0]  ( .D(
        requesterAddressIn_EAST[0]), .RN(n64), .CK(clk), .Q(
        requesterAddressInBuffer_EAST[0]) );
  DFFTRX2TS readInBuffer_SOUTH_reg ( .D(readIn_SOUTH), .RN(n390), .CK(clk), 
        .Q(n5), .QN(n96) );
  DFFTRX2TS readInBuffer_NORTH_reg ( .D(readIn_NORTH), .RN(n64), .CK(clk), .Q(
        n18), .QN(n100) );
  DFFTRX2TS readInBuffer_EAST_reg ( .D(readIn_EAST), .RN(n24), .CK(clk), .Q(
        readInBuffer_EAST) );
  DFFTRX2TS \destinationAddressInBuffer_WEST_reg[12]  ( .D(
        destinationAddressIn_WEST[12]), .RN(n51), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[12]) );
  DFFTRX2TS \destinationAddressInBuffer_WEST_reg[11]  ( .D(
        destinationAddressIn_WEST[11]), .RN(n48), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[11]) );
  DFFTRX2TS \destinationAddressInBuffer_WEST_reg[10]  ( .D(
        destinationAddressIn_WEST[10]), .RN(n38), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[10]) );
  DFFTRX2TS \destinationAddressInBuffer_WEST_reg[9]  ( .D(
        destinationAddressIn_WEST[9]), .RN(n58), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[9]) );
  DFFTRX2TS \destinationAddressInBuffer_WEST_reg[8]  ( .D(
        destinationAddressIn_WEST[8]), .RN(n20), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[8]) );
  DFFTRX2TS \destinationAddressInBuffer_WEST_reg[7]  ( .D(
        destinationAddressIn_WEST[7]), .RN(n47), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[7]) );
  DFFTRX2TS \destinationAddressInBuffer_WEST_reg[6]  ( .D(
        destinationAddressIn_WEST[6]), .RN(n387), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[6]) );
  DFFTRX2TS \destinationAddressInBuffer_WEST_reg[5]  ( .D(
        destinationAddressIn_WEST[5]), .RN(n25), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[5]) );
  DFFTRX2TS \destinationAddressInBuffer_WEST_reg[4]  ( .D(
        destinationAddressIn_WEST[4]), .RN(n33), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[4]) );
  DFFTRX2TS \destinationAddressInBuffer_WEST_reg[3]  ( .D(
        destinationAddressIn_WEST[3]), .RN(n30), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[3]) );
  DFFTRX2TS \destinationAddressInBuffer_WEST_reg[2]  ( .D(
        destinationAddressIn_WEST[2]), .RN(n42), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[2]) );
  DFFTRX2TS \destinationAddressInBuffer_WEST_reg[1]  ( .D(
        destinationAddressIn_WEST[1]), .RN(n57), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[1]) );
  DFFTRX2TS \destinationAddressInBuffer_WEST_reg[0]  ( .D(
        destinationAddressIn_WEST[0]), .RN(n44), .CK(clk), .Q(
        destinationAddressInBuffer_WEST[0]) );
  DFFTRX2TS \destinationAddressInBuffer_SOUTH_reg[13]  ( .D(
        destinationAddressIn_SOUTH[13]), .RN(n25), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[13]) );
  DFFTRX2TS \destinationAddressInBuffer_SOUTH_reg[12]  ( .D(
        destinationAddressIn_SOUTH[12]), .RN(n387), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[12]) );
  DFFTRX2TS \destinationAddressInBuffer_SOUTH_reg[11]  ( .D(
        destinationAddressIn_SOUTH[11]), .RN(n25), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[11]) );
  DFFTRX2TS \destinationAddressInBuffer_SOUTH_reg[10]  ( .D(
        destinationAddressIn_SOUTH[10]), .RN(n23), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[10]) );
  DFFTRX2TS \destinationAddressInBuffer_SOUTH_reg[9]  ( .D(
        destinationAddressIn_SOUTH[9]), .RN(n25), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[9]) );
  DFFTRX2TS \destinationAddressInBuffer_SOUTH_reg[8]  ( .D(
        destinationAddressIn_SOUTH[8]), .RN(n58), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[8]) );
  DFFTRX2TS \destinationAddressInBuffer_SOUTH_reg[7]  ( .D(
        destinationAddressIn_SOUTH[7]), .RN(n55), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[7]) );
  DFFTRX2TS \destinationAddressInBuffer_SOUTH_reg[6]  ( .D(
        destinationAddressIn_SOUTH[6]), .RN(n27), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[6]) );
  DFFTRX2TS \destinationAddressInBuffer_SOUTH_reg[5]  ( .D(
        destinationAddressIn_SOUTH[5]), .RN(n24), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[5]) );
  DFFTRX2TS \destinationAddressInBuffer_SOUTH_reg[4]  ( .D(
        destinationAddressIn_SOUTH[4]), .RN(n19), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[4]) );
  DFFTRX2TS \destinationAddressInBuffer_SOUTH_reg[3]  ( .D(
        destinationAddressIn_SOUTH[3]), .RN(n394), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[3]) );
  DFFTRX2TS \destinationAddressInBuffer_SOUTH_reg[2]  ( .D(
        destinationAddressIn_SOUTH[2]), .RN(n53), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[2]) );
  DFFTRX2TS \destinationAddressInBuffer_SOUTH_reg[1]  ( .D(
        destinationAddressIn_SOUTH[1]), .RN(n50), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[1]) );
  DFFTRX2TS \destinationAddressInBuffer_SOUTH_reg[0]  ( .D(
        destinationAddressIn_SOUTH[0]), .RN(n59), .CK(clk), .Q(
        destinationAddressInBuffer_SOUTH[0]) );
  DFFTRX2TS \destinationAddressInBuffer_NORTH_reg[13]  ( .D(
        destinationAddressIn_NORTH[13]), .RN(n35), .CK(clk), .Q(n7), .QN(n82)
         );
  DFFTRX2TS \destinationAddressInBuffer_NORTH_reg[12]  ( .D(
        destinationAddressIn_NORTH[12]), .RN(n389), .CK(clk), .Q(n6), .QN(n66)
         );
  DFFTRX2TS \destinationAddressInBuffer_NORTH_reg[11]  ( .D(
        destinationAddressIn_NORTH[11]), .RN(n392), .CK(clk), .Q(n8), .QN(n74)
         );
  DFFTRX2TS \destinationAddressInBuffer_NORTH_reg[10]  ( .D(
        destinationAddressIn_NORTH[10]), .RN(n24), .CK(clk), .Q(n9), .QN(n70)
         );
  DFFTRX2TS \destinationAddressInBuffer_NORTH_reg[9]  ( .D(
        destinationAddressIn_NORTH[9]), .RN(n26), .CK(clk), .Q(n10), .QN(n86)
         );
  DFFTRX2TS \destinationAddressInBuffer_NORTH_reg[8]  ( .D(
        destinationAddressIn_NORTH[8]), .RN(n22), .CK(clk), .Q(n11), .QN(n78)
         );
  DFFTRX2TS \destinationAddressInBuffer_NORTH_reg[7]  ( .D(
        destinationAddressIn_NORTH[7]), .RN(n21), .CK(clk), .Q(n2) );
  DFFTRX2TS \destinationAddressInBuffer_NORTH_reg[6]  ( .D(
        destinationAddressIn_NORTH[6]), .RN(n39), .CK(clk), .Q(n1) );
  DFFTRX2TS \destinationAddressInBuffer_NORTH_reg[5]  ( .D(
        destinationAddressIn_NORTH[5]), .RN(n56), .CK(clk), .Q(
        destinationAddressInBuffer_NORTH_5) );
  DFFTRX2TS \destinationAddressInBuffer_NORTH_reg[4]  ( .D(
        destinationAddressIn_NORTH[4]), .RN(n47), .CK(clk), .Q(
        destinationAddressInBuffer_NORTH_4) );
  DFFTRX2TS \destinationAddressInBuffer_NORTH_reg[3]  ( .D(
        destinationAddressIn_NORTH[3]), .RN(n45), .CK(clk), .Q(
        destinationAddressInBuffer_NORTH_3) );
  DFFTRX2TS \destinationAddressInBuffer_NORTH_reg[2]  ( .D(
        destinationAddressIn_NORTH[2]), .RN(n19), .CK(clk), .Q(
        destinationAddressInBuffer_NORTH_2) );
  DFFTRX2TS \destinationAddressInBuffer_NORTH_reg[1]  ( .D(
        destinationAddressIn_NORTH[1]), .RN(n20), .CK(clk), .Q(
        destinationAddressInBuffer_NORTH_1) );
  DFFTRX2TS \destinationAddressInBuffer_NORTH_reg[0]  ( .D(
        destinationAddressIn_NORTH[0]), .RN(n32), .CK(clk), .Q(
        destinationAddressInBuffer_NORTH_0) );
  DFFTRX2TS \destinationAddressInBuffer_EAST_reg[13]  ( .D(
        destinationAddressIn_EAST[13]), .RN(n29), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[13]) );
  DFFTRX2TS \destinationAddressInBuffer_EAST_reg[12]  ( .D(
        destinationAddressIn_EAST[12]), .RN(n41), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[12]) );
  DFFTRX2TS \destinationAddressInBuffer_EAST_reg[11]  ( .D(
        destinationAddressIn_EAST[11]), .RN(n401), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[11]) );
  DFFTRX2TS \destinationAddressInBuffer_EAST_reg[10]  ( .D(
        destinationAddressIn_EAST[10]), .RN(n44), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[10]) );
  DFFTRX2TS \destinationAddressInBuffer_EAST_reg[9]  ( .D(
        destinationAddressIn_EAST[9]), .RN(n21), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[9]) );
  DFFTRX2TS \destinationAddressInBuffer_EAST_reg[8]  ( .D(
        destinationAddressIn_EAST[8]), .RN(n44), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[8]) );
  DFFTRX2TS \destinationAddressInBuffer_EAST_reg[7]  ( .D(
        destinationAddressIn_EAST[7]), .RN(n46), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[7]) );
  DFFTRX2TS \destinationAddressInBuffer_EAST_reg[6]  ( .D(
        destinationAddressIn_EAST[6]), .RN(n51), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[6]) );
  DFFTRX2TS \destinationAddressInBuffer_EAST_reg[5]  ( .D(
        destinationAddressIn_EAST[5]), .RN(n48), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[5]) );
  DFFTRX2TS \destinationAddressInBuffer_EAST_reg[4]  ( .D(
        destinationAddressIn_EAST[4]), .RN(n56), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[4]) );
  DFFTRX2TS \destinationAddressInBuffer_EAST_reg[3]  ( .D(
        destinationAddressIn_EAST[3]), .RN(n54), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[3]) );
  DFFTRX2TS \destinationAddressInBuffer_EAST_reg[2]  ( .D(
        destinationAddressIn_EAST[2]), .RN(n29), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[2]) );
  DFFTRX2TS \destinationAddressInBuffer_EAST_reg[1]  ( .D(
        destinationAddressIn_EAST[1]), .RN(n43), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[1]) );
  DFFTRX2TS \destinationAddressInBuffer_EAST_reg[0]  ( .D(
        destinationAddressIn_EAST[0]), .RN(reset), .CK(clk), .Q(
        destinationAddressInBuffer_EAST[0]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[31]  ( .D(dataIn_WEST[31]), .RN(n393), .CK(
        clk), .Q(dataInBuffer_WEST[31]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[30]  ( .D(dataIn_WEST[30]), .RN(n38), .CK(
        clk), .Q(dataInBuffer_WEST[30]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[29]  ( .D(dataIn_WEST[29]), .RN(n32), .CK(
        clk), .Q(dataInBuffer_WEST[29]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[28]  ( .D(dataIn_WEST[28]), .RN(n57), .CK(
        clk), .Q(dataInBuffer_WEST[28]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[27]  ( .D(dataIn_WEST[27]), .RN(n36), .CK(
        clk), .Q(dataInBuffer_WEST[27]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[26]  ( .D(dataIn_WEST[26]), .RN(n27), .CK(
        clk), .Q(dataInBuffer_WEST[26]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[25]  ( .D(dataIn_WEST[25]), .RN(n405), .CK(
        clk), .Q(dataInBuffer_WEST[25]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[24]  ( .D(dataIn_WEST[24]), .RN(n30), .CK(
        clk), .Q(dataInBuffer_WEST[24]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[23]  ( .D(dataIn_WEST[23]), .RN(n45), .CK(
        clk), .Q(dataInBuffer_WEST[23]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[11]  ( .D(dataIn_WEST[11]), .RN(n51), .CK(
        clk), .Q(dataInBuffer_WEST[11]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[10]  ( .D(dataIn_WEST[10]), .RN(n48), .CK(
        clk), .Q(dataInBuffer_WEST[10]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[8]  ( .D(dataIn_WEST[8]), .RN(n38), .CK(clk), .Q(dataInBuffer_WEST[8]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[7]  ( .D(dataIn_WEST[7]), .RN(n42), .CK(clk), .Q(dataInBuffer_WEST[7]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[6]  ( .D(dataIn_WEST[6]), .RN(n20), .CK(clk), .Q(dataInBuffer_WEST[6]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[5]  ( .D(dataIn_WEST[5]), .RN(n60), .CK(clk), .Q(dataInBuffer_WEST[5]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[4]  ( .D(dataIn_WEST[4]), .RN(n391), .CK(
        clk), .Q(dataInBuffer_WEST[4]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[3]  ( .D(dataIn_WEST[3]), .RN(n43), .CK(clk), .Q(dataInBuffer_WEST[3]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[2]  ( .D(dataIn_WEST[2]), .RN(n33), .CK(clk), .Q(dataInBuffer_WEST[2]) );
  DFFTRX2TS \dataInBuffer_WEST_reg[0]  ( .D(dataIn_WEST[0]), .RN(n30), .CK(clk), .Q(dataInBuffer_WEST[0]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[31]  ( .D(dataIn_SOUTH[31]), .RN(n42), 
        .CK(clk), .Q(dataInBuffer_SOUTH[31]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[30]  ( .D(dataIn_SOUTH[30]), .RN(n59), 
        .CK(clk), .Q(dataInBuffer_SOUTH[30]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[29]  ( .D(dataIn_SOUTH[29]), .RN(n27), 
        .CK(clk), .Q(dataInBuffer_SOUTH[29]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[28]  ( .D(dataIn_SOUTH[28]), .RN(n24), 
        .CK(clk), .Q(dataInBuffer_SOUTH[28]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[27]  ( .D(dataIn_SOUTH[27]), .RN(n392), 
        .CK(clk), .Q(dataInBuffer_SOUTH[27]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[26]  ( .D(dataIn_SOUTH[26]), .RN(n49), 
        .CK(clk), .Q(dataInBuffer_SOUTH[26]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[25]  ( .D(dataIn_SOUTH[25]), .RN(n53), 
        .CK(clk), .Q(dataInBuffer_SOUTH[25]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[24]  ( .D(dataIn_SOUTH[24]), .RN(n50), 
        .CK(clk), .Q(dataInBuffer_SOUTH[24]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[23]  ( .D(dataIn_SOUTH[23]), .RN(n406), 
        .CK(clk), .Q(dataInBuffer_SOUTH[23]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[22]  ( .D(dataIn_SOUTH[22]), .RN(n55), 
        .CK(clk), .Q(dataInBuffer_SOUTH[22]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[21]  ( .D(dataIn_SOUTH[21]), .RN(reset), 
        .CK(clk), .Q(dataInBuffer_SOUTH[21]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[20]  ( .D(dataIn_SOUTH[20]), .RN(n46), 
        .CK(clk), .Q(dataInBuffer_SOUTH[20]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[19]  ( .D(dataIn_SOUTH[19]), .RN(n391), 
        .CK(clk), .Q(dataInBuffer_SOUTH[19]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[18]  ( .D(dataIn_SOUTH[18]), .RN(n390), 
        .CK(clk), .Q(dataInBuffer_SOUTH[18]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[17]  ( .D(dataIn_SOUTH[17]), .RN(n22), 
        .CK(clk), .Q(dataInBuffer_SOUTH[17]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[16]  ( .D(dataIn_SOUTH[16]), .RN(n21), 
        .CK(clk), .Q(dataInBuffer_SOUTH[16]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[15]  ( .D(dataIn_SOUTH[15]), .RN(n407), 
        .CK(clk), .Q(dataInBuffer_SOUTH[15]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[14]  ( .D(dataIn_SOUTH[14]), .RN(n35), 
        .CK(clk), .Q(dataInBuffer_SOUTH[14]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[13]  ( .D(dataIn_SOUTH[13]), .RN(n388), 
        .CK(clk), .Q(dataInBuffer_SOUTH[13]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[12]  ( .D(dataIn_SOUTH[12]), .RN(n60), 
        .CK(clk), .Q(dataInBuffer_SOUTH[12]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[11]  ( .D(dataIn_SOUTH[11]), .RN(n408), 
        .CK(clk), .Q(dataInBuffer_SOUTH[11]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[10]  ( .D(dataIn_SOUTH[10]), .RN(n60), 
        .CK(clk), .Q(dataInBuffer_SOUTH[10]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[9]  ( .D(dataIn_SOUTH[9]), .RN(n53), .CK(
        clk), .Q(dataInBuffer_SOUTH[9]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[8]  ( .D(dataIn_SOUTH[8]), .RN(n50), .CK(
        clk), .Q(dataInBuffer_SOUTH[8]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[7]  ( .D(dataIn_SOUTH[7]), .RN(n39), .CK(
        clk), .Q(dataInBuffer_SOUTH[7]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[6]  ( .D(dataIn_SOUTH[6]), .RN(n58), .CK(
        clk), .Q(dataInBuffer_SOUTH[6]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[5]  ( .D(dataIn_SOUTH[5]), .RN(n392), .CK(
        clk), .Q(dataInBuffer_SOUTH[5]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[4]  ( .D(dataIn_SOUTH[4]), .RN(n52), .CK(
        clk), .Q(dataInBuffer_SOUTH[4]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[3]  ( .D(dataIn_SOUTH[3]), .RN(n49), .CK(
        clk), .Q(dataInBuffer_SOUTH[3]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[2]  ( .D(dataIn_SOUTH[2]), .RN(n26), .CK(
        clk), .Q(dataInBuffer_SOUTH[2]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[1]  ( .D(dataIn_SOUTH[1]), .RN(n32), .CK(
        clk), .Q(dataInBuffer_SOUTH[1]) );
  DFFTRX2TS \dataInBuffer_SOUTH_reg[0]  ( .D(dataIn_SOUTH[0]), .RN(n29), .CK(
        clk), .Q(dataInBuffer_SOUTH[0]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[31]  ( .D(dataIn_NORTH[31]), .RN(n41), 
        .CK(clk), .Q(dataInBuffer_NORTH[31]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[30]  ( .D(dataIn_NORTH[30]), .RN(n57), 
        .CK(clk), .Q(dataInBuffer_NORTH[30]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[29]  ( .D(dataIn_NORTH[29]), .RN(n52), 
        .CK(clk), .Q(dataInBuffer_NORTH[29]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[28]  ( .D(dataIn_NORTH[28]), .RN(n19), 
        .CK(clk), .Q(dataInBuffer_NORTH[28]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[27]  ( .D(dataIn_NORTH[27]), .RN(n23), 
        .CK(clk), .Q(dataInBuffer_NORTH[27]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[26]  ( .D(dataIn_NORTH[26]), .RN(n52), 
        .CK(clk), .Q(dataInBuffer_NORTH[26]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[25]  ( .D(dataIn_NORTH[25]), .RN(n36), 
        .CK(clk), .Q(dataInBuffer_NORTH[25]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[24]  ( .D(dataIn_NORTH[24]), .RN(n43), 
        .CK(clk), .Q(dataInBuffer_NORTH[24]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[23]  ( .D(dataIn_NORTH[23]), .RN(n58), 
        .CK(clk), .Q(dataInBuffer_NORTH[23]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[22]  ( .D(dataIn_NORTH[22]), .RN(n54), 
        .CK(clk), .Q(dataInBuffer_NORTH[22]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[21]  ( .D(dataIn_NORTH[21]), .RN(n23), 
        .CK(clk), .Q(dataInBuffer_NORTH[21]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[20]  ( .D(dataIn_NORTH[20]), .RN(n391), 
        .CK(clk), .Q(dataInBuffer_NORTH[20]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[19]  ( .D(dataIn_NORTH[19]), .RN(reset), 
        .CK(clk), .Q(dataInBuffer_NORTH[19]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[18]  ( .D(dataIn_NORTH[18]), .RN(n26), 
        .CK(clk), .Q(dataInBuffer_NORTH[18]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[17]  ( .D(dataIn_NORTH[17]), .RN(n51), 
        .CK(clk), .Q(dataInBuffer_NORTH[17]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[16]  ( .D(dataIn_NORTH[16]), .RN(n48), 
        .CK(clk), .Q(dataInBuffer_NORTH[16]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[15]  ( .D(dataIn_NORTH[15]), .RN(n59), 
        .CK(clk), .Q(dataInBuffer_NORTH[15]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[14]  ( .D(dataIn_NORTH[14]), .RN(n36), 
        .CK(clk), .Q(dataInBuffer_NORTH[14]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[13]  ( .D(dataIn_NORTH[13]), .RN(n405), 
        .CK(clk), .Q(dataInBuffer_NORTH[13]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[12]  ( .D(dataIn_NORTH[12]), .RN(n60), 
        .CK(clk), .Q(dataInBuffer_NORTH[12]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[11]  ( .D(dataIn_NORTH[11]), .RN(n389), 
        .CK(clk), .Q(dataInBuffer_NORTH[11]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[10]  ( .D(dataIn_NORTH[10]), .RN(n64), 
        .CK(clk), .Q(dataInBuffer_NORTH[10]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[9]  ( .D(dataIn_NORTH[9]), .RN(n35), .CK(
        clk), .Q(dataInBuffer_NORTH[9]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[8]  ( .D(dataIn_NORTH[8]), .RN(n44), .CK(
        clk), .Q(dataInBuffer_NORTH[8]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[7]  ( .D(dataIn_NORTH[7]), .RN(n38), .CK(
        clk), .Q(dataInBuffer_NORTH[7]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[6]  ( .D(dataIn_NORTH[6]), .RN(n56), .CK(
        clk), .Q(dataInBuffer_NORTH[6]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[5]  ( .D(dataIn_NORTH[5]), .RN(n62), .CK(
        clk), .Q(dataInBuffer_NORTH[5]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[4]  ( .D(dataIn_NORTH[4]), .RN(n62), .CK(
        clk), .Q(dataInBuffer_NORTH[4]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[3]  ( .D(dataIn_NORTH[3]), .RN(n62), .CK(
        clk), .Q(dataInBuffer_NORTH[3]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[2]  ( .D(dataIn_NORTH[2]), .RN(n63), .CK(
        clk), .Q(dataInBuffer_NORTH[2]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[1]  ( .D(dataIn_NORTH[1]), .RN(n63), .CK(
        clk), .Q(dataInBuffer_NORTH[1]) );
  DFFTRX2TS \dataInBuffer_NORTH_reg[0]  ( .D(dataIn_NORTH[0]), .RN(n63), .CK(
        clk), .Q(dataInBuffer_NORTH[0]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[31]  ( .D(dataIn_EAST[31]), .RN(n388), .CK(
        clk), .Q(dataInBuffer_EAST[31]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[30]  ( .D(dataIn_EAST[30]), .RN(n46), .CK(
        clk), .Q(dataInBuffer_EAST[30]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[29]  ( .D(dataIn_EAST[29]), .RN(n49), .CK(
        clk), .Q(dataInBuffer_EAST[29]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[28]  ( .D(dataIn_EAST[28]), .RN(n19), .CK(
        clk), .Q(dataInBuffer_EAST[28]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[27]  ( .D(dataIn_EAST[27]), .RN(n32), .CK(
        clk), .Q(dataInBuffer_EAST[27]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[26]  ( .D(dataIn_EAST[26]), .RN(n29), .CK(
        clk), .Q(dataInBuffer_EAST[26]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[25]  ( .D(dataIn_EAST[25]), .RN(n41), .CK(
        clk), .Q(dataInBuffer_EAST[25]) );
  DFFTRX2TS \dataInBuffer_EAST_reg[24]  ( .D(dataIn_EAST[24]), .RN(n59), .CK(
        clk), .Q(dataInBuffer_EAST[24]) );
  CLKBUFX2TS U2 ( .A(localRouterAddress[3]), .Y(n12) );
  CLKBUFX2TS U3 ( .A(localRouterAddress[3]), .Y(n13) );
  CLKBUFX2TS U4 ( .A(localRouterAddress[4]), .Y(n14) );
  CLKBUFX2TS U5 ( .A(localRouterAddress[4]), .Y(n15) );
  CLKBUFX2TS U6 ( .A(localRouterAddress[5]), .Y(n16) );
  CLKBUFX2TS U7 ( .A(localRouterAddress[5]), .Y(n17) );
  INVXLTS U8 ( .A(n379), .Y(n19) );
  INVXLTS U9 ( .A(n40), .Y(n20) );
  INVXLTS U10 ( .A(n381), .Y(n21) );
  INVXLTS U11 ( .A(n386), .Y(n22) );
  INVXLTS U12 ( .A(n40), .Y(n23) );
  INVXLTS U13 ( .A(n381), .Y(n24) );
  INVXLTS U14 ( .A(n383), .Y(n25) );
  INVXLTS U15 ( .A(n34), .Y(n26) );
  INVXLTS U16 ( .A(n384), .Y(n27) );
  INVXLTS U17 ( .A(n4), .Y(n28) );
  INVXLTS U18 ( .A(n386), .Y(n29) );
  INVXLTS U19 ( .A(n386), .Y(n30) );
  INVXLTS U20 ( .A(n39), .Y(n31) );
  INVXLTS U21 ( .A(n31), .Y(n32) );
  INVXLTS U22 ( .A(n31), .Y(n33) );
  INVXLTS U23 ( .A(n54), .Y(n34) );
  INVXLTS U24 ( .A(n34), .Y(n35) );
  INVXLTS U25 ( .A(n34), .Y(n36) );
  INVXLTS U26 ( .A(n407), .Y(n37) );
  INVXLTS U27 ( .A(n37), .Y(n38) );
  INVXLTS U28 ( .A(n37), .Y(n39) );
  INVXLTS U29 ( .A(n406), .Y(n40) );
  INVXLTS U30 ( .A(n40), .Y(n41) );
  INVXLTS U31 ( .A(n40), .Y(n42) );
  INVXLTS U32 ( .A(n34), .Y(n43) );
  INVXLTS U33 ( .A(n31), .Y(n44) );
  INVXLTS U34 ( .A(n379), .Y(n45) );
  INVXLTS U35 ( .A(n380), .Y(n46) );
  INVXLTS U36 ( .A(n37), .Y(n47) );
  INVXLTS U37 ( .A(n381), .Y(n48) );
  INVXLTS U38 ( .A(n380), .Y(n49) );
  INVXLTS U39 ( .A(n380), .Y(n50) );
  INVXLTS U40 ( .A(n379), .Y(n51) );
  INVXLTS U41 ( .A(n37), .Y(n52) );
  INVXLTS U42 ( .A(n31), .Y(n53) );
  INVXLTS U43 ( .A(n383), .Y(n54) );
  INVXLTS U44 ( .A(n383), .Y(n55) );
  INVXLTS U45 ( .A(n384), .Y(n56) );
  INVXLTS U46 ( .A(n382), .Y(n57) );
  INVXLTS U47 ( .A(n384), .Y(n58) );
  INVXLTS U48 ( .A(n382), .Y(n59) );
  CLKINVX1TS U49 ( .A(n382), .Y(n60) );
  INVXLTS U50 ( .A(reset), .Y(n61) );
  INVXLTS U51 ( .A(n61), .Y(n62) );
  INVXLTS U52 ( .A(n61), .Y(n63) );
  INVX2TS U53 ( .A(n61), .Y(n64) );
  INVX2TS U54 ( .A(n66), .Y(n67) );
  INVX2TS U55 ( .A(n66), .Y(n68) );
  INVX2TS U56 ( .A(n66), .Y(n69) );
  INVX2TS U57 ( .A(n70), .Y(n71) );
  INVX2TS U58 ( .A(n70), .Y(n72) );
  INVX2TS U59 ( .A(n70), .Y(n73) );
  INVX2TS U60 ( .A(n74), .Y(n75) );
  INVX2TS U61 ( .A(n74), .Y(n76) );
  INVX2TS U62 ( .A(n74), .Y(n77) );
  INVX2TS U63 ( .A(n78), .Y(n79) );
  INVX2TS U64 ( .A(n78), .Y(n80) );
  INVX2TS U65 ( .A(n78), .Y(n81) );
  INVX2TS U66 ( .A(n82), .Y(n83) );
  INVX2TS U67 ( .A(n82), .Y(n84) );
  INVX2TS U68 ( .A(n82), .Y(n85) );
  INVX2TS U69 ( .A(n86), .Y(n87) );
  INVX2TS U70 ( .A(n86), .Y(n88) );
  INVX2TS U71 ( .A(n86), .Y(n89) );
  CLKBUFX2TS U72 ( .A(n1), .Y(n90) );
  CLKBUFX2TS U73 ( .A(n1), .Y(n91) );
  CLKBUFX2TS U74 ( .A(n1), .Y(n92) );
  CLKBUFX2TS U75 ( .A(n2), .Y(n93) );
  CLKBUFX2TS U76 ( .A(n2), .Y(n94) );
  CLKBUFX2TS U77 ( .A(n2), .Y(n95) );
  INVX2TS U78 ( .A(n96), .Y(n97) );
  INVX2TS U79 ( .A(n96), .Y(n98) );
  INVX2TS U80 ( .A(n96), .Y(n99) );
  INVX2TS U81 ( .A(n100), .Y(n101) );
  INVX2TS U82 ( .A(n100), .Y(n102) );
  INVX2TS U83 ( .A(n100), .Y(n103) );
  CLKBUFX2TS U84 ( .A(dataInBuffer_EAST[30]), .Y(n307) );
  CLKBUFX2TS U85 ( .A(dataInBuffer_EAST[28]), .Y(n303) );
  CLKBUFX2TS U86 ( .A(dataInBuffer_EAST[27]), .Y(n301) );
  CLKBUFX2TS U87 ( .A(dataInBuffer_EAST[26]), .Y(n299) );
  CLKBUFX2TS U88 ( .A(dataInBuffer_EAST[25]), .Y(n297) );
  CLKBUFX2TS U89 ( .A(dataInBuffer_EAST[24]), .Y(n295) );
  CLKBUFX2TS U90 ( .A(dataInBuffer_EAST[23]), .Y(n293) );
  CLKBUFX2TS U91 ( .A(dataInBuffer_EAST[18]), .Y(n283) );
  CLKBUFX2TS U92 ( .A(dataInBuffer_EAST[13]), .Y(n273) );
  CLKBUFX2TS U93 ( .A(dataInBuffer_EAST[9]), .Y(n265) );
  CLKBUFX2TS U94 ( .A(dataInBuffer_EAST[7]), .Y(n261) );
  CLKBUFX2TS U95 ( .A(dataInBuffer_EAST[5]), .Y(n257) );
  CLKBUFX2TS U96 ( .A(dataInBuffer_EAST[4]), .Y(n255) );
  CLKBUFX2TS U97 ( .A(dataInBuffer_EAST[2]), .Y(n251) );
  CLKBUFX2TS U98 ( .A(dataInBuffer_EAST[31]), .Y(n309) );
  CLKBUFX2TS U99 ( .A(dataInBuffer_EAST[29]), .Y(n305) );
  CLKBUFX2TS U100 ( .A(dataInBuffer_EAST[22]), .Y(n291) );
  CLKBUFX2TS U101 ( .A(dataInBuffer_EAST[21]), .Y(n289) );
  CLKBUFX2TS U102 ( .A(dataInBuffer_EAST[20]), .Y(n287) );
  CLKBUFX2TS U103 ( .A(dataInBuffer_EAST[19]), .Y(n285) );
  CLKBUFX2TS U104 ( .A(dataInBuffer_EAST[16]), .Y(n279) );
  CLKBUFX2TS U105 ( .A(dataInBuffer_EAST[12]), .Y(n271) );
  CLKBUFX2TS U106 ( .A(dataInBuffer_EAST[11]), .Y(n269) );
  CLKBUFX2TS U107 ( .A(dataInBuffer_EAST[10]), .Y(n267) );
  CLKBUFX2TS U108 ( .A(dataInBuffer_EAST[8]), .Y(n263) );
  CLKBUFX2TS U109 ( .A(dataInBuffer_EAST[6]), .Y(n259) );
  CLKBUFX2TS U110 ( .A(dataInBuffer_EAST[1]), .Y(n249) );
  CLKBUFX2TS U111 ( .A(dataInBuffer_EAST[0]), .Y(n247) );
  CLKBUFX2TS U112 ( .A(dataInBuffer_EAST[17]), .Y(n281) );
  CLKBUFX2TS U113 ( .A(dataInBuffer_EAST[15]), .Y(n277) );
  CLKBUFX2TS U114 ( .A(dataInBuffer_EAST[14]), .Y(n275) );
  CLKBUFX2TS U115 ( .A(dataInBuffer_EAST[3]), .Y(n253) );
  CLKBUFX2TS U116 ( .A(destinationAddressInBuffer_EAST[7]), .Y(n111) );
  CLKBUFX2TS U117 ( .A(destinationAddressInBuffer_EAST[6]), .Y(n110) );
  CLKBUFX2TS U118 ( .A(destinationAddressInBuffer_EAST[2]), .Y(n106) );
  CLKBUFX2TS U119 ( .A(destinationAddressInBuffer_EAST[5]), .Y(n109) );
  CLKBUFX2TS U120 ( .A(destinationAddressInBuffer_EAST[4]), .Y(n108) );
  CLKBUFX2TS U121 ( .A(destinationAddressInBuffer_EAST[3]), .Y(n107) );
  CLKBUFX2TS U122 ( .A(destinationAddressInBuffer_EAST[1]), .Y(n105) );
  CLKBUFX2TS U123 ( .A(destinationAddressInBuffer_EAST[0]), .Y(n104) );
  CLKBUFX2TS U124 ( .A(requesterAddressInBuffer_WEST[3]), .Y(n135) );
  CLKBUFX2TS U125 ( .A(requesterAddressInBuffer_WEST[2]), .Y(n133) );
  CLKBUFX2TS U126 ( .A(requesterAddressInBuffer_WEST[1]), .Y(n131) );
  CLKBUFX2TS U127 ( .A(requesterAddressInBuffer_WEST[0]), .Y(n129) );
  CLKBUFX2TS U128 ( .A(requesterAddressInBuffer_WEST[5]), .Y(n139) );
  CLKBUFX2TS U129 ( .A(requesterAddressInBuffer_WEST[4]), .Y(n137) );
  CLKBUFX2TS U130 ( .A(requesterAddressInBuffer_EAST[4]), .Y(n188) );
  CLKBUFX2TS U131 ( .A(requesterAddressInBuffer_EAST[1]), .Y(n185) );
  CLKBUFX2TS U132 ( .A(requesterAddressInBuffer_EAST[0]), .Y(n184) );
  CLKBUFX2TS U133 ( .A(requesterAddressInBuffer_EAST[5]), .Y(n189) );
  CLKBUFX2TS U134 ( .A(requesterAddressInBuffer_EAST[3]), .Y(n187) );
  CLKBUFX2TS U135 ( .A(requesterAddressInBuffer_EAST[2]), .Y(n186) );
  CLKBUFX2TS U136 ( .A(destinationAddressInBuffer_WEST[5]), .Y(n117) );
  CLKBUFX2TS U137 ( .A(destinationAddressInBuffer_WEST[4]), .Y(n116) );
  CLKBUFX2TS U138 ( .A(destinationAddressInBuffer_WEST[3]), .Y(n115) );
  CLKBUFX2TS U139 ( .A(destinationAddressInBuffer_WEST[2]), .Y(n114) );
  CLKBUFX2TS U140 ( .A(destinationAddressInBuffer_WEST[1]), .Y(n113) );
  CLKBUFX2TS U141 ( .A(destinationAddressInBuffer_WEST[0]), .Y(n112) );
  CLKBUFX2TS U142 ( .A(dataInBuffer_WEST[30]), .Y(n245) );
  CLKBUFX2TS U143 ( .A(dataInBuffer_WEST[28]), .Y(n243) );
  CLKBUFX2TS U144 ( .A(dataInBuffer_WEST[27]), .Y(n242) );
  CLKBUFX2TS U145 ( .A(dataInBuffer_WEST[26]), .Y(n241) );
  CLKBUFX2TS U146 ( .A(dataInBuffer_WEST[25]), .Y(n240) );
  CLKBUFX2TS U147 ( .A(dataInBuffer_WEST[24]), .Y(n239) );
  CLKBUFX2TS U148 ( .A(dataInBuffer_WEST[23]), .Y(n238) );
  CLKBUFX2TS U149 ( .A(dataInBuffer_WEST[18]), .Y(n233) );
  CLKBUFX2TS U150 ( .A(dataInBuffer_WEST[13]), .Y(n228) );
  CLKBUFX2TS U151 ( .A(dataInBuffer_WEST[9]), .Y(n224) );
  CLKBUFX2TS U152 ( .A(dataInBuffer_WEST[7]), .Y(n222) );
  CLKBUFX2TS U153 ( .A(dataInBuffer_WEST[5]), .Y(n220) );
  CLKBUFX2TS U154 ( .A(dataInBuffer_WEST[4]), .Y(n219) );
  CLKBUFX2TS U155 ( .A(dataInBuffer_WEST[2]), .Y(n217) );
  CLKBUFX2TS U156 ( .A(dataInBuffer_WEST[31]), .Y(n246) );
  CLKBUFX2TS U157 ( .A(dataInBuffer_WEST[29]), .Y(n244) );
  CLKBUFX2TS U158 ( .A(dataInBuffer_WEST[22]), .Y(n237) );
  CLKBUFX2TS U159 ( .A(dataInBuffer_WEST[21]), .Y(n236) );
  CLKBUFX2TS U160 ( .A(dataInBuffer_WEST[20]), .Y(n235) );
  CLKBUFX2TS U161 ( .A(dataInBuffer_WEST[19]), .Y(n234) );
  CLKBUFX2TS U162 ( .A(dataInBuffer_WEST[16]), .Y(n231) );
  CLKBUFX2TS U163 ( .A(dataInBuffer_WEST[12]), .Y(n227) );
  CLKBUFX2TS U164 ( .A(dataInBuffer_WEST[11]), .Y(n226) );
  CLKBUFX2TS U165 ( .A(dataInBuffer_WEST[10]), .Y(n225) );
  CLKBUFX2TS U166 ( .A(dataInBuffer_WEST[8]), .Y(n223) );
  CLKBUFX2TS U167 ( .A(dataInBuffer_WEST[6]), .Y(n221) );
  CLKBUFX2TS U168 ( .A(dataInBuffer_WEST[1]), .Y(n216) );
  CLKBUFX2TS U169 ( .A(dataInBuffer_WEST[0]), .Y(n215) );
  CLKBUFX2TS U170 ( .A(dataInBuffer_WEST[17]), .Y(n232) );
  CLKBUFX2TS U171 ( .A(dataInBuffer_WEST[15]), .Y(n230) );
  CLKBUFX2TS U172 ( .A(dataInBuffer_WEST[14]), .Y(n229) );
  CLKBUFX2TS U173 ( .A(dataInBuffer_WEST[3]), .Y(n218) );
  INVX2TS U174 ( .A(n387), .Y(n386) );
  INVX2TS U175 ( .A(n394), .Y(n379) );
  INVX2TS U176 ( .A(n393), .Y(n380) );
  INVX2TS U177 ( .A(n392), .Y(n381) );
  INVX2TS U178 ( .A(n388), .Y(n385) );
  INVX2TS U179 ( .A(n390), .Y(n383) );
  INVX2TS U180 ( .A(n391), .Y(n382) );
  INVX2TS U181 ( .A(n389), .Y(n384) );
  CLKBUFX2TS U182 ( .A(n401), .Y(n400) );
  CLKBUFX2TS U183 ( .A(n401), .Y(n399) );
  CLKBUFX2TS U184 ( .A(n402), .Y(n398) );
  CLKBUFX2TS U185 ( .A(n402), .Y(n397) );
  CLKBUFX2TS U186 ( .A(n402), .Y(n396) );
  CLKBUFX2TS U187 ( .A(n402), .Y(n395) );
  CLKBUFX2TS U188 ( .A(n403), .Y(n394) );
  CLKBUFX2TS U189 ( .A(n403), .Y(n393) );
  CLKBUFX2TS U190 ( .A(n403), .Y(n392) );
  CLKBUFX2TS U191 ( .A(n404), .Y(n388) );
  CLKBUFX2TS U192 ( .A(n404), .Y(n387) );
  CLKBUFX2TS U193 ( .A(n403), .Y(n391) );
  CLKBUFX2TS U194 ( .A(n404), .Y(n390) );
  CLKBUFX2TS U195 ( .A(n404), .Y(n389) );
  CLKBUFX2TS U196 ( .A(n406), .Y(n401) );
  CLKBUFX2TS U197 ( .A(n406), .Y(n402) );
  CLKBUFX2TS U198 ( .A(n405), .Y(n403) );
  CLKBUFX2TS U199 ( .A(n405), .Y(n404) );
  CLKBUFX2TS U200 ( .A(n407), .Y(n406) );
  CLKBUFX2TS U201 ( .A(n408), .Y(n405) );
  CLKBUFX2TS U202 ( .A(n62), .Y(n408) );
  CLKBUFX2TS U203 ( .A(n63), .Y(n407) );
  CLKBUFX2TS U204 ( .A(destinationAddressInBuffer_SOUTH[7]), .Y(n202) );
  CLKBUFX2TS U205 ( .A(destinationAddressInBuffer_SOUTH[6]), .Y(n201) );
  CLKBUFX2TS U206 ( .A(dataInBuffer_EAST[0]), .Y(n248) );
  CLKBUFX2TS U207 ( .A(dataInBuffer_EAST[1]), .Y(n250) );
  CLKBUFX2TS U208 ( .A(dataInBuffer_EAST[2]), .Y(n252) );
  CLKBUFX2TS U209 ( .A(dataInBuffer_EAST[3]), .Y(n254) );
  CLKBUFX2TS U210 ( .A(dataInBuffer_EAST[4]), .Y(n256) );
  CLKBUFX2TS U211 ( .A(dataInBuffer_EAST[5]), .Y(n258) );
  CLKBUFX2TS U212 ( .A(dataInBuffer_EAST[6]), .Y(n260) );
  CLKBUFX2TS U213 ( .A(dataInBuffer_EAST[7]), .Y(n262) );
  CLKBUFX2TS U214 ( .A(dataInBuffer_EAST[8]), .Y(n264) );
  CLKBUFX2TS U215 ( .A(dataInBuffer_EAST[9]), .Y(n266) );
  CLKBUFX2TS U216 ( .A(dataInBuffer_EAST[10]), .Y(n268) );
  CLKBUFX2TS U217 ( .A(dataInBuffer_EAST[11]), .Y(n270) );
  CLKBUFX2TS U218 ( .A(dataInBuffer_EAST[12]), .Y(n272) );
  CLKBUFX2TS U219 ( .A(dataInBuffer_EAST[13]), .Y(n274) );
  CLKBUFX2TS U220 ( .A(dataInBuffer_EAST[14]), .Y(n276) );
  CLKBUFX2TS U221 ( .A(dataInBuffer_EAST[15]), .Y(n278) );
  CLKBUFX2TS U222 ( .A(dataInBuffer_EAST[16]), .Y(n280) );
  CLKBUFX2TS U223 ( .A(dataInBuffer_EAST[17]), .Y(n282) );
  CLKBUFX2TS U224 ( .A(dataInBuffer_EAST[18]), .Y(n284) );
  CLKBUFX2TS U225 ( .A(dataInBuffer_EAST[19]), .Y(n286) );
  CLKBUFX2TS U226 ( .A(dataInBuffer_EAST[20]), .Y(n288) );
  CLKBUFX2TS U227 ( .A(dataInBuffer_EAST[21]), .Y(n290) );
  CLKBUFX2TS U228 ( .A(dataInBuffer_EAST[22]), .Y(n292) );
  CLKBUFX2TS U229 ( .A(dataInBuffer_EAST[23]), .Y(n294) );
  CLKBUFX2TS U230 ( .A(dataInBuffer_EAST[24]), .Y(n296) );
  CLKBUFX2TS U231 ( .A(dataInBuffer_EAST[25]), .Y(n298) );
  CLKBUFX2TS U232 ( .A(dataInBuffer_EAST[26]), .Y(n300) );
  CLKBUFX2TS U233 ( .A(dataInBuffer_EAST[27]), .Y(n302) );
  CLKBUFX2TS U234 ( .A(dataInBuffer_EAST[28]), .Y(n304) );
  CLKBUFX2TS U235 ( .A(dataInBuffer_EAST[29]), .Y(n306) );
  CLKBUFX2TS U236 ( .A(dataInBuffer_EAST[30]), .Y(n308) );
  CLKBUFX2TS U237 ( .A(dataInBuffer_EAST[31]), .Y(n310) );
  CLKBUFX2TS U238 ( .A(destinationAddressInBuffer_WEST[13]), .Y(n127) );
  CLKBUFX2TS U239 ( .A(destinationAddressInBuffer_WEST[11]), .Y(n125) );
  CLKBUFX2TS U240 ( .A(destinationAddressInBuffer_WEST[9]), .Y(n122) );
  CLKBUFX2TS U241 ( .A(destinationAddressInBuffer_WEST[12]), .Y(n126) );
  CLKBUFX2TS U242 ( .A(destinationAddressInBuffer_WEST[10]), .Y(n124) );
  CLKBUFX2TS U243 ( .A(requesterAddressInBuffer_SOUTH[4]), .Y(n375) );
  CLKBUFX2TS U244 ( .A(requesterAddressInBuffer_SOUTH[1]), .Y(n369) );
  CLKBUFX2TS U245 ( .A(requesterAddressInBuffer_SOUTH[5]), .Y(n377) );
  CLKBUFX2TS U246 ( .A(requesterAddressInBuffer_SOUTH[3]), .Y(n373) );
  CLKBUFX2TS U247 ( .A(requesterAddressInBuffer_SOUTH[2]), .Y(n371) );
  CLKBUFX2TS U248 ( .A(destinationAddressInBuffer_SOUTH[4]), .Y(n198) );
  CLKBUFX2TS U249 ( .A(destinationAddressInBuffer_SOUTH[3]), .Y(n196) );
  CLKBUFX2TS U250 ( .A(destinationAddressInBuffer_SOUTH[0]), .Y(n192) );
  CLKBUFX2TS U251 ( .A(dataInBuffer_SOUTH[30]), .Y(n364) );
  CLKBUFX2TS U252 ( .A(dataInBuffer_SOUTH[28]), .Y(n360) );
  CLKBUFX2TS U253 ( .A(dataInBuffer_SOUTH[27]), .Y(n358) );
  CLKBUFX2TS U254 ( .A(dataInBuffer_SOUTH[25]), .Y(n355) );
  CLKBUFX2TS U255 ( .A(dataInBuffer_SOUTH[24]), .Y(n353) );
  CLKBUFX2TS U256 ( .A(dataInBuffer_SOUTH[18]), .Y(n343) );
  CLKBUFX2TS U257 ( .A(dataInBuffer_SOUTH[13]), .Y(n335) );
  CLKBUFX2TS U258 ( .A(dataInBuffer_SOUTH[7]), .Y(n324) );
  CLKBUFX2TS U259 ( .A(dataInBuffer_SOUTH[5]), .Y(n320) );
  CLKBUFX2TS U260 ( .A(dataInBuffer_SOUTH[2]), .Y(n315) );
  CLKBUFX2TS U261 ( .A(dataInBuffer_SOUTH[31]), .Y(n366) );
  CLKBUFX2TS U262 ( .A(dataInBuffer_SOUTH[29]), .Y(n362) );
  CLKBUFX2TS U263 ( .A(dataInBuffer_SOUTH[22]), .Y(n350) );
  CLKBUFX2TS U264 ( .A(dataInBuffer_SOUTH[21]), .Y(n348) );
  CLKBUFX2TS U265 ( .A(dataInBuffer_SOUTH[19]), .Y(n345) );
  CLKBUFX2TS U266 ( .A(dataInBuffer_SOUTH[12]), .Y(n333) );
  CLKBUFX2TS U267 ( .A(dataInBuffer_SOUTH[11]), .Y(n331) );
  CLKBUFX2TS U268 ( .A(dataInBuffer_SOUTH[10]), .Y(n329) );
  CLKBUFX2TS U269 ( .A(dataInBuffer_SOUTH[8]), .Y(n326) );
  CLKBUFX2TS U270 ( .A(dataInBuffer_SOUTH[6]), .Y(n322) );
  CLKBUFX2TS U271 ( .A(dataInBuffer_SOUTH[1]), .Y(n313) );
  CLKBUFX2TS U272 ( .A(dataInBuffer_SOUTH[0]), .Y(n311) );
  CLKBUFX2TS U273 ( .A(dataInBuffer_SOUTH[17]), .Y(n341) );
  CLKBUFX2TS U274 ( .A(dataInBuffer_SOUTH[15]), .Y(n338) );
  CLKBUFX2TS U275 ( .A(dataInBuffer_SOUTH[3]), .Y(n317) );
  CLKBUFX2TS U276 ( .A(destinationAddressInBuffer_WEST[9]), .Y(n121) );
  CLKBUFX2TS U277 ( .A(destinationAddressInBuffer_WEST[7]), .Y(n119) );
  CLKBUFX2TS U278 ( .A(destinationAddressInBuffer_WEST[10]), .Y(n123) );
  CLKBUFX2TS U279 ( .A(destinationAddressInBuffer_WEST[8]), .Y(n120) );
  CLKBUFX2TS U280 ( .A(destinationAddressInBuffer_WEST[6]), .Y(n118) );
  CLKBUFX2TS U281 ( .A(requesterAddressInBuffer_SOUTH[0]), .Y(n368) );
  CLKBUFX2TS U282 ( .A(requesterAddressInBuffer_SOUTH[1]), .Y(n370) );
  CLKBUFX2TS U283 ( .A(requesterAddressInBuffer_SOUTH[2]), .Y(n372) );
  CLKBUFX2TS U284 ( .A(requesterAddressInBuffer_SOUTH[3]), .Y(n374) );
  CLKBUFX2TS U285 ( .A(requesterAddressInBuffer_SOUTH[4]), .Y(n376) );
  CLKBUFX2TS U286 ( .A(requesterAddressInBuffer_SOUTH[5]), .Y(n378) );
  CLKBUFX2TS U287 ( .A(dataInBuffer_SOUTH[0]), .Y(n312) );
  CLKBUFX2TS U288 ( .A(dataInBuffer_SOUTH[1]), .Y(n314) );
  CLKBUFX2TS U289 ( .A(dataInBuffer_SOUTH[2]), .Y(n316) );
  CLKBUFX2TS U290 ( .A(dataInBuffer_SOUTH[3]), .Y(n318) );
  CLKBUFX2TS U291 ( .A(dataInBuffer_SOUTH[4]), .Y(n319) );
  CLKBUFX2TS U292 ( .A(dataInBuffer_SOUTH[5]), .Y(n321) );
  CLKBUFX2TS U293 ( .A(dataInBuffer_SOUTH[6]), .Y(n323) );
  CLKBUFX2TS U294 ( .A(dataInBuffer_SOUTH[7]), .Y(n325) );
  CLKBUFX2TS U295 ( .A(dataInBuffer_SOUTH[8]), .Y(n327) );
  CLKBUFX2TS U296 ( .A(dataInBuffer_SOUTH[9]), .Y(n328) );
  CLKBUFX2TS U297 ( .A(dataInBuffer_SOUTH[10]), .Y(n330) );
  CLKBUFX2TS U298 ( .A(dataInBuffer_SOUTH[11]), .Y(n332) );
  CLKBUFX2TS U299 ( .A(dataInBuffer_SOUTH[12]), .Y(n334) );
  CLKBUFX2TS U300 ( .A(dataInBuffer_SOUTH[13]), .Y(n336) );
  CLKBUFX2TS U301 ( .A(dataInBuffer_SOUTH[14]), .Y(n337) );
  CLKBUFX2TS U302 ( .A(dataInBuffer_SOUTH[15]), .Y(n339) );
  CLKBUFX2TS U303 ( .A(dataInBuffer_SOUTH[16]), .Y(n340) );
  CLKBUFX2TS U304 ( .A(dataInBuffer_SOUTH[17]), .Y(n342) );
  CLKBUFX2TS U305 ( .A(dataInBuffer_SOUTH[18]), .Y(n344) );
  CLKBUFX2TS U306 ( .A(dataInBuffer_SOUTH[19]), .Y(n346) );
  CLKBUFX2TS U307 ( .A(dataInBuffer_SOUTH[20]), .Y(n347) );
  CLKBUFX2TS U308 ( .A(dataInBuffer_SOUTH[21]), .Y(n349) );
  CLKBUFX2TS U309 ( .A(dataInBuffer_SOUTH[22]), .Y(n351) );
  CLKBUFX2TS U310 ( .A(dataInBuffer_SOUTH[23]), .Y(n352) );
  CLKBUFX2TS U311 ( .A(dataInBuffer_SOUTH[24]), .Y(n354) );
  CLKBUFX2TS U312 ( .A(dataInBuffer_SOUTH[25]), .Y(n356) );
  CLKBUFX2TS U313 ( .A(dataInBuffer_SOUTH[26]), .Y(n357) );
  CLKBUFX2TS U314 ( .A(dataInBuffer_SOUTH[27]), .Y(n359) );
  CLKBUFX2TS U315 ( .A(dataInBuffer_SOUTH[28]), .Y(n361) );
  CLKBUFX2TS U316 ( .A(dataInBuffer_SOUTH[29]), .Y(n363) );
  CLKBUFX2TS U317 ( .A(dataInBuffer_SOUTH[30]), .Y(n365) );
  CLKBUFX2TS U318 ( .A(dataInBuffer_SOUTH[31]), .Y(n367) );
  CLKBUFX2TS U319 ( .A(destinationAddressInBuffer_SOUTH[0]), .Y(n193) );
  CLKBUFX2TS U320 ( .A(destinationAddressInBuffer_SOUTH[1]), .Y(n194) );
  CLKBUFX2TS U321 ( .A(destinationAddressInBuffer_SOUTH[2]), .Y(n195) );
  CLKBUFX2TS U322 ( .A(destinationAddressInBuffer_SOUTH[3]), .Y(n197) );
  CLKBUFX2TS U323 ( .A(destinationAddressInBuffer_SOUTH[4]), .Y(n199) );
  CLKBUFX2TS U324 ( .A(destinationAddressInBuffer_SOUTH[5]), .Y(n200) );
  CLKBUFX2TS U325 ( .A(writeInBuffer_SOUTH), .Y(n190) );
  CLKBUFX2TS U326 ( .A(destinationAddressInBuffer_SOUTH[13]), .Y(n214) );
  CLKBUFX2TS U327 ( .A(destinationAddressInBuffer_SOUTH[11]), .Y(n210) );
  CLKBUFX2TS U328 ( .A(destinationAddressInBuffer_SOUTH[9]), .Y(n206) );
  CLKBUFX2TS U329 ( .A(destinationAddressInBuffer_SOUTH[12]), .Y(n212) );
  CLKBUFX2TS U330 ( .A(destinationAddressInBuffer_SOUTH[10]), .Y(n208) );
  CLKBUFX2TS U331 ( .A(destinationAddressInBuffer_SOUTH[8]), .Y(n204) );
  CLKBUFX2TS U332 ( .A(writeInBuffer_SOUTH), .Y(n191) );
  CLKBUFX2TS U333 ( .A(destinationAddressInBuffer_SOUTH[13]), .Y(n213) );
  CLKBUFX2TS U334 ( .A(destinationAddressInBuffer_SOUTH[11]), .Y(n209) );
  CLKBUFX2TS U335 ( .A(destinationAddressInBuffer_SOUTH[9]), .Y(n205) );
  CLKBUFX2TS U336 ( .A(destinationAddressInBuffer_SOUTH[12]), .Y(n211) );
  CLKBUFX2TS U337 ( .A(destinationAddressInBuffer_SOUTH[10]), .Y(n207) );
  CLKBUFX2TS U338 ( .A(destinationAddressInBuffer_SOUTH[8]), .Y(n203) );
  CLKBUFX2TS U339 ( .A(requesterAddressInBuffer_WEST[0]), .Y(n128) );
  CLKBUFX2TS U340 ( .A(requesterAddressInBuffer_WEST[1]), .Y(n130) );
  CLKBUFX2TS U341 ( .A(requesterAddressInBuffer_WEST[2]), .Y(n132) );
  CLKBUFX2TS U342 ( .A(requesterAddressInBuffer_WEST[3]), .Y(n134) );
  CLKBUFX2TS U343 ( .A(requesterAddressInBuffer_WEST[4]), .Y(n136) );
  CLKBUFX2TS U344 ( .A(requesterAddressInBuffer_WEST[5]), .Y(n138) );
  CLKBUFX2TS U345 ( .A(requesterAddressInBuffer_NORTH[4]), .Y(n150) );
  CLKBUFX2TS U346 ( .A(requesterAddressInBuffer_NORTH[1]), .Y(n147) );
  CLKBUFX2TS U347 ( .A(requesterAddressInBuffer_NORTH[0]), .Y(n146) );
  CLKBUFX2TS U348 ( .A(requesterAddressInBuffer_NORTH[3]), .Y(n149) );
  CLKBUFX2TS U349 ( .A(requesterAddressInBuffer_NORTH[2]), .Y(n148) );
  CLKBUFX2TS U350 ( .A(destinationAddressInBuffer_NORTH_4), .Y(n144) );
  CLKBUFX2TS U351 ( .A(destinationAddressInBuffer_NORTH_2), .Y(n142) );
  CLKBUFX2TS U352 ( .A(destinationAddressInBuffer_NORTH_1), .Y(n141) );
  CLKBUFX2TS U353 ( .A(dataInBuffer_NORTH[30]), .Y(n182) );
  CLKBUFX2TS U354 ( .A(dataInBuffer_NORTH[28]), .Y(n180) );
  CLKBUFX2TS U355 ( .A(dataInBuffer_NORTH[26]), .Y(n178) );
  CLKBUFX2TS U356 ( .A(dataInBuffer_NORTH[25]), .Y(n177) );
  CLKBUFX2TS U357 ( .A(dataInBuffer_NORTH[24]), .Y(n176) );
  CLKBUFX2TS U358 ( .A(dataInBuffer_NORTH[23]), .Y(n175) );
  CLKBUFX2TS U359 ( .A(dataInBuffer_NORTH[18]), .Y(n170) );
  CLKBUFX2TS U360 ( .A(dataInBuffer_NORTH[13]), .Y(n165) );
  CLKBUFX2TS U361 ( .A(dataInBuffer_NORTH[7]), .Y(n159) );
  CLKBUFX2TS U362 ( .A(dataInBuffer_NORTH[4]), .Y(n156) );
  CLKBUFX2TS U363 ( .A(dataInBuffer_NORTH[2]), .Y(n154) );
  CLKBUFX2TS U364 ( .A(dataInBuffer_NORTH[29]), .Y(n181) );
  CLKBUFX2TS U365 ( .A(dataInBuffer_NORTH[22]), .Y(n174) );
  CLKBUFX2TS U366 ( .A(dataInBuffer_NORTH[21]), .Y(n173) );
  CLKBUFX2TS U367 ( .A(dataInBuffer_NORTH[20]), .Y(n172) );
  CLKBUFX2TS U368 ( .A(dataInBuffer_NORTH[19]), .Y(n171) );
  CLKBUFX2TS U369 ( .A(dataInBuffer_NORTH[16]), .Y(n168) );
  CLKBUFX2TS U370 ( .A(dataInBuffer_NORTH[12]), .Y(n164) );
  CLKBUFX2TS U371 ( .A(dataInBuffer_NORTH[11]), .Y(n163) );
  CLKBUFX2TS U372 ( .A(dataInBuffer_NORTH[10]), .Y(n162) );
  CLKBUFX2TS U373 ( .A(dataInBuffer_NORTH[8]), .Y(n160) );
  CLKBUFX2TS U374 ( .A(dataInBuffer_NORTH[6]), .Y(n158) );
  CLKBUFX2TS U375 ( .A(dataInBuffer_NORTH[0]), .Y(n152) );
  CLKBUFX2TS U376 ( .A(dataInBuffer_NORTH[17]), .Y(n169) );
  CLKBUFX2TS U377 ( .A(dataInBuffer_NORTH[15]), .Y(n167) );
  CLKBUFX2TS U378 ( .A(dataInBuffer_NORTH[14]), .Y(n166) );
  CLKBUFX2TS U379 ( .A(dataInBuffer_NORTH[3]), .Y(n155) );
  CLKBUFX2TS U380 ( .A(destinationAddressInBuffer_NORTH_0), .Y(n140) );
  CLKBUFX2TS U381 ( .A(destinationAddressInBuffer_NORTH_3), .Y(n143) );
  CLKBUFX2TS U382 ( .A(dataInBuffer_NORTH[9]), .Y(n161) );
  CLKBUFX2TS U383 ( .A(dataInBuffer_NORTH[5]), .Y(n157) );
  CLKBUFX2TS U384 ( .A(dataInBuffer_NORTH[1]), .Y(n153) );
  CLKBUFX2TS U385 ( .A(requesterAddressInBuffer_NORTH[5]), .Y(n151) );
  CLKBUFX2TS U386 ( .A(destinationAddressInBuffer_NORTH_5), .Y(n145) );
  CLKBUFX2TS U387 ( .A(dataInBuffer_NORTH[27]), .Y(n179) );
  CLKBUFX2TS U388 ( .A(dataInBuffer_NORTH[31]), .Y(n183) );
endmodule


module Node ( clk, reset, localRouterAddress, destinationAddressIn_NORTH, 
        requesterAddressIn_NORTH, readIn_NORTH, writeIn_NORTH, dataIn_NORTH, 
        destinationAddressOut_NORTH, requesterAddressOut_NORTH, readOut_NORTH, 
        writeOut_NORTH, dataOut_NORTH, destinationAddressIn_SOUTH, 
        requesterAddressIn_SOUTH, readIn_SOUTH, writeIn_SOUTH, dataIn_SOUTH, 
        destinationAddressOut_SOUTH, requesterAddressOut_SOUTH, readOut_SOUTH, 
        writeOut_SOUTH, dataOut_SOUTH, destinationAddressIn_EAST, 
        requesterAddressIn_EAST, readIn_EAST, writeIn_EAST, dataIn_EAST, 
        destinationAddressOut_EAST, requesterAddressOut_EAST, readOut_EAST, 
        writeOut_EAST, dataOut_EAST, destinationAddressIn_WEST, 
        requesterAddressIn_WEST, readIn_WEST, writeIn_WEST, dataIn_WEST, 
        destinationAddressOut_WEST, requesterAddressOut_WEST, readOut_WEST, 
        writeOut_WEST, dataOut_WEST );
  input [5:0] localRouterAddress;
  input [13:0] destinationAddressIn_NORTH;
  input [5:0] requesterAddressIn_NORTH;
  input [31:0] dataIn_NORTH;
  output [13:0] destinationAddressOut_NORTH;
  output [5:0] requesterAddressOut_NORTH;
  output [31:0] dataOut_NORTH;
  input [13:0] destinationAddressIn_SOUTH;
  input [5:0] requesterAddressIn_SOUTH;
  input [31:0] dataIn_SOUTH;
  output [13:0] destinationAddressOut_SOUTH;
  output [5:0] requesterAddressOut_SOUTH;
  output [31:0] dataOut_SOUTH;
  input [13:0] destinationAddressIn_EAST;
  input [5:0] requesterAddressIn_EAST;
  input [31:0] dataIn_EAST;
  output [13:0] destinationAddressOut_EAST;
  output [5:0] requesterAddressOut_EAST;
  output [31:0] dataOut_EAST;
  input [13:0] destinationAddressIn_WEST;
  input [5:0] requesterAddressIn_WEST;
  input [31:0] dataIn_WEST;
  output [13:0] destinationAddressOut_WEST;
  output [5:0] requesterAddressOut_WEST;
  output [31:0] dataOut_WEST;
  input clk, reset, readIn_NORTH, writeIn_NORTH, readIn_SOUTH, writeIn_SOUTH,
         readIn_EAST, writeIn_EAST, readIn_WEST, writeIn_WEST;
  output readOut_NORTH, writeOut_NORTH, readOut_SOUTH, writeOut_SOUTH,
         readOut_EAST, writeOut_EAST, readOut_WEST, writeOut_WEST;
  wire   memWrite_A, memWrite_B, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69;
  wire   [31:0] cacheDataIn_A;
  wire   [7:0] cacheAddressIn_A;
  wire   [31:0] cacheDataOut_A;
  wire   [31:0] cacheDataIn_B;
  wire   [7:0] cacheAddressIn_B;
  wire   [31:0] cacheDataOut_B;

  router rtr ( .clk(clk), .localRouterAddress({n65, n69, n67, n45, n43, n55}), 
        .destinationAddressIn_NORTH({n9, destinationAddressIn_NORTH[12], n17, 
        n63, n53, n41, destinationAddressIn_NORTH[7:0]}), 
        .requesterAddressIn_NORTH(requesterAddressIn_NORTH), .readIn_NORTH(n33), .writeIn_NORTH(n25), .dataIn_NORTH(dataIn_NORTH), 
        .destinationAddressOut_NORTH(destinationAddressOut_NORTH), 
        .requesterAddressOut_NORTH(requesterAddressOut_NORTH), .readOut_NORTH(
        readOut_NORTH), .writeOut_NORTH(writeOut_NORTH), .dataOut_NORTH(
        dataOut_NORTH), .destinationAddressIn_SOUTH({n7, 
        destinationAddressIn_SOUTH[12], n15, n61, n51, n39, 
        destinationAddressIn_SOUTH[7:0]}), .requesterAddressIn_SOUTH(
        requesterAddressIn_SOUTH), .readIn_SOUTH(n31), .writeIn_SOUTH(n23), 
        .dataIn_SOUTH(dataIn_SOUTH), .destinationAddressOut_SOUTH(
        destinationAddressOut_SOUTH), .requesterAddressOut_SOUTH(
        requesterAddressOut_SOUTH), .readOut_SOUTH(readOut_SOUTH), 
        .writeOut_SOUTH(writeOut_SOUTH), .dataOut_SOUTH(dataOut_SOUTH), 
        .destinationAddressIn_EAST({n5, destinationAddressIn_EAST[12], n13, 
        n59, n49, n37, destinationAddressIn_EAST[7:0]}), 
        .requesterAddressIn_EAST(requesterAddressIn_EAST), .readIn_EAST(n29), 
        .writeIn_EAST(n21), .dataIn_EAST(dataIn_EAST), 
        .destinationAddressOut_EAST(destinationAddressOut_EAST), 
        .requesterAddressOut_EAST(requesterAddressOut_EAST), .readOut_EAST(
        readOut_EAST), .writeOut_EAST(writeOut_EAST), .dataOut_EAST(
        dataOut_EAST), .destinationAddressIn_WEST({n3, 
        destinationAddressIn_WEST[12], n11, n57, n47, n35, 
        destinationAddressIn_WEST[7:0]}), .requesterAddressIn_WEST(
        requesterAddressIn_WEST), .readIn_WEST(n27), .writeIn_WEST(n19), 
        .dataIn_WEST(dataIn_WEST), .destinationAddressOut_WEST(
        destinationAddressOut_WEST), .requesterAddressOut_WEST(
        requesterAddressOut_WEST), .readOut_WEST(readOut_WEST), 
        .writeOut_WEST(writeOut_WEST), .dataOut_WEST(dataOut_WEST), 
        .cacheDataIn_A(cacheDataIn_A), .cacheAddressIn_A(cacheAddressIn_A), 
        .cacheDataOut_A(cacheDataOut_A), .memWrite_A(memWrite_A), 
        .portA_writtenTo(1'b0), .cacheDataIn_B(cacheDataIn_B), 
        .cacheAddressIn_B(cacheAddressIn_B), .cacheDataOut_B(cacheDataOut_B), 
        .memWrite_B(memWrite_B), .portB_writtenTo(1'b0), .reset_BAR(n1) );
  cacheBank localCacheBank ( .clk(clk), .reset(reset), .cacheDataIn_A(
        cacheDataIn_A), .cacheAddressIn_A(cacheAddressIn_A), .memWrite_A(
        memWrite_A), .cacheDataOut_A(cacheDataOut_A), .cacheDataIn_B(
        cacheDataIn_B), .cacheAddressIn_B(cacheAddressIn_B), .memWrite_B(
        memWrite_B), .cacheDataOut_B(cacheDataOut_B) );
  INVXLTS U1 ( .A(reset), .Y(n1) );
  INVXLTS U2 ( .A(destinationAddressIn_WEST[13]), .Y(n2) );
  INVXLTS U3 ( .A(n2), .Y(n3) );
  INVXLTS U4 ( .A(destinationAddressIn_EAST[13]), .Y(n4) );
  INVXLTS U5 ( .A(n4), .Y(n5) );
  INVXLTS U6 ( .A(destinationAddressIn_SOUTH[13]), .Y(n6) );
  INVXLTS U7 ( .A(n6), .Y(n7) );
  INVXLTS U8 ( .A(destinationAddressIn_NORTH[13]), .Y(n8) );
  INVXLTS U9 ( .A(n8), .Y(n9) );
  INVXLTS U10 ( .A(destinationAddressIn_WEST[11]), .Y(n10) );
  INVXLTS U11 ( .A(n10), .Y(n11) );
  INVXLTS U12 ( .A(destinationAddressIn_EAST[11]), .Y(n12) );
  INVXLTS U13 ( .A(n12), .Y(n13) );
  INVXLTS U14 ( .A(destinationAddressIn_SOUTH[11]), .Y(n14) );
  INVXLTS U15 ( .A(n14), .Y(n15) );
  INVXLTS U16 ( .A(destinationAddressIn_NORTH[11]), .Y(n16) );
  INVXLTS U17 ( .A(n16), .Y(n17) );
  INVXLTS U18 ( .A(writeIn_WEST), .Y(n18) );
  INVXLTS U19 ( .A(n18), .Y(n19) );
  INVXLTS U20 ( .A(writeIn_EAST), .Y(n20) );
  INVXLTS U21 ( .A(n20), .Y(n21) );
  INVXLTS U22 ( .A(writeIn_SOUTH), .Y(n22) );
  INVXLTS U23 ( .A(n22), .Y(n23) );
  INVXLTS U24 ( .A(writeIn_NORTH), .Y(n24) );
  INVXLTS U25 ( .A(n24), .Y(n25) );
  INVXLTS U26 ( .A(readIn_WEST), .Y(n26) );
  INVXLTS U27 ( .A(n26), .Y(n27) );
  INVXLTS U28 ( .A(readIn_EAST), .Y(n28) );
  INVXLTS U29 ( .A(n28), .Y(n29) );
  INVXLTS U30 ( .A(readIn_SOUTH), .Y(n30) );
  INVXLTS U31 ( .A(n30), .Y(n31) );
  INVXLTS U32 ( .A(readIn_NORTH), .Y(n32) );
  INVXLTS U33 ( .A(n32), .Y(n33) );
  INVXLTS U34 ( .A(destinationAddressIn_WEST[8]), .Y(n34) );
  INVXLTS U35 ( .A(n34), .Y(n35) );
  INVXLTS U36 ( .A(destinationAddressIn_EAST[8]), .Y(n36) );
  INVXLTS U37 ( .A(n36), .Y(n37) );
  INVXLTS U38 ( .A(destinationAddressIn_SOUTH[8]), .Y(n38) );
  INVXLTS U39 ( .A(n38), .Y(n39) );
  INVXLTS U40 ( .A(destinationAddressIn_NORTH[8]), .Y(n40) );
  INVXLTS U41 ( .A(n40), .Y(n41) );
  INVXLTS U42 ( .A(localRouterAddress[1]), .Y(n42) );
  INVXLTS U43 ( .A(n42), .Y(n43) );
  INVXLTS U44 ( .A(localRouterAddress[2]), .Y(n44) );
  INVXLTS U45 ( .A(n44), .Y(n45) );
  INVXLTS U46 ( .A(destinationAddressIn_WEST[9]), .Y(n46) );
  INVXLTS U47 ( .A(n46), .Y(n47) );
  INVXLTS U48 ( .A(destinationAddressIn_EAST[9]), .Y(n48) );
  INVXLTS U49 ( .A(n48), .Y(n49) );
  INVXLTS U50 ( .A(destinationAddressIn_SOUTH[9]), .Y(n50) );
  INVXLTS U51 ( .A(n50), .Y(n51) );
  INVXLTS U52 ( .A(destinationAddressIn_NORTH[9]), .Y(n52) );
  INVXLTS U53 ( .A(n52), .Y(n53) );
  INVXLTS U54 ( .A(localRouterAddress[0]), .Y(n54) );
  INVXLTS U55 ( .A(n54), .Y(n55) );
  INVXLTS U56 ( .A(destinationAddressIn_WEST[10]), .Y(n56) );
  INVXLTS U57 ( .A(n56), .Y(n57) );
  INVXLTS U58 ( .A(destinationAddressIn_EAST[10]), .Y(n58) );
  INVXLTS U59 ( .A(n58), .Y(n59) );
  INVXLTS U60 ( .A(destinationAddressIn_SOUTH[10]), .Y(n60) );
  INVXLTS U61 ( .A(n60), .Y(n61) );
  INVXLTS U62 ( .A(destinationAddressIn_NORTH[10]), .Y(n62) );
  INVXLTS U63 ( .A(n62), .Y(n63) );
  INVXLTS U64 ( .A(localRouterAddress[5]), .Y(n64) );
  INVXLTS U65 ( .A(n64), .Y(n65) );
  INVXLTS U66 ( .A(localRouterAddress[3]), .Y(n66) );
  INVXLTS U67 ( .A(n66), .Y(n67) );
  INVXLTS U68 ( .A(localRouterAddress[4]), .Y(n68) );
  INVXLTS U69 ( .A(n68), .Y(n69) );
endmodule

